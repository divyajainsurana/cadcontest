//
// Conformal-LEC Version 19.20-d255 (16-Apr-2020)
//
module top(\s[31] ,\s[30] ,\s[29] ,\s[28] ,\s[27] ,\s[26] ,\s[25] ,\s[24] ,\s[23] ,
        \s[22] ,\s[21] ,\s[20] ,\s[19] ,\s[18] ,\s[17] ,\s[16] ,\s[15] ,\s[14] ,\s[13] ,
        \s[12] ,\s[11] ,\s[10] ,\s[9] ,\s[8] ,\s[7] ,\s[6] ,\s[5] ,\s[4] ,\s[3] ,
        \s[2] ,\s[1] ,\s[0] ,\a[31] ,\a[30] ,\a[29] ,\a[28] ,\a[27] ,\a[26] ,\a[25] ,
        \a[24] ,\a[23] ,\a[22] ,\a[21] ,\a[20] ,\a[19] ,\a[18] ,\a[17] ,\a[16] ,\a[15] ,
        \a[14] ,\a[13] ,\a[12] ,\a[11] ,\a[10] ,\a[9] ,\a[8] ,\a[7] ,\a[6] ,\a[5] ,
        \a[4] ,\a[3] ,\a[2] ,\a[1] ,\a[0] ,\b[31] ,\b[30] ,\b[29] ,\b[28] ,\b[27] ,
        \b[26] ,\b[25] ,\b[24] ,\b[23] ,\b[22] ,\b[21] ,\b[20] ,\b[19] ,\b[18] ,\b[17] ,
        \b[16] ,\b[15] ,\b[14] ,\b[13] ,\b[12] ,\b[11] ,\b[10] ,\b[9] ,\b[8] ,\b[7] ,
        \b[6] ,\b[5] ,\b[4] ,\b[3] ,\b[2] ,\b[1] ,\b[0] ,\c[31] ,\c[30] ,\c[29] ,
        \c[28] ,\c[27] ,\c[26] ,\c[25] ,\c[24] ,\c[23] ,\c[22] ,\c[21] ,\c[20] ,\c[19] ,
        \c[18] ,\c[17] ,\c[16] ,\c[15] ,\c[14] ,\c[13] ,\c[12] ,\c[11] ,\c[10] ,\c[9] ,
        \c[8] ,\c[7] ,\c[6] ,\c[5] ,\c[4] ,\c[3] ,\c[2] ,\c[1] ,\c[0] ,\d[31] ,
        \d[30] ,\d[29] ,\d[28] ,\d[27] ,\d[26] ,\d[25] ,\d[24] ,\d[23] ,\d[22] ,\d[21] ,
        \d[20] ,\d[19] ,\d[18] ,\d[17] ,\d[16] ,\d[15] ,\d[14] ,\d[13] ,\d[12] ,\d[11] ,
        \d[10] ,\d[9] ,\d[8] ,\d[7] ,\d[6] ,\d[5] ,\d[4] ,\d[3] ,\d[2] ,\d[1] ,
        \d[0] ,\o[31] ,\o[30] ,\o[29] ,\o[28] ,\o[27] ,\o[26] ,\o[25] ,\o[24] ,\o[23] ,
        \o[22] ,\o[21] ,\o[20] ,\o[19] ,\o[18] ,\o[17] ,\o[16] ,\o[15] ,\o[14] ,\o[13] ,
        \o[12] ,\o[11] ,\o[10] ,\o[9] ,\o[8] ,\o[7] ,\o[6] ,\o[5] ,\o[4] ,\o[3] ,
        \o[2] ,\o[1] ,\o[0] );
input \s[31] ,\s[30] ,\s[29] ,\s[28] ,\s[27] ,\s[26] ,\s[25] ,\s[24] ,\s[23] ,
        \s[22] ,\s[21] ,\s[20] ,\s[19] ,\s[18] ,\s[17] ,\s[16] ,\s[15] ,\s[14] ,\s[13] ,
        \s[12] ,\s[11] ,\s[10] ,\s[9] ,\s[8] ,\s[7] ,\s[6] ,\s[5] ,\s[4] ,\s[3] ,
        \s[2] ,\s[1] ,\s[0] ,\a[31] ,\a[30] ,\a[29] ,\a[28] ,\a[27] ,\a[26] ,\a[25] ,
        \a[24] ,\a[23] ,\a[22] ,\a[21] ,\a[20] ,\a[19] ,\a[18] ,\a[17] ,\a[16] ,\a[15] ,
        \a[14] ,\a[13] ,\a[12] ,\a[11] ,\a[10] ,\a[9] ,\a[8] ,\a[7] ,\a[6] ,\a[5] ,
        \a[4] ,\a[3] ,\a[2] ,\a[1] ,\a[0] ,\b[31] ,\b[30] ,\b[29] ,\b[28] ,\b[27] ,
        \b[26] ,\b[25] ,\b[24] ,\b[23] ,\b[22] ,\b[21] ,\b[20] ,\b[19] ,\b[18] ,\b[17] ,
        \b[16] ,\b[15] ,\b[14] ,\b[13] ,\b[12] ,\b[11] ,\b[10] ,\b[9] ,\b[8] ,\b[7] ,
        \b[6] ,\b[5] ,\b[4] ,\b[3] ,\b[2] ,\b[1] ,\b[0] ,\c[31] ,\c[30] ,\c[29] ,
        \c[28] ,\c[27] ,\c[26] ,\c[25] ,\c[24] ,\c[23] ,\c[22] ,\c[21] ,\c[20] ,\c[19] ,
        \c[18] ,\c[17] ,\c[16] ,\c[15] ,\c[14] ,\c[13] ,\c[12] ,\c[11] ,\c[10] ,\c[9] ,
        \c[8] ,\c[7] ,\c[6] ,\c[5] ,\c[4] ,\c[3] ,\c[2] ,\c[1] ,\c[0] ,\d[31] ,
        \d[30] ,\d[29] ,\d[28] ,\d[27] ,\d[26] ,\d[25] ,\d[24] ,\d[23] ,\d[22] ,\d[21] ,
        \d[20] ,\d[19] ,\d[18] ,\d[17] ,\d[16] ,\d[15] ,\d[14] ,\d[13] ,\d[12] ,\d[11] ,
        \d[10] ,\d[9] ,\d[8] ,\d[7] ,\d[6] ,\d[5] ,\d[4] ,\d[3] ,\d[2] ,\d[1] ,
        \d[0] ;
output \o[31] ,\o[30] ,\o[29] ,\o[28] ,\o[27] ,\o[26] ,\o[25] ,\o[24] ,\o[23] ,
        \o[22] ,\o[21] ,\o[20] ,\o[19] ,\o[18] ,\o[17] ,\o[16] ,\o[15] ,\o[14] ,\o[13] ,
        \o[12] ,\o[11] ,\o[10] ,\o[9] ,\o[8] ,\o[7] ,\o[6] ,\o[5] ,\o[4] ,\o[3] ,
        \o[2] ,\o[1] ,\o[0] ;

wire \193_ZERO , \194 , \195 , \196 , \197 , \198 , \199 , \200 , \201 ,
         \202 , \203 , \204_ONE , \205_n5[0] , \206 , \207_A[0] , \208_B[0] , \209 , \210_SUM[0] , \211 ,
         \212 , \213 , \214 , \215 , \216 , \217 , \218 , \219 , \220 , \221 ,
         \222 , \223 , \224 , \225 , \226 , \227 , \228 , \229 , \230 , \231 ,
         \232 , \233 , \234 , \235 , \236 , \237 , \238 , \239 , \240 , \241 ,
         \242 , \243_A[0] , \244_B[0] , \245 , \246_SUM[0] , \247 , \248 , \249 , \250 , \251 ,
         \252 , \253 , \254 , \255 , \256 , \257 , \258 , \259 , \260 , \261 ,
         \262 , \263 , \264 , \265 , \266 , \267 , \268 , \269 , \270 , \271 ,
         \272 , \273 , \274 , \275 , \276 , \277 , \278 , \279_n5[1] , \280 , \281_A[1] ,
         \282_B[1] , \283 , \284 , \285 , \286 , \287 , \288_SUM[1] , \289 , \290_A[1] , \291_B[1] ,
         \292 , \293 , \294 , \295_SUM[1] , \296 , \297_n5[2] , \298 , \299_A[2] , \300_B[2] , \301 ,
         \302 , \303 , \304 , \305 , \306 , \307 , \308_SUM[2] , \309 , \310_A[2] , \311_B[2] ,
         \312 , \313 , \314 , \315 , \316 , \317 , \318_SUM[2] , \319 , \320_n5[3] , \321 ,
         \322_A[3] , \323_B[3] , \324 , \325 , \326 , \327 , \328 , \329 , \330 , \331_SUM[3] ,
         \332 , \333_A[3] , \334_B[3] , \335 , \336 , \337 , \338 , \339 , \340 , \341_SUM[3] ,
         \342 , \343_n5[4] , \344 , \345_A[4] , \346_B[4] , \347 , \348 , \349 , \350 , \351 ,
         \352 , \353 , \354_SUM[4] , \355 , \356_A[4] , \357_B[4] , \358 , \359 , \360 , \361 ,
         \362 , \363 , \364_SUM[4] , \365 , \366_n5[5] , \367 , \368_A[5] , \369_B[5] , \370 , \371 ,
         \372 , \373 , \374 , \375 , \376 , \377_SUM[5] , \378 , \379_A[5] , \380_B[5] , \381 ,
         \382 , \383 , \384 , \385 , \386 , \387_SUM[5] , \388 , \389_n5[6] , \390 , \391_A[6] ,
         \392_B[6] , \393 , \394 , \395 , \396 , \397 , \398 , \399 , \400_SUM[6] , \401 ,
         \402_A[6] , \403_B[6] , \404 , \405 , \406 , \407 , \408 , \409 , \410_SUM[6] , \411 ,
         \412_n5[7] , \413 , \414_A[7] , \415_B[7] , \416 , \417 , \418 , \419 , \420 , \421 ,
         \422 , \423_SUM[7] , \424 , \425_A[7] , \426_B[7] , \427 , \428 , \429 , \430 , \431 ,
         \432 , \433_SUM[7] , \434 , \435_n5[8] , \436 , \437_A[8] , \438_B[8] , \439 , \440 , \441 ,
         \442 , \443 , \444 , \445 , \446_SUM[8] , \447 , \448_A[8] , \449_B[8] , \450 , \451 ,
         \452 , \453 , \454 , \455 , \456_SUM[8] , \457 , \458_n5[9] , \459 , \460_A[9] , \461_B[9] ,
         \462 , \463 , \464 , \465 , \466 , \467 , \468 , \469_SUM[9] , \470 , \471_A[9] ,
         \472_B[9] , \473 , \474 , \475 , \476 , \477 , \478 , \479_SUM[9] , \480 , \481_n5[10] ,
         \482 , \483_A[10] , \484_B[10] , \485 , \486 , \487 , \488 , \489 , \490 , \491 ,
         \492_SUM[10] , \493 , \494_A[10] , \495_B[10] , \496 , \497 , \498 , \499 , \500 , \501 ,
         \502_SUM[10] , \503 , \504_n5[11] , \505 , \506_A[11] , \507_B[11] , \508 , \509 , \510 , \511 ,
         \512 , \513 , \514 , \515_SUM[11] , \516 , \517_A[11] , \518_B[11] , \519 , \520 , \521 ,
         \522 , \523 , \524 , \525_SUM[11] , \526 , \527_n5[12] , \528 , \529_A[12] , \530_B[12] , \531 ,
         \532 , \533 , \534 , \535 , \536 , \537 , \538_SUM[12] , \539 , \540_A[12] , \541_B[12] ,
         \542 , \543 , \544 , \545 , \546 , \547 , \548_SUM[12] , \549 , \550_n5[13] , \551 ,
         \552_A[13] , \553_B[13] , \554 , \555 , \556 , \557 , \558 , \559 , \560 , \561_SUM[13] ,
         \562 , \563_A[13] , \564_B[13] , \565 , \566 , \567 , \568 , \569 , \570 , \571_SUM[13] ,
         \572 , \573_n5[14] , \574 , \575_A[14] , \576_B[14] , \577 , \578 , \579 , \580 , \581 ,
         \582 , \583 , \584_SUM[14] , \585 , \586_A[14] , \587_B[14] , \588 , \589 , \590 , \591 ,
         \592 , \593 , \594_SUM[14] , \595 , \596_n5[15] , \597 , \598_A[15] , \599_B[15] , \600 , \601 ,
         \602 , \603 , \604 , \605 , \606 , \607_SUM[15] , \608 , \609_A[15] , \610_B[15] , \611 ,
         \612 , \613 , \614 , \615 , \616 , \617_SUM[15] , \618 , \619_n5[16] , \620 , \621_A[16] ,
         \622_B[16] , \623 , \624 , \625 , \626 , \627 , \628 , \629 , \630_SUM[16] , \631 ,
         \632_A[16] , \633_B[16] , \634 , \635 , \636 , \637 , \638 , \639 , \640_SUM[16] , \641 ,
         \642_n5[17] , \643 , \644_A[17] , \645_B[17] , \646 , \647 , \648 , \649 , \650 , \651 ,
         \652 , \653_SUM[17] , \654 , \655_A[17] , \656_B[17] , \657 , \658 , \659 , \660 , \661 ,
         \662 , \663_SUM[17] , \664 , \665_n5[18] , \666 , \667_A[18] , \668_B[18] , \669 , \670 , \671 ,
         \672 , \673 , \674 , \675 , \676_SUM[18] , \677 , \678_A[18] , \679_B[18] , \680 , \681 ,
         \682 , \683 , \684 , \685 , \686_SUM[18] , \687 , \688_n5[19] , \689 , \690_A[19] , \691_B[19] ,
         \692 , \693 , \694 , \695 , \696 , \697 , \698 , \699_SUM[19] , \700 , \701_A[19] ,
         \702_B[19] , \703 , \704 , \705 , \706 , \707 , \708 , \709_SUM[19] , \710 , \711_n5[20] ,
         \712 , \713_A[20] , \714_B[20] , \715 , \716 , \717 , \718 , \719 , \720 , \721 ,
         \722_SUM[20] , \723 , \724_A[20] , \725_B[20] , \726 , \727 , \728 , \729 , \730 , \731 ,
         \732_SUM[20] , \733 , \734_n5[21] , \735 , \736_A[21] , \737_B[21] , \738 , \739 , \740 , \741 ,
         \742 , \743 , \744 , \745_SUM[21] , \746 , \747_A[21] , \748_B[21] , \749 , \750 , \751 ,
         \752 , \753 , \754 , \755_SUM[21] , \756 , \757_n5[22] , \758 , \759_A[22] , \760_B[22] , \761 ,
         \762 , \763 , \764 , \765 , \766 , \767 , \768_SUM[22] , \769 , \770_A[22] , \771_B[22] ,
         \772 , \773 , \774 , \775 , \776 , \777 , \778_SUM[22] , \779 , \780_n5[23] , \781 ,
         \782_A[23] , \783_B[23] , \784 , \785 , \786 , \787 , \788 , \789 , \790 , \791_SUM[23] ,
         \792 , \793_A[23] , \794_B[23] , \795 , \796 , \797 , \798 , \799 , \800 , \801_SUM[23] ,
         \802 , \803_n5[24] , \804 , \805_A[24] , \806_B[24] , \807 , \808 , \809 , \810 , \811 ,
         \812 , \813 , \814_SUM[24] , \815 , \816_A[24] , \817_B[24] , \818 , \819 , \820 , \821 ,
         \822 , \823 , \824_SUM[24] , \825 , \826_n5[25] , \827 , \828_A[25] , \829_B[25] , \830 , \831 ,
         \832 , \833 , \834 , \835 , \836 , \837_SUM[25] , \838 , \839_A[25] , \840_B[25] , \841 ,
         \842 , \843 , \844 , \845 , \846 , \847_SUM[25] , \848 , \849_n5[26] , \850 , \851_A[26] ,
         \852_B[26] , \853 , \854 , \855 , \856 , \857 , \858 , \859 , \860_SUM[26] , \861 ,
         \862_A[26] , \863_B[26] , \864 , \865 , \866 , \867 , \868 , \869 , \870_SUM[26] , \871 ,
         \872_n5[27] , \873 , \874_A[27] , \875_B[27] , \876 , \877 , \878 , \879 , \880 , \881 ,
         \882 , \883_SUM[27] , \884 , \885_A[27] , \886_B[27] , \887 , \888 , \889 , \890 , \891 ,
         \892 , \893_SUM[27] , \894 , \895_n5[28] , \896 , \897_A[28] , \898_B[28] , \899 , \900 , \901 ,
         \902 , \903 , \904 , \905 , \906_SUM[28] , \907 , \908_A[28] , \909_B[28] , \910 , \911 ,
         \912 , \913 , \914 , \915 , \916_SUM[28] , \917 , \918_n5[29] , \919 , \920_A[29] , \921_B[29] ,
         \922 , \923 , \924 , \925 , \926 , \927 , \928 , \929_SUM[29] , \930 , \931_A[29] ,
         \932_B[29] , \933 , \934 , \935 , \936 , \937 , \938 , \939_SUM[29] , \940 , \941_n5[30] ,
         \942 , \943_A[30] , \944_B[30] , \945 , \946 , \947 , \948 , \949 , \950 , \951 ,
         \952_SUM[30] , \953 , \954_A[30] , \955_B[30] , \956 , \957 , \958 , \959 , \960 , \961 ,
         \962_SUM[30] , \963 , \964_n5[31] , \965 , \966_A[31] , \967_B[31] , \968 , \969 , \970 , \971 ,
         \972 , \973 , \974 , \975_SUM[31] , \976 , \977_A[31] , \978_B[31] , \979 , \980 , \981 ,
         \982 , \983 , \984 , \985_SUM[31] , \986 , \987_A[31] , \988_B[31] , \989 , \990_A[30] , \991_B[30] ,
         \992 , \993_A[29] , \994_B[29] , \995 , \996_A[28] , \997_B[28] , \998 , \999_A[27] , \1000_B[27] , \1001 ,
         \1002_A[26] , \1003_B[26] , \1004 , \1005_A[25] , \1006_B[25] , \1007 , \1008_A[24] , \1009_B[24] , \1010 , \1011_A[23] ,
         \1012_B[23] , \1013 , \1014_A[22] , \1015_B[22] , \1016 , \1017_A[21] , \1018_B[21] , \1019 , \1020_A[20] , \1021_B[20] ,
         \1022 , \1023_A[19] , \1024_B[19] , \1025 , \1026_A[18] , \1027_B[18] , \1028 , \1029_A[17] , \1030_B[17] , \1031 ,
         \1032_A[16] , \1033_B[16] , \1034 , \1035_A[15] , \1036_B[15] , \1037 , \1038_A[14] , \1039_B[14] , \1040 , \1041_A[13] ,
         \1042_B[13] , \1043 , \1044_A[12] , \1045_B[12] , \1046 , \1047_A[11] , \1048_B[11] , \1049 , \1050_A[10] , \1051_B[10] ,
         \1052 , \1053_A[9] , \1054_B[9] , \1055 , \1056_A[8] , \1057_B[8] , \1058 , \1059_A[7] , \1060_B[7] , \1061 ,
         \1062_A[6] , \1063_B[6] , \1064 , \1065_A[5] , \1066_B[5] , \1067 , \1068_A[4] , \1069_B[4] , \1070 , \1071_A[3] ,
         \1072_B[3] , \1073 , \1074_A[2] , \1075_B[2] , \1076 , \1077_A[1] , \1078_B[1] , \1079 , \1080_A[0] , \1081_B[0] ,
         \1082 , \1083 , \1084 , \1085 , \1086 , \1087 , \1088 , \1089 , \1090 , \1091 ,
         \1092 , \1093 , \1094 , \1095 , \1096 , \1097 , \1098 , \1099 , \1100 , \1101 ,
         \1102 , \1103 , \1104 , \1105 , \1106 , \1107 , \1108 , \1109 , \1110 , \1111 ,
         \1112 , \1113 , \1114 , \1115 , \1116 , \1117 , \1118 , \1119 , \1120 , \1121 ,
         \1122 , \1123 , \1124 , \1125 , \1126 , \1127 , \1128 , \1129 , \1130 , \1131 ,
         \1132 , \1133 , \1134 , \1135 , \1136 , \1137 , \1138 , \1139 , \1140 , \1141 ,
         \1142 , \1143 , \1144 , \1145 , \1146 , \1147 , \1148 , \1149 , \1150 , \1151 ,
         \1152 , \1153 , \1154 , \1155 , \1156 , \1157 , \1158 , \1159 , \1160 , \1161 ,
         \1162 , \1163 , \1164 , \1165 , \1166 , \1167 , \1168 , \1169 , \1170 , \1171 ,
         \1172 , \1173 , \1174_SUM[31] , \1175_A[31] , \1176 , \1177 , \1178_SUM[30] , \1179_A[30] , \1180 , \1181 ,
         \1182_SUM[29] , \1183_A[29] , \1184 , \1185 , \1186_SUM[28] , \1187_A[28] , \1188 , \1189 , \1190_SUM[27] , \1191_A[27] ,
         \1192 , \1193 , \1194_SUM[26] , \1195_A[26] , \1196 , \1197 , \1198_SUM[25] , \1199_A[25] , \1200 , \1201 ,
         \1202_SUM[24] , \1203_A[24] , \1204 , \1205 , \1206_SUM[23] , \1207_A[23] , \1208 , \1209 , \1210_SUM[22] , \1211_A[22] ,
         \1212 , \1213 , \1214_SUM[21] , \1215_A[21] , \1216 , \1217 , \1218_SUM[20] , \1219_A[20] , \1220 , \1221 ,
         \1222_SUM[19] , \1223_A[19] , \1224 , \1225 , \1226_SUM[18] , \1227_A[18] , \1228 , \1229 , \1230_SUM[17] , \1231_A[17] ,
         \1232 , \1233 , \1234_SUM[16] , \1235_A[16] , \1236 , \1237 , \1238_SUM[15] , \1239_A[15] , \1240 , \1241 ,
         \1242_SUM[14] , \1243_A[14] , \1244 , \1245 , \1246_SUM[13] , \1247_A[13] , \1248 , \1249 , \1250_SUM[12] , \1251_A[12] ,
         \1252 , \1253 , \1254_SUM[11] , \1255_A[11] , \1256 , \1257 , \1258_SUM[10] , \1259_A[10] , \1260 , \1261 ,
         \1262_SUM[9] , \1263_A[9] , \1264 , \1265 , \1266_SUM[8] , \1267_A[8] , \1268 , \1269 , \1270_SUM[7] , \1271_A[7] ,
         \1272 , \1273 , \1274_SUM[6] , \1275_A[6] , \1276 , \1277 , \1278_SUM[5] , \1279_A[5] , \1280 , \1281 ,
         \1282_SUM[4] , \1283_A[4] , \1284 , \1285 , \1286_SUM[3] , \1287_A[3] , \1288 , \1289 , \1290_SUM[2] , \1291_A[2] ,
         \1292 , \1293 , \1294_SUM[1] , \1295_A[1] , \1296 , \1297_SUM[0] , \1298_A[0] , \1299_B[31] , \1300_B[30] , \1301_B[29] ,
         \1302_B[28] , \1303_B[27] , \1304_B[26] , \1305_B[25] , \1306_B[24] , \1307_B[23] , \1308_B[22] , \1309_B[21] , \1310_B[20] , \1311_B[19] ,
         \1312_B[18] , \1313_B[17] , \1314_B[16] , \1315_B[15] , \1316_B[14] , \1317_B[13] , \1318_B[12] , \1319_B[11] , \1320_B[10] , \1321_B[9] ,
         \1322_B[8] , \1323_B[7] , \1324_B[6] , \1325_B[5] , \1326_B[4] , \1327_B[3] , \1328_B[2] , \1329_B[1] , \1330_B[0] , \1331 ,
         \1332 , \1333 , \1334 , \1335 , \1336 , \1337 , \1338 , \1339 , \1340 , \1341 ,
         \1342 , \1343 , \1344 , \1345 , \1346 , \1347 , \1348 , \1349 , \1350 , \1351 ,
         \1352 , \1353 , \1354 , \1355 , \1356 , \1357 , \1358 , \1359 , \1360 , \1361 ,
         \1362 , \1363 , \1364 , \1365 , \1366 , \1367 , \1368 , \1369 , \1370 , \1371 ,
         \1372 , \1373 , \1374 , \1375 , \1376 , \1377 , \1378 , \1379 , \1380 , \1381 ,
         \1382 , \1383 , \1384 , \1385 , \1386 , \1387 , \1388 , \1389 , \1390 , \1391 ,
         \1392 , \1393 , \1394 , \1395 , \1396 , \1397 , \1398 , \1399 , \1400 , \1401 ,
         \1402 , \1403 , \1404 , \1405 , \1406 , \1407 , \1408 , \1409 , \1410 , \1411 ,
         \1412 , \1413 , \1414 , \1415 , \1416 , \1417 , \1418 , \1419 , \1420 , \1421 ,
         \1422 , \1423 , \1424 , \1425 , \1426 , \1427 , \1428 , \1429 , \1430 , \1431 ,
         \1432 , \1433 , \1434 , \1435 , \1436 , \1437 , \1438 , \1439 , \1440 , \1441 ,
         \1442 , \1443 , \1444 , \1445 , \1446 , \1447 , \1448 , \1449 , \1450 , \1451 ,
         \1452 , \1453 , \1454 , \1455 , \1456 , \1457 , \1458 , \1459 , \1460 , \1461 ,
         \1462 , \1463 , \1464 , \1465 , \1466 , \1467 , \1468 , \1469 , \1470 , \1471 ,
         \1472 , \1473 , \1474 , \1475 , \1476 , \1477 , \1478 , \1479 , \1480 , \1481 ,
         \1482 , \1483 , \1484 , \1485 , \1486 , \1487 , \1488 , \1489 , \1490 , \1491 ,
         \1492 , \1493 , \1494 , \1495 , \1496 , \1497 , \1498 , \1499 , \1500 , \1501 ,
         \1502 , \1503 , \1504 , \1505 , \1506 , \1507 , \1508 , \1509 , \1510 , \1511 ,
         \1512 , \1513 , \1514 , \1515 , \1516 , \1517 , \1518 , \1519 , \1520 , \1521 ,
         \1522 , \1523 , \1524 , \1525 , \1526 , \1527 , \1528 , \1529 , \1530 , \1531 ,
         \1532 , \1533 , \1534 , \1535 , \1536 , \1537 , \1538 , \1539 , \1540 , \1541 ,
         \1542 , \1543 , \1544 , \1545 , \1546 , \1547 , \1548 , \1549 , \1550 , \1551 ,
         \1552 , \1553 , \1554 , \1555 , \1556 , \1557 , \1558 , \1559 , \1560 , \1561 ,
         \1562 , \1563 , \1564 , \1565 , \1566 , \1567 , \1568 , \1569 , \1570 , \1571 ,
         \1572 , \1573 , \1574 , \1575 , \1576 , \1577 , \1578 , \1579 , \1580 , \1581 ,
         \1582 , \1583 , \1584 , \1585 , \1586 , \1587 , \1588 , \1589 , \1590 , \1591 ,
         \1592 , \1593 , \1594 , \1595 , \1596 , \1597 , \1598 , \1599 , \1600 , \1601 ,
         \1602 , \1603 , \1604 , \1605 , \1606 , \1607 , \1608 , \1609 , \1610 , \1611 ,
         \1612 , \1613 , \1614 , \1615 , \1616 , \1617 , \1618 , \1619 , \1620 , \1621 ,
         \1622 , \1623 , \1624 , \1625 , \1626 , \1627 , \1628 , \1629 , \1630 , \1631 ,
         \1632 , \1633 , \1634 , \1635 , \1636 , \1637 , \1638 , \1639 , \1640 , \1641 ,
         \1642 , \1643 , \1644 , \1645 , \1646 , \1647 , \1648 , \1649 , \1650 , \1651 ,
         \1652 , \1653 , \1654 , \1655 , \1656 , \1657 , \1658 , \1659 , \1660 , \1661 ,
         \1662 , \1663 , \1664 , \1665 , \1666 , \1667 , \1668 , \1669 , \1670 , \1671 ,
         \1672 , \1673 , \1674 , \1675 , \1676 , \1677 , \1678 , \1679 , \1680 , \1681 ,
         \1682 , \1683 , \1684 , \1685 , \1686 , \1687 , \1688 , \1689 , \1690 , \1691 ,
         \1692 , \1693 , \1694 , \1695 , \1696 , \1697 , \1698 , \1699 , \1700 , \1701 ,
         \1702 , \1703 , \1704 , \1705 , \1706 , \1707 , \1708 , \1709 , \1710 , \1711 ,
         \1712 , \1713 , \1714 , \1715 , \1716 , \1717 , \1718 , \1719 , \1720 , \1721 ,
         \1722 , \1723 , \1724 , \1725 , \1726 , \1727 , \1728 , \1729 , \1730 , \1731 ,
         \1732 , \1733 , \1734 , \1735 , \1736 , \1737 , \1738 , \1739 , \1740 , \1741 ,
         \1742 , \1743 , \1744 , \1745 , \1746 , \1747 , \1748 , \1749 , \1750 , \1751 ,
         \1752 , \1753 , \1754 , \1755 , \1756 , \1757 , \1758 , \1759 , \1760 , \1761 ,
         \1762 , \1763 , \1764 , \1765 , \1766 , \1767 , \1768 , \1769 , \1770 , \1771 ,
         \1772 , \1773 , \1774 , \1775 , \1776 , \1777 , \1778 , \1779 , \1780 , \1781 ,
         \1782 , \1783 , \1784 , \1785 , \1786 , \1787 , \1788 , \1789 , \1790 , \1791 ,
         \1792 , \1793 , \1794 , \1795 , \1796 , \1797 , \1798 , \1799 , \1800 , \1801 ,
         \1802 , \1803 , \1804 , \1805 , \1806 , \1807 , \1808 , \1809 , \1810 , \1811 ,
         \1812 , \1813 , \1814 , \1815 , \1816 , \1817 , \1818 , \1819 , \1820 , \1821 ,
         \1822 , \1823 , \1824 , \1825 , \1826 , \1827 , \1828 , \1829 , \1830 , \1831 ,
         \1832 , \1833 , \1834 , \1835 , \1836 , \1837 , \1838 , \1839 , \1840 , \1841 ,
         \1842 , \1843 , \1844 , \1845 , \1846 , \1847 , \1848 , \1849 , \1850 , \1851 ,
         \1852 , \1853 , \1854 , \1855 , \1856 , \1857 , \1858 , \1859 , \1860 , \1861 ,
         \1862 , \1863 , \1864 , \1865 , \1866 , \1867 , \1868 , \1869 , \1870 , \1871 ,
         \1872 , \1873 , \1874 , \1875 , \1876 , \1877 , \1878 , \1879 , \1880 , \1881 ,
         \1882 , \1883 , \1884 , \1885 , \1886 , \1887 , \1888 , \1889 , \1890 , \1891 ,
         \1892 , \1893 , \1894 , \1895 , \1896 , \1897 , \1898 , \1899 , \1900 , \1901 ,
         \1902 , \1903 , \1904 , \1905 , \1906 , \1907 , \1908 , \1909 , \1910 , \1911 ,
         \1912 , \1913 , \1914 , \1915 , \1916 , \1917 , \1918 , \1919 , \1920 , \1921 ,
         \1922 , \1923 , \1924 , \1925 , \1926 , \1927 , \1928 , \1929 , \1930 , \1931 ,
         \1932 , \1933 , \1934 , \1935 , \1936 , \1937 , \1938 , \1939 , \1940 , \1941 ,
         \1942 , \1943 , \1944 , \1945 , \1946 , \1947 , \1948 , \1949 , \1950 , \1951 ,
         \1952 , \1953 , \1954 , \1955 , \1956 , \1957 , \1958 , \1959 , \1960 , \1961 ,
         \1962 , \1963 , \1964 , \1965 , \1966 , \1967 , \1968 , \1969 , \1970 , \1971 ,
         \1972 , \1973 , \1974 , \1975 , \1976 , \1977 , \1978 , \1979 , \1980 , \1981 ,
         \1982 , \1983 , \1984 , \1985 , \1986 , \1987 , \1988 , \1989 , \1990 , \1991 ,
         \1992 , \1993 , \1994 , \1995 , \1996 , \1997 , \1998 , \1999 , \2000 , \2001 ,
         \2002 , \2003 , \2004 , \2005 , \2006 , \2007 , \2008 , \2009 , \2010 , \2011 ,
         \2012 , \2013 , \2014 , \2015 , \2016 , \2017 , \2018 , \2019 , \2020 , \2021 ,
         \2022 , \2023 , \2024 , \2025 , \2026 , \2027 , \2028 , \2029 , \2030 , \2031 ,
         \2032 , \2033 , \2034 , \2035 , \2036 , \2037 , \2038 , \2039 , \2040 , \2041 ,
         \2042 , \2043 , \2044 , \2045 , \2046 , \2047 , \2048 , \2049 , \2050 , \2051 ,
         \2052 , \2053 , \2054 , \2055 , \2056 , \2057 , \2058 , \2059 , \2060 , \2061 ,
         \2062 , \2063 , \2064 , \2065 , \2066 , \2067 , \2068 , \2069 , \2070 , \2071 ,
         \2072 , \2073 , \2074 , \2075 , \2076 , \2077 , \2078 , \2079 , \2080 , \2081 ,
         \2082 , \2083 , \2084 , \2085 , \2086 , \2087 , \2088 , \2089 , \2090 , \2091 ,
         \2092 , \2093 , \2094 , \2095 , \2096 , \2097 , \2098 , \2099 , \2100 , \2101 ,
         \2102 , \2103 , \2104 , \2105 , \2106 , \2107 , \2108 , \2109 , \2110 , \2111 ,
         \2112 , \2113 , \2114 , \2115 , \2116 , \2117 , \2118 , \2119 , \2120 , \2121 ,
         \2122 , \2123 , \2124 , \2125 , \2126 , \2127 , \2128 , \2129 , \2130 , \2131 ,
         \2132 , \2133 , \2134 , \2135 , \2136 , \2137 , \2138 , \2139 , \2140 , \2141 ,
         \2142 , \2143 , \2144 , \2145 , \2146 , \2147 , \2148 , \2149 , \2150 , \2151 ,
         \2152 , \2153 , \2154 , \2155 , \2156 , \2157 , \2158 , \2159 , \2160 , \2161 ,
         \2162 , \2163 , \2164 , \2165 , \2166 , \2167 , \2168 , \2169 , \2170 , \2171 ,
         \2172 , \2173 , \2174 , \2175 , \2176 , \2177 , \2178 , \2179 , \2180 , \2181 ,
         \2182 , \2183 , \2184 , \2185 , \2186 , \2187 , \2188 , \2189 , \2190 , \2191 ,
         \2192 , \2193 , \2194 , \2195 , \2196 , \2197 , \2198 , \2199 , \2200 , \2201 ,
         \2202 , \2203 , \2204 , \2205 , \2206 , \2207 , \2208 , \2209 , \2210 , \2211 ,
         \2212 , \2213 , \2214 , \2215 , \2216 , \2217 , \2218 , \2219 , \2220 , \2221 ,
         \2222 , \2223 , \2224 , \2225 , \2226 , \2227 , \2228 , \2229 , \2230 , \2231 ,
         \2232 , \2233 , \2234 , \2235 , \2236 , \2237 , \2238 , \2239 , \2240 , \2241 ,
         \2242 , \2243 , \2244 , \2245 , \2246 , \2247 , \2248 , \2249 , \2250 , \2251 ,
         \2252 , \2253 , \2254 , \2255 , \2256 , \2257 , \2258 , \2259 , \2260 , \2261 ,
         \2262 , \2263 , \2264 , \2265 , \2266 , \2267 , \2268 , \2269 , \2270 , \2271 ,
         \2272 , \2273 , \2274 , \2275 , \2276 , \2277 , \2278 , \2279 , \2280 , \2281 ,
         \2282 , \2283 , \2284 , \2285 , \2286 , \2287 , \2288 , \2289 , \2290 , \2291 ,
         \2292 , \2293 , \2294 , \2295 , \2296 , \2297 , \2298 , \2299 , \2300 , \2301 ,
         \2302 , \2303 , \2304 , \2305 , \2306 , \2307 , \2308 , \2309 , \2310 , \2311 ,
         \2312 , \2313 , \2314 , \2315 , \2316 , \2317 , \2318 , \2319 , \2320 , \2321 ,
         \2322 , \2323 , \2324 , \2325 , \2326 , \2327 , \2328 , \2329 , \2330 , \2331 ,
         \2332 , \2333 , \2334 , \2335 , \2336 , \2337 , \2338 , \2339 , \2340 , \2341 ,
         \2342 , \2343 , \2344 , \2345 , \2346 , \2347 , \2348 , \2349 , \2350 , \2351 ,
         \2352 , \2353 , \2354 , \2355 , \2356 , \2357 , \2358 , \2359 , \2360 , \2361 ,
         \2362 , \2363 , \2364 , \2365 , \2366 , \2367 , \2368 , \2369 , \2370 , \2371 ,
         \2372 , \2373 , \2374 , \2375 , \2376 , \2377 , \2378 , \2379 , \2380 , \2381 ,
         \2382 , \2383 , \2384 , \2385 , \2386 , \2387 , \2388 , \2389 , \2390 , \2391 ,
         \2392 , \2393 , \2394 , \2395 , \2396 , \2397 , \2398 , \2399 , \2400 , \2401 ,
         \2402 , \2403 , \2404 , \2405 , \2406 , \2407 , \2408 , \2409 , \2410 , \2411 ,
         \2412 , \2413 , \2414 , \2415 , \2416 , \2417 , \2418 , \2419 , \2420 , \2421 ,
         \2422 , \2423 , \2424 , \2425 , \2426 , \2427 , \2428 , \2429 , \2430 , \2431 ,
         \2432 , \2433 , \2434 , \2435 , \2436 , \2437 , \2438 , \2439 , \2440 , \2441 ,
         \2442 , \2443 , \2444 , \2445 , \2446 , \2447 , \2448 , \2449 , \2450 , \2451 ,
         \2452 , \2453 , \2454 , \2455 , \2456 , \2457 , \2458 , \2459 , \2460 , \2461 ,
         \2462 , \2463 , \2464 , \2465 , \2466 , \2467 , \2468 , \2469 , \2470 , \2471 ,
         \2472 , \2473 , \2474 , \2475 , \2476 , \2477 , \2478 , \2479 , \2480 , \2481 ,
         \2482 , \2483 , \2484 , \2485 , \2486 , \2487 , \2488 , \2489 , \2490 , \2491 ,
         \2492 , \2493 , \2494 , \2495 , \2496 , \2497 , \2498 , \2499 , \2500 , \2501 ,
         \2502 , \2503 , \2504 , \2505 , \2506 , \2507 , \2508 , \2509 , \2510 , \2511 ,
         \2512 , \2513 , \2514 , \2515 , \2516 , \2517 , \2518 , \2519 , \2520 , \2521 ,
         \2522 , \2523 , \2524 , \2525 , \2526 , \2527 , \2528 , \2529 , \2530 , \2531 ,
         \2532 , \2533 , \2534 , \2535 , \2536 , \2537 , \2538 , \2539 , \2540 , \2541 ,
         \2542 , \2543 , \2544 , \2545 , \2546 , \2547 , \2548 , \2549 , \2550 , \2551 ,
         \2552 , \2553 , \2554 , \2555 , \2556 , \2557 , \2558 , \2559 , \2560 , \2561 ,
         \2562 , \2563 , \2564 , \2565 , \2566 , \2567 , \2568 , \2569 , \2570 , \2571 ,
         \2572 , \2573 , \2574 , \2575 , \2576 , \2577 , \2578 , \2579 , \2580 , \2581 ,
         \2582 , \2583 , \2584 , \2585 , \2586 , \2587 , \2588 , \2589 , \2590 , \2591 ,
         \2592 , \2593 , \2594 , \2595 , \2596 , \2597 , \2598 , \2599 , \2600 , \2601 ,
         \2602 , \2603 , \2604 , \2605 , \2606 , \2607 , \2608 , \2609 , \2610 , \2611 ,
         \2612 , \2613 , \2614 , \2615 , \2616 , \2617 , \2618 , \2619 , \2620 , \2621 ,
         \2622 , \2623 , \2624 , \2625 , \2626 , \2627 , \2628 , \2629 , \2630 , \2631 ,
         \2632 , \2633 , \2634 , \2635 , \2636 , \2637 , \2638 , \2639 , \2640 , \2641 ,
         \2642 , \2643 , \2644 , \2645 , \2646 , \2647 , \2648 , \2649 , \2650 , \2651 ,
         \2652 , \2653 , \2654 , \2655 , \2656 , \2657 , \2658 , \2659 , \2660 , \2661 ,
         \2662 , \2663 , \2664 , \2665 , \2666 , \2667 , \2668 , \2669 , \2670 , \2671 ,
         \2672 , \2673 , \2674 , \2675 , \2676 , \2677 , \2678 , \2679 , \2680 , \2681 ,
         \2682 , \2683 , \2684 , \2685 , \2686 , \2687 , \2688 , \2689 , \2690 , \2691 ,
         \2692 , \2693 , \2694 , \2695 , \2696 , \2697 , \2698 , \2699 , \2700 , \2701 ,
         \2702 , \2703 , \2704 , \2705 , \2706 , \2707 , \2708 , \2709 , \2710 , \2711 ,
         \2712 , \2713 , \2714 , \2715 , \2716 , \2717 , \2718 , \2719 , \2720 , \2721 ,
         \2722 , \2723 , \2724 , \2725 , \2726 , \2727 , \2728 , \2729 , \2730 , \2731 ,
         \2732 , \2733 , \2734 , \2735 , \2736 , \2737 , \2738 , \2739 , \2740 , \2741 ,
         \2742 , \2743 , \2744 , \2745 , \2746 , \2747 , \2748 , \2749 , \2750 , \2751 ,
         \2752 , \2753 , \2754 , \2755 , \2756 , \2757 , \2758 , \2759 , \2760 , \2761 ,
         \2762 , \2763 , \2764 , \2765 , \2766 , \2767 , \2768 , \2769 , \2770 , \2771 ,
         \2772 , \2773 , \2774 , \2775 , \2776 , \2777 , \2778 , \2779 , \2780 , \2781 ,
         \2782 , \2783 , \2784 , \2785 , \2786 , \2787 , \2788 , \2789 , \2790 , \2791 ,
         \2792 , \2793 , \2794 , \2795 , \2796 , \2797 , \2798 , \2799 , \2800 , \2801 ,
         \2802 , \2803 , \2804 , \2805 , \2806 , \2807 , \2808 , \2809 , \2810 , \2811 ,
         \2812 , \2813 , \2814 , \2815 , \2816 , \2817 , \2818 , \2819 , \2820 , \2821 ,
         \2822 , \2823 , \2824 , \2825 , \2826 , \2827 , \2828 , \2829 , \2830 , \2831 ,
         \2832 , \2833 , \2834 , \2835 , \2836 , \2837 , \2838 , \2839 , \2840 , \2841 ,
         \2842 , \2843 , \2844 , \2845 , \2846 , \2847 , \2848 , \2849 , \2850 , \2851 ,
         \2852 , \2853 , \2854 , \2855 , \2856 , \2857 , \2858 , \2859 , \2860 , \2861 ,
         \2862 , \2863 , \2864 , \2865 , \2866 , \2867 , \2868 , \2869 , \2870 , \2871 ,
         \2872 , \2873 , \2874 , \2875 , \2876 , \2877 , \2878 , \2879 , \2880 , \2881 ,
         \2882 , \2883 , \2884 , \2885 , \2886 , \2887 , \2888 , \2889 , \2890 , \2891 ,
         \2892 , \2893 , \2894 , \2895 , \2896 , \2897 , \2898 , \2899 , \2900 , \2901 ,
         \2902 , \2903 , \2904 , \2905 , \2906 , \2907 , \2908 , \2909 , \2910 , \2911 ,
         \2912 , \2913 , \2914 , \2915 , \2916 , \2917 , \2918 , \2919 , \2920 , \2921 ,
         \2922 , \2923 , \2924 , \2925 , \2926 , \2927 , \2928 , \2929 , \2930 , \2931 ,
         \2932 , \2933 , \2934 , \2935 , \2936 , \2937 , \2938 , \2939 , \2940 , \2941 ,
         \2942 , \2943 , \2944 , \2945 , \2946 , \2947 , \2948 , \2949 , \2950 , \2951 ,
         \2952 , \2953 , \2954 , \2955 , \2956 , \2957 , \2958 , \2959 , \2960 , \2961 ,
         \2962 , \2963 , \2964 , \2965 , \2966 , \2967 , \2968 , \2969 , \2970 , \2971 ,
         \2972 , \2973 , \2974 , \2975 , \2976 , \2977 , \2978 , \2979 , \2980 , \2981 ,
         \2982 , \2983 , \2984 , \2985 , \2986 , \2987 , \2988 , \2989 , \2990 , \2991 ,
         \2992 , \2993 , \2994 , \2995 , \2996 , \2997 , \2998 , \2999 , \3000 , \3001 ,
         \3002 , \3003 , \3004 , \3005 , \3006 , \3007 , \3008 , \3009 , \3010 , \3011 ,
         \3012 , \3013 , \3014 , \3015 , \3016 , \3017 , \3018 , \3019 , \3020 , \3021 ,
         \3022 , \3023 , \3024 , \3025 , \3026 , \3027 , \3028 , \3029 , \3030 , \3031 ,
         \3032 , \3033 , \3034 , \3035 , \3036 , \3037 , \3038 , \3039 , \3040 , \3041 ,
         \3042 , \3043 , \3044 , \3045 , \3046 , \3047 , \3048 , \3049 , \3050 , \3051 ,
         \3052 , \3053 , \3054 , \3055 , \3056 , \3057 , \3058 , \3059 , \3060 , \3061 ,
         \3062 , \3063 , \3064 , \3065 , \3066 , \3067 , \3068 , \3069 , \3070 , \3071 ,
         \3072 , \3073 , \3074 , \3075 , \3076 , \3077 , \3078 , \3079 , \3080 , \3081 ,
         \3082 , \3083 , \3084 , \3085 , \3086 , \3087 , \3088 , \3089 , \3090 , \3091 ,
         \3092 , \3093 , \3094 , \3095 , \3096 , \3097 , \3098 , \3099 , \3100 , \3101 ,
         \3102 , \3103 , \3104 , \3105 , \3106 , \3107 , \3108 , \3109 , \3110 , \3111 ,
         \3112 , \3113 , \3114 , \3115 , \3116 , \3117 , \3118 , \3119 , \3120 , \3121 ,
         \3122 , \3123 , \3124 , \3125 , \3126 , \3127 , \3128 , \3129 , \3130 , \3131 ,
         \3132 , \3133 , \3134 , \3135 , \3136 , \3137 , \3138 , \3139 , \3140 , \3141 ,
         \3142 , \3143 , \3144 , \3145 , \3146 , \3147 , \3148 , \3149 , \3150 , \3151 ,
         \3152 , \3153 , \3154 , \3155 , \3156 , \3157 , \3158 , \3159 , \3160 , \3161 ,
         \3162 , \3163 , \3164 , \3165 , \3166 , \3167 , \3168 , \3169 , \3170 , \3171 ,
         \3172 , \3173 , \3174 , \3175 , \3176 , \3177 , \3178 , \3179 , \3180 , \3181 ,
         \3182 , \3183 , \3184 , \3185 , \3186 , \3187 , \3188 , \3189 , \3190 , \3191 ,
         \3192 , \3193 , \3194 , \3195 , \3196 , \3197 , \3198 , \3199 , \3200 , \3201 ,
         \3202 , \3203 , \3204 , \3205 , \3206 , \3207 , \3208 , \3209 , \3210 , \3211 ,
         \3212 , \3213 , \3214 , \3215 , \3216 , \3217 , \3218 , \3219 , \3220 , \3221 ,
         \3222 , \3223 , \3224 , \3225 , \3226 , \3227 , \3228 , \3229 , \3230 , \3231 ,
         \3232 , \3233 , \3234 , \3235 , \3236 , \3237 , \3238 , \3239 , \3240 , \3241 ,
         \3242 , \3243 , \3244 , \3245 , \3246 , \3247 , \3248 , \3249 , \3250 , \3251 ,
         \3252 , \3253 , \3254 , \3255 , \3256 , \3257 , \3258 , \3259 , \3260 , \3261 ,
         \3262 , \3263 , \3264 , \3265 , \3266 , \3267 , \3268 , \3269 , \3270 , \3271 ,
         \3272 , \3273 , \3274 , \3275 , \3276 , \3277 , \3278 , \3279 , \3280 , \3281 ,
         \3282 , \3283 , \3284 , \3285 , \3286 , \3287 , \3288 , \3289 , \3290 , \3291 ,
         \3292 , \3293 , \3294 , \3295 , \3296 , \3297 , \3298 , \3299 , \3300 , \3301 ,
         \3302 , \3303 , \3304 , \3305 , \3306 , \3307 , \3308 , \3309 , \3310 , \3311 ,
         \3312 , \3313 , \3314 , \3315 , \3316 , \3317 , \3318 , \3319 , \3320 , \3321 ,
         \3322 , \3323 , \3324 , \3325 , \3326 , \3327 , \3328 , \3329 , \3330 , \3331 ,
         \3332 , \3333 , \3334 , \3335 , \3336 , \3337 , \3338 , \3339 , \3340 , \3341 ,
         \3342 , \3343 , \3344 , \3345 , \3346 , \3347 , \3348 , \3349 , \3350 , \3351 ,
         \3352 , \3353 , \3354 , \3355 , \3356 , \3357 , \3358 , \3359 , \3360 , \3361 ,
         \3362 , \3363 , \3364 , \3365 , \3366 , \3367 , \3368 , \3369 , \3370 , \3371 ,
         \3372 , \3373 , \3374 , \3375 , \3376 , \3377 , \3378 , \3379 , \3380 , \3381 ,
         \3382 , \3383 , \3384 , \3385 , \3386 , \3387 , \3388 , \3389 , \3390 , \3391 ,
         \3392 , \3393 , \3394 , \3395 , \3396 , \3397 , \3398 , \3399 , \3400 , \3401 ,
         \3402 , \3403 , \3404 , \3405 , \3406 , \3407 , \3408 , \3409 , \3410 , \3411 ,
         \3412 , \3413 , \3414 , \3415 , \3416 , \3417 , \3418 , \3419 , \3420 , \3421 ,
         \3422 , \3423 , \3424 , \3425 , \3426 , \3427 , \3428 , \3429 , \3430 , \3431 ,
         \3432 , \3433 , \3434 , \3435 , \3436 , \3437 , \3438 , \3439 , \3440 , \3441 ,
         \3442 , \3443 , \3444 , \3445 , \3446 , \3447 , \3448 , \3449 , \3450 , \3451 ,
         \3452 , \3453 , \3454 , \3455 , \3456 , \3457 , \3458 , \3459 , \3460 , \3461 ,
         \3462 , \3463 , \3464 , \3465 , \3466 , \3467 , \3468 , \3469 , \3470 , \3471 ,
         \3472 , \3473 , \3474 , \3475 , \3476 , \3477 , \3478 , \3479 , \3480 , \3481 ,
         \3482 , \3483 , \3484 , \3485 , \3486 , \3487 , \3488 , \3489 , \3490 , \3491 ,
         \3492 , \3493 , \3494 , \3495 , \3496 , \3497 , \3498 , \3499 , \3500 , \3501 ,
         \3502 , \3503 , \3504 , \3505 , \3506 , \3507 , \3508 , \3509 , \3510 , \3511 ,
         \3512 , \3513 , \3514 , \3515 , \3516 , \3517 , \3518 , \3519 , \3520 , \3521 ,
         \3522 , \3523 , \3524 , \3525 , \3526 , \3527 , \3528 , \3529 , \3530 , \3531 ,
         \3532 , \3533 , \3534 , \3535 , \3536 , \3537 , \3538 , \3539 , \3540 , \3541 ,
         \3542 , \3543 , \3544 , \3545 , \3546 , \3547 , \3548 , \3549 , \3550 , \3551 ,
         \3552 , \3553 , \3554 , \3555 , \3556 , \3557 , \3558 , \3559 , \3560 , \3561 ,
         \3562 , \3563 , \3564 , \3565 , \3566 , \3567 , \3568 , \3569 , \3570 , \3571 ,
         \3572 , \3573 , \3574 , \3575 , \3576 , \3577 , \3578 , \3579 , \3580 , \3581 ,
         \3582 , \3583 , \3584 , \3585 , \3586 , \3587 , \3588 , \3589 , \3590 , \3591 ,
         \3592 , \3593 , \3594 , \3595 , \3596 , \3597 , \3598 , \3599 , \3600 , \3601 ,
         \3602 , \3603 , \3604 , \3605 , \3606 , \3607 , \3608 , \3609 , \3610 , \3611 ,
         \3612 , \3613 , \3614 , \3615 , \3616 , \3617 , \3618 , \3619 , \3620 , \3621 ,
         \3622 , \3623 , \3624 , \3625 , \3626 , \3627 , \3628 , \3629 , \3630 , \3631 ,
         \3632 , \3633 , \3634 , \3635 , \3636 , \3637 , \3638 , \3639 , \3640 , \3641 ,
         \3642 , \3643 , \3644 , \3645 , \3646 , \3647 , \3648 , \3649 , \3650 , \3651 ,
         \3652 , \3653 , \3654 , \3655 , \3656 , \3657 , \3658 , \3659 , \3660 , \3661 ,
         \3662 , \3663 , \3664 , \3665 , \3666 , \3667 , \3668 , \3669 , \3670 , \3671 ,
         \3672 , \3673 , \3674 , \3675 , \3676 , \3677 , \3678 , \3679 , \3680 , \3681 ,
         \3682 , \3683 , \3684 , \3685 , \3686 , \3687 , \3688 , \3689 , \3690 , \3691 ,
         \3692 , \3693 , \3694 , \3695 , \3696 , \3697 , \3698 , \3699 , \3700 , \3701 ,
         \3702 , \3703 , \3704 , \3705 , \3706 , \3707 , \3708 , \3709 , \3710 , \3711 ,
         \3712 , \3713 , \3714 , \3715 , \3716 , \3717 , \3718 , \3719 , \3720 , \3721 ,
         \3722 , \3723 , \3724 , \3725 , \3726 , \3727 , \3728 , \3729 , \3730 , \3731 ,
         \3732 , \3733 , \3734 , \3735 , \3736 , \3737 , \3738 , \3739 , \3740 , \3741 ,
         \3742 , \3743 , \3744 , \3745 , \3746 , \3747 , \3748 , \3749 , \3750 , \3751 ,
         \3752 , \3753 , \3754 , \3755 , \3756 , \3757 , \3758 , \3759 , \3760 , \3761 ,
         \3762 , \3763 , \3764 , \3765 , \3766 , \3767 , \3768 , \3769 , \3770 , \3771 ,
         \3772 , \3773 , \3774 , \3775 , \3776 , \3777 , \3778 , \3779 , \3780 , \3781 ,
         \3782 , \3783 , \3784 , \3785 , \3786 , \3787 , \3788 , \3789 , \3790 , \3791 ,
         \3792 , \3793 , \3794 , \3795 , \3796 , \3797 , \3798 , \3799 , \3800 , \3801 ,
         \3802 , \3803 , \3804 , \3805 , \3806 , \3807 , \3808 , \3809 , \3810 , \3811 ,
         \3812 , \3813 , \3814 , \3815 , \3816 , \3817 , \3818 , \3819 , \3820 , \3821 ,
         \3822 , \3823 , \3824 , \3825 , \3826 , \3827 , \3828 , \3829 , \3830 , \3831 ,
         \3832 , \3833 , \3834 , \3835 , \3836 , \3837 , \3838 , \3839 , \3840 , \3841 ,
         \3842 , \3843 , \3844 , \3845 , \3846 , \3847 , \3848 , \3849 , \3850 , \3851 ,
         \3852 , \3853 , \3854 , \3855 , \3856 , \3857 , \3858 , \3859 , \3860 , \3861 ,
         \3862 , \3863 , \3864 , \3865 , \3866 , \3867 , \3868 , \3869 , \3870 , \3871 ,
         \3872 , \3873 , \3874 , \3875 , \3876 , \3877 , \3878 , \3879 , \3880 , \3881 ,
         \3882 , \3883 , \3884 , \3885 , \3886 , \3887 , \3888 , \3889 , \3890 , \3891 ,
         \3892 , \3893 , \3894 , \3895 , \3896 , \3897 , \3898 , \3899 , \3900 , \3901 ,
         \3902 , \3903 , \3904 , \3905 , \3906 , \3907 , \3908 , \3909 , \3910 , \3911 ,
         \3912 , \3913 , \3914 , \3915 , \3916 , \3917 , \3918 , \3919 , \3920 , \3921 ,
         \3922 , \3923 , \3924 , \3925 , \3926 , \3927_Z[31] , \3928 , \3929_Z[30] , \3930 , \3931_Z[29] ,
         \3932 , \3933_Z[28] , \3934 , \3935_Z[27] , \3936 , \3937_Z[26] , \3938 , \3939_Z[25] , \3940 , \3941_Z[24] ,
         \3942 , \3943_Z[23] , \3944 , \3945_Z[22] , \3946 , \3947_Z[21] , \3948 , \3949_Z[20] , \3950 , \3951_Z[19] ,
         \3952 , \3953_Z[18] , \3954 , \3955_Z[17] , \3956 , \3957_Z[16] , \3958 , \3959_Z[15] , \3960 , \3961_Z[14] ,
         \3962 , \3963_Z[13] , \3964 , \3965_Z[12] , \3966 , \3967_Z[11] , \3968 , \3969_Z[10] , \3970 , \3971_Z[9] ,
         \3972 , \3973_Z[8] , \3974 , \3975_Z[7] , \3976 , \3977_Z[6] , \3978 , \3979_Z[5] , \3980 , \3981_Z[4] ,
         \3982 , \3983_Z[3] , \3984 , \3985_Z[2] , \3986 , \3987_Z[1] , \3988 , \3989_Z[0] ;
buf \U$labaj426 ( \o[31] , \3927_Z[31] );
buf \U$labaj427 ( \o[30] , \3929_Z[30] );
buf \U$labaj428 ( \o[29] , \3931_Z[29] );
buf \U$labaj429 ( \o[28] , \3933_Z[28] );
buf \U$labaj430 ( \o[27] , \3935_Z[27] );
buf \U$labaj431 ( \o[26] , \3937_Z[26] );
buf \U$labaj432 ( \o[25] , \3939_Z[25] );
buf \U$labaj433 ( \o[24] , \3941_Z[24] );
buf \U$labaj434 ( \o[23] , \3943_Z[23] );
buf \U$labaj435 ( \o[22] , \3945_Z[22] );
buf \U$labaj436 ( \o[21] , \3947_Z[21] );
buf \U$labaj437 ( \o[20] , \3949_Z[20] );
buf \U$labaj438 ( \o[19] , \3951_Z[19] );
buf \U$labaj439 ( \o[18] , \3953_Z[18] );
buf \U$labaj440 ( \o[17] , \3955_Z[17] );
buf \U$labaj441 ( \o[16] , \3957_Z[16] );
buf \U$labaj442 ( \o[15] , \3959_Z[15] );
buf \U$labaj443 ( \o[14] , \3961_Z[14] );
buf \U$labaj444 ( \o[13] , \3963_Z[13] );
buf \U$labaj445 ( \o[12] , \3965_Z[12] );
buf \U$labaj446 ( \o[11] , \3967_Z[11] );
buf \U$labaj447 ( \o[10] , \3969_Z[10] );
buf \U$labaj448 ( \o[9] , \3971_Z[9] );
buf \U$labaj449 ( \o[8] , \3973_Z[8] );
buf \U$labaj450 ( \o[7] , \3975_Z[7] );
buf \U$labaj451 ( \o[6] , \3977_Z[6] );
buf \U$labaj452 ( \o[5] , \3979_Z[5] );
buf \U$labaj453 ( \o[4] , \3981_Z[4] );
buf \U$labaj454 ( \o[3] , \3983_Z[3] );
buf \U$labaj455 ( \o[2] , \3985_Z[2] );
buf \U$labaj456 ( \o[1] , \3987_Z[1] );
buf \U$labaj457 ( \o[0] , \3989_Z[0] );
_DC \n5[0] ( \205_n5[0] , 1'b0 , 1'b1 );
or \U$5/U$1 ( \206 , \b[0] , \205_n5[0] );
buf \sub_5_33/A[0] ( \207_A[0] , \c[0] );
buf \sub_5_33/B[0] ( \208_B[0] , \d[0] );
xor \sub_5_33/U$215 ( \209 , \207_A[0] , \208_B[0] );
buf \sub_5_33/SUM[0] ( \210_SUM[0] , \209 );
xor \U$4 ( \211 , \a[31] , \a[30] );
xor \U$4_g1 ( \212 , \a[29] , \a[28] );
xor \U$4_g2 ( \213 , \211 , \212 );
xor \U$4_g3 ( \214 , \a[27] , \a[26] );
xor \U$4_g4 ( \215 , \a[25] , \a[24] );
xor \U$4_g5 ( \216 , \214 , \215 );
xor \U$4_g6 ( \217 , \213 , \216 );
xor \U$4_g7 ( \218 , \a[23] , \a[22] );
xor \U$4_g8 ( \219 , \a[21] , \a[20] );
xor \U$4_g9 ( \220 , \218 , \219 );
xor \U$4_g10 ( \221 , \a[19] , \a[18] );
xor \U$4_g11 ( \222 , \a[17] , \a[16] );
xor \U$4_g12 ( \223 , \221 , \222 );
xor \U$4_g13 ( \224 , \220 , \223 );
xor \U$4_g14 ( \225 , \217 , \224 );
xor \U$4_g15 ( \226 , \a[15] , \a[14] );
xor \U$4_g16 ( \227 , \a[13] , \a[12] );
xor \U$4_g17 ( \228 , \226 , \227 );
xor \U$4_g18 ( \229 , \a[11] , \a[10] );
xor \U$4_g19 ( \230 , \a[9] , \a[8] );
xor \U$4_g20 ( \231 , \229 , \230 );
xor \U$4_g21 ( \232 , \228 , \231 );
xor \U$4_g22 ( \233 , \a[7] , \a[6] );
xor \U$4_g23 ( \234 , \a[5] , \a[4] );
xor \U$4_g24 ( \235 , \233 , \234 );
xor \U$4_g25 ( \236 , \a[3] , \a[2] );
xor \U$4_g26 ( \237 , \a[1] , \a[0] );
xor \U$4_g27 ( \238 , \236 , \237 );
xor \U$4_g28 ( \239 , \235 , \238 );
xor \U$4_g29 ( \240 , \232 , \239 );
xor \U$4_g30 ( \241 , \225 , \240 );
_HMUX \U$3/U$1 ( \242 , \206 , \210_SUM[0] , \241 );
buf \add_5_20/A[0] ( \243_A[0] , \c[0] );
buf \add_5_20/B[0] ( \244_B[0] , \d[0] );
xor \add_5_20/U$184 ( \245 , \243_A[0] , \244_B[0] );
buf \add_5_20/SUM[0] ( \246_SUM[0] , \245 );
xor \U$2 ( \247 , \s[31] , \s[30] );
xor \U$2_g1 ( \248 , \s[29] , \s[28] );
xor \U$2_g2 ( \249 , \247 , \248 );
xor \U$2_g3 ( \250 , \s[27] , \s[26] );
xor \U$2_g4 ( \251 , \s[25] , \s[24] );
xor \U$2_g5 ( \252 , \250 , \251 );
xor \U$2_g6 ( \253 , \249 , \252 );
xor \U$2_g7 ( \254 , \s[23] , \s[22] );
xor \U$2_g8 ( \255 , \s[21] , \s[20] );
xor \U$2_g9 ( \256 , \254 , \255 );
xor \U$2_g10 ( \257 , \s[19] , \s[18] );
xor \U$2_g11 ( \258 , \s[17] , \s[16] );
xor \U$2_g12 ( \259 , \257 , \258 );
xor \U$2_g13 ( \260 , \256 , \259 );
xor \U$2_g14 ( \261 , \253 , \260 );
xor \U$2_g15 ( \262 , \s[15] , \s[14] );
xor \U$2_g16 ( \263 , \s[13] , \s[12] );
xor \U$2_g17 ( \264 , \262 , \263 );
xor \U$2_g18 ( \265 , \s[11] , \s[10] );
xor \U$2_g19 ( \266 , \s[9] , \s[8] );
xor \U$2_g20 ( \267 , \265 , \266 );
xor \U$2_g21 ( \268 , \264 , \267 );
xor \U$2_g22 ( \269 , \s[7] , \s[6] );
xor \U$2_g23 ( \270 , \s[5] , \s[4] );
xor \U$2_g24 ( \271 , \269 , \270 );
xor \U$2_g25 ( \272 , \s[3] , \s[2] );
xor \U$2_g26 ( \273 , \s[1] , \s[0] );
xor \U$2_g27 ( \274 , \272 , \273 );
xor \U$2_g28 ( \275 , \271 , \274 );
xor \U$2_g29 ( \276 , \268 , \275 );
xor \U$2_g30 ( \277 , \261 , \276 );
_HMUX \U$1/U$1 ( \278 , \242 , \246_SUM[0] , \277 );
_DC \n5[1] ( \279_n5[1] , 1'b0 , 1'b1 );
or \U$5/U$2 ( \280 , \b[1] , \279_n5[1] );
buf \sub_5_33/A[1] ( \281_A[1] , \c[1] );
buf \sub_5_33/B[1] ( \282_B[1] , \d[1] );
not \sub_5_33/U$213 ( \283 , \282_B[1] );
xor \sub_5_33/U$212 ( \284 , \281_A[1] , \283 );
not \sub_5_33/U$216 ( \285 , \208_B[0] );
or \sub_5_33/U$214 ( \286 , \207_A[0] , \285 );
xor \sub_5_33/U$211 ( \287 , \284 , \286 );
buf \sub_5_33/SUM[1] ( \288_SUM[1] , \287 );
_HMUX \U$3/U$2 ( \289 , \280 , \288_SUM[1] , \241 );
buf \add_5_20/A[1] ( \290_A[1] , \c[1] );
buf \add_5_20/B[1] ( \291_B[1] , \d[1] );
xor \add_5_20/U$182 ( \292 , \290_A[1] , \291_B[1] );
and \add_5_20/U$183 ( \293 , \243_A[0] , \244_B[0] );
xor \add_5_20/U$181 ( \294 , \292 , \293 );
buf \add_5_20/SUM[1] ( \295_SUM[1] , \294 );
_HMUX \U$1/U$2 ( \296 , \289 , \295_SUM[1] , \277 );
_DC \n5[2] ( \297_n5[2] , 1'b0 , 1'b1 );
or \U$5/U$3 ( \298 , \b[2] , \297_n5[2] );
buf \sub_5_33/A[2] ( \299_A[2] , \c[2] );
buf \sub_5_33/B[2] ( \300_B[2] , \d[2] );
not \sub_5_33/U$206 ( \301 , \300_B[2] );
xor \sub_5_33/U$205 ( \302 , \299_A[2] , \301 );
and \sub_5_33/U$210 ( \303 , \281_A[1] , \283 );
and \sub_5_33/U$209 ( \304 , \283 , \286 );
and \sub_5_33/U$208 ( \305 , \281_A[1] , \286 );
or \sub_5_33/U$207 ( \306 , \303 , \304 , \305 );
xor \sub_5_33/U$204 ( \307 , \302 , \306 );
buf \sub_5_33/SUM[2] ( \308_SUM[2] , \307 );
_HMUX \U$3/U$3 ( \309 , \298 , \308_SUM[2] , \241 );
buf \add_5_20/A[2] ( \310_A[2] , \c[2] );
buf \add_5_20/B[2] ( \311_B[2] , \d[2] );
xor \add_5_20/U$176 ( \312 , \310_A[2] , \311_B[2] );
and \add_5_20/U$180 ( \313 , \290_A[1] , \291_B[1] );
and \add_5_20/U$179 ( \314 , \291_B[1] , \293 );
and \add_5_20/U$178 ( \315 , \290_A[1] , \293 );
or \add_5_20/U$177 ( \316 , \313 , \314 , \315 );
xor \add_5_20/U$175 ( \317 , \312 , \316 );
buf \add_5_20/SUM[2] ( \318_SUM[2] , \317 );
_HMUX \U$1/U$3 ( \319 , \309 , \318_SUM[2] , \277 );
_DC \n5[3] ( \320_n5[3] , 1'b0 , 1'b1 );
or \U$5/U$4 ( \321 , \b[3] , \320_n5[3] );
buf \sub_5_33/A[3] ( \322_A[3] , \c[3] );
buf \sub_5_33/B[3] ( \323_B[3] , \d[3] );
not \sub_5_33/U$199 ( \324 , \323_B[3] );
xor \sub_5_33/U$198 ( \325 , \322_A[3] , \324 );
and \sub_5_33/U$203 ( \326 , \299_A[2] , \301 );
and \sub_5_33/U$202 ( \327 , \301 , \306 );
and \sub_5_33/U$201 ( \328 , \299_A[2] , \306 );
or \sub_5_33/U$200 ( \329 , \326 , \327 , \328 );
xor \sub_5_33/U$197 ( \330 , \325 , \329 );
buf \sub_5_33/SUM[3] ( \331_SUM[3] , \330 );
_HMUX \U$3/U$4 ( \332 , \321 , \331_SUM[3] , \241 );
buf \add_5_20/A[3] ( \333_A[3] , \c[3] );
buf \add_5_20/B[3] ( \334_B[3] , \d[3] );
xor \add_5_20/U$170 ( \335 , \333_A[3] , \334_B[3] );
and \add_5_20/U$174 ( \336 , \310_A[2] , \311_B[2] );
and \add_5_20/U$173 ( \337 , \311_B[2] , \316 );
and \add_5_20/U$172 ( \338 , \310_A[2] , \316 );
or \add_5_20/U$171 ( \339 , \336 , \337 , \338 );
xor \add_5_20/U$169 ( \340 , \335 , \339 );
buf \add_5_20/SUM[3] ( \341_SUM[3] , \340 );
_HMUX \U$1/U$4 ( \342 , \332 , \341_SUM[3] , \277 );
_DC \n5[4] ( \343_n5[4] , 1'b0 , 1'b1 );
or \U$5/U$5 ( \344 , \b[4] , \343_n5[4] );
buf \sub_5_33/A[4] ( \345_A[4] , \c[4] );
buf \sub_5_33/B[4] ( \346_B[4] , \d[4] );
not \sub_5_33/U$192 ( \347 , \346_B[4] );
xor \sub_5_33/U$191 ( \348 , \345_A[4] , \347 );
and \sub_5_33/U$196 ( \349 , \322_A[3] , \324 );
and \sub_5_33/U$195 ( \350 , \324 , \329 );
and \sub_5_33/U$194 ( \351 , \322_A[3] , \329 );
or \sub_5_33/U$193 ( \352 , \349 , \350 , \351 );
xor \sub_5_33/U$190 ( \353 , \348 , \352 );
buf \sub_5_33/SUM[4] ( \354_SUM[4] , \353 );
_HMUX \U$3/U$5 ( \355 , \344 , \354_SUM[4] , \241 );
buf \add_5_20/A[4] ( \356_A[4] , \c[4] );
buf \add_5_20/B[4] ( \357_B[4] , \d[4] );
xor \add_5_20/U$164 ( \358 , \356_A[4] , \357_B[4] );
and \add_5_20/U$168 ( \359 , \333_A[3] , \334_B[3] );
and \add_5_20/U$167 ( \360 , \334_B[3] , \339 );
and \add_5_20/U$166 ( \361 , \333_A[3] , \339 );
or \add_5_20/U$165 ( \362 , \359 , \360 , \361 );
xor \add_5_20/U$163 ( \363 , \358 , \362 );
buf \add_5_20/SUM[4] ( \364_SUM[4] , \363 );
_HMUX \U$1/U$5 ( \365 , \355 , \364_SUM[4] , \277 );
_DC \n5[5] ( \366_n5[5] , 1'b0 , 1'b1 );
or \U$5/U$6 ( \367 , \b[5] , \366_n5[5] );
buf \sub_5_33/A[5] ( \368_A[5] , \c[5] );
buf \sub_5_33/B[5] ( \369_B[5] , \d[5] );
not \sub_5_33/U$185 ( \370 , \369_B[5] );
xor \sub_5_33/U$184 ( \371 , \368_A[5] , \370 );
and \sub_5_33/U$189 ( \372 , \345_A[4] , \347 );
and \sub_5_33/U$188 ( \373 , \347 , \352 );
and \sub_5_33/U$187 ( \374 , \345_A[4] , \352 );
or \sub_5_33/U$186 ( \375 , \372 , \373 , \374 );
xor \sub_5_33/U$183 ( \376 , \371 , \375 );
buf \sub_5_33/SUM[5] ( \377_SUM[5] , \376 );
_HMUX \U$3/U$6 ( \378 , \367 , \377_SUM[5] , \241 );
buf \add_5_20/A[5] ( \379_A[5] , \c[5] );
buf \add_5_20/B[5] ( \380_B[5] , \d[5] );
xor \add_5_20/U$158 ( \381 , \379_A[5] , \380_B[5] );
and \add_5_20/U$162 ( \382 , \356_A[4] , \357_B[4] );
and \add_5_20/U$161 ( \383 , \357_B[4] , \362 );
and \add_5_20/U$160 ( \384 , \356_A[4] , \362 );
or \add_5_20/U$159 ( \385 , \382 , \383 , \384 );
xor \add_5_20/U$157 ( \386 , \381 , \385 );
buf \add_5_20/SUM[5] ( \387_SUM[5] , \386 );
_HMUX \U$1/U$6 ( \388 , \378 , \387_SUM[5] , \277 );
_DC \n5[6] ( \389_n5[6] , 1'b0 , 1'b1 );
or \U$5/U$7 ( \390 , \b[6] , \389_n5[6] );
buf \sub_5_33/A[6] ( \391_A[6] , \c[6] );
buf \sub_5_33/B[6] ( \392_B[6] , \d[6] );
not \sub_5_33/U$178 ( \393 , \392_B[6] );
xor \sub_5_33/U$177 ( \394 , \391_A[6] , \393 );
and \sub_5_33/U$182 ( \395 , \368_A[5] , \370 );
and \sub_5_33/U$181 ( \396 , \370 , \375 );
and \sub_5_33/U$180 ( \397 , \368_A[5] , \375 );
or \sub_5_33/U$179 ( \398 , \395 , \396 , \397 );
xor \sub_5_33/U$176 ( \399 , \394 , \398 );
buf \sub_5_33/SUM[6] ( \400_SUM[6] , \399 );
_HMUX \U$3/U$7 ( \401 , \390 , \400_SUM[6] , \241 );
buf \add_5_20/A[6] ( \402_A[6] , \c[6] );
buf \add_5_20/B[6] ( \403_B[6] , \d[6] );
xor \add_5_20/U$152 ( \404 , \402_A[6] , \403_B[6] );
and \add_5_20/U$156 ( \405 , \379_A[5] , \380_B[5] );
and \add_5_20/U$155 ( \406 , \380_B[5] , \385 );
and \add_5_20/U$154 ( \407 , \379_A[5] , \385 );
or \add_5_20/U$153 ( \408 , \405 , \406 , \407 );
xor \add_5_20/U$151 ( \409 , \404 , \408 );
buf \add_5_20/SUM[6] ( \410_SUM[6] , \409 );
_HMUX \U$1/U$7 ( \411 , \401 , \410_SUM[6] , \277 );
_DC \n5[7] ( \412_n5[7] , 1'b0 , 1'b1 );
or \U$5/U$8 ( \413 , \b[7] , \412_n5[7] );
buf \sub_5_33/A[7] ( \414_A[7] , \c[7] );
buf \sub_5_33/B[7] ( \415_B[7] , \d[7] );
not \sub_5_33/U$171 ( \416 , \415_B[7] );
xor \sub_5_33/U$170 ( \417 , \414_A[7] , \416 );
and \sub_5_33/U$175 ( \418 , \391_A[6] , \393 );
and \sub_5_33/U$174 ( \419 , \393 , \398 );
and \sub_5_33/U$173 ( \420 , \391_A[6] , \398 );
or \sub_5_33/U$172 ( \421 , \418 , \419 , \420 );
xor \sub_5_33/U$169 ( \422 , \417 , \421 );
buf \sub_5_33/SUM[7] ( \423_SUM[7] , \422 );
_HMUX \U$3/U$8 ( \424 , \413 , \423_SUM[7] , \241 );
buf \add_5_20/A[7] ( \425_A[7] , \c[7] );
buf \add_5_20/B[7] ( \426_B[7] , \d[7] );
xor \add_5_20/U$146 ( \427 , \425_A[7] , \426_B[7] );
and \add_5_20/U$150 ( \428 , \402_A[6] , \403_B[6] );
and \add_5_20/U$149 ( \429 , \403_B[6] , \408 );
and \add_5_20/U$148 ( \430 , \402_A[6] , \408 );
or \add_5_20/U$147 ( \431 , \428 , \429 , \430 );
xor \add_5_20/U$145 ( \432 , \427 , \431 );
buf \add_5_20/SUM[7] ( \433_SUM[7] , \432 );
_HMUX \U$1/U$8 ( \434 , \424 , \433_SUM[7] , \277 );
_DC \n5[8] ( \435_n5[8] , 1'b0 , 1'b1 );
or \U$5/U$9 ( \436 , \b[8] , \435_n5[8] );
buf \sub_5_33/A[8] ( \437_A[8] , \c[8] );
buf \sub_5_33/B[8] ( \438_B[8] , \d[8] );
not \sub_5_33/U$164 ( \439 , \438_B[8] );
xor \sub_5_33/U$163 ( \440 , \437_A[8] , \439 );
and \sub_5_33/U$168 ( \441 , \414_A[7] , \416 );
and \sub_5_33/U$167 ( \442 , \416 , \421 );
and \sub_5_33/U$166 ( \443 , \414_A[7] , \421 );
or \sub_5_33/U$165 ( \444 , \441 , \442 , \443 );
xor \sub_5_33/U$162 ( \445 , \440 , \444 );
buf \sub_5_33/SUM[8] ( \446_SUM[8] , \445 );
_HMUX \U$3/U$9 ( \447 , \436 , \446_SUM[8] , \241 );
buf \add_5_20/A[8] ( \448_A[8] , \c[8] );
buf \add_5_20/B[8] ( \449_B[8] , \d[8] );
xor \add_5_20/U$140 ( \450 , \448_A[8] , \449_B[8] );
and \add_5_20/U$144 ( \451 , \425_A[7] , \426_B[7] );
and \add_5_20/U$143 ( \452 , \426_B[7] , \431 );
and \add_5_20/U$142 ( \453 , \425_A[7] , \431 );
or \add_5_20/U$141 ( \454 , \451 , \452 , \453 );
xor \add_5_20/U$139 ( \455 , \450 , \454 );
buf \add_5_20/SUM[8] ( \456_SUM[8] , \455 );
_HMUX \U$1/U$9 ( \457 , \447 , \456_SUM[8] , \277 );
_DC \n5[9] ( \458_n5[9] , 1'b0 , 1'b1 );
or \U$5/U$10 ( \459 , \b[9] , \458_n5[9] );
buf \sub_5_33/A[9] ( \460_A[9] , \c[9] );
buf \sub_5_33/B[9] ( \461_B[9] , \d[9] );
not \sub_5_33/U$157 ( \462 , \461_B[9] );
xor \sub_5_33/U$156 ( \463 , \460_A[9] , \462 );
and \sub_5_33/U$161 ( \464 , \437_A[8] , \439 );
and \sub_5_33/U$160 ( \465 , \439 , \444 );
and \sub_5_33/U$159 ( \466 , \437_A[8] , \444 );
or \sub_5_33/U$158 ( \467 , \464 , \465 , \466 );
xor \sub_5_33/U$155 ( \468 , \463 , \467 );
buf \sub_5_33/SUM[9] ( \469_SUM[9] , \468 );
_HMUX \U$3/U$10 ( \470 , \459 , \469_SUM[9] , \241 );
buf \add_5_20/A[9] ( \471_A[9] , \c[9] );
buf \add_5_20/B[9] ( \472_B[9] , \d[9] );
xor \add_5_20/U$134 ( \473 , \471_A[9] , \472_B[9] );
and \add_5_20/U$138 ( \474 , \448_A[8] , \449_B[8] );
and \add_5_20/U$137 ( \475 , \449_B[8] , \454 );
and \add_5_20/U$136 ( \476 , \448_A[8] , \454 );
or \add_5_20/U$135 ( \477 , \474 , \475 , \476 );
xor \add_5_20/U$133 ( \478 , \473 , \477 );
buf \add_5_20/SUM[9] ( \479_SUM[9] , \478 );
_HMUX \U$1/U$10 ( \480 , \470 , \479_SUM[9] , \277 );
_DC \n5[10] ( \481_n5[10] , 1'b0 , 1'b1 );
or \U$5/U$11 ( \482 , \b[10] , \481_n5[10] );
buf \sub_5_33/A[10] ( \483_A[10] , \c[10] );
buf \sub_5_33/B[10] ( \484_B[10] , \d[10] );
not \sub_5_33/U$150 ( \485 , \484_B[10] );
xor \sub_5_33/U$149 ( \486 , \483_A[10] , \485 );
and \sub_5_33/U$154 ( \487 , \460_A[9] , \462 );
and \sub_5_33/U$153 ( \488 , \462 , \467 );
and \sub_5_33/U$152 ( \489 , \460_A[9] , \467 );
or \sub_5_33/U$151 ( \490 , \487 , \488 , \489 );
xor \sub_5_33/U$148 ( \491 , \486 , \490 );
buf \sub_5_33/SUM[10] ( \492_SUM[10] , \491 );
_HMUX \U$3/U$11 ( \493 , \482 , \492_SUM[10] , \241 );
buf \add_5_20/A[10] ( \494_A[10] , \c[10] );
buf \add_5_20/B[10] ( \495_B[10] , \d[10] );
xor \add_5_20/U$128 ( \496 , \494_A[10] , \495_B[10] );
and \add_5_20/U$132 ( \497 , \471_A[9] , \472_B[9] );
and \add_5_20/U$131 ( \498 , \472_B[9] , \477 );
and \add_5_20/U$130 ( \499 , \471_A[9] , \477 );
or \add_5_20/U$129 ( \500 , \497 , \498 , \499 );
xor \add_5_20/U$127 ( \501 , \496 , \500 );
buf \add_5_20/SUM[10] ( \502_SUM[10] , \501 );
_HMUX \U$1/U$11 ( \503 , \493 , \502_SUM[10] , \277 );
_DC \n5[11] ( \504_n5[11] , 1'b0 , 1'b1 );
or \U$5/U$12 ( \505 , \b[11] , \504_n5[11] );
buf \sub_5_33/A[11] ( \506_A[11] , \c[11] );
buf \sub_5_33/B[11] ( \507_B[11] , \d[11] );
not \sub_5_33/U$143 ( \508 , \507_B[11] );
xor \sub_5_33/U$142 ( \509 , \506_A[11] , \508 );
and \sub_5_33/U$147 ( \510 , \483_A[10] , \485 );
and \sub_5_33/U$146 ( \511 , \485 , \490 );
and \sub_5_33/U$145 ( \512 , \483_A[10] , \490 );
or \sub_5_33/U$144 ( \513 , \510 , \511 , \512 );
xor \sub_5_33/U$141 ( \514 , \509 , \513 );
buf \sub_5_33/SUM[11] ( \515_SUM[11] , \514 );
_HMUX \U$3/U$12 ( \516 , \505 , \515_SUM[11] , \241 );
buf \add_5_20/A[11] ( \517_A[11] , \c[11] );
buf \add_5_20/B[11] ( \518_B[11] , \d[11] );
xor \add_5_20/U$122 ( \519 , \517_A[11] , \518_B[11] );
and \add_5_20/U$126 ( \520 , \494_A[10] , \495_B[10] );
and \add_5_20/U$125 ( \521 , \495_B[10] , \500 );
and \add_5_20/U$124 ( \522 , \494_A[10] , \500 );
or \add_5_20/U$123 ( \523 , \520 , \521 , \522 );
xor \add_5_20/U$121 ( \524 , \519 , \523 );
buf \add_5_20/SUM[11] ( \525_SUM[11] , \524 );
_HMUX \U$1/U$12 ( \526 , \516 , \525_SUM[11] , \277 );
_DC \n5[12] ( \527_n5[12] , 1'b0 , 1'b1 );
or \U$5/U$13 ( \528 , \b[12] , \527_n5[12] );
buf \sub_5_33/A[12] ( \529_A[12] , \c[12] );
buf \sub_5_33/B[12] ( \530_B[12] , \d[12] );
not \sub_5_33/U$136 ( \531 , \530_B[12] );
xor \sub_5_33/U$135 ( \532 , \529_A[12] , \531 );
and \sub_5_33/U$140 ( \533 , \506_A[11] , \508 );
and \sub_5_33/U$139 ( \534 , \508 , \513 );
and \sub_5_33/U$138 ( \535 , \506_A[11] , \513 );
or \sub_5_33/U$137 ( \536 , \533 , \534 , \535 );
xor \sub_5_33/U$134 ( \537 , \532 , \536 );
buf \sub_5_33/SUM[12] ( \538_SUM[12] , \537 );
_HMUX \U$3/U$13 ( \539 , \528 , \538_SUM[12] , \241 );
buf \add_5_20/A[12] ( \540_A[12] , \c[12] );
buf \add_5_20/B[12] ( \541_B[12] , \d[12] );
xor \add_5_20/U$116 ( \542 , \540_A[12] , \541_B[12] );
and \add_5_20/U$120 ( \543 , \517_A[11] , \518_B[11] );
and \add_5_20/U$119 ( \544 , \518_B[11] , \523 );
and \add_5_20/U$118 ( \545 , \517_A[11] , \523 );
or \add_5_20/U$117 ( \546 , \543 , \544 , \545 );
xor \add_5_20/U$115 ( \547 , \542 , \546 );
buf \add_5_20/SUM[12] ( \548_SUM[12] , \547 );
_HMUX \U$1/U$13 ( \549 , \539 , \548_SUM[12] , \277 );
_DC \n5[13] ( \550_n5[13] , 1'b0 , 1'b1 );
or \U$5/U$14 ( \551 , \b[13] , \550_n5[13] );
buf \sub_5_33/A[13] ( \552_A[13] , \c[13] );
buf \sub_5_33/B[13] ( \553_B[13] , \d[13] );
not \sub_5_33/U$129 ( \554 , \553_B[13] );
xor \sub_5_33/U$128 ( \555 , \552_A[13] , \554 );
and \sub_5_33/U$133 ( \556 , \529_A[12] , \531 );
and \sub_5_33/U$132 ( \557 , \531 , \536 );
and \sub_5_33/U$131 ( \558 , \529_A[12] , \536 );
or \sub_5_33/U$130 ( \559 , \556 , \557 , \558 );
xor \sub_5_33/U$127 ( \560 , \555 , \559 );
buf \sub_5_33/SUM[13] ( \561_SUM[13] , \560 );
_HMUX \U$3/U$14 ( \562 , \551 , \561_SUM[13] , \241 );
buf \add_5_20/A[13] ( \563_A[13] , \c[13] );
buf \add_5_20/B[13] ( \564_B[13] , \d[13] );
xor \add_5_20/U$110 ( \565 , \563_A[13] , \564_B[13] );
and \add_5_20/U$114 ( \566 , \540_A[12] , \541_B[12] );
and \add_5_20/U$113 ( \567 , \541_B[12] , \546 );
and \add_5_20/U$112 ( \568 , \540_A[12] , \546 );
or \add_5_20/U$111 ( \569 , \566 , \567 , \568 );
xor \add_5_20/U$109 ( \570 , \565 , \569 );
buf \add_5_20/SUM[13] ( \571_SUM[13] , \570 );
_HMUX \U$1/U$14 ( \572 , \562 , \571_SUM[13] , \277 );
_DC \n5[14] ( \573_n5[14] , 1'b0 , 1'b1 );
or \U$5/U$15 ( \574 , \b[14] , \573_n5[14] );
buf \sub_5_33/A[14] ( \575_A[14] , \c[14] );
buf \sub_5_33/B[14] ( \576_B[14] , \d[14] );
not \sub_5_33/U$122 ( \577 , \576_B[14] );
xor \sub_5_33/U$121 ( \578 , \575_A[14] , \577 );
and \sub_5_33/U$126 ( \579 , \552_A[13] , \554 );
and \sub_5_33/U$125 ( \580 , \554 , \559 );
and \sub_5_33/U$124 ( \581 , \552_A[13] , \559 );
or \sub_5_33/U$123 ( \582 , \579 , \580 , \581 );
xor \sub_5_33/U$120 ( \583 , \578 , \582 );
buf \sub_5_33/SUM[14] ( \584_SUM[14] , \583 );
_HMUX \U$3/U$15 ( \585 , \574 , \584_SUM[14] , \241 );
buf \add_5_20/A[14] ( \586_A[14] , \c[14] );
buf \add_5_20/B[14] ( \587_B[14] , \d[14] );
xor \add_5_20/U$104 ( \588 , \586_A[14] , \587_B[14] );
and \add_5_20/U$108 ( \589 , \563_A[13] , \564_B[13] );
and \add_5_20/U$107 ( \590 , \564_B[13] , \569 );
and \add_5_20/U$106 ( \591 , \563_A[13] , \569 );
or \add_5_20/U$105 ( \592 , \589 , \590 , \591 );
xor \add_5_20/U$103 ( \593 , \588 , \592 );
buf \add_5_20/SUM[14] ( \594_SUM[14] , \593 );
_HMUX \U$1/U$15 ( \595 , \585 , \594_SUM[14] , \277 );
_DC \n5[15] ( \596_n5[15] , 1'b0 , 1'b1 );
or \U$5/U$16 ( \597 , \b[15] , \596_n5[15] );
buf \sub_5_33/A[15] ( \598_A[15] , \c[15] );
buf \sub_5_33/B[15] ( \599_B[15] , \d[15] );
not \sub_5_33/U$115 ( \600 , \599_B[15] );
xor \sub_5_33/U$114 ( \601 , \598_A[15] , \600 );
and \sub_5_33/U$119 ( \602 , \575_A[14] , \577 );
and \sub_5_33/U$118 ( \603 , \577 , \582 );
and \sub_5_33/U$117 ( \604 , \575_A[14] , \582 );
or \sub_5_33/U$116 ( \605 , \602 , \603 , \604 );
xor \sub_5_33/U$113 ( \606 , \601 , \605 );
buf \sub_5_33/SUM[15] ( \607_SUM[15] , \606 );
_HMUX \U$3/U$16 ( \608 , \597 , \607_SUM[15] , \241 );
buf \add_5_20/A[15] ( \609_A[15] , \c[15] );
buf \add_5_20/B[15] ( \610_B[15] , \d[15] );
xor \add_5_20/U$98 ( \611 , \609_A[15] , \610_B[15] );
and \add_5_20/U$102 ( \612 , \586_A[14] , \587_B[14] );
and \add_5_20/U$101 ( \613 , \587_B[14] , \592 );
and \add_5_20/U$100 ( \614 , \586_A[14] , \592 );
or \add_5_20/U$99 ( \615 , \612 , \613 , \614 );
xor \add_5_20/U$97 ( \616 , \611 , \615 );
buf \add_5_20/SUM[15] ( \617_SUM[15] , \616 );
_HMUX \U$1/U$16 ( \618 , \608 , \617_SUM[15] , \277 );
_DC \n5[16] ( \619_n5[16] , 1'b0 , 1'b1 );
or \U$5/U$17 ( \620 , \b[16] , \619_n5[16] );
buf \sub_5_33/A[16] ( \621_A[16] , \c[16] );
buf \sub_5_33/B[16] ( \622_B[16] , \d[16] );
not \sub_5_33/U$108 ( \623 , \622_B[16] );
xor \sub_5_33/U$107 ( \624 , \621_A[16] , \623 );
and \sub_5_33/U$112 ( \625 , \598_A[15] , \600 );
and \sub_5_33/U$111 ( \626 , \600 , \605 );
and \sub_5_33/U$110 ( \627 , \598_A[15] , \605 );
or \sub_5_33/U$109 ( \628 , \625 , \626 , \627 );
xor \sub_5_33/U$106 ( \629 , \624 , \628 );
buf \sub_5_33/SUM[16] ( \630_SUM[16] , \629 );
_HMUX \U$3/U$17 ( \631 , \620 , \630_SUM[16] , \241 );
buf \add_5_20/A[16] ( \632_A[16] , \c[16] );
buf \add_5_20/B[16] ( \633_B[16] , \d[16] );
xor \add_5_20/U$92 ( \634 , \632_A[16] , \633_B[16] );
and \add_5_20/U$96 ( \635 , \609_A[15] , \610_B[15] );
and \add_5_20/U$95 ( \636 , \610_B[15] , \615 );
and \add_5_20/U$94 ( \637 , \609_A[15] , \615 );
or \add_5_20/U$93 ( \638 , \635 , \636 , \637 );
xor \add_5_20/U$91 ( \639 , \634 , \638 );
buf \add_5_20/SUM[16] ( \640_SUM[16] , \639 );
_HMUX \U$1/U$17 ( \641 , \631 , \640_SUM[16] , \277 );
_DC \n5[17] ( \642_n5[17] , 1'b0 , 1'b1 );
or \U$5/U$18 ( \643 , \b[17] , \642_n5[17] );
buf \sub_5_33/A[17] ( \644_A[17] , \c[17] );
buf \sub_5_33/B[17] ( \645_B[17] , \d[17] );
not \sub_5_33/U$101 ( \646 , \645_B[17] );
xor \sub_5_33/U$100 ( \647 , \644_A[17] , \646 );
and \sub_5_33/U$105 ( \648 , \621_A[16] , \623 );
and \sub_5_33/U$104 ( \649 , \623 , \628 );
and \sub_5_33/U$103 ( \650 , \621_A[16] , \628 );
or \sub_5_33/U$102 ( \651 , \648 , \649 , \650 );
xor \sub_5_33/U$99 ( \652 , \647 , \651 );
buf \sub_5_33/SUM[17] ( \653_SUM[17] , \652 );
_HMUX \U$3/U$18 ( \654 , \643 , \653_SUM[17] , \241 );
buf \add_5_20/A[17] ( \655_A[17] , \c[17] );
buf \add_5_20/B[17] ( \656_B[17] , \d[17] );
xor \add_5_20/U$86 ( \657 , \655_A[17] , \656_B[17] );
and \add_5_20/U$90 ( \658 , \632_A[16] , \633_B[16] );
and \add_5_20/U$89 ( \659 , \633_B[16] , \638 );
and \add_5_20/U$88 ( \660 , \632_A[16] , \638 );
or \add_5_20/U$87 ( \661 , \658 , \659 , \660 );
xor \add_5_20/U$85 ( \662 , \657 , \661 );
buf \add_5_20/SUM[17] ( \663_SUM[17] , \662 );
_HMUX \U$1/U$18 ( \664 , \654 , \663_SUM[17] , \277 );
_DC \n5[18] ( \665_n5[18] , 1'b0 , 1'b1 );
or \U$5/U$19 ( \666 , \b[18] , \665_n5[18] );
buf \sub_5_33/A[18] ( \667_A[18] , \c[18] );
buf \sub_5_33/B[18] ( \668_B[18] , \d[18] );
not \sub_5_33/U$94 ( \669 , \668_B[18] );
xor \sub_5_33/U$93 ( \670 , \667_A[18] , \669 );
and \sub_5_33/U$98 ( \671 , \644_A[17] , \646 );
and \sub_5_33/U$97 ( \672 , \646 , \651 );
and \sub_5_33/U$96 ( \673 , \644_A[17] , \651 );
or \sub_5_33/U$95 ( \674 , \671 , \672 , \673 );
xor \sub_5_33/U$92 ( \675 , \670 , \674 );
buf \sub_5_33/SUM[18] ( \676_SUM[18] , \675 );
_HMUX \U$3/U$19 ( \677 , \666 , \676_SUM[18] , \241 );
buf \add_5_20/A[18] ( \678_A[18] , \c[18] );
buf \add_5_20/B[18] ( \679_B[18] , \d[18] );
xor \add_5_20/U$80 ( \680 , \678_A[18] , \679_B[18] );
and \add_5_20/U$84 ( \681 , \655_A[17] , \656_B[17] );
and \add_5_20/U$83 ( \682 , \656_B[17] , \661 );
and \add_5_20/U$82 ( \683 , \655_A[17] , \661 );
or \add_5_20/U$81 ( \684 , \681 , \682 , \683 );
xor \add_5_20/U$79 ( \685 , \680 , \684 );
buf \add_5_20/SUM[18] ( \686_SUM[18] , \685 );
_HMUX \U$1/U$19 ( \687 , \677 , \686_SUM[18] , \277 );
_DC \n5[19] ( \688_n5[19] , 1'b0 , 1'b1 );
or \U$5/U$20 ( \689 , \b[19] , \688_n5[19] );
buf \sub_5_33/A[19] ( \690_A[19] , \c[19] );
buf \sub_5_33/B[19] ( \691_B[19] , \d[19] );
not \sub_5_33/U$87 ( \692 , \691_B[19] );
xor \sub_5_33/U$86 ( \693 , \690_A[19] , \692 );
and \sub_5_33/U$91 ( \694 , \667_A[18] , \669 );
and \sub_5_33/U$90 ( \695 , \669 , \674 );
and \sub_5_33/U$89 ( \696 , \667_A[18] , \674 );
or \sub_5_33/U$88 ( \697 , \694 , \695 , \696 );
xor \sub_5_33/U$85 ( \698 , \693 , \697 );
buf \sub_5_33/SUM[19] ( \699_SUM[19] , \698 );
_HMUX \U$3/U$20 ( \700 , \689 , \699_SUM[19] , \241 );
buf \add_5_20/A[19] ( \701_A[19] , \c[19] );
buf \add_5_20/B[19] ( \702_B[19] , \d[19] );
xor \add_5_20/U$74 ( \703 , \701_A[19] , \702_B[19] );
and \add_5_20/U$78 ( \704 , \678_A[18] , \679_B[18] );
and \add_5_20/U$77 ( \705 , \679_B[18] , \684 );
and \add_5_20/U$76 ( \706 , \678_A[18] , \684 );
or \add_5_20/U$75 ( \707 , \704 , \705 , \706 );
xor \add_5_20/U$73 ( \708 , \703 , \707 );
buf \add_5_20/SUM[19] ( \709_SUM[19] , \708 );
_HMUX \U$1/U$20 ( \710 , \700 , \709_SUM[19] , \277 );
_DC \n5[20] ( \711_n5[20] , 1'b0 , 1'b1 );
or \U$5/U$21 ( \712 , \b[20] , \711_n5[20] );
buf \sub_5_33/A[20] ( \713_A[20] , \c[20] );
buf \sub_5_33/B[20] ( \714_B[20] , \d[20] );
not \sub_5_33/U$80 ( \715 , \714_B[20] );
xor \sub_5_33/U$79 ( \716 , \713_A[20] , \715 );
and \sub_5_33/U$84 ( \717 , \690_A[19] , \692 );
and \sub_5_33/U$83 ( \718 , \692 , \697 );
and \sub_5_33/U$82 ( \719 , \690_A[19] , \697 );
or \sub_5_33/U$81 ( \720 , \717 , \718 , \719 );
xor \sub_5_33/U$78 ( \721 , \716 , \720 );
buf \sub_5_33/SUM[20] ( \722_SUM[20] , \721 );
_HMUX \U$3/U$21 ( \723 , \712 , \722_SUM[20] , \241 );
buf \add_5_20/A[20] ( \724_A[20] , \c[20] );
buf \add_5_20/B[20] ( \725_B[20] , \d[20] );
xor \add_5_20/U$68 ( \726 , \724_A[20] , \725_B[20] );
and \add_5_20/U$72 ( \727 , \701_A[19] , \702_B[19] );
and \add_5_20/U$71 ( \728 , \702_B[19] , \707 );
and \add_5_20/U$70 ( \729 , \701_A[19] , \707 );
or \add_5_20/U$69 ( \730 , \727 , \728 , \729 );
xor \add_5_20/U$67 ( \731 , \726 , \730 );
buf \add_5_20/SUM[20] ( \732_SUM[20] , \731 );
_HMUX \U$1/U$21 ( \733 , \723 , \732_SUM[20] , \277 );
_DC \n5[21] ( \734_n5[21] , 1'b0 , 1'b1 );
or \U$5/U$22 ( \735 , \b[21] , \734_n5[21] );
buf \sub_5_33/A[21] ( \736_A[21] , \c[21] );
buf \sub_5_33/B[21] ( \737_B[21] , \d[21] );
not \sub_5_33/U$73 ( \738 , \737_B[21] );
xor \sub_5_33/U$72 ( \739 , \736_A[21] , \738 );
and \sub_5_33/U$77 ( \740 , \713_A[20] , \715 );
and \sub_5_33/U$76 ( \741 , \715 , \720 );
and \sub_5_33/U$75 ( \742 , \713_A[20] , \720 );
or \sub_5_33/U$74 ( \743 , \740 , \741 , \742 );
xor \sub_5_33/U$71 ( \744 , \739 , \743 );
buf \sub_5_33/SUM[21] ( \745_SUM[21] , \744 );
_HMUX \U$3/U$22 ( \746 , \735 , \745_SUM[21] , \241 );
buf \add_5_20/A[21] ( \747_A[21] , \c[21] );
buf \add_5_20/B[21] ( \748_B[21] , \d[21] );
xor \add_5_20/U$62 ( \749 , \747_A[21] , \748_B[21] );
and \add_5_20/U$66 ( \750 , \724_A[20] , \725_B[20] );
and \add_5_20/U$65 ( \751 , \725_B[20] , \730 );
and \add_5_20/U$64 ( \752 , \724_A[20] , \730 );
or \add_5_20/U$63 ( \753 , \750 , \751 , \752 );
xor \add_5_20/U$61 ( \754 , \749 , \753 );
buf \add_5_20/SUM[21] ( \755_SUM[21] , \754 );
_HMUX \U$1/U$22 ( \756 , \746 , \755_SUM[21] , \277 );
_DC \n5[22] ( \757_n5[22] , 1'b0 , 1'b1 );
or \U$5/U$23 ( \758 , \b[22] , \757_n5[22] );
buf \sub_5_33/A[22] ( \759_A[22] , \c[22] );
buf \sub_5_33/B[22] ( \760_B[22] , \d[22] );
not \sub_5_33/U$66 ( \761 , \760_B[22] );
xor \sub_5_33/U$65 ( \762 , \759_A[22] , \761 );
and \sub_5_33/U$70 ( \763 , \736_A[21] , \738 );
and \sub_5_33/U$69 ( \764 , \738 , \743 );
and \sub_5_33/U$68 ( \765 , \736_A[21] , \743 );
or \sub_5_33/U$67 ( \766 , \763 , \764 , \765 );
xor \sub_5_33/U$64 ( \767 , \762 , \766 );
buf \sub_5_33/SUM[22] ( \768_SUM[22] , \767 );
_HMUX \U$3/U$23 ( \769 , \758 , \768_SUM[22] , \241 );
buf \add_5_20/A[22] ( \770_A[22] , \c[22] );
buf \add_5_20/B[22] ( \771_B[22] , \d[22] );
xor \add_5_20/U$56 ( \772 , \770_A[22] , \771_B[22] );
and \add_5_20/U$60 ( \773 , \747_A[21] , \748_B[21] );
and \add_5_20/U$59 ( \774 , \748_B[21] , \753 );
and \add_5_20/U$58 ( \775 , \747_A[21] , \753 );
or \add_5_20/U$57 ( \776 , \773 , \774 , \775 );
xor \add_5_20/U$55 ( \777 , \772 , \776 );
buf \add_5_20/SUM[22] ( \778_SUM[22] , \777 );
_HMUX \U$1/U$23 ( \779 , \769 , \778_SUM[22] , \277 );
_DC \n5[23] ( \780_n5[23] , 1'b0 , 1'b1 );
or \U$5/U$24 ( \781 , \b[23] , \780_n5[23] );
buf \sub_5_33/A[23] ( \782_A[23] , \c[23] );
buf \sub_5_33/B[23] ( \783_B[23] , \d[23] );
not \sub_5_33/U$59 ( \784 , \783_B[23] );
xor \sub_5_33/U$58 ( \785 , \782_A[23] , \784 );
and \sub_5_33/U$63 ( \786 , \759_A[22] , \761 );
and \sub_5_33/U$62 ( \787 , \761 , \766 );
and \sub_5_33/U$61 ( \788 , \759_A[22] , \766 );
or \sub_5_33/U$60 ( \789 , \786 , \787 , \788 );
xor \sub_5_33/U$57 ( \790 , \785 , \789 );
buf \sub_5_33/SUM[23] ( \791_SUM[23] , \790 );
_HMUX \U$3/U$24 ( \792 , \781 , \791_SUM[23] , \241 );
buf \add_5_20/A[23] ( \793_A[23] , \c[23] );
buf \add_5_20/B[23] ( \794_B[23] , \d[23] );
xor \add_5_20/U$50 ( \795 , \793_A[23] , \794_B[23] );
and \add_5_20/U$54 ( \796 , \770_A[22] , \771_B[22] );
and \add_5_20/U$53 ( \797 , \771_B[22] , \776 );
and \add_5_20/U$52 ( \798 , \770_A[22] , \776 );
or \add_5_20/U$51 ( \799 , \796 , \797 , \798 );
xor \add_5_20/U$49 ( \800 , \795 , \799 );
buf \add_5_20/SUM[23] ( \801_SUM[23] , \800 );
_HMUX \U$1/U$24 ( \802 , \792 , \801_SUM[23] , \277 );
_DC \n5[24] ( \803_n5[24] , 1'b0 , 1'b1 );
or \U$5/U$25 ( \804 , \b[24] , \803_n5[24] );
buf \sub_5_33/A[24] ( \805_A[24] , \c[24] );
buf \sub_5_33/B[24] ( \806_B[24] , \d[24] );
not \sub_5_33/U$52 ( \807 , \806_B[24] );
xor \sub_5_33/U$51 ( \808 , \805_A[24] , \807 );
and \sub_5_33/U$56 ( \809 , \782_A[23] , \784 );
and \sub_5_33/U$55 ( \810 , \784 , \789 );
and \sub_5_33/U$54 ( \811 , \782_A[23] , \789 );
or \sub_5_33/U$53 ( \812 , \809 , \810 , \811 );
xor \sub_5_33/U$50 ( \813 , \808 , \812 );
buf \sub_5_33/SUM[24] ( \814_SUM[24] , \813 );
_HMUX \U$3/U$25 ( \815 , \804 , \814_SUM[24] , \241 );
buf \add_5_20/A[24] ( \816_A[24] , \c[24] );
buf \add_5_20/B[24] ( \817_B[24] , \d[24] );
xor \add_5_20/U$44 ( \818 , \816_A[24] , \817_B[24] );
and \add_5_20/U$48 ( \819 , \793_A[23] , \794_B[23] );
and \add_5_20/U$47 ( \820 , \794_B[23] , \799 );
and \add_5_20/U$46 ( \821 , \793_A[23] , \799 );
or \add_5_20/U$45 ( \822 , \819 , \820 , \821 );
xor \add_5_20/U$43 ( \823 , \818 , \822 );
buf \add_5_20/SUM[24] ( \824_SUM[24] , \823 );
_HMUX \U$1/U$25 ( \825 , \815 , \824_SUM[24] , \277 );
_DC \n5[25] ( \826_n5[25] , 1'b0 , 1'b1 );
or \U$5/U$26 ( \827 , \b[25] , \826_n5[25] );
buf \sub_5_33/A[25] ( \828_A[25] , \c[25] );
buf \sub_5_33/B[25] ( \829_B[25] , \d[25] );
not \sub_5_33/U$45 ( \830 , \829_B[25] );
xor \sub_5_33/U$44 ( \831 , \828_A[25] , \830 );
and \sub_5_33/U$49 ( \832 , \805_A[24] , \807 );
and \sub_5_33/U$48 ( \833 , \807 , \812 );
and \sub_5_33/U$47 ( \834 , \805_A[24] , \812 );
or \sub_5_33/U$46 ( \835 , \832 , \833 , \834 );
xor \sub_5_33/U$43 ( \836 , \831 , \835 );
buf \sub_5_33/SUM[25] ( \837_SUM[25] , \836 );
_HMUX \U$3/U$26 ( \838 , \827 , \837_SUM[25] , \241 );
buf \add_5_20/A[25] ( \839_A[25] , \c[25] );
buf \add_5_20/B[25] ( \840_B[25] , \d[25] );
xor \add_5_20/U$38 ( \841 , \839_A[25] , \840_B[25] );
and \add_5_20/U$42 ( \842 , \816_A[24] , \817_B[24] );
and \add_5_20/U$41 ( \843 , \817_B[24] , \822 );
and \add_5_20/U$40 ( \844 , \816_A[24] , \822 );
or \add_5_20/U$39 ( \845 , \842 , \843 , \844 );
xor \add_5_20/U$37 ( \846 , \841 , \845 );
buf \add_5_20/SUM[25] ( \847_SUM[25] , \846 );
_HMUX \U$1/U$26 ( \848 , \838 , \847_SUM[25] , \277 );
_DC \n5[26] ( \849_n5[26] , 1'b0 , 1'b1 );
or \U$5/U$27 ( \850 , \b[26] , \849_n5[26] );
buf \sub_5_33/A[26] ( \851_A[26] , \c[26] );
buf \sub_5_33/B[26] ( \852_B[26] , \d[26] );
not \sub_5_33/U$38 ( \853 , \852_B[26] );
xor \sub_5_33/U$37 ( \854 , \851_A[26] , \853 );
and \sub_5_33/U$42 ( \855 , \828_A[25] , \830 );
and \sub_5_33/U$41 ( \856 , \830 , \835 );
and \sub_5_33/U$40 ( \857 , \828_A[25] , \835 );
or \sub_5_33/U$39 ( \858 , \855 , \856 , \857 );
xor \sub_5_33/U$36 ( \859 , \854 , \858 );
buf \sub_5_33/SUM[26] ( \860_SUM[26] , \859 );
_HMUX \U$3/U$27 ( \861 , \850 , \860_SUM[26] , \241 );
buf \add_5_20/A[26] ( \862_A[26] , \c[26] );
buf \add_5_20/B[26] ( \863_B[26] , \d[26] );
xor \add_5_20/U$32 ( \864 , \862_A[26] , \863_B[26] );
and \add_5_20/U$36 ( \865 , \839_A[25] , \840_B[25] );
and \add_5_20/U$35 ( \866 , \840_B[25] , \845 );
and \add_5_20/U$34 ( \867 , \839_A[25] , \845 );
or \add_5_20/U$33 ( \868 , \865 , \866 , \867 );
xor \add_5_20/U$31 ( \869 , \864 , \868 );
buf \add_5_20/SUM[26] ( \870_SUM[26] , \869 );
_HMUX \U$1/U$27 ( \871 , \861 , \870_SUM[26] , \277 );
_DC \n5[27] ( \872_n5[27] , 1'b0 , 1'b1 );
or \U$5/U$28 ( \873 , \b[27] , \872_n5[27] );
buf \sub_5_33/A[27] ( \874_A[27] , \c[27] );
buf \sub_5_33/B[27] ( \875_B[27] , \d[27] );
not \sub_5_33/U$31 ( \876 , \875_B[27] );
xor \sub_5_33/U$30 ( \877 , \874_A[27] , \876 );
and \sub_5_33/U$35 ( \878 , \851_A[26] , \853 );
and \sub_5_33/U$34 ( \879 , \853 , \858 );
and \sub_5_33/U$33 ( \880 , \851_A[26] , \858 );
or \sub_5_33/U$32 ( \881 , \878 , \879 , \880 );
xor \sub_5_33/U$29 ( \882 , \877 , \881 );
buf \sub_5_33/SUM[27] ( \883_SUM[27] , \882 );
_HMUX \U$3/U$28 ( \884 , \873 , \883_SUM[27] , \241 );
buf \add_5_20/A[27] ( \885_A[27] , \c[27] );
buf \add_5_20/B[27] ( \886_B[27] , \d[27] );
xor \add_5_20/U$26 ( \887 , \885_A[27] , \886_B[27] );
and \add_5_20/U$30 ( \888 , \862_A[26] , \863_B[26] );
and \add_5_20/U$29 ( \889 , \863_B[26] , \868 );
and \add_5_20/U$28 ( \890 , \862_A[26] , \868 );
or \add_5_20/U$27 ( \891 , \888 , \889 , \890 );
xor \add_5_20/U$25 ( \892 , \887 , \891 );
buf \add_5_20/SUM[27] ( \893_SUM[27] , \892 );
_HMUX \U$1/U$28 ( \894 , \884 , \893_SUM[27] , \277 );
_DC \n5[28] ( \895_n5[28] , 1'b0 , 1'b1 );
or \U$5/U$29 ( \896 , \b[28] , \895_n5[28] );
buf \sub_5_33/A[28] ( \897_A[28] , \c[28] );
buf \sub_5_33/B[28] ( \898_B[28] , \d[28] );
not \sub_5_33/U$24 ( \899 , \898_B[28] );
xor \sub_5_33/U$23 ( \900 , \897_A[28] , \899 );
and \sub_5_33/U$28 ( \901 , \874_A[27] , \876 );
and \sub_5_33/U$27 ( \902 , \876 , \881 );
and \sub_5_33/U$26 ( \903 , \874_A[27] , \881 );
or \sub_5_33/U$25 ( \904 , \901 , \902 , \903 );
xor \sub_5_33/U$22 ( \905 , \900 , \904 );
buf \sub_5_33/SUM[28] ( \906_SUM[28] , \905 );
_HMUX \U$3/U$29 ( \907 , \896 , \906_SUM[28] , \241 );
buf \add_5_20/A[28] ( \908_A[28] , \c[28] );
buf \add_5_20/B[28] ( \909_B[28] , \d[28] );
xor \add_5_20/U$20 ( \910 , \908_A[28] , \909_B[28] );
and \add_5_20/U$24 ( \911 , \885_A[27] , \886_B[27] );
and \add_5_20/U$23 ( \912 , \886_B[27] , \891 );
and \add_5_20/U$22 ( \913 , \885_A[27] , \891 );
or \add_5_20/U$21 ( \914 , \911 , \912 , \913 );
xor \add_5_20/U$19 ( \915 , \910 , \914 );
buf \add_5_20/SUM[28] ( \916_SUM[28] , \915 );
_HMUX \U$1/U$29 ( \917 , \907 , \916_SUM[28] , \277 );
_DC \n5[29] ( \918_n5[29] , 1'b0 , 1'b1 );
or \U$5/U$30 ( \919 , \b[29] , \918_n5[29] );
buf \sub_5_33/A[29] ( \920_A[29] , \c[29] );
buf \sub_5_33/B[29] ( \921_B[29] , \d[29] );
not \sub_5_33/U$17 ( \922 , \921_B[29] );
xor \sub_5_33/U$16 ( \923 , \920_A[29] , \922 );
and \sub_5_33/U$21 ( \924 , \897_A[28] , \899 );
and \sub_5_33/U$20 ( \925 , \899 , \904 );
and \sub_5_33/U$19 ( \926 , \897_A[28] , \904 );
or \sub_5_33/U$18 ( \927 , \924 , \925 , \926 );
xor \sub_5_33/U$15 ( \928 , \923 , \927 );
buf \sub_5_33/SUM[29] ( \929_SUM[29] , \928 );
_HMUX \U$3/U$30 ( \930 , \919 , \929_SUM[29] , \241 );
buf \add_5_20/A[29] ( \931_A[29] , \c[29] );
buf \add_5_20/B[29] ( \932_B[29] , \d[29] );
xor \add_5_20/U$14 ( \933 , \931_A[29] , \932_B[29] );
and \add_5_20/U$18 ( \934 , \908_A[28] , \909_B[28] );
and \add_5_20/U$17 ( \935 , \909_B[28] , \914 );
and \add_5_20/U$16 ( \936 , \908_A[28] , \914 );
or \add_5_20/U$15 ( \937 , \934 , \935 , \936 );
xor \add_5_20/U$13 ( \938 , \933 , \937 );
buf \add_5_20/SUM[29] ( \939_SUM[29] , \938 );
_HMUX \U$1/U$30 ( \940 , \930 , \939_SUM[29] , \277 );
_DC \n5[30] ( \941_n5[30] , 1'b0 , 1'b1 );
or \U$5/U$31 ( \942 , \b[30] , \941_n5[30] );
buf \sub_5_33/A[30] ( \943_A[30] , \c[30] );
buf \sub_5_33/B[30] ( \944_B[30] , \d[30] );
not \sub_5_33/U$10 ( \945 , \944_B[30] );
xor \sub_5_33/U$9 ( \946 , \943_A[30] , \945 );
and \sub_5_33/U$14 ( \947 , \920_A[29] , \922 );
and \sub_5_33/U$13 ( \948 , \922 , \927 );
and \sub_5_33/U$12 ( \949 , \920_A[29] , \927 );
or \sub_5_33/U$11 ( \950 , \947 , \948 , \949 );
xor \sub_5_33/U$8 ( \951 , \946 , \950 );
buf \sub_5_33/SUM[30] ( \952_SUM[30] , \951 );
_HMUX \U$3/U$31 ( \953 , \942 , \952_SUM[30] , \241 );
buf \add_5_20/A[30] ( \954_A[30] , \c[30] );
buf \add_5_20/B[30] ( \955_B[30] , \d[30] );
xor \add_5_20/U$8 ( \956 , \954_A[30] , \955_B[30] );
and \add_5_20/U$12 ( \957 , \931_A[29] , \932_B[29] );
and \add_5_20/U$11 ( \958 , \932_B[29] , \937 );
and \add_5_20/U$10 ( \959 , \931_A[29] , \937 );
or \add_5_20/U$9 ( \960 , \957 , \958 , \959 );
xor \add_5_20/U$7 ( \961 , \956 , \960 );
buf \add_5_20/SUM[30] ( \962_SUM[30] , \961 );
_HMUX \U$1/U$31 ( \963 , \953 , \962_SUM[30] , \277 );
_DC \n5[31] ( \964_n5[31] , 1'b0 , 1'b1 );
or \U$5/U$32 ( \965 , \b[31] , \964_n5[31] );
buf \sub_5_33/A[31] ( \966_A[31] , \c[31] );
buf \sub_5_33/B[31] ( \967_B[31] , \d[31] );
not \sub_5_33/U$3 ( \968 , \967_B[31] );
xor \sub_5_33/U$2 ( \969 , \966_A[31] , \968 );
and \sub_5_33/U$7 ( \970 , \943_A[30] , \945 );
and \sub_5_33/U$6 ( \971 , \945 , \950 );
and \sub_5_33/U$5 ( \972 , \943_A[30] , \950 );
or \sub_5_33/U$4 ( \973 , \970 , \971 , \972 );
xor \sub_5_33/U$1 ( \974 , \969 , \973 );
buf \sub_5_33/SUM[31] ( \975_SUM[31] , \974 );
_HMUX \U$3/U$32 ( \976 , \965 , \975_SUM[31] , \241 );
buf \add_5_20/A[31] ( \977_A[31] , \c[31] );
buf \add_5_20/B[31] ( \978_B[31] , \d[31] );
xor \add_5_20/U$2 ( \979 , \977_A[31] , \978_B[31] );
and \add_5_20/U$6 ( \980 , \954_A[30] , \955_B[30] );
and \add_5_20/U$5 ( \981 , \955_B[30] , \960 );
and \add_5_20/U$4 ( \982 , \954_A[30] , \960 );
or \add_5_20/U$3 ( \983 , \980 , \981 , \982 );
xor \add_5_20/U$1 ( \984 , \979 , \983 );
buf \add_5_20/SUM[31] ( \985_SUM[31] , \984 );
_HMUX \U$1/U$32 ( \986 , \976 , \985_SUM[31] , \277 );
buf \add_6_14/A[31] ( \987_A[31] , \a[31] );
buf \add_6_14/B[31] ( \988_B[31] , \b[31] );
xor \add_6_14/U$2 ( \989 , \987_A[31] , \988_B[31] );
buf \add_6_14/A[30] ( \990_A[30] , \a[30] );
buf \add_6_14/B[30] ( \991_B[30] , \b[30] );
and \add_6_14/U$6 ( \992 , \990_A[30] , \991_B[30] );
buf \add_6_14/A[29] ( \993_A[29] , \a[29] );
buf \add_6_14/B[29] ( \994_B[29] , \b[29] );
and \add_6_14/U$12 ( \995 , \993_A[29] , \994_B[29] );
buf \add_6_14/A[28] ( \996_A[28] , \a[28] );
buf \add_6_14/B[28] ( \997_B[28] , \b[28] );
and \add_6_14/U$18 ( \998 , \996_A[28] , \997_B[28] );
buf \add_6_14/A[27] ( \999_A[27] , \a[27] );
buf \add_6_14/B[27] ( \1000_B[27] , \b[27] );
and \add_6_14/U$24 ( \1001 , \999_A[27] , \1000_B[27] );
buf \add_6_14/A[26] ( \1002_A[26] , \a[26] );
buf \add_6_14/B[26] ( \1003_B[26] , \b[26] );
and \add_6_14/U$30 ( \1004 , \1002_A[26] , \1003_B[26] );
buf \add_6_14/A[25] ( \1005_A[25] , \a[25] );
buf \add_6_14/B[25] ( \1006_B[25] , \b[25] );
and \add_6_14/U$36 ( \1007 , \1005_A[25] , \1006_B[25] );
buf \add_6_14/A[24] ( \1008_A[24] , \a[24] );
buf \add_6_14/B[24] ( \1009_B[24] , \b[24] );
and \add_6_14/U$42 ( \1010 , \1008_A[24] , \1009_B[24] );
buf \add_6_14/A[23] ( \1011_A[23] , \a[23] );
buf \add_6_14/B[23] ( \1012_B[23] , \b[23] );
and \add_6_14/U$48 ( \1013 , \1011_A[23] , \1012_B[23] );
buf \add_6_14/A[22] ( \1014_A[22] , \a[22] );
buf \add_6_14/B[22] ( \1015_B[22] , \b[22] );
and \add_6_14/U$54 ( \1016 , \1014_A[22] , \1015_B[22] );
buf \add_6_14/A[21] ( \1017_A[21] , \a[21] );
buf \add_6_14/B[21] ( \1018_B[21] , \b[21] );
and \add_6_14/U$60 ( \1019 , \1017_A[21] , \1018_B[21] );
buf \add_6_14/A[20] ( \1020_A[20] , \a[20] );
buf \add_6_14/B[20] ( \1021_B[20] , \b[20] );
and \add_6_14/U$66 ( \1022 , \1020_A[20] , \1021_B[20] );
buf \add_6_14/A[19] ( \1023_A[19] , \a[19] );
buf \add_6_14/B[19] ( \1024_B[19] , \b[19] );
and \add_6_14/U$72 ( \1025 , \1023_A[19] , \1024_B[19] );
buf \add_6_14/A[18] ( \1026_A[18] , \a[18] );
buf \add_6_14/B[18] ( \1027_B[18] , \b[18] );
and \add_6_14/U$78 ( \1028 , \1026_A[18] , \1027_B[18] );
buf \add_6_14/A[17] ( \1029_A[17] , \a[17] );
buf \add_6_14/B[17] ( \1030_B[17] , \b[17] );
and \add_6_14/U$84 ( \1031 , \1029_A[17] , \1030_B[17] );
buf \add_6_14/A[16] ( \1032_A[16] , \a[16] );
buf \add_6_14/B[16] ( \1033_B[16] , \b[16] );
and \add_6_14/U$90 ( \1034 , \1032_A[16] , \1033_B[16] );
buf \add_6_14/A[15] ( \1035_A[15] , \a[15] );
buf \add_6_14/B[15] ( \1036_B[15] , \b[15] );
and \add_6_14/U$96 ( \1037 , \1035_A[15] , \1036_B[15] );
buf \add_6_14/A[14] ( \1038_A[14] , \a[14] );
buf \add_6_14/B[14] ( \1039_B[14] , \b[14] );
and \add_6_14/U$102 ( \1040 , \1038_A[14] , \1039_B[14] );
buf \add_6_14/A[13] ( \1041_A[13] , \a[13] );
buf \add_6_14/B[13] ( \1042_B[13] , \b[13] );
and \add_6_14/U$108 ( \1043 , \1041_A[13] , \1042_B[13] );
buf \add_6_14/A[12] ( \1044_A[12] , \a[12] );
buf \add_6_14/B[12] ( \1045_B[12] , \b[12] );
and \add_6_14/U$114 ( \1046 , \1044_A[12] , \1045_B[12] );
buf \add_6_14/A[11] ( \1047_A[11] , \a[11] );
buf \add_6_14/B[11] ( \1048_B[11] , \b[11] );
and \add_6_14/U$120 ( \1049 , \1047_A[11] , \1048_B[11] );
buf \add_6_14/A[10] ( \1050_A[10] , \a[10] );
buf \add_6_14/B[10] ( \1051_B[10] , \b[10] );
and \add_6_14/U$126 ( \1052 , \1050_A[10] , \1051_B[10] );
buf \add_6_14/A[9] ( \1053_A[9] , \a[9] );
buf \add_6_14/B[9] ( \1054_B[9] , \b[9] );
and \add_6_14/U$132 ( \1055 , \1053_A[9] , \1054_B[9] );
buf \add_6_14/A[8] ( \1056_A[8] , \a[8] );
buf \add_6_14/B[8] ( \1057_B[8] , \b[8] );
and \add_6_14/U$138 ( \1058 , \1056_A[8] , \1057_B[8] );
buf \add_6_14/A[7] ( \1059_A[7] , \a[7] );
buf \add_6_14/B[7] ( \1060_B[7] , \b[7] );
and \add_6_14/U$144 ( \1061 , \1059_A[7] , \1060_B[7] );
buf \add_6_14/A[6] ( \1062_A[6] , \a[6] );
buf \add_6_14/B[6] ( \1063_B[6] , \b[6] );
and \add_6_14/U$150 ( \1064 , \1062_A[6] , \1063_B[6] );
buf \add_6_14/A[5] ( \1065_A[5] , \a[5] );
buf \add_6_14/B[5] ( \1066_B[5] , \b[5] );
and \add_6_14/U$156 ( \1067 , \1065_A[5] , \1066_B[5] );
buf \add_6_14/A[4] ( \1068_A[4] , \a[4] );
buf \add_6_14/B[4] ( \1069_B[4] , \b[4] );
and \add_6_14/U$162 ( \1070 , \1068_A[4] , \1069_B[4] );
buf \add_6_14/A[3] ( \1071_A[3] , \a[3] );
buf \add_6_14/B[3] ( \1072_B[3] , \b[3] );
and \add_6_14/U$168 ( \1073 , \1071_A[3] , \1072_B[3] );
buf \add_6_14/A[2] ( \1074_A[2] , \a[2] );
buf \add_6_14/B[2] ( \1075_B[2] , \b[2] );
and \add_6_14/U$174 ( \1076 , \1074_A[2] , \1075_B[2] );
buf \add_6_14/A[1] ( \1077_A[1] , \a[1] );
buf \add_6_14/B[1] ( \1078_B[1] , \b[1] );
and \add_6_14/U$180 ( \1079 , \1077_A[1] , \1078_B[1] );
buf \add_6_14/A[0] ( \1080_A[0] , \a[0] );
buf \add_6_14/B[0] ( \1081_B[0] , \b[0] );
and \add_6_14/U$183 ( \1082 , \1080_A[0] , \1081_B[0] );
and \add_6_14/U$179 ( \1083 , \1078_B[1] , \1082 );
and \add_6_14/U$178 ( \1084 , \1077_A[1] , \1082 );
or \add_6_14/U$177 ( \1085 , \1079 , \1083 , \1084 );
and \add_6_14/U$173 ( \1086 , \1075_B[2] , \1085 );
and \add_6_14/U$172 ( \1087 , \1074_A[2] , \1085 );
or \add_6_14/U$171 ( \1088 , \1076 , \1086 , \1087 );
and \add_6_14/U$167 ( \1089 , \1072_B[3] , \1088 );
and \add_6_14/U$166 ( \1090 , \1071_A[3] , \1088 );
or \add_6_14/U$165 ( \1091 , \1073 , \1089 , \1090 );
and \add_6_14/U$161 ( \1092 , \1069_B[4] , \1091 );
and \add_6_14/U$160 ( \1093 , \1068_A[4] , \1091 );
or \add_6_14/U$159 ( \1094 , \1070 , \1092 , \1093 );
and \add_6_14/U$155 ( \1095 , \1066_B[5] , \1094 );
and \add_6_14/U$154 ( \1096 , \1065_A[5] , \1094 );
or \add_6_14/U$153 ( \1097 , \1067 , \1095 , \1096 );
and \add_6_14/U$149 ( \1098 , \1063_B[6] , \1097 );
and \add_6_14/U$148 ( \1099 , \1062_A[6] , \1097 );
or \add_6_14/U$147 ( \1100 , \1064 , \1098 , \1099 );
and \add_6_14/U$143 ( \1101 , \1060_B[7] , \1100 );
and \add_6_14/U$142 ( \1102 , \1059_A[7] , \1100 );
or \add_6_14/U$141 ( \1103 , \1061 , \1101 , \1102 );
and \add_6_14/U$137 ( \1104 , \1057_B[8] , \1103 );
and \add_6_14/U$136 ( \1105 , \1056_A[8] , \1103 );
or \add_6_14/U$135 ( \1106 , \1058 , \1104 , \1105 );
and \add_6_14/U$131 ( \1107 , \1054_B[9] , \1106 );
and \add_6_14/U$130 ( \1108 , \1053_A[9] , \1106 );
or \add_6_14/U$129 ( \1109 , \1055 , \1107 , \1108 );
and \add_6_14/U$125 ( \1110 , \1051_B[10] , \1109 );
and \add_6_14/U$124 ( \1111 , \1050_A[10] , \1109 );
or \add_6_14/U$123 ( \1112 , \1052 , \1110 , \1111 );
and \add_6_14/U$119 ( \1113 , \1048_B[11] , \1112 );
and \add_6_14/U$118 ( \1114 , \1047_A[11] , \1112 );
or \add_6_14/U$117 ( \1115 , \1049 , \1113 , \1114 );
and \add_6_14/U$113 ( \1116 , \1045_B[12] , \1115 );
and \add_6_14/U$112 ( \1117 , \1044_A[12] , \1115 );
or \add_6_14/U$111 ( \1118 , \1046 , \1116 , \1117 );
and \add_6_14/U$107 ( \1119 , \1042_B[13] , \1118 );
and \add_6_14/U$106 ( \1120 , \1041_A[13] , \1118 );
or \add_6_14/U$105 ( \1121 , \1043 , \1119 , \1120 );
and \add_6_14/U$101 ( \1122 , \1039_B[14] , \1121 );
and \add_6_14/U$100 ( \1123 , \1038_A[14] , \1121 );
or \add_6_14/U$99 ( \1124 , \1040 , \1122 , \1123 );
and \add_6_14/U$95 ( \1125 , \1036_B[15] , \1124 );
and \add_6_14/U$94 ( \1126 , \1035_A[15] , \1124 );
or \add_6_14/U$93 ( \1127 , \1037 , \1125 , \1126 );
and \add_6_14/U$89 ( \1128 , \1033_B[16] , \1127 );
and \add_6_14/U$88 ( \1129 , \1032_A[16] , \1127 );
or \add_6_14/U$87 ( \1130 , \1034 , \1128 , \1129 );
and \add_6_14/U$83 ( \1131 , \1030_B[17] , \1130 );
and \add_6_14/U$82 ( \1132 , \1029_A[17] , \1130 );
or \add_6_14/U$81 ( \1133 , \1031 , \1131 , \1132 );
and \add_6_14/U$77 ( \1134 , \1027_B[18] , \1133 );
and \add_6_14/U$76 ( \1135 , \1026_A[18] , \1133 );
or \add_6_14/U$75 ( \1136 , \1028 , \1134 , \1135 );
and \add_6_14/U$71 ( \1137 , \1024_B[19] , \1136 );
and \add_6_14/U$70 ( \1138 , \1023_A[19] , \1136 );
or \add_6_14/U$69 ( \1139 , \1025 , \1137 , \1138 );
and \add_6_14/U$65 ( \1140 , \1021_B[20] , \1139 );
and \add_6_14/U$64 ( \1141 , \1020_A[20] , \1139 );
or \add_6_14/U$63 ( \1142 , \1022 , \1140 , \1141 );
and \add_6_14/U$59 ( \1143 , \1018_B[21] , \1142 );
and \add_6_14/U$58 ( \1144 , \1017_A[21] , \1142 );
or \add_6_14/U$57 ( \1145 , \1019 , \1143 , \1144 );
and \add_6_14/U$53 ( \1146 , \1015_B[22] , \1145 );
and \add_6_14/U$52 ( \1147 , \1014_A[22] , \1145 );
or \add_6_14/U$51 ( \1148 , \1016 , \1146 , \1147 );
and \add_6_14/U$47 ( \1149 , \1012_B[23] , \1148 );
and \add_6_14/U$46 ( \1150 , \1011_A[23] , \1148 );
or \add_6_14/U$45 ( \1151 , \1013 , \1149 , \1150 );
and \add_6_14/U$41 ( \1152 , \1009_B[24] , \1151 );
and \add_6_14/U$40 ( \1153 , \1008_A[24] , \1151 );
or \add_6_14/U$39 ( \1154 , \1010 , \1152 , \1153 );
and \add_6_14/U$35 ( \1155 , \1006_B[25] , \1154 );
and \add_6_14/U$34 ( \1156 , \1005_A[25] , \1154 );
or \add_6_14/U$33 ( \1157 , \1007 , \1155 , \1156 );
and \add_6_14/U$29 ( \1158 , \1003_B[26] , \1157 );
and \add_6_14/U$28 ( \1159 , \1002_A[26] , \1157 );
or \add_6_14/U$27 ( \1160 , \1004 , \1158 , \1159 );
and \add_6_14/U$23 ( \1161 , \1000_B[27] , \1160 );
and \add_6_14/U$22 ( \1162 , \999_A[27] , \1160 );
or \add_6_14/U$21 ( \1163 , \1001 , \1161 , \1162 );
and \add_6_14/U$17 ( \1164 , \997_B[28] , \1163 );
and \add_6_14/U$16 ( \1165 , \996_A[28] , \1163 );
or \add_6_14/U$15 ( \1166 , \998 , \1164 , \1165 );
and \add_6_14/U$11 ( \1167 , \994_B[29] , \1166 );
and \add_6_14/U$10 ( \1168 , \993_A[29] , \1166 );
or \add_6_14/U$9 ( \1169 , \995 , \1167 , \1168 );
and \add_6_14/U$5 ( \1170 , \991_B[30] , \1169 );
and \add_6_14/U$4 ( \1171 , \990_A[30] , \1169 );
or \add_6_14/U$3 ( \1172 , \992 , \1170 , \1171 );
xor \add_6_14/U$1 ( \1173 , \989 , \1172 );
buf \add_6_14/SUM[31] ( \1174_SUM[31] , \1173 );
buf \mul_6_18/A[31] ( \1175_A[31] , \1174_SUM[31] );
xor \add_6_14/U$8 ( \1176 , \990_A[30] , \991_B[30] );
xor \add_6_14/U$7 ( \1177 , \1176 , \1169 );
buf \add_6_14/SUM[30] ( \1178_SUM[30] , \1177 );
buf \mul_6_18/A[30] ( \1179_A[30] , \1178_SUM[30] );
xor \add_6_14/U$14 ( \1180 , \993_A[29] , \994_B[29] );
xor \add_6_14/U$13 ( \1181 , \1180 , \1166 );
buf \add_6_14/SUM[29] ( \1182_SUM[29] , \1181 );
buf \mul_6_18/A[29] ( \1183_A[29] , \1182_SUM[29] );
xor \add_6_14/U$20 ( \1184 , \996_A[28] , \997_B[28] );
xor \add_6_14/U$19 ( \1185 , \1184 , \1163 );
buf \add_6_14/SUM[28] ( \1186_SUM[28] , \1185 );
buf \mul_6_18/A[28] ( \1187_A[28] , \1186_SUM[28] );
xor \add_6_14/U$26 ( \1188 , \999_A[27] , \1000_B[27] );
xor \add_6_14/U$25 ( \1189 , \1188 , \1160 );
buf \add_6_14/SUM[27] ( \1190_SUM[27] , \1189 );
buf \mul_6_18/A[27] ( \1191_A[27] , \1190_SUM[27] );
xor \add_6_14/U$32 ( \1192 , \1002_A[26] , \1003_B[26] );
xor \add_6_14/U$31 ( \1193 , \1192 , \1157 );
buf \add_6_14/SUM[26] ( \1194_SUM[26] , \1193 );
buf \mul_6_18/A[26] ( \1195_A[26] , \1194_SUM[26] );
xor \add_6_14/U$38 ( \1196 , \1005_A[25] , \1006_B[25] );
xor \add_6_14/U$37 ( \1197 , \1196 , \1154 );
buf \add_6_14/SUM[25] ( \1198_SUM[25] , \1197 );
buf \mul_6_18/A[25] ( \1199_A[25] , \1198_SUM[25] );
xor \add_6_14/U$44 ( \1200 , \1008_A[24] , \1009_B[24] );
xor \add_6_14/U$43 ( \1201 , \1200 , \1151 );
buf \add_6_14/SUM[24] ( \1202_SUM[24] , \1201 );
buf \mul_6_18/A[24] ( \1203_A[24] , \1202_SUM[24] );
xor \add_6_14/U$50 ( \1204 , \1011_A[23] , \1012_B[23] );
xor \add_6_14/U$49 ( \1205 , \1204 , \1148 );
buf \add_6_14/SUM[23] ( \1206_SUM[23] , \1205 );
buf \mul_6_18/A[23] ( \1207_A[23] , \1206_SUM[23] );
xor \add_6_14/U$56 ( \1208 , \1014_A[22] , \1015_B[22] );
xor \add_6_14/U$55 ( \1209 , \1208 , \1145 );
buf \add_6_14/SUM[22] ( \1210_SUM[22] , \1209 );
buf \mul_6_18/A[22] ( \1211_A[22] , \1210_SUM[22] );
xor \add_6_14/U$62 ( \1212 , \1017_A[21] , \1018_B[21] );
xor \add_6_14/U$61 ( \1213 , \1212 , \1142 );
buf \add_6_14/SUM[21] ( \1214_SUM[21] , \1213 );
buf \mul_6_18/A[21] ( \1215_A[21] , \1214_SUM[21] );
xor \add_6_14/U$68 ( \1216 , \1020_A[20] , \1021_B[20] );
xor \add_6_14/U$67 ( \1217 , \1216 , \1139 );
buf \add_6_14/SUM[20] ( \1218_SUM[20] , \1217 );
buf \mul_6_18/A[20] ( \1219_A[20] , \1218_SUM[20] );
xor \add_6_14/U$74 ( \1220 , \1023_A[19] , \1024_B[19] );
xor \add_6_14/U$73 ( \1221 , \1220 , \1136 );
buf \add_6_14/SUM[19] ( \1222_SUM[19] , \1221 );
buf \mul_6_18/A[19] ( \1223_A[19] , \1222_SUM[19] );
xor \add_6_14/U$80 ( \1224 , \1026_A[18] , \1027_B[18] );
xor \add_6_14/U$79 ( \1225 , \1224 , \1133 );
buf \add_6_14/SUM[18] ( \1226_SUM[18] , \1225 );
buf \mul_6_18/A[18] ( \1227_A[18] , \1226_SUM[18] );
xor \add_6_14/U$86 ( \1228 , \1029_A[17] , \1030_B[17] );
xor \add_6_14/U$85 ( \1229 , \1228 , \1130 );
buf \add_6_14/SUM[17] ( \1230_SUM[17] , \1229 );
buf \mul_6_18/A[17] ( \1231_A[17] , \1230_SUM[17] );
xor \add_6_14/U$92 ( \1232 , \1032_A[16] , \1033_B[16] );
xor \add_6_14/U$91 ( \1233 , \1232 , \1127 );
buf \add_6_14/SUM[16] ( \1234_SUM[16] , \1233 );
buf \mul_6_18/A[16] ( \1235_A[16] , \1234_SUM[16] );
xor \add_6_14/U$98 ( \1236 , \1035_A[15] , \1036_B[15] );
xor \add_6_14/U$97 ( \1237 , \1236 , \1124 );
buf \add_6_14/SUM[15] ( \1238_SUM[15] , \1237 );
buf \mul_6_18/A[15] ( \1239_A[15] , \1238_SUM[15] );
xor \add_6_14/U$104 ( \1240 , \1038_A[14] , \1039_B[14] );
xor \add_6_14/U$103 ( \1241 , \1240 , \1121 );
buf \add_6_14/SUM[14] ( \1242_SUM[14] , \1241 );
buf \mul_6_18/A[14] ( \1243_A[14] , \1242_SUM[14] );
xor \add_6_14/U$110 ( \1244 , \1041_A[13] , \1042_B[13] );
xor \add_6_14/U$109 ( \1245 , \1244 , \1118 );
buf \add_6_14/SUM[13] ( \1246_SUM[13] , \1245 );
buf \mul_6_18/A[13] ( \1247_A[13] , \1246_SUM[13] );
xor \add_6_14/U$116 ( \1248 , \1044_A[12] , \1045_B[12] );
xor \add_6_14/U$115 ( \1249 , \1248 , \1115 );
buf \add_6_14/SUM[12] ( \1250_SUM[12] , \1249 );
buf \mul_6_18/A[12] ( \1251_A[12] , \1250_SUM[12] );
xor \add_6_14/U$122 ( \1252 , \1047_A[11] , \1048_B[11] );
xor \add_6_14/U$121 ( \1253 , \1252 , \1112 );
buf \add_6_14/SUM[11] ( \1254_SUM[11] , \1253 );
buf \mul_6_18/A[11] ( \1255_A[11] , \1254_SUM[11] );
xor \add_6_14/U$128 ( \1256 , \1050_A[10] , \1051_B[10] );
xor \add_6_14/U$127 ( \1257 , \1256 , \1109 );
buf \add_6_14/SUM[10] ( \1258_SUM[10] , \1257 );
buf \mul_6_18/A[10] ( \1259_A[10] , \1258_SUM[10] );
xor \add_6_14/U$134 ( \1260 , \1053_A[9] , \1054_B[9] );
xor \add_6_14/U$133 ( \1261 , \1260 , \1106 );
buf \add_6_14/SUM[9] ( \1262_SUM[9] , \1261 );
buf \mul_6_18/A[9] ( \1263_A[9] , \1262_SUM[9] );
xor \add_6_14/U$140 ( \1264 , \1056_A[8] , \1057_B[8] );
xor \add_6_14/U$139 ( \1265 , \1264 , \1103 );
buf \add_6_14/SUM[8] ( \1266_SUM[8] , \1265 );
buf \mul_6_18/A[8] ( \1267_A[8] , \1266_SUM[8] );
xor \add_6_14/U$146 ( \1268 , \1059_A[7] , \1060_B[7] );
xor \add_6_14/U$145 ( \1269 , \1268 , \1100 );
buf \add_6_14/SUM[7] ( \1270_SUM[7] , \1269 );
buf \mul_6_18/A[7] ( \1271_A[7] , \1270_SUM[7] );
xor \add_6_14/U$152 ( \1272 , \1062_A[6] , \1063_B[6] );
xor \add_6_14/U$151 ( \1273 , \1272 , \1097 );
buf \add_6_14/SUM[6] ( \1274_SUM[6] , \1273 );
buf \mul_6_18/A[6] ( \1275_A[6] , \1274_SUM[6] );
xor \add_6_14/U$158 ( \1276 , \1065_A[5] , \1066_B[5] );
xor \add_6_14/U$157 ( \1277 , \1276 , \1094 );
buf \add_6_14/SUM[5] ( \1278_SUM[5] , \1277 );
buf \mul_6_18/A[5] ( \1279_A[5] , \1278_SUM[5] );
xor \add_6_14/U$164 ( \1280 , \1068_A[4] , \1069_B[4] );
xor \add_6_14/U$163 ( \1281 , \1280 , \1091 );
buf \add_6_14/SUM[4] ( \1282_SUM[4] , \1281 );
buf \mul_6_18/A[4] ( \1283_A[4] , \1282_SUM[4] );
xor \add_6_14/U$170 ( \1284 , \1071_A[3] , \1072_B[3] );
xor \add_6_14/U$169 ( \1285 , \1284 , \1088 );
buf \add_6_14/SUM[3] ( \1286_SUM[3] , \1285 );
buf \mul_6_18/A[3] ( \1287_A[3] , \1286_SUM[3] );
xor \add_6_14/U$176 ( \1288 , \1074_A[2] , \1075_B[2] );
xor \add_6_14/U$175 ( \1289 , \1288 , \1085 );
buf \add_6_14/SUM[2] ( \1290_SUM[2] , \1289 );
buf \mul_6_18/A[2] ( \1291_A[2] , \1290_SUM[2] );
xor \add_6_14/U$182 ( \1292 , \1077_A[1] , \1078_B[1] );
xor \add_6_14/U$181 ( \1293 , \1292 , \1082 );
buf \add_6_14/SUM[1] ( \1294_SUM[1] , \1293 );
buf \mul_6_18/A[1] ( \1295_A[1] , \1294_SUM[1] );
xor \add_6_14/U$184 ( \1296 , \1080_A[0] , \1081_B[0] );
buf \add_6_14/SUM[0] ( \1297_SUM[0] , \1296 );
buf \mul_6_18/A[0] ( \1298_A[0] , \1297_SUM[0] );
buf \mul_6_18/B[31] ( \1299_B[31] , \986 );
buf \mul_6_18/B[30] ( \1300_B[30] , \963 );
buf \mul_6_18/B[29] ( \1301_B[29] , \940 );
buf \mul_6_18/B[28] ( \1302_B[28] , \917 );
buf \mul_6_18/B[27] ( \1303_B[27] , \894 );
buf \mul_6_18/B[26] ( \1304_B[26] , \871 );
buf \mul_6_18/B[25] ( \1305_B[25] , \848 );
buf \mul_6_18/B[24] ( \1306_B[24] , \825 );
buf \mul_6_18/B[23] ( \1307_B[23] , \802 );
buf \mul_6_18/B[22] ( \1308_B[22] , \779 );
buf \mul_6_18/B[21] ( \1309_B[21] , \756 );
buf \mul_6_18/B[20] ( \1310_B[20] , \733 );
buf \mul_6_18/B[19] ( \1311_B[19] , \710 );
buf \mul_6_18/B[18] ( \1312_B[18] , \687 );
buf \mul_6_18/B[17] ( \1313_B[17] , \664 );
buf \mul_6_18/B[16] ( \1314_B[16] , \641 );
buf \mul_6_18/B[15] ( \1315_B[15] , \618 );
buf \mul_6_18/B[14] ( \1316_B[14] , \595 );
buf \mul_6_18/B[13] ( \1317_B[13] , \572 );
buf \mul_6_18/B[12] ( \1318_B[12] , \549 );
buf \mul_6_18/B[11] ( \1319_B[11] , \526 );
buf \mul_6_18/B[10] ( \1320_B[10] , \503 );
buf \mul_6_18/B[9] ( \1321_B[9] , \480 );
buf \mul_6_18/B[8] ( \1322_B[8] , \457 );
buf \mul_6_18/B[7] ( \1323_B[7] , \434 );
buf \mul_6_18/B[6] ( \1324_B[6] , \411 );
buf \mul_6_18/B[5] ( \1325_B[5] , \388 );
buf \mul_6_18/B[4] ( \1326_B[4] , \365 );
buf \mul_6_18/B[3] ( \1327_B[3] , \342 );
buf \mul_6_18/B[2] ( \1328_B[2] , \319 );
buf \mul_6_18/B[1] ( \1329_B[1] , \296 );
buf \mul_6_18/B[0] ( \1330_B[0] , \278 );
buf mul_6_18( \1331 , \1191_A[27] );
buf mul_6_18_g1( \1332 , \1329_B[1] );
buf mul_6_18_g2( \1333 , \1330_B[0] );
xor mul_6_18_g3( \1334 , \1332 , \1333 );
not mul_6_18_g4( \1335 , \1333 );
and mul_6_18_g5( \1336 , \1334 , \1335 );
and mul_6_18_g6( \1337 , \1331 , \1336 );
buf mul_6_18_g7( \1338 , \1187_A[28] );
and mul_6_18_g8( \1339 , \1338 , \1333 );
nor mul_6_18_g9( \1340 , \1337 , \1339 );
xnor mul_6_18_g10( \1341 , \1340 , \1332 );
buf mul_6_18_g11( \1342 , \1215_A[21] );
buf mul_6_18_g12( \1343 , \1323_B[7] );
buf mul_6_18_g13( \1344 , \1324_B[6] );
xor mul_6_18_g14( \1345 , \1343 , \1344 );
buf mul_6_18_g15( \1346 , \1325_B[5] );
xor mul_6_18_g16( \1347 , \1344 , \1346 );
not mul_6_18_g17( \1348 , \1347 );
and mul_6_18_g18( \1349 , \1345 , \1348 );
and mul_6_18_g19( \1350 , \1342 , \1349 );
buf mul_6_18_g20( \1351 , \1211_A[22] );
and mul_6_18_g21( \1352 , \1351 , \1347 );
nor mul_6_18_g22( \1353 , \1350 , \1352 );
and mul_6_18_g23( \1354 , \1344 , \1346 );
not mul_6_18_g24( \1355 , \1354 );
and mul_6_18_g25( \1356 , \1343 , \1355 );
xnor mul_6_18_g26( \1357 , \1353 , \1356 );
xor mul_6_18_g27( \1358 , \1341 , \1357 );
buf mul_6_18_g28( \1359 , \1247_A[13] );
buf mul_6_18_g29( \1360 , \1315_B[15] );
buf mul_6_18_g30( \1361 , \1316_B[14] );
xor mul_6_18_g31( \1362 , \1360 , \1361 );
buf mul_6_18_g32( \1363 , \1317_B[13] );
xor mul_6_18_g33( \1364 , \1361 , \1363 );
not mul_6_18_g34( \1365 , \1364 );
and mul_6_18_g35( \1366 , \1362 , \1365 );
and mul_6_18_g36( \1367 , \1359 , \1366 );
buf mul_6_18_g37( \1368 , \1243_A[14] );
and mul_6_18_g38( \1369 , \1368 , \1364 );
nor mul_6_18_g39( \1370 , \1367 , \1369 );
and mul_6_18_g40( \1371 , \1361 , \1363 );
not mul_6_18_g41( \1372 , \1371 );
and mul_6_18_g42( \1373 , \1360 , \1372 );
xnor mul_6_18_g43( \1374 , \1370 , \1373 );
xor mul_6_18_g44( \1375 , \1358 , \1374 );
buf mul_6_18_g45( \1376 , \1223_A[19] );
buf mul_6_18_g46( \1377 , \1321_B[9] );
buf mul_6_18_g47( \1378 , \1322_B[8] );
xor mul_6_18_g48( \1379 , \1377 , \1378 );
xor mul_6_18_g49( \1380 , \1378 , \1343 );
not mul_6_18_g50( \1381 , \1380 );
and mul_6_18_g51( \1382 , \1379 , \1381 );
and mul_6_18_g52( \1383 , \1376 , \1382 );
buf mul_6_18_g53( \1384 , \1219_A[20] );
and mul_6_18_g54( \1385 , \1384 , \1380 );
nor mul_6_18_g55( \1386 , \1383 , \1385 );
and mul_6_18_g56( \1387 , \1378 , \1343 );
not mul_6_18_g57( \1388 , \1387 );
and mul_6_18_g58( \1389 , \1377 , \1388 );
xnor mul_6_18_g59( \1390 , \1386 , \1389 );
buf mul_6_18_g60( \1391 , \1255_A[11] );
buf mul_6_18_g61( \1392 , \1313_B[17] );
buf mul_6_18_g62( \1393 , \1314_B[16] );
xor mul_6_18_g63( \1394 , \1392 , \1393 );
xor mul_6_18_g64( \1395 , \1393 , \1360 );
not mul_6_18_g65( \1396 , \1395 );
and mul_6_18_g66( \1397 , \1394 , \1396 );
and mul_6_18_g67( \1398 , \1391 , \1397 );
buf mul_6_18_g68( \1399 , \1251_A[12] );
and mul_6_18_g69( \1400 , \1399 , \1395 );
nor mul_6_18_g70( \1401 , \1398 , \1400 );
and mul_6_18_g71( \1402 , \1393 , \1360 );
not mul_6_18_g72( \1403 , \1402 );
and mul_6_18_g73( \1404 , \1392 , \1403 );
xnor mul_6_18_g74( \1405 , \1401 , \1404 );
xor mul_6_18_g75( \1406 , \1390 , \1405 );
buf mul_6_18_g76( \1407 , \1271_A[7] );
buf mul_6_18_g77( \1408 , \1309_B[21] );
buf mul_6_18_g78( \1409 , \1310_B[20] );
xor mul_6_18_g79( \1410 , \1408 , \1409 );
buf mul_6_18_g80( \1411 , \1311_B[19] );
xor mul_6_18_g81( \1412 , \1409 , \1411 );
not mul_6_18_g82( \1413 , \1412 );
and mul_6_18_g83( \1414 , \1410 , \1413 );
and mul_6_18_g84( \1415 , \1407 , \1414 );
buf mul_6_18_g85( \1416 , \1267_A[8] );
and mul_6_18_g86( \1417 , \1416 , \1412 );
nor mul_6_18_g87( \1418 , \1415 , \1417 );
and mul_6_18_g88( \1419 , \1409 , \1411 );
not mul_6_18_g89( \1420 , \1419 );
and mul_6_18_g90( \1421 , \1408 , \1420 );
xnor mul_6_18_g91( \1422 , \1418 , \1421 );
xor mul_6_18_g92( \1423 , \1406 , \1422 );
and mul_6_18_g93( \1424 , \1375 , \1423 );
buf mul_6_18_g94( \1425 , \1203_A[24] );
buf mul_6_18_g95( \1426 , \1327_B[3] );
buf mul_6_18_g96( \1427 , \1328_B[2] );
xor mul_6_18_g97( \1428 , \1426 , \1427 );
xor mul_6_18_g98( \1429 , \1427 , \1332 );
not mul_6_18_g99( \1430 , \1429 );
and mul_6_18_g100( \1431 , \1428 , \1430 );
and mul_6_18_g101( \1432 , \1425 , \1431 );
buf mul_6_18_g102( \1433 , \1199_A[25] );
and mul_6_18_g103( \1434 , \1433 , \1429 );
nor mul_6_18_g104( \1435 , \1432 , \1434 );
and mul_6_18_g105( \1436 , \1427 , \1332 );
not mul_6_18_g106( \1437 , \1436 );
and mul_6_18_g107( \1438 , \1426 , \1437 );
xnor mul_6_18_g108( \1439 , \1435 , \1438 );
buf mul_6_18_g109( \1440 , \1326_B[4] );
xor mul_6_18_g110( \1441 , \1346 , \1440 );
xor mul_6_18_g111( \1442 , \1440 , \1426 );
not mul_6_18_g112( \1443 , \1442 );
and mul_6_18_g113( \1444 , \1441 , \1443 );
and mul_6_18_g114( \1445 , \1351 , \1444 );
buf mul_6_18_g115( \1446 , \1207_A[23] );
and mul_6_18_g116( \1447 , \1446 , \1442 );
nor mul_6_18_g117( \1448 , \1445 , \1447 );
and mul_6_18_g118( \1449 , \1440 , \1426 );
not mul_6_18_g119( \1450 , \1449 );
and mul_6_18_g120( \1451 , \1346 , \1450 );
xnor mul_6_18_g121( \1452 , \1448 , \1451 );
and mul_6_18_g122( \1453 , \1439 , \1452 );
buf mul_6_18_g123( \1454 , \1231_A[17] );
buf mul_6_18_g124( \1455 , \1319_B[11] );
buf mul_6_18_g125( \1456 , \1320_B[10] );
xor mul_6_18_g126( \1457 , \1455 , \1456 );
xor mul_6_18_g127( \1458 , \1456 , \1377 );
not mul_6_18_g128( \1459 , \1458 );
and mul_6_18_g129( \1460 , \1457 , \1459 );
and mul_6_18_g130( \1461 , \1454 , \1460 );
buf mul_6_18_g131( \1462 , \1227_A[18] );
and mul_6_18_g132( \1463 , \1462 , \1458 );
nor mul_6_18_g133( \1464 , \1461 , \1463 );
and mul_6_18_g134( \1465 , \1456 , \1377 );
not mul_6_18_g135( \1466 , \1465 );
and mul_6_18_g136( \1467 , \1455 , \1466 );
xnor mul_6_18_g137( \1468 , \1464 , \1467 );
xor mul_6_18_g138( \1469 , \1453 , \1468 );
buf mul_6_18_g139( \1470 , \1239_A[15] );
buf mul_6_18_g140( \1471 , \1318_B[12] );
xor mul_6_18_g141( \1472 , \1363 , \1471 );
xor mul_6_18_g142( \1473 , \1471 , \1455 );
not mul_6_18_g143( \1474 , \1473 );
and mul_6_18_g144( \1475 , \1472 , \1474 );
and mul_6_18_g145( \1476 , \1470 , \1475 );
buf mul_6_18_g146( \1477 , \1235_A[16] );
and mul_6_18_g147( \1478 , \1477 , \1473 );
nor mul_6_18_g148( \1479 , \1476 , \1478 );
and mul_6_18_g149( \1480 , \1471 , \1455 );
not mul_6_18_g150( \1481 , \1480 );
and mul_6_18_g151( \1482 , \1363 , \1481 );
xnor mul_6_18_g152( \1483 , \1479 , \1482 );
xor mul_6_18_g153( \1484 , \1469 , \1483 );
and mul_6_18_g154( \1485 , \1423 , \1484 );
and mul_6_18_g155( \1486 , \1375 , \1484 );
or mul_6_18_g156( \1487 , \1424 , \1485 , \1486 );
and mul_6_18_g157( \1488 , \1433 , \1431 );
buf mul_6_18_g158( \1489 , \1195_A[26] );
and mul_6_18_g159( \1490 , \1489 , \1429 );
nor mul_6_18_g160( \1491 , \1488 , \1490 );
xnor mul_6_18_g161( \1492 , \1491 , \1438 );
and mul_6_18_g162( \1493 , \1446 , \1444 );
and mul_6_18_g163( \1494 , \1425 , \1442 );
nor mul_6_18_g164( \1495 , \1493 , \1494 );
xnor mul_6_18_g165( \1496 , \1495 , \1451 );
and mul_6_18_g166( \1497 , \1492 , \1496 );
buf mul_6_18_g167( \1498 , \1298_A[0] );
buf mul_6_18_g168( \1499 , \1302_B[28] );
buf mul_6_18_g169( \1500 , \1303_B[27] );
xor mul_6_18_g170( \1501 , \1499 , \1500 );
and mul_6_18_g171( \1502 , \1498 , \1501 );
and mul_6_18_g172( \1503 , \1496 , \1502 );
and mul_6_18_g173( \1504 , \1492 , \1502 );
or mul_6_18_g174( \1505 , \1497 , \1503 , \1504 );
and mul_6_18_g175( \1506 , \1341 , \1357 );
and mul_6_18_g176( \1507 , \1357 , \1374 );
and mul_6_18_g177( \1508 , \1341 , \1374 );
or mul_6_18_g178( \1509 , \1506 , \1507 , \1508 );
xor mul_6_18_g179( \1510 , \1505 , \1509 );
and mul_6_18_g180( \1511 , \1390 , \1405 );
and mul_6_18_g181( \1512 , \1405 , \1422 );
and mul_6_18_g182( \1513 , \1390 , \1422 );
or mul_6_18_g183( \1514 , \1511 , \1512 , \1513 );
xor mul_6_18_g184( \1515 , \1510 , \1514 );
and mul_6_18_g185( \1516 , \1487 , \1515 );
buf mul_6_18_g186( \1517 , \1283_A[4] );
buf mul_6_18_g187( \1518 , \1305_B[25] );
buf mul_6_18_g188( \1519 , \1306_B[24] );
xor mul_6_18_g189( \1520 , \1518 , \1519 );
buf mul_6_18_g190( \1521 , \1307_B[23] );
xor mul_6_18_g191( \1522 , \1519 , \1521 );
not mul_6_18_g192( \1523 , \1522 );
and mul_6_18_g193( \1524 , \1520 , \1523 );
and mul_6_18_g194( \1525 , \1517 , \1524 );
buf mul_6_18_g195( \1526 , \1279_A[5] );
and mul_6_18_g196( \1527 , \1526 , \1522 );
nor mul_6_18_g197( \1528 , \1525 , \1527 );
and mul_6_18_g198( \1529 , \1519 , \1521 );
not mul_6_18_g199( \1530 , \1529 );
and mul_6_18_g200( \1531 , \1518 , \1530 );
xnor mul_6_18_g201( \1532 , \1528 , \1531 );
buf mul_6_18_g202( \1533 , \1291_A[2] );
buf mul_6_18_g203( \1534 , \1304_B[26] );
xor mul_6_18_g204( \1535 , \1500 , \1534 );
xor mul_6_18_g205( \1536 , \1534 , \1518 );
not mul_6_18_g206( \1537 , \1536 );
and mul_6_18_g207( \1538 , \1535 , \1537 );
and mul_6_18_g208( \1539 , \1533 , \1538 );
buf mul_6_18_g209( \1540 , \1287_A[3] );
and mul_6_18_g210( \1541 , \1540 , \1536 );
nor mul_6_18_g211( \1542 , \1539 , \1541 );
and mul_6_18_g212( \1543 , \1534 , \1518 );
not mul_6_18_g213( \1544 , \1543 );
and mul_6_18_g214( \1545 , \1500 , \1544 );
xnor mul_6_18_g215( \1546 , \1542 , \1545 );
xor mul_6_18_g216( \1547 , \1532 , \1546 );
buf mul_6_18_g217( \1548 , \1301_B[29] );
xor mul_6_18_g218( \1549 , \1548 , \1499 );
not mul_6_18_g219( \1550 , \1501 );
and mul_6_18_g220( \1551 , \1549 , \1550 );
and mul_6_18_g221( \1552 , \1498 , \1551 );
buf mul_6_18_g222( \1553 , \1295_A[1] );
and mul_6_18_g223( \1554 , \1553 , \1501 );
nor mul_6_18_g224( \1555 , \1552 , \1554 );
and mul_6_18_g225( \1556 , \1499 , \1500 );
not mul_6_18_g226( \1557 , \1556 );
and mul_6_18_g227( \1558 , \1548 , \1557 );
xnor mul_6_18_g228( \1559 , \1555 , \1558 );
xor mul_6_18_g229( \1560 , \1547 , \1559 );
and mul_6_18_g230( \1561 , \1384 , \1382 );
and mul_6_18_g231( \1562 , \1342 , \1380 );
nor mul_6_18_g232( \1563 , \1561 , \1562 );
xnor mul_6_18_g233( \1564 , \1563 , \1389 );
and mul_6_18_g234( \1565 , \1368 , \1366 );
and mul_6_18_g235( \1566 , \1470 , \1364 );
nor mul_6_18_g236( \1567 , \1565 , \1566 );
xnor mul_6_18_g237( \1568 , \1567 , \1373 );
xor mul_6_18_g238( \1569 , \1564 , \1568 );
and mul_6_18_g239( \1570 , \1399 , \1397 );
and mul_6_18_g240( \1571 , \1359 , \1395 );
nor mul_6_18_g241( \1572 , \1570 , \1571 );
xnor mul_6_18_g242( \1573 , \1572 , \1404 );
xor mul_6_18_g243( \1574 , \1569 , \1573 );
xor mul_6_18_g244( \1575 , \1560 , \1574 );
and mul_6_18_g245( \1576 , \1462 , \1460 );
and mul_6_18_g246( \1577 , \1376 , \1458 );
nor mul_6_18_g247( \1578 , \1576 , \1577 );
xnor mul_6_18_g248( \1579 , \1578 , \1467 );
and mul_6_18_g249( \1580 , \1477 , \1475 );
and mul_6_18_g250( \1581 , \1454 , \1473 );
nor mul_6_18_g251( \1582 , \1580 , \1581 );
xnor mul_6_18_g252( \1583 , \1582 , \1482 );
xor mul_6_18_g253( \1584 , \1579 , \1583 );
and mul_6_18_g254( \1585 , \1416 , \1414 );
buf mul_6_18_g255( \1586 , \1263_A[9] );
and mul_6_18_g256( \1587 , \1586 , \1412 );
nor mul_6_18_g257( \1588 , \1585 , \1587 );
xnor mul_6_18_g258( \1589 , \1588 , \1421 );
xor mul_6_18_g259( \1590 , \1584 , \1589 );
xor mul_6_18_g260( \1591 , \1575 , \1590 );
and mul_6_18_g261( \1592 , \1515 , \1591 );
and mul_6_18_g262( \1593 , \1487 , \1591 );
or mul_6_18_g263( \1594 , \1516 , \1592 , \1593 );
and mul_6_18_g264( \1595 , \1433 , \1336 );
and mul_6_18_g265( \1596 , \1489 , \1333 );
nor mul_6_18_g266( \1597 , \1595 , \1596 );
xnor mul_6_18_g267( \1598 , \1597 , \1332 );
and mul_6_18_g268( \1599 , \1376 , \1349 );
and mul_6_18_g269( \1600 , \1384 , \1347 );
nor mul_6_18_g270( \1601 , \1599 , \1600 );
xnor mul_6_18_g271( \1602 , \1601 , \1356 );
and mul_6_18_g272( \1603 , \1598 , \1602 );
and mul_6_18_g273( \1604 , \1391 , \1366 );
and mul_6_18_g274( \1605 , \1399 , \1364 );
nor mul_6_18_g275( \1606 , \1604 , \1605 );
xnor mul_6_18_g276( \1607 , \1606 , \1373 );
and mul_6_18_g277( \1608 , \1602 , \1607 );
and mul_6_18_g278( \1609 , \1598 , \1607 );
or mul_6_18_g279( \1610 , \1603 , \1608 , \1609 );
and mul_6_18_g280( \1611 , \1454 , \1382 );
and mul_6_18_g281( \1612 , \1462 , \1380 );
nor mul_6_18_g282( \1613 , \1611 , \1612 );
xnor mul_6_18_g283( \1614 , \1613 , \1389 );
and mul_6_18_g284( \1615 , \1586 , \1397 );
buf mul_6_18_g285( \1616 , \1259_A[10] );
and mul_6_18_g286( \1617 , \1616 , \1395 );
nor mul_6_18_g287( \1618 , \1615 , \1617 );
xnor mul_6_18_g288( \1619 , \1618 , \1404 );
and mul_6_18_g289( \1620 , \1614 , \1619 );
and mul_6_18_g290( \1621 , \1526 , \1414 );
buf mul_6_18_g291( \1622 , \1275_A[6] );
and mul_6_18_g292( \1623 , \1622 , \1412 );
nor mul_6_18_g293( \1624 , \1621 , \1623 );
xnor mul_6_18_g294( \1625 , \1624 , \1421 );
and mul_6_18_g295( \1626 , \1619 , \1625 );
and mul_6_18_g296( \1627 , \1614 , \1625 );
or mul_6_18_g297( \1628 , \1620 , \1626 , \1627 );
and mul_6_18_g298( \1629 , \1610 , \1628 );
and mul_6_18_g299( \1630 , \1351 , \1431 );
and mul_6_18_g300( \1631 , \1446 , \1429 );
nor mul_6_18_g301( \1632 , \1630 , \1631 );
xnor mul_6_18_g302( \1633 , \1632 , \1438 );
and mul_6_18_g303( \1634 , \1384 , \1444 );
and mul_6_18_g304( \1635 , \1342 , \1442 );
nor mul_6_18_g305( \1636 , \1634 , \1635 );
xnor mul_6_18_g306( \1637 , \1636 , \1451 );
and mul_6_18_g307( \1638 , \1633 , \1637 );
buf mul_6_18_g308( \1639 , \1308_B[22] );
xor mul_6_18_g309( \1640 , \1521 , \1639 );
xor mul_6_18_g310( \1641 , \1639 , \1408 );
not mul_6_18_g311( \1642 , \1641 );
and mul_6_18_g312( \1643 , \1640 , \1642 );
and mul_6_18_g313( \1644 , \1540 , \1643 );
and mul_6_18_g314( \1645 , \1517 , \1641 );
nor mul_6_18_g315( \1646 , \1644 , \1645 );
and mul_6_18_g316( \1647 , \1639 , \1408 );
not mul_6_18_g317( \1648 , \1647 );
and mul_6_18_g318( \1649 , \1521 , \1648 );
xnor mul_6_18_g319( \1650 , \1646 , \1649 );
and mul_6_18_g320( \1651 , \1638 , \1650 );
and mul_6_18_g321( \1652 , \1553 , \1524 );
and mul_6_18_g322( \1653 , \1533 , \1522 );
nor mul_6_18_g323( \1654 , \1652 , \1653 );
xnor mul_6_18_g324( \1655 , \1654 , \1531 );
and mul_6_18_g325( \1656 , \1650 , \1655 );
and mul_6_18_g326( \1657 , \1638 , \1655 );
or mul_6_18_g327( \1658 , \1651 , \1656 , \1657 );
and mul_6_18_g328( \1659 , \1628 , \1658 );
and mul_6_18_g329( \1660 , \1610 , \1658 );
or mul_6_18_g330( \1661 , \1629 , \1659 , \1660 );
and mul_6_18_g331( \1662 , \1470 , \1460 );
and mul_6_18_g332( \1663 , \1477 , \1458 );
nor mul_6_18_g333( \1664 , \1662 , \1663 );
xnor mul_6_18_g334( \1665 , \1664 , \1467 );
and mul_6_18_g335( \1666 , \1359 , \1475 );
and mul_6_18_g336( \1667 , \1368 , \1473 );
nor mul_6_18_g337( \1668 , \1666 , \1667 );
xnor mul_6_18_g338( \1669 , \1668 , \1482 );
and mul_6_18_g339( \1670 , \1665 , \1669 );
buf mul_6_18_g340( \1671 , \1312_B[18] );
xor mul_6_18_g341( \1672 , \1411 , \1671 );
xor mul_6_18_g342( \1673 , \1671 , \1392 );
not mul_6_18_g343( \1674 , \1673 );
and mul_6_18_g344( \1675 , \1672 , \1674 );
and mul_6_18_g345( \1676 , \1407 , \1675 );
and mul_6_18_g346( \1677 , \1416 , \1673 );
nor mul_6_18_g347( \1678 , \1676 , \1677 );
and mul_6_18_g348( \1679 , \1671 , \1392 );
not mul_6_18_g349( \1680 , \1679 );
and mul_6_18_g350( \1681 , \1411 , \1680 );
xnor mul_6_18_g351( \1682 , \1678 , \1681 );
and mul_6_18_g352( \1683 , \1669 , \1682 );
and mul_6_18_g353( \1684 , \1665 , \1682 );
or mul_6_18_g354( \1685 , \1670 , \1683 , \1684 );
and mul_6_18_g355( \1686 , \1462 , \1382 );
and mul_6_18_g356( \1687 , \1376 , \1380 );
nor mul_6_18_g357( \1688 , \1686 , \1687 );
xnor mul_6_18_g358( \1689 , \1688 , \1389 );
and mul_6_18_g359( \1690 , \1399 , \1366 );
and mul_6_18_g360( \1691 , \1359 , \1364 );
nor mul_6_18_g361( \1692 , \1690 , \1691 );
xnor mul_6_18_g362( \1693 , \1692 , \1373 );
xor mul_6_18_g363( \1694 , \1689 , \1693 );
and mul_6_18_g364( \1695 , \1616 , \1397 );
and mul_6_18_g365( \1696 , \1391 , \1395 );
nor mul_6_18_g366( \1697 , \1695 , \1696 );
xnor mul_6_18_g367( \1698 , \1697 , \1404 );
xor mul_6_18_g368( \1699 , \1694 , \1698 );
and mul_6_18_g369( \1700 , \1685 , \1699 );
and mul_6_18_g370( \1701 , \1477 , \1460 );
and mul_6_18_g371( \1702 , \1454 , \1458 );
nor mul_6_18_g372( \1703 , \1701 , \1702 );
xnor mul_6_18_g373( \1704 , \1703 , \1467 );
and mul_6_18_g374( \1705 , \1368 , \1475 );
and mul_6_18_g375( \1706 , \1470 , \1473 );
nor mul_6_18_g376( \1707 , \1705 , \1706 );
xnor mul_6_18_g377( \1708 , \1707 , \1482 );
xor mul_6_18_g378( \1709 , \1704 , \1708 );
and mul_6_18_g379( \1710 , \1622 , \1414 );
and mul_6_18_g380( \1711 , \1407 , \1412 );
nor mul_6_18_g381( \1712 , \1710 , \1711 );
xnor mul_6_18_g382( \1713 , \1712 , \1421 );
xor mul_6_18_g383( \1714 , \1709 , \1713 );
and mul_6_18_g384( \1715 , \1699 , \1714 );
and mul_6_18_g385( \1716 , \1685 , \1714 );
or mul_6_18_g386( \1717 , \1700 , \1715 , \1716 );
and mul_6_18_g387( \1718 , \1661 , \1717 );
and mul_6_18_g388( \1719 , \1689 , \1693 );
and mul_6_18_g389( \1720 , \1693 , \1698 );
and mul_6_18_g390( \1721 , \1689 , \1698 );
or mul_6_18_g391( \1722 , \1719 , \1720 , \1721 );
and mul_6_18_g392( \1723 , \1704 , \1708 );
and mul_6_18_g393( \1724 , \1708 , \1713 );
and mul_6_18_g394( \1725 , \1704 , \1713 );
or mul_6_18_g395( \1726 , \1723 , \1724 , \1725 );
xor mul_6_18_g396( \1727 , \1722 , \1726 );
xor mul_6_18_g397( \1728 , \1439 , \1452 );
and mul_6_18_g398( \1729 , \1416 , \1675 );
and mul_6_18_g399( \1730 , \1586 , \1673 );
nor mul_6_18_g400( \1731 , \1729 , \1730 );
xnor mul_6_18_g401( \1732 , \1731 , \1681 );
and mul_6_18_g402( \1733 , \1728 , \1732 );
and mul_6_18_g403( \1734 , \1517 , \1643 );
and mul_6_18_g404( \1735 , \1526 , \1641 );
nor mul_6_18_g405( \1736 , \1734 , \1735 );
xnor mul_6_18_g406( \1737 , \1736 , \1649 );
and mul_6_18_g407( \1738 , \1732 , \1737 );
and mul_6_18_g408( \1739 , \1728 , \1737 );
or mul_6_18_g409( \1740 , \1733 , \1738 , \1739 );
xor mul_6_18_g410( \1741 , \1727 , \1740 );
and mul_6_18_g411( \1742 , \1717 , \1741 );
and mul_6_18_g412( \1743 , \1661 , \1741 );
or mul_6_18_g413( \1744 , \1718 , \1742 , \1743 );
and mul_6_18_g414( \1745 , \1446 , \1431 );
and mul_6_18_g415( \1746 , \1425 , \1429 );
nor mul_6_18_g416( \1747 , \1745 , \1746 );
xnor mul_6_18_g417( \1748 , \1747 , \1438 );
and mul_6_18_g418( \1749 , \1342 , \1444 );
and mul_6_18_g419( \1750 , \1351 , \1442 );
nor mul_6_18_g420( \1751 , \1749 , \1750 );
xnor mul_6_18_g421( \1752 , \1751 , \1451 );
and mul_6_18_g422( \1753 , \1748 , \1752 );
and mul_6_18_g423( \1754 , \1498 , \1536 );
and mul_6_18_g424( \1755 , \1752 , \1754 );
and mul_6_18_g425( \1756 , \1748 , \1754 );
or mul_6_18_g426( \1757 , \1753 , \1755 , \1756 );
and mul_6_18_g427( \1758 , \1533 , \1524 );
and mul_6_18_g428( \1759 , \1540 , \1522 );
nor mul_6_18_g429( \1760 , \1758 , \1759 );
xnor mul_6_18_g430( \1761 , \1760 , \1531 );
and mul_6_18_g431( \1762 , \1757 , \1761 );
and mul_6_18_g432( \1763 , \1498 , \1538 );
and mul_6_18_g433( \1764 , \1553 , \1536 );
nor mul_6_18_g434( \1765 , \1763 , \1764 );
xnor mul_6_18_g435( \1766 , \1765 , \1545 );
and mul_6_18_g436( \1767 , \1761 , \1766 );
and mul_6_18_g437( \1768 , \1757 , \1766 );
or mul_6_18_g438( \1769 , \1762 , \1767 , \1768 );
and mul_6_18_g439( \1770 , \1586 , \1675 );
and mul_6_18_g440( \1771 , \1616 , \1673 );
nor mul_6_18_g441( \1772 , \1770 , \1771 );
xnor mul_6_18_g442( \1773 , \1772 , \1681 );
and mul_6_18_g443( \1774 , \1526 , \1643 );
and mul_6_18_g444( \1775 , \1622 , \1641 );
nor mul_6_18_g445( \1776 , \1774 , \1775 );
xnor mul_6_18_g446( \1777 , \1776 , \1649 );
xor mul_6_18_g447( \1778 , \1773 , \1777 );
and mul_6_18_g448( \1779 , \1540 , \1524 );
and mul_6_18_g449( \1780 , \1517 , \1522 );
nor mul_6_18_g450( \1781 , \1779 , \1780 );
xnor mul_6_18_g451( \1782 , \1781 , \1531 );
xor mul_6_18_g452( \1783 , \1778 , \1782 );
and mul_6_18_g453( \1784 , \1769 , \1783 );
and mul_6_18_g454( \1785 , \1489 , \1336 );
and mul_6_18_g455( \1786 , \1331 , \1333 );
nor mul_6_18_g456( \1787 , \1785 , \1786 );
xnor mul_6_18_g457( \1788 , \1787 , \1332 );
and mul_6_18_g458( \1789 , \1384 , \1349 );
and mul_6_18_g459( \1790 , \1342 , \1347 );
nor mul_6_18_g460( \1791 , \1789 , \1790 );
xnor mul_6_18_g461( \1792 , \1791 , \1356 );
and mul_6_18_g462( \1793 , \1788 , \1792 );
not mul_6_18_g463( \1794 , \1754 );
and mul_6_18_g464( \1795 , \1794 , \1545 );
and mul_6_18_g465( \1796 , \1792 , \1795 );
and mul_6_18_g466( \1797 , \1788 , \1795 );
or mul_6_18_g467( \1798 , \1793 , \1796 , \1797 );
and mul_6_18_g468( \1799 , \1553 , \1538 );
and mul_6_18_g469( \1800 , \1533 , \1536 );
nor mul_6_18_g470( \1801 , \1799 , \1800 );
xnor mul_6_18_g471( \1802 , \1801 , \1545 );
xor mul_6_18_g472( \1803 , \1798 , \1802 );
xor mul_6_18_g473( \1804 , \1492 , \1496 );
xor mul_6_18_g474( \1805 , \1804 , \1502 );
xor mul_6_18_g475( \1806 , \1803 , \1805 );
and mul_6_18_g476( \1807 , \1783 , \1806 );
and mul_6_18_g477( \1808 , \1769 , \1806 );
or mul_6_18_g478( \1809 , \1784 , \1807 , \1808 );
and mul_6_18_g479( \1810 , \1744 , \1809 );
and mul_6_18_g480( \1811 , \1773 , \1777 );
and mul_6_18_g481( \1812 , \1777 , \1782 );
and mul_6_18_g482( \1813 , \1773 , \1782 );
or mul_6_18_g483( \1814 , \1811 , \1812 , \1813 );
and mul_6_18_g484( \1815 , \1453 , \1468 );
and mul_6_18_g485( \1816 , \1468 , \1483 );
and mul_6_18_g486( \1817 , \1453 , \1483 );
or mul_6_18_g487( \1818 , \1815 , \1816 , \1817 );
xor mul_6_18_g488( \1819 , \1814 , \1818 );
and mul_6_18_g489( \1820 , \1338 , \1336 );
buf mul_6_18_g490( \1821 , \1183_A[29] );
and mul_6_18_g491( \1822 , \1821 , \1333 );
nor mul_6_18_g492( \1823 , \1820 , \1822 );
xnor mul_6_18_g493( \1824 , \1823 , \1332 );
and mul_6_18_g494( \1825 , \1425 , \1444 );
and mul_6_18_g495( \1826 , \1433 , \1442 );
nor mul_6_18_g496( \1827 , \1825 , \1826 );
xnor mul_6_18_g497( \1828 , \1827 , \1451 );
xor mul_6_18_g498( \1829 , \1824 , \1828 );
and mul_6_18_g499( \1830 , \1351 , \1349 );
and mul_6_18_g500( \1831 , \1446 , \1347 );
nor mul_6_18_g501( \1832 , \1830 , \1831 );
xnor mul_6_18_g502( \1833 , \1832 , \1356 );
xor mul_6_18_g503( \1834 , \1829 , \1833 );
xor mul_6_18_g504( \1835 , \1819 , \1834 );
and mul_6_18_g505( \1836 , \1809 , \1835 );
and mul_6_18_g506( \1837 , \1744 , \1835 );
or mul_6_18_g507( \1838 , \1810 , \1836 , \1837 );
and mul_6_18_g508( \1839 , \1594 , \1838 );
and mul_6_18_g509( \1840 , \1560 , \1574 );
and mul_6_18_g510( \1841 , \1574 , \1590 );
and mul_6_18_g511( \1842 , \1560 , \1590 );
or mul_6_18_g512( \1843 , \1840 , \1841 , \1842 );
and mul_6_18_g513( \1844 , \1814 , \1818 );
and mul_6_18_g514( \1845 , \1818 , \1834 );
and mul_6_18_g515( \1846 , \1814 , \1834 );
or mul_6_18_g516( \1847 , \1844 , \1845 , \1846 );
xor mul_6_18_g517( \1848 , \1843 , \1847 );
and mul_6_18_g518( \1849 , \1489 , \1431 );
and mul_6_18_g519( \1850 , \1331 , \1429 );
nor mul_6_18_g520( \1851 , \1849 , \1850 );
xnor mul_6_18_g521( \1852 , \1851 , \1438 );
not mul_6_18_g522( \1853 , \1502 );
and mul_6_18_g523( \1854 , \1853 , \1558 );
xor mul_6_18_g524( \1855 , \1852 , \1854 );
and mul_6_18_g525( \1856 , \1616 , \1675 );
and mul_6_18_g526( \1857 , \1391 , \1673 );
nor mul_6_18_g527( \1858 , \1856 , \1857 );
xnor mul_6_18_g528( \1859 , \1858 , \1681 );
and mul_6_18_g529( \1860 , \1855 , \1859 );
and mul_6_18_g530( \1861 , \1622 , \1643 );
and mul_6_18_g531( \1862 , \1407 , \1641 );
nor mul_6_18_g532( \1863 , \1861 , \1862 );
xnor mul_6_18_g533( \1864 , \1863 , \1649 );
and mul_6_18_g534( \1865 , \1859 , \1864 );
and mul_6_18_g535( \1866 , \1855 , \1864 );
or mul_6_18_g536( \1867 , \1860 , \1865 , \1866 );
and mul_6_18_g537( \1868 , \1342 , \1382 );
and mul_6_18_g538( \1869 , \1351 , \1380 );
nor mul_6_18_g539( \1870 , \1868 , \1869 );
xnor mul_6_18_g540( \1871 , \1870 , \1389 );
and mul_6_18_g541( \1872 , \1359 , \1397 );
and mul_6_18_g542( \1873 , \1368 , \1395 );
nor mul_6_18_g543( \1874 , \1872 , \1873 );
xnor mul_6_18_g544( \1875 , \1874 , \1404 );
xor mul_6_18_g545( \1876 , \1871 , \1875 );
and mul_6_18_g546( \1877 , \1586 , \1414 );
and mul_6_18_g547( \1878 , \1616 , \1412 );
nor mul_6_18_g548( \1879 , \1877 , \1878 );
xnor mul_6_18_g549( \1880 , \1879 , \1421 );
xor mul_6_18_g550( \1881 , \1876 , \1880 );
xor mul_6_18_g551( \1882 , \1867 , \1881 );
and mul_6_18_g552( \1883 , \1391 , \1675 );
and mul_6_18_g553( \1884 , \1399 , \1673 );
nor mul_6_18_g554( \1885 , \1883 , \1884 );
xnor mul_6_18_g555( \1886 , \1885 , \1681 );
and mul_6_18_g556( \1887 , \1407 , \1643 );
and mul_6_18_g557( \1888 , \1416 , \1641 );
nor mul_6_18_g558( \1889 , \1887 , \1888 );
xnor mul_6_18_g559( \1890 , \1889 , \1649 );
xor mul_6_18_g560( \1891 , \1886 , \1890 );
and mul_6_18_g561( \1892 , \1526 , \1524 );
and mul_6_18_g562( \1893 , \1622 , \1522 );
nor mul_6_18_g563( \1894 , \1892 , \1893 );
xnor mul_6_18_g564( \1895 , \1894 , \1531 );
xor mul_6_18_g565( \1896 , \1891 , \1895 );
xor mul_6_18_g566( \1897 , \1882 , \1896 );
xor mul_6_18_g567( \1898 , \1848 , \1897 );
and mul_6_18_g568( \1899 , \1838 , \1898 );
and mul_6_18_g569( \1900 , \1594 , \1898 );
or mul_6_18_g570( \1901 , \1839 , \1899 , \1900 );
xor mul_6_18_g571( \1902 , \1788 , \1792 );
xor mul_6_18_g572( \1903 , \1902 , \1795 );
xor mul_6_18_g573( \1904 , \1757 , \1761 );
xor mul_6_18_g574( \1905 , \1904 , \1766 );
and mul_6_18_g575( \1906 , \1903 , \1905 );
xor mul_6_18_g576( \1907 , \1728 , \1732 );
xor mul_6_18_g577( \1908 , \1907 , \1737 );
and mul_6_18_g578( \1909 , \1905 , \1908 );
and mul_6_18_g579( \1910 , \1903 , \1908 );
or mul_6_18_g580( \1911 , \1906 , \1909 , \1910 );
and mul_6_18_g581( \1912 , \1425 , \1336 );
and mul_6_18_g582( \1913 , \1433 , \1333 );
nor mul_6_18_g583( \1914 , \1912 , \1913 );
xnor mul_6_18_g584( \1915 , \1914 , \1332 );
and mul_6_18_g585( \1916 , \1462 , \1349 );
and mul_6_18_g586( \1917 , \1376 , \1347 );
nor mul_6_18_g587( \1918 , \1916 , \1917 );
xnor mul_6_18_g588( \1919 , \1918 , \1356 );
and mul_6_18_g589( \1920 , \1915 , \1919 );
and mul_6_18_g590( \1921 , \1498 , \1522 );
not mul_6_18_g591( \1922 , \1921 );
and mul_6_18_g592( \1923 , \1922 , \1531 );
and mul_6_18_g593( \1924 , \1919 , \1923 );
and mul_6_18_g594( \1925 , \1915 , \1923 );
or mul_6_18_g595( \1926 , \1920 , \1924 , \1925 );
and mul_6_18_g596( \1927 , \1368 , \1460 );
and mul_6_18_g597( \1928 , \1470 , \1458 );
nor mul_6_18_g598( \1929 , \1927 , \1928 );
xnor mul_6_18_g599( \1930 , \1929 , \1467 );
and mul_6_18_g600( \1931 , \1399 , \1475 );
and mul_6_18_g601( \1932 , \1359 , \1473 );
nor mul_6_18_g602( \1933 , \1931 , \1932 );
xnor mul_6_18_g603( \1934 , \1933 , \1482 );
and mul_6_18_g604( \1935 , \1930 , \1934 );
and mul_6_18_g605( \1936 , \1517 , \1414 );
and mul_6_18_g606( \1937 , \1526 , \1412 );
nor mul_6_18_g607( \1938 , \1936 , \1937 );
xnor mul_6_18_g608( \1939 , \1938 , \1421 );
and mul_6_18_g609( \1940 , \1934 , \1939 );
and mul_6_18_g610( \1941 , \1930 , \1939 );
or mul_6_18_g611( \1942 , \1935 , \1940 , \1941 );
and mul_6_18_g612( \1943 , \1926 , \1942 );
and mul_6_18_g613( \1944 , \1477 , \1382 );
and mul_6_18_g614( \1945 , \1454 , \1380 );
nor mul_6_18_g615( \1946 , \1944 , \1945 );
xnor mul_6_18_g616( \1947 , \1946 , \1389 );
and mul_6_18_g617( \1948 , \1616 , \1366 );
and mul_6_18_g618( \1949 , \1391 , \1364 );
nor mul_6_18_g619( \1950 , \1948 , \1949 );
xnor mul_6_18_g620( \1951 , \1950 , \1373 );
and mul_6_18_g621( \1952 , \1947 , \1951 );
and mul_6_18_g622( \1953 , \1416 , \1397 );
and mul_6_18_g623( \1954 , \1586 , \1395 );
nor mul_6_18_g624( \1955 , \1953 , \1954 );
xnor mul_6_18_g625( \1956 , \1955 , \1404 );
and mul_6_18_g626( \1957 , \1951 , \1956 );
and mul_6_18_g627( \1958 , \1947 , \1956 );
or mul_6_18_g628( \1959 , \1952 , \1957 , \1958 );
and mul_6_18_g629( \1960 , \1942 , \1959 );
and mul_6_18_g630( \1961 , \1926 , \1959 );
or mul_6_18_g631( \1962 , \1943 , \1960 , \1961 );
xor mul_6_18_g632( \1963 , \1633 , \1637 );
and mul_6_18_g633( \1964 , \1622 , \1675 );
and mul_6_18_g634( \1965 , \1407 , \1673 );
nor mul_6_18_g635( \1966 , \1964 , \1965 );
xnor mul_6_18_g636( \1967 , \1966 , \1681 );
and mul_6_18_g637( \1968 , \1963 , \1967 );
and mul_6_18_g638( \1969 , \1533 , \1643 );
and mul_6_18_g639( \1970 , \1540 , \1641 );
nor mul_6_18_g640( \1971 , \1969 , \1970 );
xnor mul_6_18_g641( \1972 , \1971 , \1649 );
and mul_6_18_g642( \1973 , \1967 , \1972 );
and mul_6_18_g643( \1974 , \1963 , \1972 );
or mul_6_18_g644( \1975 , \1968 , \1973 , \1974 );
xor mul_6_18_g645( \1976 , \1748 , \1752 );
xor mul_6_18_g646( \1977 , \1976 , \1754 );
and mul_6_18_g647( \1978 , \1975 , \1977 );
xor mul_6_18_g648( \1979 , \1598 , \1602 );
xor mul_6_18_g649( \1980 , \1979 , \1607 );
and mul_6_18_g650( \1981 , \1977 , \1980 );
and mul_6_18_g651( \1982 , \1975 , \1980 );
or mul_6_18_g652( \1983 , \1978 , \1981 , \1982 );
and mul_6_18_g653( \1984 , \1962 , \1983 );
xor mul_6_18_g654( \1985 , \1610 , \1628 );
xor mul_6_18_g655( \1986 , \1985 , \1658 );
and mul_6_18_g656( \1987 , \1983 , \1986 );
and mul_6_18_g657( \1988 , \1962 , \1986 );
or mul_6_18_g658( \1989 , \1984 , \1987 , \1988 );
and mul_6_18_g659( \1990 , \1911 , \1989 );
xor mul_6_18_g660( \1991 , \1375 , \1423 );
xor mul_6_18_g661( \1992 , \1991 , \1484 );
and mul_6_18_g662( \1993 , \1989 , \1992 );
and mul_6_18_g663( \1994 , \1911 , \1992 );
or mul_6_18_g664( \1995 , \1990 , \1993 , \1994 );
and mul_6_18_g665( \1996 , \1722 , \1726 );
and mul_6_18_g666( \1997 , \1726 , \1740 );
and mul_6_18_g667( \1998 , \1722 , \1740 );
or mul_6_18_g668( \1999 , \1996 , \1997 , \1998 );
and mul_6_18_g669( \2000 , \1798 , \1802 );
and mul_6_18_g670( \2001 , \1802 , \1805 );
and mul_6_18_g671( \2002 , \1798 , \1805 );
or mul_6_18_g672( \2003 , \2000 , \2001 , \2002 );
xor mul_6_18_g673( \2004 , \1999 , \2003 );
xor mul_6_18_g674( \2005 , \1855 , \1859 );
xor mul_6_18_g675( \2006 , \2005 , \1864 );
xor mul_6_18_g676( \2007 , \2004 , \2006 );
and mul_6_18_g677( \2008 , \1995 , \2007 );
xor mul_6_18_g678( \2009 , \1487 , \1515 );
xor mul_6_18_g679( \2010 , \2009 , \1591 );
and mul_6_18_g680( \2011 , \2007 , \2010 );
and mul_6_18_g681( \2012 , \1995 , \2010 );
or mul_6_18_g682( \2013 , \2008 , \2011 , \2012 );
and mul_6_18_g683( \2014 , \1999 , \2003 );
and mul_6_18_g684( \2015 , \2003 , \2006 );
and mul_6_18_g685( \2016 , \1999 , \2006 );
or mul_6_18_g686( \2017 , \2014 , \2015 , \2016 );
and mul_6_18_g687( \2018 , \1532 , \1546 );
and mul_6_18_g688( \2019 , \1546 , \1559 );
and mul_6_18_g689( \2020 , \1532 , \1559 );
or mul_6_18_g690( \2021 , \2018 , \2019 , \2020 );
and mul_6_18_g691( \2022 , \1821 , \1336 );
buf mul_6_18_g692( \2023 , \1179_A[30] );
and mul_6_18_g693( \2024 , \2023 , \1333 );
nor mul_6_18_g694( \2025 , \2022 , \2024 );
xnor mul_6_18_g695( \2026 , \2025 , \1332 );
and mul_6_18_g696( \2027 , \1446 , \1349 );
and mul_6_18_g697( \2028 , \1425 , \1347 );
nor mul_6_18_g698( \2029 , \2027 , \2028 );
xnor mul_6_18_g699( \2030 , \2029 , \1356 );
xor mul_6_18_g700( \2031 , \2026 , \2030 );
and mul_6_18_g701( \2032 , \1470 , \1366 );
and mul_6_18_g702( \2033 , \1477 , \1364 );
nor mul_6_18_g703( \2034 , \2032 , \2033 );
xnor mul_6_18_g704( \2035 , \2034 , \1373 );
xor mul_6_18_g705( \2036 , \2031 , \2035 );
xor mul_6_18_g706( \2037 , \2021 , \2036 );
and mul_6_18_g707( \2038 , \1852 , \1854 );
and mul_6_18_g708( \2039 , \1376 , \1460 );
and mul_6_18_g709( \2040 , \1384 , \1458 );
nor mul_6_18_g710( \2041 , \2039 , \2040 );
xnor mul_6_18_g711( \2042 , \2041 , \1467 );
xor mul_6_18_g712( \2043 , \2038 , \2042 );
and mul_6_18_g713( \2044 , \1454 , \1475 );
and mul_6_18_g714( \2045 , \1462 , \1473 );
nor mul_6_18_g715( \2046 , \2044 , \2045 );
xnor mul_6_18_g716( \2047 , \2046 , \1482 );
xor mul_6_18_g717( \2048 , \2043 , \2047 );
xor mul_6_18_g718( \2049 , \2037 , \2048 );
xor mul_6_18_g719( \2050 , \2017 , \2049 );
and mul_6_18_g720( \2051 , \1505 , \1509 );
and mul_6_18_g721( \2052 , \1509 , \1514 );
and mul_6_18_g722( \2053 , \1505 , \1514 );
or mul_6_18_g723( \2054 , \2051 , \2052 , \2053 );
and mul_6_18_g724( \2055 , \1564 , \1568 );
and mul_6_18_g725( \2056 , \1568 , \1573 );
and mul_6_18_g726( \2057 , \1564 , \1573 );
or mul_6_18_g727( \2058 , \2055 , \2056 , \2057 );
and mul_6_18_g728( \2059 , \1579 , \1583 );
and mul_6_18_g729( \2060 , \1583 , \1589 );
and mul_6_18_g730( \2061 , \1579 , \1589 );
or mul_6_18_g731( \2062 , \2059 , \2060 , \2061 );
xor mul_6_18_g732( \2063 , \2058 , \2062 );
and mul_6_18_g733( \2064 , \1824 , \1828 );
and mul_6_18_g734( \2065 , \1828 , \1833 );
and mul_6_18_g735( \2066 , \1824 , \1833 );
or mul_6_18_g736( \2067 , \2064 , \2065 , \2066 );
xor mul_6_18_g737( \2068 , \2063 , \2067 );
xor mul_6_18_g738( \2069 , \2054 , \2068 );
and mul_6_18_g739( \2070 , \1540 , \1538 );
and mul_6_18_g740( \2071 , \1517 , \1536 );
nor mul_6_18_g741( \2072 , \2070 , \2071 );
xnor mul_6_18_g742( \2073 , \2072 , \1545 );
and mul_6_18_g743( \2074 , \1553 , \1551 );
and mul_6_18_g744( \2075 , \1533 , \1501 );
nor mul_6_18_g745( \2076 , \2074 , \2075 );
xnor mul_6_18_g746( \2077 , \2076 , \1558 );
xor mul_6_18_g747( \2078 , \2073 , \2077 );
and mul_6_18_g748( \2079 , \1331 , \1431 );
and mul_6_18_g749( \2080 , \1338 , \1429 );
nor mul_6_18_g750( \2081 , \2079 , \2080 );
xnor mul_6_18_g751( \2082 , \2081 , \1438 );
and mul_6_18_g752( \2083 , \1433 , \1444 );
and mul_6_18_g753( \2084 , \1489 , \1442 );
nor mul_6_18_g754( \2085 , \2083 , \2084 );
xnor mul_6_18_g755( \2086 , \2085 , \1451 );
xor mul_6_18_g756( \2087 , \2082 , \2086 );
buf mul_6_18_g757( \2088 , \1300_B[30] );
xor mul_6_18_g758( \2089 , \2088 , \1548 );
and mul_6_18_g759( \2090 , \1498 , \2089 );
xor mul_6_18_g760( \2091 , \2087 , \2090 );
xor mul_6_18_g761( \2092 , \2078 , \2091 );
xor mul_6_18_g762( \2093 , \2069 , \2092 );
xor mul_6_18_g763( \2094 , \2050 , \2093 );
and mul_6_18_g764( \2095 , \2013 , \2094 );
xor mul_6_18_g765( \2096 , \1594 , \1838 );
xor mul_6_18_g766( \2097 , \2096 , \1898 );
and mul_6_18_g767( \2098 , \2094 , \2097 );
and mul_6_18_g768( \2099 , \2013 , \2097 );
or mul_6_18_g769( \2100 , \2095 , \2098 , \2099 );
xor mul_6_18_g770( \2101 , \1901 , \2100 );
and mul_6_18_g771( \2102 , \2017 , \2049 );
and mul_6_18_g772( \2103 , \2049 , \2093 );
and mul_6_18_g773( \2104 , \2017 , \2093 );
or mul_6_18_g774( \2105 , \2102 , \2103 , \2104 );
and mul_6_18_g775( \2106 , \2054 , \2068 );
and mul_6_18_g776( \2107 , \2068 , \2092 );
and mul_6_18_g777( \2108 , \2054 , \2092 );
or mul_6_18_g778( \2109 , \2106 , \2107 , \2108 );
and mul_6_18_g779( \2110 , \1871 , \1875 );
and mul_6_18_g780( \2111 , \1875 , \1880 );
and mul_6_18_g781( \2112 , \1871 , \1880 );
or mul_6_18_g782( \2113 , \2110 , \2111 , \2112 );
and mul_6_18_g783( \2114 , \2073 , \2077 );
and mul_6_18_g784( \2115 , \2077 , \2091 );
and mul_6_18_g785( \2116 , \2073 , \2091 );
or mul_6_18_g786( \2117 , \2114 , \2115 , \2116 );
xor mul_6_18_g787( \2118 , \2113 , \2117 );
and mul_6_18_g788( \2119 , \1399 , \1675 );
and mul_6_18_g789( \2120 , \1359 , \1673 );
nor mul_6_18_g790( \2121 , \2119 , \2120 );
xnor mul_6_18_g791( \2122 , \2121 , \1681 );
and mul_6_18_g792( \2123 , \1517 , \1538 );
and mul_6_18_g793( \2124 , \1526 , \1536 );
nor mul_6_18_g794( \2125 , \2123 , \2124 );
xnor mul_6_18_g795( \2126 , \2125 , \1545 );
xor mul_6_18_g796( \2127 , \2122 , \2126 );
and mul_6_18_g797( \2128 , \1533 , \1551 );
and mul_6_18_g798( \2129 , \1540 , \1501 );
nor mul_6_18_g799( \2130 , \2128 , \2129 );
xnor mul_6_18_g800( \2131 , \2130 , \1558 );
xor mul_6_18_g801( \2132 , \2127 , \2131 );
xor mul_6_18_g802( \2133 , \2118 , \2132 );
xor mul_6_18_g803( \2134 , \2109 , \2133 );
and mul_6_18_g804( \2135 , \1886 , \1890 );
and mul_6_18_g805( \2136 , \1890 , \1895 );
and mul_6_18_g806( \2137 , \1886 , \1895 );
or mul_6_18_g807( \2138 , \2135 , \2136 , \2137 );
and mul_6_18_g808( \2139 , \2038 , \2042 );
and mul_6_18_g809( \2140 , \2042 , \2047 );
and mul_6_18_g810( \2141 , \2038 , \2047 );
or mul_6_18_g811( \2142 , \2139 , \2140 , \2141 );
xor mul_6_18_g812( \2143 , \2138 , \2142 );
and mul_6_18_g813( \2144 , \1338 , \1431 );
and mul_6_18_g814( \2145 , \1821 , \1429 );
nor mul_6_18_g815( \2146 , \2144 , \2145 );
xnor mul_6_18_g816( \2147 , \2146 , \1438 );
and mul_6_18_g817( \2148 , \1489 , \1444 );
and mul_6_18_g818( \2149 , \1331 , \1442 );
nor mul_6_18_g819( \2150 , \2148 , \2149 );
xnor mul_6_18_g820( \2151 , \2150 , \1451 );
xor mul_6_18_g821( \2152 , \2147 , \2151 );
and mul_6_18_g822( \2153 , \1616 , \1414 );
and mul_6_18_g823( \2154 , \1391 , \1412 );
nor mul_6_18_g824( \2155 , \2153 , \2154 );
xnor mul_6_18_g825( \2156 , \2155 , \1421 );
xor mul_6_18_g826( \2157 , \2152 , \2156 );
and mul_6_18_g827( \2158 , \1622 , \1524 );
and mul_6_18_g828( \2159 , \1407 , \1522 );
nor mul_6_18_g829( \2160 , \2158 , \2159 );
xnor mul_6_18_g830( \2161 , \2160 , \1531 );
xor mul_6_18_g831( \2162 , \2157 , \2161 );
xor mul_6_18_g832( \2163 , \2143 , \2162 );
and mul_6_18_g833( \2164 , \1425 , \1349 );
and mul_6_18_g834( \2165 , \1433 , \1347 );
nor mul_6_18_g835( \2166 , \2164 , \2165 );
xnor mul_6_18_g836( \2167 , \2166 , \1356 );
and mul_6_18_g837( \2168 , \1462 , \1475 );
and mul_6_18_g838( \2169 , \1376 , \1473 );
nor mul_6_18_g839( \2170 , \2168 , \2169 );
xnor mul_6_18_g840( \2171 , \2170 , \1482 );
xor mul_6_18_g841( \2172 , \2167 , \2171 );
and mul_6_18_g842( \2173 , \1477 , \1366 );
and mul_6_18_g843( \2174 , \1454 , \1364 );
nor mul_6_18_g844( \2175 , \2173 , \2174 );
xnor mul_6_18_g845( \2176 , \2175 , \1373 );
xor mul_6_18_g846( \2177 , \2172 , \2176 );
and mul_6_18_g847( \2178 , \1368 , \1397 );
and mul_6_18_g848( \2179 , \1470 , \1395 );
nor mul_6_18_g849( \2180 , \2178 , \2179 );
xnor mul_6_18_g850( \2181 , \2180 , \1404 );
xor mul_6_18_g851( \2182 , \2177 , \2181 );
xor mul_6_18_g852( \2183 , \2163 , \2182 );
xor mul_6_18_g853( \2184 , \2134 , \2183 );
xor mul_6_18_g854( \2185 , \2105 , \2184 );
and mul_6_18_g855( \2186 , \2058 , \2062 );
and mul_6_18_g856( \2187 , \2062 , \2067 );
and mul_6_18_g857( \2188 , \2058 , \2067 );
or mul_6_18_g858( \2189 , \2186 , \2187 , \2188 );
and mul_6_18_g859( \2190 , \2021 , \2036 );
and mul_6_18_g860( \2191 , \2036 , \2048 );
and mul_6_18_g861( \2192 , \2021 , \2048 );
or mul_6_18_g862( \2193 , \2190 , \2191 , \2192 );
xor mul_6_18_g863( \2194 , \2189 , \2193 );
and mul_6_18_g864( \2195 , \1867 , \1881 );
and mul_6_18_g865( \2196 , \1881 , \1896 );
and mul_6_18_g866( \2197 , \1867 , \1896 );
or mul_6_18_g867( \2198 , \2195 , \2196 , \2197 );
and mul_6_18_g868( \2199 , \1843 , \1847 );
and mul_6_18_g869( \2200 , \1847 , \1897 );
and mul_6_18_g870( \2201 , \1843 , \1897 );
or mul_6_18_g871( \2202 , \2199 , \2200 , \2201 );
xor mul_6_18_g872( \2203 , \2198 , \2202 );
and mul_6_18_g873( \2204 , \2026 , \2030 );
and mul_6_18_g874( \2205 , \2030 , \2035 );
and mul_6_18_g875( \2206 , \2026 , \2035 );
or mul_6_18_g876( \2207 , \2204 , \2205 , \2206 );
and mul_6_18_g877( \2208 , \2082 , \2086 );
and mul_6_18_g878( \2209 , \2086 , \2090 );
and mul_6_18_g879( \2210 , \2082 , \2090 );
or mul_6_18_g880( \2211 , \2208 , \2209 , \2210 );
xor mul_6_18_g881( \2212 , \2207 , \2211 );
and mul_6_18_g882( \2213 , \1351 , \1382 );
and mul_6_18_g883( \2214 , \1446 , \1380 );
nor mul_6_18_g884( \2215 , \2213 , \2214 );
xnor mul_6_18_g885( \2216 , \2215 , \1389 );
and mul_6_18_g886( \2217 , \1384 , \1460 );
and mul_6_18_g887( \2218 , \1342 , \1458 );
nor mul_6_18_g888( \2219 , \2217 , \2218 );
xnor mul_6_18_g889( \2220 , \2219 , \1467 );
xor mul_6_18_g890( \2221 , \2216 , \2220 );
and mul_6_18_g891( \2222 , \1416 , \1643 );
and mul_6_18_g892( \2223 , \1586 , \1641 );
nor mul_6_18_g893( \2224 , \2222 , \2223 );
xnor mul_6_18_g894( \2225 , \2224 , \1649 );
xor mul_6_18_g895( \2226 , \2221 , \2225 );
and mul_6_18_g896( \2227 , \2023 , \1336 );
buf mul_6_18_g897( \2228 , \1175_A[31] );
and mul_6_18_g898( \2229 , \2228 , \1333 );
nor mul_6_18_g899( \2230 , \2227 , \2229 );
xnor mul_6_18_g900( \2231 , \2230 , \1332 );
not mul_6_18_g901( \2232 , \2090 );
buf mul_6_18_g902( \2233 , \1299_B[31] );
and mul_6_18_g903( \2234 , \2088 , \1548 );
not mul_6_18_g904( \2235 , \2234 );
and mul_6_18_g905( \2236 , \2233 , \2235 );
and mul_6_18_g906( \2237 , \2232 , \2236 );
xor mul_6_18_g907( \2238 , \2231 , \2237 );
xor mul_6_18_g908( \2239 , \2233 , \2088 );
not mul_6_18_g909( \2240 , \2089 );
and mul_6_18_g910( \2241 , \2239 , \2240 );
and mul_6_18_g911( \2242 , \1498 , \2241 );
and mul_6_18_g912( \2243 , \1553 , \2089 );
nor mul_6_18_g913( \2244 , \2242 , \2243 );
xnor mul_6_18_g914( \2245 , \2244 , \2236 );
xor mul_6_18_g915( \2246 , \2238 , \2245 );
xor mul_6_18_g916( \2247 , \2226 , \2246 );
xor mul_6_18_g917( \2248 , \2212 , \2247 );
xor mul_6_18_g918( \2249 , \2203 , \2248 );
xor mul_6_18_g919( \2250 , \2194 , \2249 );
xor mul_6_18_g920( \2251 , \2185 , \2250 );
xor mul_6_18_g921( \2252 , \2101 , \2251 );
xor mul_6_18_g922( \2253 , \2013 , \2094 );
xor mul_6_18_g923( \2254 , \2253 , \2097 );
xor mul_6_18_g924( \2255 , \1665 , \1669 );
xor mul_6_18_g925( \2256 , \2255 , \1682 );
xor mul_6_18_g926( \2257 , \1614 , \1619 );
xor mul_6_18_g927( \2258 , \2257 , \1625 );
and mul_6_18_g928( \2259 , \2256 , \2258 );
xor mul_6_18_g929( \2260 , \1638 , \1650 );
xor mul_6_18_g930( \2261 , \2260 , \1655 );
and mul_6_18_g931( \2262 , \2258 , \2261 );
and mul_6_18_g932( \2263 , \2256 , \2261 );
or mul_6_18_g933( \2264 , \2259 , \2262 , \2263 );
xor mul_6_18_g934( \2265 , \1685 , \1699 );
xor mul_6_18_g935( \2266 , \2265 , \1714 );
and mul_6_18_g936( \2267 , \2264 , \2266 );
xor mul_6_18_g937( \2268 , \1903 , \1905 );
xor mul_6_18_g938( \2269 , \2268 , \1908 );
and mul_6_18_g939( \2270 , \2266 , \2269 );
and mul_6_18_g940( \2271 , \2264 , \2269 );
or mul_6_18_g941( \2272 , \2267 , \2270 , \2271 );
xor mul_6_18_g942( \2273 , \1661 , \1717 );
xor mul_6_18_g943( \2274 , \2273 , \1741 );
and mul_6_18_g944( \2275 , \2272 , \2274 );
xor mul_6_18_g945( \2276 , \1769 , \1783 );
xor mul_6_18_g946( \2277 , \2276 , \1806 );
and mul_6_18_g947( \2278 , \2274 , \2277 );
and mul_6_18_g948( \2279 , \2272 , \2277 );
or mul_6_18_g949( \2280 , \2275 , \2278 , \2279 );
xor mul_6_18_g950( \2281 , \1744 , \1809 );
xor mul_6_18_g951( \2282 , \2281 , \1835 );
and mul_6_18_g952( \2283 , \2280 , \2282 );
xor mul_6_18_g953( \2284 , \1995 , \2007 );
xor mul_6_18_g954( \2285 , \2284 , \2010 );
and mul_6_18_g955( \2286 , \2282 , \2285 );
and mul_6_18_g956( \2287 , \2280 , \2285 );
or mul_6_18_g957( \2288 , \2283 , \2286 , \2287 );
and mul_6_18_g958( \2289 , \2254 , \2288 );
xor mul_6_18_g959( \2290 , \2254 , \2288 );
and mul_6_18_g960( \2291 , \1342 , \1431 );
and mul_6_18_g961( \2292 , \1351 , \1429 );
nor mul_6_18_g962( \2293 , \2291 , \2292 );
xnor mul_6_18_g963( \2294 , \2293 , \1438 );
and mul_6_18_g964( \2295 , \1376 , \1444 );
and mul_6_18_g965( \2296 , \1384 , \1442 );
nor mul_6_18_g966( \2297 , \2295 , \2296 );
xnor mul_6_18_g967( \2298 , \2297 , \1451 );
and mul_6_18_g968( \2299 , \2294 , \2298 );
and mul_6_18_g969( \2300 , \2298 , \1921 );
and mul_6_18_g970( \2301 , \2294 , \1921 );
or mul_6_18_g971( \2302 , \2299 , \2300 , \2301 );
and mul_6_18_g972( \2303 , \1446 , \1336 );
and mul_6_18_g973( \2304 , \1425 , \1333 );
nor mul_6_18_g974( \2305 , \2303 , \2304 );
xnor mul_6_18_g975( \2306 , \2305 , \1332 );
and mul_6_18_g976( \2307 , \1454 , \1349 );
and mul_6_18_g977( \2308 , \1462 , \1347 );
nor mul_6_18_g978( \2309 , \2307 , \2308 );
xnor mul_6_18_g979( \2310 , \2309 , \1356 );
and mul_6_18_g980( \2311 , \2306 , \2310 );
and mul_6_18_g981( \2312 , \1586 , \1366 );
and mul_6_18_g982( \2313 , \1616 , \1364 );
nor mul_6_18_g983( \2314 , \2312 , \2313 );
xnor mul_6_18_g984( \2315 , \2314 , \1373 );
and mul_6_18_g985( \2316 , \2310 , \2315 );
and mul_6_18_g986( \2317 , \2306 , \2315 );
or mul_6_18_g987( \2318 , \2311 , \2316 , \2317 );
and mul_6_18_g988( \2319 , \2302 , \2318 );
and mul_6_18_g989( \2320 , \1498 , \1524 );
and mul_6_18_g990( \2321 , \1553 , \1522 );
nor mul_6_18_g991( \2322 , \2320 , \2321 );
xnor mul_6_18_g992( \2323 , \2322 , \1531 );
and mul_6_18_g993( \2324 , \2318 , \2323 );
and mul_6_18_g994( \2325 , \2302 , \2323 );
or mul_6_18_g995( \2326 , \2319 , \2324 , \2325 );
and mul_6_18_g996( \2327 , \1470 , \1382 );
and mul_6_18_g997( \2328 , \1477 , \1380 );
nor mul_6_18_g998( \2329 , \2327 , \2328 );
xnor mul_6_18_g999( \2330 , \2329 , \1389 );
and mul_6_18_g1000( \2331 , \1407 , \1397 );
and mul_6_18_g1001( \2332 , \1416 , \1395 );
nor mul_6_18_g1002( \2333 , \2331 , \2332 );
xnor mul_6_18_g1003( \2334 , \2333 , \1404 );
and mul_6_18_g1004( \2335 , \2330 , \2334 );
and mul_6_18_g1005( \2336 , \1540 , \1414 );
and mul_6_18_g1006( \2337 , \1517 , \1412 );
nor mul_6_18_g1007( \2338 , \2336 , \2337 );
xnor mul_6_18_g1008( \2339 , \2338 , \1421 );
and mul_6_18_g1009( \2340 , \2334 , \2339 );
and mul_6_18_g1010( \2341 , \2330 , \2339 );
or mul_6_18_g1011( \2342 , \2335 , \2340 , \2341 );
and mul_6_18_g1012( \2343 , \1359 , \1460 );
and mul_6_18_g1013( \2344 , \1368 , \1458 );
nor mul_6_18_g1014( \2345 , \2343 , \2344 );
xnor mul_6_18_g1015( \2346 , \2345 , \1467 );
and mul_6_18_g1016( \2347 , \1391 , \1475 );
and mul_6_18_g1017( \2348 , \1399 , \1473 );
nor mul_6_18_g1018( \2349 , \2347 , \2348 );
xnor mul_6_18_g1019( \2350 , \2349 , \1482 );
and mul_6_18_g1020( \2351 , \2346 , \2350 );
and mul_6_18_g1021( \2352 , \1526 , \1675 );
and mul_6_18_g1022( \2353 , \1622 , \1673 );
nor mul_6_18_g1023( \2354 , \2352 , \2353 );
xnor mul_6_18_g1024( \2355 , \2354 , \1681 );
and mul_6_18_g1025( \2356 , \2350 , \2355 );
and mul_6_18_g1026( \2357 , \2346 , \2355 );
or mul_6_18_g1027( \2358 , \2351 , \2356 , \2357 );
and mul_6_18_g1028( \2359 , \2342 , \2358 );
xor mul_6_18_g1029( \2360 , \1915 , \1919 );
xor mul_6_18_g1030( \2361 , \2360 , \1923 );
and mul_6_18_g1031( \2362 , \2358 , \2361 );
and mul_6_18_g1032( \2363 , \2342 , \2361 );
or mul_6_18_g1033( \2364 , \2359 , \2362 , \2363 );
and mul_6_18_g1034( \2365 , \2326 , \2364 );
xor mul_6_18_g1035( \2366 , \1926 , \1942 );
xor mul_6_18_g1036( \2367 , \2366 , \1959 );
and mul_6_18_g1037( \2368 , \2364 , \2367 );
and mul_6_18_g1038( \2369 , \2326 , \2367 );
or mul_6_18_g1039( \2370 , \2365 , \2368 , \2369 );
xor mul_6_18_g1040( \2371 , \1930 , \1934 );
xor mul_6_18_g1041( \2372 , \2371 , \1939 );
xor mul_6_18_g1042( \2373 , \1947 , \1951 );
xor mul_6_18_g1043( \2374 , \2373 , \1956 );
and mul_6_18_g1044( \2375 , \2372 , \2374 );
xor mul_6_18_g1045( \2376 , \1963 , \1967 );
xor mul_6_18_g1046( \2377 , \2376 , \1972 );
and mul_6_18_g1047( \2378 , \2374 , \2377 );
and mul_6_18_g1048( \2379 , \2372 , \2377 );
or mul_6_18_g1049( \2380 , \2375 , \2378 , \2379 );
xor mul_6_18_g1050( \2381 , \2256 , \2258 );
xor mul_6_18_g1051( \2382 , \2381 , \2261 );
and mul_6_18_g1052( \2383 , \2380 , \2382 );
xor mul_6_18_g1053( \2384 , \1975 , \1977 );
xor mul_6_18_g1054( \2385 , \2384 , \1980 );
and mul_6_18_g1055( \2386 , \2382 , \2385 );
and mul_6_18_g1056( \2387 , \2380 , \2385 );
or mul_6_18_g1057( \2388 , \2383 , \2386 , \2387 );
and mul_6_18_g1058( \2389 , \2370 , \2388 );
xor mul_6_18_g1059( \2390 , \1962 , \1983 );
xor mul_6_18_g1060( \2391 , \2390 , \1986 );
and mul_6_18_g1061( \2392 , \2388 , \2391 );
and mul_6_18_g1062( \2393 , \2370 , \2391 );
or mul_6_18_g1063( \2394 , \2389 , \2392 , \2393 );
xor mul_6_18_g1064( \2395 , \1911 , \1989 );
xor mul_6_18_g1065( \2396 , \2395 , \1992 );
and mul_6_18_g1066( \2397 , \2394 , \2396 );
xor mul_6_18_g1067( \2398 , \2272 , \2274 );
xor mul_6_18_g1068( \2399 , \2398 , \2277 );
and mul_6_18_g1069( \2400 , \2396 , \2399 );
and mul_6_18_g1070( \2401 , \2394 , \2399 );
or mul_6_18_g1071( \2402 , \2397 , \2400 , \2401 );
xor mul_6_18_g1072( \2403 , \2280 , \2282 );
xor mul_6_18_g1073( \2404 , \2403 , \2285 );
and mul_6_18_g1074( \2405 , \2402 , \2404 );
xor mul_6_18_g1075( \2406 , \2402 , \2404 );
xor mul_6_18_g1076( \2407 , \2394 , \2396 );
xor mul_6_18_g1077( \2408 , \2407 , \2399 );
and mul_6_18_g1078( \2409 , \1368 , \1382 );
and mul_6_18_g1079( \2410 , \1470 , \1380 );
nor mul_6_18_g1080( \2411 , \2409 , \2410 );
xnor mul_6_18_g1081( \2412 , \2411 , \1389 );
and mul_6_18_g1082( \2413 , \1416 , \1366 );
and mul_6_18_g1083( \2414 , \1586 , \1364 );
nor mul_6_18_g1084( \2415 , \2413 , \2414 );
xnor mul_6_18_g1085( \2416 , \2415 , \1373 );
and mul_6_18_g1086( \2417 , \2412 , \2416 );
and mul_6_18_g1087( \2418 , \1622 , \1397 );
and mul_6_18_g1088( \2419 , \1407 , \1395 );
nor mul_6_18_g1089( \2420 , \2418 , \2419 );
xnor mul_6_18_g1090( \2421 , \2420 , \1404 );
and mul_6_18_g1091( \2422 , \2416 , \2421 );
and mul_6_18_g1092( \2423 , \2412 , \2421 );
or mul_6_18_g1093( \2424 , \2417 , \2422 , \2423 );
and mul_6_18_g1094( \2425 , \1384 , \1431 );
and mul_6_18_g1095( \2426 , \1342 , \1429 );
nor mul_6_18_g1096( \2427 , \2425 , \2426 );
xnor mul_6_18_g1097( \2428 , \2427 , \1438 );
and mul_6_18_g1098( \2429 , \1462 , \1444 );
and mul_6_18_g1099( \2430 , \1376 , \1442 );
nor mul_6_18_g1100( \2431 , \2429 , \2430 );
xnor mul_6_18_g1101( \2432 , \2431 , \1451 );
and mul_6_18_g1102( \2433 , \2428 , \2432 );
and mul_6_18_g1103( \2434 , \2424 , \2433 );
and mul_6_18_g1104( \2435 , \1553 , \1643 );
and mul_6_18_g1105( \2436 , \1533 , \1641 );
nor mul_6_18_g1106( \2437 , \2435 , \2436 );
xnor mul_6_18_g1107( \2438 , \2437 , \1649 );
and mul_6_18_g1108( \2439 , \2433 , \2438 );
and mul_6_18_g1109( \2440 , \2424 , \2438 );
or mul_6_18_g1110( \2441 , \2434 , \2439 , \2440 );
and mul_6_18_g1111( \2442 , \1399 , \1460 );
and mul_6_18_g1112( \2443 , \1359 , \1458 );
nor mul_6_18_g1113( \2444 , \2442 , \2443 );
xnor mul_6_18_g1114( \2445 , \2444 , \1467 );
and mul_6_18_g1115( \2446 , \1616 , \1475 );
and mul_6_18_g1116( \2447 , \1391 , \1473 );
nor mul_6_18_g1117( \2448 , \2446 , \2447 );
xnor mul_6_18_g1118( \2449 , \2448 , \1482 );
and mul_6_18_g1119( \2450 , \2445 , \2449 );
and mul_6_18_g1120( \2451 , \1533 , \1414 );
and mul_6_18_g1121( \2452 , \1540 , \1412 );
nor mul_6_18_g1122( \2453 , \2451 , \2452 );
xnor mul_6_18_g1123( \2454 , \2453 , \1421 );
and mul_6_18_g1124( \2455 , \2449 , \2454 );
and mul_6_18_g1125( \2456 , \2445 , \2454 );
or mul_6_18_g1126( \2457 , \2450 , \2455 , \2456 );
and mul_6_18_g1127( \2458 , \1351 , \1336 );
and mul_6_18_g1128( \2459 , \1446 , \1333 );
nor mul_6_18_g1129( \2460 , \2458 , \2459 );
xnor mul_6_18_g1130( \2461 , \2460 , \1332 );
and mul_6_18_g1131( \2462 , \1477 , \1349 );
and mul_6_18_g1132( \2463 , \1454 , \1347 );
nor mul_6_18_g1133( \2464 , \2462 , \2463 );
xnor mul_6_18_g1134( \2465 , \2464 , \1356 );
and mul_6_18_g1135( \2466 , \2461 , \2465 );
and mul_6_18_g1136( \2467 , \1498 , \1641 );
not mul_6_18_g1137( \2468 , \2467 );
and mul_6_18_g1138( \2469 , \2468 , \1649 );
and mul_6_18_g1139( \2470 , \2465 , \2469 );
and mul_6_18_g1140( \2471 , \2461 , \2469 );
or mul_6_18_g1141( \2472 , \2466 , \2470 , \2471 );
and mul_6_18_g1142( \2473 , \2457 , \2472 );
xor mul_6_18_g1143( \2474 , \2294 , \2298 );
xor mul_6_18_g1144( \2475 , \2474 , \1921 );
and mul_6_18_g1145( \2476 , \2472 , \2475 );
and mul_6_18_g1146( \2477 , \2457 , \2475 );
or mul_6_18_g1147( \2478 , \2473 , \2476 , \2477 );
and mul_6_18_g1148( \2479 , \2441 , \2478 );
xor mul_6_18_g1149( \2480 , \2302 , \2318 );
xor mul_6_18_g1150( \2481 , \2480 , \2323 );
and mul_6_18_g1151( \2482 , \2478 , \2481 );
and mul_6_18_g1152( \2483 , \2441 , \2481 );
or mul_6_18_g1153( \2484 , \2479 , \2482 , \2483 );
xor mul_6_18_g1154( \2485 , \2306 , \2310 );
xor mul_6_18_g1155( \2486 , \2485 , \2315 );
xor mul_6_18_g1156( \2487 , \2330 , \2334 );
xor mul_6_18_g1157( \2488 , \2487 , \2339 );
and mul_6_18_g1158( \2489 , \2486 , \2488 );
xor mul_6_18_g1159( \2490 , \2346 , \2350 );
xor mul_6_18_g1160( \2491 , \2490 , \2355 );
and mul_6_18_g1161( \2492 , \2488 , \2491 );
and mul_6_18_g1162( \2493 , \2486 , \2491 );
or mul_6_18_g1163( \2494 , \2489 , \2492 , \2493 );
xor mul_6_18_g1164( \2495 , \2342 , \2358 );
xor mul_6_18_g1165( \2496 , \2495 , \2361 );
and mul_6_18_g1166( \2497 , \2494 , \2496 );
xor mul_6_18_g1167( \2498 , \2372 , \2374 );
xor mul_6_18_g1168( \2499 , \2498 , \2377 );
and mul_6_18_g1169( \2500 , \2496 , \2499 );
and mul_6_18_g1170( \2501 , \2494 , \2499 );
or mul_6_18_g1171( \2502 , \2497 , \2500 , \2501 );
and mul_6_18_g1172( \2503 , \2484 , \2502 );
xor mul_6_18_g1173( \2504 , \2326 , \2364 );
xor mul_6_18_g1174( \2505 , \2504 , \2367 );
and mul_6_18_g1175( \2506 , \2502 , \2505 );
and mul_6_18_g1176( \2507 , \2484 , \2505 );
or mul_6_18_g1177( \2508 , \2503 , \2506 , \2507 );
xor mul_6_18_g1178( \2509 , \2264 , \2266 );
xor mul_6_18_g1179( \2510 , \2509 , \2269 );
and mul_6_18_g1180( \2511 , \2508 , \2510 );
xor mul_6_18_g1181( \2512 , \2370 , \2388 );
xor mul_6_18_g1182( \2513 , \2512 , \2391 );
and mul_6_18_g1183( \2514 , \2510 , \2513 );
and mul_6_18_g1184( \2515 , \2508 , \2513 );
or mul_6_18_g1185( \2516 , \2511 , \2514 , \2515 );
and mul_6_18_g1186( \2517 , \2408 , \2516 );
xor mul_6_18_g1187( \2518 , \2408 , \2516 );
xor mul_6_18_g1188( \2519 , \2508 , \2510 );
xor mul_6_18_g1189( \2520 , \2519 , \2513 );
and mul_6_18_g1190( \2521 , \1376 , \1431 );
and mul_6_18_g1191( \2522 , \1384 , \1429 );
nor mul_6_18_g1192( \2523 , \2521 , \2522 );
xnor mul_6_18_g1193( \2524 , \2523 , \1438 );
and mul_6_18_g1194( \2525 , \1454 , \1444 );
and mul_6_18_g1195( \2526 , \1462 , \1442 );
nor mul_6_18_g1196( \2527 , \2525 , \2526 );
xnor mul_6_18_g1197( \2528 , \2527 , \1451 );
and mul_6_18_g1198( \2529 , \2524 , \2528 );
and mul_6_18_g1199( \2530 , \2528 , \2467 );
and mul_6_18_g1200( \2531 , \2524 , \2467 );
or mul_6_18_g1201( \2532 , \2529 , \2530 , \2531 );
and mul_6_18_g1202( \2533 , \1359 , \1382 );
and mul_6_18_g1203( \2534 , \1368 , \1380 );
nor mul_6_18_g1204( \2535 , \2533 , \2534 );
xnor mul_6_18_g1205( \2536 , \2535 , \1389 );
and mul_6_18_g1206( \2537 , \1526 , \1397 );
and mul_6_18_g1207( \2538 , \1622 , \1395 );
nor mul_6_18_g1208( \2539 , \2537 , \2538 );
xnor mul_6_18_g1209( \2540 , \2539 , \1404 );
and mul_6_18_g1210( \2541 , \2536 , \2540 );
and mul_6_18_g1211( \2542 , \1553 , \1414 );
and mul_6_18_g1212( \2543 , \1533 , \1412 );
nor mul_6_18_g1213( \2544 , \2542 , \2543 );
xnor mul_6_18_g1214( \2545 , \2544 , \1421 );
and mul_6_18_g1215( \2546 , \2540 , \2545 );
and mul_6_18_g1216( \2547 , \2536 , \2545 );
or mul_6_18_g1217( \2548 , \2541 , \2546 , \2547 );
and mul_6_18_g1218( \2549 , \2532 , \2548 );
and mul_6_18_g1219( \2550 , \1342 , \1336 );
and mul_6_18_g1220( \2551 , \1351 , \1333 );
nor mul_6_18_g1221( \2552 , \2550 , \2551 );
xnor mul_6_18_g1222( \2553 , \2552 , \1332 );
and mul_6_18_g1223( \2554 , \1470 , \1349 );
and mul_6_18_g1224( \2555 , \1477 , \1347 );
nor mul_6_18_g1225( \2556 , \2554 , \2555 );
xnor mul_6_18_g1226( \2557 , \2556 , \1356 );
and mul_6_18_g1227( \2558 , \2553 , \2557 );
and mul_6_18_g1228( \2559 , \1407 , \1366 );
and mul_6_18_g1229( \2560 , \1416 , \1364 );
nor mul_6_18_g1230( \2561 , \2559 , \2560 );
xnor mul_6_18_g1231( \2562 , \2561 , \1373 );
and mul_6_18_g1232( \2563 , \2557 , \2562 );
and mul_6_18_g1233( \2564 , \2553 , \2562 );
or mul_6_18_g1234( \2565 , \2558 , \2563 , \2564 );
and mul_6_18_g1235( \2566 , \2548 , \2565 );
and mul_6_18_g1236( \2567 , \2532 , \2565 );
or mul_6_18_g1237( \2568 , \2549 , \2566 , \2567 );
xor mul_6_18_g1238( \2569 , \2428 , \2432 );
and mul_6_18_g1239( \2570 , \1517 , \1675 );
and mul_6_18_g1240( \2571 , \1526 , \1673 );
nor mul_6_18_g1241( \2572 , \2570 , \2571 );
xnor mul_6_18_g1242( \2573 , \2572 , \1681 );
and mul_6_18_g1243( \2574 , \2569 , \2573 );
and mul_6_18_g1244( \2575 , \1498 , \1643 );
and mul_6_18_g1245( \2576 , \1553 , \1641 );
nor mul_6_18_g1246( \2577 , \2575 , \2576 );
xnor mul_6_18_g1247( \2578 , \2577 , \1649 );
and mul_6_18_g1248( \2579 , \2573 , \2578 );
and mul_6_18_g1249( \2580 , \2569 , \2578 );
or mul_6_18_g1250( \2581 , \2574 , \2579 , \2580 );
and mul_6_18_g1251( \2582 , \2568 , \2581 );
xor mul_6_18_g1252( \2583 , \2424 , \2433 );
xor mul_6_18_g1253( \2584 , \2583 , \2438 );
and mul_6_18_g1254( \2585 , \2581 , \2584 );
and mul_6_18_g1255( \2586 , \2568 , \2584 );
or mul_6_18_g1256( \2587 , \2582 , \2585 , \2586 );
and mul_6_18_g1257( \2588 , \1391 , \1460 );
and mul_6_18_g1258( \2589 , \1399 , \1458 );
nor mul_6_18_g1259( \2590 , \2588 , \2589 );
xnor mul_6_18_g1260( \2591 , \2590 , \1467 );
and mul_6_18_g1261( \2592 , \1586 , \1475 );
and mul_6_18_g1262( \2593 , \1616 , \1473 );
nor mul_6_18_g1263( \2594 , \2592 , \2593 );
xnor mul_6_18_g1264( \2595 , \2594 , \1482 );
and mul_6_18_g1265( \2596 , \2591 , \2595 );
and mul_6_18_g1266( \2597 , \1540 , \1675 );
and mul_6_18_g1267( \2598 , \1517 , \1673 );
nor mul_6_18_g1268( \2599 , \2597 , \2598 );
xnor mul_6_18_g1269( \2600 , \2599 , \1681 );
and mul_6_18_g1270( \2601 , \2595 , \2600 );
and mul_6_18_g1271( \2602 , \2591 , \2600 );
or mul_6_18_g1272( \2603 , \2596 , \2601 , \2602 );
xor mul_6_18_g1273( \2604 , \2412 , \2416 );
xor mul_6_18_g1274( \2605 , \2604 , \2421 );
and mul_6_18_g1275( \2606 , \2603 , \2605 );
xor mul_6_18_g1276( \2607 , \2445 , \2449 );
xor mul_6_18_g1277( \2608 , \2607 , \2454 );
and mul_6_18_g1278( \2609 , \2605 , \2608 );
and mul_6_18_g1279( \2610 , \2603 , \2608 );
or mul_6_18_g1280( \2611 , \2606 , \2609 , \2610 );
xor mul_6_18_g1281( \2612 , \2457 , \2472 );
xor mul_6_18_g1282( \2613 , \2612 , \2475 );
and mul_6_18_g1283( \2614 , \2611 , \2613 );
xor mul_6_18_g1284( \2615 , \2486 , \2488 );
xor mul_6_18_g1285( \2616 , \2615 , \2491 );
and mul_6_18_g1286( \2617 , \2613 , \2616 );
and mul_6_18_g1287( \2618 , \2611 , \2616 );
or mul_6_18_g1288( \2619 , \2614 , \2617 , \2618 );
and mul_6_18_g1289( \2620 , \2587 , \2619 );
xor mul_6_18_g1290( \2621 , \2441 , \2478 );
xor mul_6_18_g1291( \2622 , \2621 , \2481 );
and mul_6_18_g1292( \2623 , \2619 , \2622 );
and mul_6_18_g1293( \2624 , \2587 , \2622 );
or mul_6_18_g1294( \2625 , \2620 , \2623 , \2624 );
xor mul_6_18_g1295( \2626 , \2380 , \2382 );
xor mul_6_18_g1296( \2627 , \2626 , \2385 );
and mul_6_18_g1297( \2628 , \2625 , \2627 );
xor mul_6_18_g1298( \2629 , \2484 , \2502 );
xor mul_6_18_g1299( \2630 , \2629 , \2505 );
and mul_6_18_g1300( \2631 , \2627 , \2630 );
and mul_6_18_g1301( \2632 , \2625 , \2630 );
or mul_6_18_g1302( \2633 , \2628 , \2631 , \2632 );
and mul_6_18_g1303( \2634 , \2520 , \2633 );
xor mul_6_18_g1304( \2635 , \2520 , \2633 );
xor mul_6_18_g1305( \2636 , \2625 , \2627 );
xor mul_6_18_g1306( \2637 , \2636 , \2630 );
and mul_6_18_g1307( \2638 , \1616 , \1460 );
and mul_6_18_g1308( \2639 , \1391 , \1458 );
nor mul_6_18_g1309( \2640 , \2638 , \2639 );
xnor mul_6_18_g1310( \2641 , \2640 , \1467 );
and mul_6_18_g1311( \2642 , \1416 , \1475 );
and mul_6_18_g1312( \2643 , \1586 , \1473 );
nor mul_6_18_g1313( \2644 , \2642 , \2643 );
xnor mul_6_18_g1314( \2645 , \2644 , \1482 );
and mul_6_18_g1315( \2646 , \2641 , \2645 );
and mul_6_18_g1316( \2647 , \1498 , \1414 );
and mul_6_18_g1317( \2648 , \1553 , \1412 );
nor mul_6_18_g1318( \2649 , \2647 , \2648 );
xnor mul_6_18_g1319( \2650 , \2649 , \1421 );
and mul_6_18_g1320( \2651 , \2645 , \2650 );
and mul_6_18_g1321( \2652 , \2641 , \2650 );
or mul_6_18_g1322( \2653 , \2646 , \2651 , \2652 );
and mul_6_18_g1323( \2654 , \1399 , \1382 );
and mul_6_18_g1324( \2655 , \1359 , \1380 );
nor mul_6_18_g1325( \2656 , \2654 , \2655 );
xnor mul_6_18_g1326( \2657 , \2656 , \1389 );
and mul_6_18_g1327( \2658 , \1622 , \1366 );
and mul_6_18_g1328( \2659 , \1407 , \1364 );
nor mul_6_18_g1329( \2660 , \2658 , \2659 );
xnor mul_6_18_g1330( \2661 , \2660 , \1373 );
and mul_6_18_g1331( \2662 , \2657 , \2661 );
and mul_6_18_g1332( \2663 , \1517 , \1397 );
and mul_6_18_g1333( \2664 , \1526 , \1395 );
nor mul_6_18_g1334( \2665 , \2663 , \2664 );
xnor mul_6_18_g1335( \2666 , \2665 , \1404 );
and mul_6_18_g1336( \2667 , \2661 , \2666 );
and mul_6_18_g1337( \2668 , \2657 , \2666 );
or mul_6_18_g1338( \2669 , \2662 , \2667 , \2668 );
and mul_6_18_g1339( \2670 , \2653 , \2669 );
and mul_6_18_g1340( \2671 , \1462 , \1431 );
and mul_6_18_g1341( \2672 , \1376 , \1429 );
nor mul_6_18_g1342( \2673 , \2671 , \2672 );
xnor mul_6_18_g1343( \2674 , \2673 , \1438 );
and mul_6_18_g1344( \2675 , \1498 , \1412 );
not mul_6_18_g1345( \2676 , \2675 );
and mul_6_18_g1346( \2677 , \2676 , \1421 );
and mul_6_18_g1347( \2678 , \2674 , \2677 );
and mul_6_18_g1348( \2679 , \2669 , \2678 );
and mul_6_18_g1349( \2680 , \2653 , \2678 );
or mul_6_18_g1350( \2681 , \2670 , \2679 , \2680 );
xor mul_6_18_g1351( \2682 , \2461 , \2465 );
xor mul_6_18_g1352( \2683 , \2682 , \2469 );
and mul_6_18_g1353( \2684 , \2681 , \2683 );
xor mul_6_18_g1354( \2685 , \2569 , \2573 );
xor mul_6_18_g1355( \2686 , \2685 , \2578 );
and mul_6_18_g1356( \2687 , \2683 , \2686 );
and mul_6_18_g1357( \2688 , \2681 , \2686 );
or mul_6_18_g1358( \2689 , \2684 , \2687 , \2688 );
and mul_6_18_g1359( \2690 , \1384 , \1336 );
and mul_6_18_g1360( \2691 , \1342 , \1333 );
nor mul_6_18_g1361( \2692 , \2690 , \2691 );
xnor mul_6_18_g1362( \2693 , \2692 , \1332 );
and mul_6_18_g1363( \2694 , \1477 , \1444 );
and mul_6_18_g1364( \2695 , \1454 , \1442 );
nor mul_6_18_g1365( \2696 , \2694 , \2695 );
xnor mul_6_18_g1366( \2697 , \2696 , \1451 );
and mul_6_18_g1367( \2698 , \2693 , \2697 );
and mul_6_18_g1368( \2699 , \1368 , \1349 );
and mul_6_18_g1369( \2700 , \1470 , \1347 );
nor mul_6_18_g1370( \2701 , \2699 , \2700 );
xnor mul_6_18_g1371( \2702 , \2701 , \1356 );
and mul_6_18_g1372( \2703 , \2697 , \2702 );
and mul_6_18_g1373( \2704 , \2693 , \2702 );
or mul_6_18_g1374( \2705 , \2698 , \2703 , \2704 );
xor mul_6_18_g1375( \2706 , \2524 , \2528 );
xor mul_6_18_g1376( \2707 , \2706 , \2467 );
and mul_6_18_g1377( \2708 , \2705 , \2707 );
xor mul_6_18_g1378( \2709 , \2536 , \2540 );
xor mul_6_18_g1379( \2710 , \2709 , \2545 );
and mul_6_18_g1380( \2711 , \2707 , \2710 );
and mul_6_18_g1381( \2712 , \2705 , \2710 );
or mul_6_18_g1382( \2713 , \2708 , \2711 , \2712 );
xor mul_6_18_g1383( \2714 , \2674 , \2677 );
and mul_6_18_g1384( \2715 , \1454 , \1431 );
and mul_6_18_g1385( \2716 , \1462 , \1429 );
nor mul_6_18_g1386( \2717 , \2715 , \2716 );
xnor mul_6_18_g1387( \2718 , \2717 , \1438 );
and mul_6_18_g1388( \2719 , \1470 , \1444 );
and mul_6_18_g1389( \2720 , \1477 , \1442 );
nor mul_6_18_g1390( \2721 , \2719 , \2720 );
xnor mul_6_18_g1391( \2722 , \2721 , \1451 );
and mul_6_18_g1392( \2723 , \2718 , \2722 );
and mul_6_18_g1393( \2724 , \2722 , \2675 );
and mul_6_18_g1394( \2725 , \2718 , \2675 );
or mul_6_18_g1395( \2726 , \2723 , \2724 , \2725 );
and mul_6_18_g1396( \2727 , \2714 , \2726 );
and mul_6_18_g1397( \2728 , \1533 , \1675 );
and mul_6_18_g1398( \2729 , \1540 , \1673 );
nor mul_6_18_g1399( \2730 , \2728 , \2729 );
xnor mul_6_18_g1400( \2731 , \2730 , \1681 );
and mul_6_18_g1401( \2732 , \2726 , \2731 );
and mul_6_18_g1402( \2733 , \2714 , \2731 );
or mul_6_18_g1403( \2734 , \2727 , \2732 , \2733 );
xor mul_6_18_g1404( \2735 , \2591 , \2595 );
xor mul_6_18_g1405( \2736 , \2735 , \2600 );
and mul_6_18_g1406( \2737 , \2734 , \2736 );
xor mul_6_18_g1407( \2738 , \2553 , \2557 );
xor mul_6_18_g1408( \2739 , \2738 , \2562 );
and mul_6_18_g1409( \2740 , \2736 , \2739 );
and mul_6_18_g1410( \2741 , \2734 , \2739 );
or mul_6_18_g1411( \2742 , \2737 , \2740 , \2741 );
and mul_6_18_g1412( \2743 , \2713 , \2742 );
xor mul_6_18_g1413( \2744 , \2532 , \2548 );
xor mul_6_18_g1414( \2745 , \2744 , \2565 );
and mul_6_18_g1415( \2746 , \2742 , \2745 );
and mul_6_18_g1416( \2747 , \2713 , \2745 );
or mul_6_18_g1417( \2748 , \2743 , \2746 , \2747 );
and mul_6_18_g1418( \2749 , \2689 , \2748 );
xor mul_6_18_g1419( \2750 , \2568 , \2581 );
xor mul_6_18_g1420( \2751 , \2750 , \2584 );
and mul_6_18_g1421( \2752 , \2748 , \2751 );
and mul_6_18_g1422( \2753 , \2689 , \2751 );
or mul_6_18_g1423( \2754 , \2749 , \2752 , \2753 );
xor mul_6_18_g1424( \2755 , \2494 , \2496 );
xor mul_6_18_g1425( \2756 , \2755 , \2499 );
and mul_6_18_g1426( \2757 , \2754 , \2756 );
xor mul_6_18_g1427( \2758 , \2587 , \2619 );
xor mul_6_18_g1428( \2759 , \2758 , \2622 );
and mul_6_18_g1429( \2760 , \2756 , \2759 );
and mul_6_18_g1430( \2761 , \2754 , \2759 );
or mul_6_18_g1431( \2762 , \2757 , \2760 , \2761 );
and mul_6_18_g1432( \2763 , \2637 , \2762 );
xor mul_6_18_g1433( \2764 , \2637 , \2762 );
xor mul_6_18_g1434( \2765 , \2754 , \2756 );
xor mul_6_18_g1435( \2766 , \2765 , \2759 );
and mul_6_18_g1436( \2767 , \1376 , \1336 );
and mul_6_18_g1437( \2768 , \1384 , \1333 );
nor mul_6_18_g1438( \2769 , \2767 , \2768 );
xnor mul_6_18_g1439( \2770 , \2769 , \1332 );
and mul_6_18_g1440( \2771 , \1391 , \1382 );
and mul_6_18_g1441( \2772 , \1399 , \1380 );
nor mul_6_18_g1442( \2773 , \2771 , \2772 );
xnor mul_6_18_g1443( \2774 , \2773 , \1389 );
and mul_6_18_g1444( \2775 , \2770 , \2774 );
and mul_6_18_g1445( \2776 , \1586 , \1460 );
and mul_6_18_g1446( \2777 , \1616 , \1458 );
nor mul_6_18_g1447( \2778 , \2776 , \2777 );
xnor mul_6_18_g1448( \2779 , \2778 , \1467 );
and mul_6_18_g1449( \2780 , \2774 , \2779 );
and mul_6_18_g1450( \2781 , \2770 , \2779 );
or mul_6_18_g1451( \2782 , \2775 , \2780 , \2781 );
and mul_6_18_g1452( \2783 , \1359 , \1349 );
and mul_6_18_g1453( \2784 , \1368 , \1347 );
nor mul_6_18_g1454( \2785 , \2783 , \2784 );
xnor mul_6_18_g1455( \2786 , \2785 , \1356 );
and mul_6_18_g1456( \2787 , \1526 , \1366 );
and mul_6_18_g1457( \2788 , \1622 , \1364 );
nor mul_6_18_g1458( \2789 , \2787 , \2788 );
xnor mul_6_18_g1459( \2790 , \2789 , \1373 );
and mul_6_18_g1460( \2791 , \2786 , \2790 );
and mul_6_18_g1461( \2792 , \1540 , \1397 );
and mul_6_18_g1462( \2793 , \1517 , \1395 );
nor mul_6_18_g1463( \2794 , \2792 , \2793 );
xnor mul_6_18_g1464( \2795 , \2794 , \1404 );
and mul_6_18_g1465( \2796 , \2790 , \2795 );
and mul_6_18_g1466( \2797 , \2786 , \2795 );
or mul_6_18_g1467( \2798 , \2791 , \2796 , \2797 );
and mul_6_18_g1468( \2799 , \2782 , \2798 );
xor mul_6_18_g1469( \2800 , \2641 , \2645 );
xor mul_6_18_g1470( \2801 , \2800 , \2650 );
and mul_6_18_g1471( \2802 , \2798 , \2801 );
and mul_6_18_g1472( \2803 , \2782 , \2801 );
or mul_6_18_g1473( \2804 , \2799 , \2802 , \2803 );
and mul_6_18_g1474( \2805 , \1477 , \1431 );
and mul_6_18_g1475( \2806 , \1454 , \1429 );
nor mul_6_18_g1476( \2807 , \2805 , \2806 );
xnor mul_6_18_g1477( \2808 , \2807 , \1438 );
and mul_6_18_g1478( \2809 , \1498 , \1673 );
not mul_6_18_g1479( \2810 , \2809 );
and mul_6_18_g1480( \2811 , \2810 , \1681 );
and mul_6_18_g1481( \2812 , \2808 , \2811 );
and mul_6_18_g1482( \2813 , \1407 , \1475 );
and mul_6_18_g1483( \2814 , \1416 , \1473 );
nor mul_6_18_g1484( \2815 , \2813 , \2814 );
xnor mul_6_18_g1485( \2816 , \2815 , \1482 );
and mul_6_18_g1486( \2817 , \2812 , \2816 );
and mul_6_18_g1487( \2818 , \1553 , \1675 );
and mul_6_18_g1488( \2819 , \1533 , \1673 );
nor mul_6_18_g1489( \2820 , \2818 , \2819 );
xnor mul_6_18_g1490( \2821 , \2820 , \1681 );
and mul_6_18_g1491( \2822 , \2816 , \2821 );
and mul_6_18_g1492( \2823 , \2812 , \2821 );
or mul_6_18_g1493( \2824 , \2817 , \2822 , \2823 );
xor mul_6_18_g1494( \2825 , \2693 , \2697 );
xor mul_6_18_g1495( \2826 , \2825 , \2702 );
and mul_6_18_g1496( \2827 , \2824 , \2826 );
xor mul_6_18_g1497( \2828 , \2657 , \2661 );
xor mul_6_18_g1498( \2829 , \2828 , \2666 );
and mul_6_18_g1499( \2830 , \2826 , \2829 );
and mul_6_18_g1500( \2831 , \2824 , \2829 );
or mul_6_18_g1501( \2832 , \2827 , \2830 , \2831 );
and mul_6_18_g1502( \2833 , \2804 , \2832 );
xor mul_6_18_g1503( \2834 , \2653 , \2669 );
xor mul_6_18_g1504( \2835 , \2834 , \2678 );
and mul_6_18_g1505( \2836 , \2832 , \2835 );
and mul_6_18_g1506( \2837 , \2804 , \2835 );
or mul_6_18_g1507( \2838 , \2833 , \2836 , \2837 );
xor mul_6_18_g1508( \2839 , \2603 , \2605 );
xor mul_6_18_g1509( \2840 , \2839 , \2608 );
and mul_6_18_g1510( \2841 , \2838 , \2840 );
xor mul_6_18_g1511( \2842 , \2681 , \2683 );
xor mul_6_18_g1512( \2843 , \2842 , \2686 );
and mul_6_18_g1513( \2844 , \2840 , \2843 );
and mul_6_18_g1514( \2845 , \2838 , \2843 );
or mul_6_18_g1515( \2846 , \2841 , \2844 , \2845 );
xor mul_6_18_g1516( \2847 , \2611 , \2613 );
xor mul_6_18_g1517( \2848 , \2847 , \2616 );
and mul_6_18_g1518( \2849 , \2846 , \2848 );
xor mul_6_18_g1519( \2850 , \2689 , \2748 );
xor mul_6_18_g1520( \2851 , \2850 , \2751 );
and mul_6_18_g1521( \2852 , \2848 , \2851 );
and mul_6_18_g1522( \2853 , \2846 , \2851 );
or mul_6_18_g1523( \2854 , \2849 , \2852 , \2853 );
and mul_6_18_g1524( \2855 , \2766 , \2854 );
xor mul_6_18_g1525( \2856 , \2766 , \2854 );
xor mul_6_18_g1526( \2857 , \2846 , \2848 );
xor mul_6_18_g1527( \2858 , \2857 , \2851 );
and mul_6_18_g1528( \2859 , \1462 , \1336 );
and mul_6_18_g1529( \2860 , \1376 , \1333 );
nor mul_6_18_g1530( \2861 , \2859 , \2860 );
xnor mul_6_18_g1531( \2862 , \2861 , \1332 );
and mul_6_18_g1532( \2863 , \1616 , \1382 );
and mul_6_18_g1533( \2864 , \1391 , \1380 );
nor mul_6_18_g1534( \2865 , \2863 , \2864 );
xnor mul_6_18_g1535( \2866 , \2865 , \1389 );
and mul_6_18_g1536( \2867 , \2862 , \2866 );
and mul_6_18_g1537( \2868 , \1533 , \1397 );
and mul_6_18_g1538( \2869 , \1540 , \1395 );
nor mul_6_18_g1539( \2870 , \2868 , \2869 );
xnor mul_6_18_g1540( \2871 , \2870 , \1404 );
and mul_6_18_g1541( \2872 , \2866 , \2871 );
and mul_6_18_g1542( \2873 , \2862 , \2871 );
or mul_6_18_g1543( \2874 , \2867 , \2872 , \2873 );
and mul_6_18_g1544( \2875 , \1368 , \1444 );
and mul_6_18_g1545( \2876 , \1470 , \1442 );
nor mul_6_18_g1546( \2877 , \2875 , \2876 );
xnor mul_6_18_g1547( \2878 , \2877 , \1451 );
and mul_6_18_g1548( \2879 , \1399 , \1349 );
and mul_6_18_g1549( \2880 , \1359 , \1347 );
nor mul_6_18_g1550( \2881 , \2879 , \2880 );
xnor mul_6_18_g1551( \2882 , \2881 , \1356 );
and mul_6_18_g1552( \2883 , \2878 , \2882 );
and mul_6_18_g1553( \2884 , \1517 , \1366 );
and mul_6_18_g1554( \2885 , \1526 , \1364 );
nor mul_6_18_g1555( \2886 , \2884 , \2885 );
xnor mul_6_18_g1556( \2887 , \2886 , \1373 );
and mul_6_18_g1557( \2888 , \2882 , \2887 );
and mul_6_18_g1558( \2889 , \2878 , \2887 );
or mul_6_18_g1559( \2890 , \2883 , \2888 , \2889 );
and mul_6_18_g1560( \2891 , \2874 , \2890 );
xor mul_6_18_g1561( \2892 , \2718 , \2722 );
xor mul_6_18_g1562( \2893 , \2892 , \2675 );
and mul_6_18_g1563( \2894 , \2890 , \2893 );
and mul_6_18_g1564( \2895 , \2874 , \2893 );
or mul_6_18_g1565( \2896 , \2891 , \2894 , \2895 );
xor mul_6_18_g1566( \2897 , \2714 , \2726 );
xor mul_6_18_g1567( \2898 , \2897 , \2731 );
and mul_6_18_g1568( \2899 , \2896 , \2898 );
xor mul_6_18_g1569( \2900 , \2782 , \2798 );
xor mul_6_18_g1570( \2901 , \2900 , \2801 );
and mul_6_18_g1571( \2902 , \2898 , \2901 );
and mul_6_18_g1572( \2903 , \2896 , \2901 );
or mul_6_18_g1573( \2904 , \2899 , \2902 , \2903 );
xor mul_6_18_g1574( \2905 , \2705 , \2707 );
xor mul_6_18_g1575( \2906 , \2905 , \2710 );
and mul_6_18_g1576( \2907 , \2904 , \2906 );
xor mul_6_18_g1577( \2908 , \2734 , \2736 );
xor mul_6_18_g1578( \2909 , \2908 , \2739 );
and mul_6_18_g1579( \2910 , \2906 , \2909 );
and mul_6_18_g1580( \2911 , \2904 , \2909 );
or mul_6_18_g1581( \2912 , \2907 , \2910 , \2911 );
xor mul_6_18_g1582( \2913 , \2713 , \2742 );
xor mul_6_18_g1583( \2914 , \2913 , \2745 );
and mul_6_18_g1584( \2915 , \2912 , \2914 );
xor mul_6_18_g1585( \2916 , \2838 , \2840 );
xor mul_6_18_g1586( \2917 , \2916 , \2843 );
and mul_6_18_g1587( \2918 , \2914 , \2917 );
and mul_6_18_g1588( \2919 , \2912 , \2917 );
or mul_6_18_g1589( \2920 , \2915 , \2918 , \2919 );
and mul_6_18_g1590( \2921 , \2858 , \2920 );
xor mul_6_18_g1591( \2922 , \2858 , \2920 );
xor mul_6_18_g1592( \2923 , \2808 , \2811 );
and mul_6_18_g1593( \2924 , \1416 , \1460 );
and mul_6_18_g1594( \2925 , \1586 , \1458 );
nor mul_6_18_g1595( \2926 , \2924 , \2925 );
xnor mul_6_18_g1596( \2927 , \2926 , \1467 );
and mul_6_18_g1597( \2928 , \2923 , \2927 );
and mul_6_18_g1598( \2929 , \1622 , \1475 );
and mul_6_18_g1599( \2930 , \1407 , \1473 );
nor mul_6_18_g1600( \2931 , \2929 , \2930 );
xnor mul_6_18_g1601( \2932 , \2931 , \1482 );
and mul_6_18_g1602( \2933 , \2927 , \2932 );
and mul_6_18_g1603( \2934 , \2923 , \2932 );
or mul_6_18_g1604( \2935 , \2928 , \2933 , \2934 );
xor mul_6_18_g1605( \2936 , \2770 , \2774 );
xor mul_6_18_g1606( \2937 , \2936 , \2779 );
and mul_6_18_g1607( \2938 , \2935 , \2937 );
xor mul_6_18_g1608( \2939 , \2786 , \2790 );
xor mul_6_18_g1609( \2940 , \2939 , \2795 );
and mul_6_18_g1610( \2941 , \2937 , \2940 );
and mul_6_18_g1611( \2942 , \2935 , \2940 );
or mul_6_18_g1612( \2943 , \2938 , \2941 , \2942 );
and mul_6_18_g1613( \2944 , \1470 , \1431 );
and mul_6_18_g1614( \2945 , \1477 , \1429 );
nor mul_6_18_g1615( \2946 , \2944 , \2945 );
xnor mul_6_18_g1616( \2947 , \2946 , \1438 );
and mul_6_18_g1617( \2948 , \1359 , \1444 );
and mul_6_18_g1618( \2949 , \1368 , \1442 );
nor mul_6_18_g1619( \2950 , \2948 , \2949 );
xnor mul_6_18_g1620( \2951 , \2950 , \1451 );
and mul_6_18_g1621( \2952 , \2947 , \2951 );
and mul_6_18_g1622( \2953 , \2951 , \2809 );
and mul_6_18_g1623( \2954 , \2947 , \2809 );
or mul_6_18_g1624( \2955 , \2952 , \2953 , \2954 );
and mul_6_18_g1625( \2956 , \1391 , \1349 );
and mul_6_18_g1626( \2957 , \1399 , \1347 );
nor mul_6_18_g1627( \2958 , \2956 , \2957 );
xnor mul_6_18_g1628( \2959 , \2958 , \1356 );
and mul_6_18_g1629( \2960 , \1540 , \1366 );
and mul_6_18_g1630( \2961 , \1517 , \1364 );
nor mul_6_18_g1631( \2962 , \2960 , \2961 );
xnor mul_6_18_g1632( \2963 , \2962 , \1373 );
and mul_6_18_g1633( \2964 , \2959 , \2963 );
and mul_6_18_g1634( \2965 , \1553 , \1397 );
and mul_6_18_g1635( \2966 , \1533 , \1395 );
nor mul_6_18_g1636( \2967 , \2965 , \2966 );
xnor mul_6_18_g1637( \2968 , \2967 , \1404 );
and mul_6_18_g1638( \2969 , \2963 , \2968 );
and mul_6_18_g1639( \2970 , \2959 , \2968 );
or mul_6_18_g1640( \2971 , \2964 , \2969 , \2970 );
and mul_6_18_g1641( \2972 , \2955 , \2971 );
and mul_6_18_g1642( \2973 , \1498 , \1675 );
and mul_6_18_g1643( \2974 , \1553 , \1673 );
nor mul_6_18_g1644( \2975 , \2973 , \2974 );
xnor mul_6_18_g1645( \2976 , \2975 , \1681 );
and mul_6_18_g1646( \2977 , \2971 , \2976 );
and mul_6_18_g1647( \2978 , \2955 , \2976 );
or mul_6_18_g1648( \2979 , \2972 , \2977 , \2978 );
xor mul_6_18_g1649( \2980 , \2812 , \2816 );
xor mul_6_18_g1650( \2981 , \2980 , \2821 );
and mul_6_18_g1651( \2982 , \2979 , \2981 );
xor mul_6_18_g1652( \2983 , \2874 , \2890 );
xor mul_6_18_g1653( \2984 , \2983 , \2893 );
and mul_6_18_g1654( \2985 , \2981 , \2984 );
and mul_6_18_g1655( \2986 , \2979 , \2984 );
or mul_6_18_g1656( \2987 , \2982 , \2985 , \2986 );
and mul_6_18_g1657( \2988 , \2943 , \2987 );
xor mul_6_18_g1658( \2989 , \2824 , \2826 );
xor mul_6_18_g1659( \2990 , \2989 , \2829 );
and mul_6_18_g1660( \2991 , \2987 , \2990 );
and mul_6_18_g1661( \2992 , \2943 , \2990 );
or mul_6_18_g1662( \2993 , \2988 , \2991 , \2992 );
xor mul_6_18_g1663( \2994 , \2804 , \2832 );
xor mul_6_18_g1664( \2995 , \2994 , \2835 );
and mul_6_18_g1665( \2996 , \2993 , \2995 );
xor mul_6_18_g1666( \2997 , \2904 , \2906 );
xor mul_6_18_g1667( \2998 , \2997 , \2909 );
and mul_6_18_g1668( \2999 , \2995 , \2998 );
and mul_6_18_g1669( \3000 , \2993 , \2998 );
or mul_6_18_g1670( \3001 , \2996 , \2999 , \3000 );
xor mul_6_18_g1671( \3002 , \2912 , \2914 );
xor mul_6_18_g1672( \3003 , \3002 , \2917 );
and mul_6_18_g1673( \3004 , \3001 , \3003 );
xor mul_6_18_g1674( \3005 , \3001 , \3003 );
xor mul_6_18_g1675( \3006 , \2993 , \2995 );
xor mul_6_18_g1676( \3007 , \3006 , \2998 );
and mul_6_18_g1677( \3008 , \1454 , \1336 );
and mul_6_18_g1678( \3009 , \1462 , \1333 );
nor mul_6_18_g1679( \3010 , \3008 , \3009 );
xnor mul_6_18_g1680( \3011 , \3010 , \1332 );
and mul_6_18_g1681( \3012 , \1586 , \1382 );
and mul_6_18_g1682( \3013 , \1616 , \1380 );
nor mul_6_18_g1683( \3014 , \3012 , \3013 );
xnor mul_6_18_g1684( \3015 , \3014 , \1389 );
and mul_6_18_g1685( \3016 , \3011 , \3015 );
and mul_6_18_g1686( \3017 , \1407 , \1460 );
and mul_6_18_g1687( \3018 , \1416 , \1458 );
nor mul_6_18_g1688( \3019 , \3017 , \3018 );
xnor mul_6_18_g1689( \3020 , \3019 , \1467 );
and mul_6_18_g1690( \3021 , \3015 , \3020 );
and mul_6_18_g1691( \3022 , \3011 , \3020 );
or mul_6_18_g1692( \3023 , \3016 , \3021 , \3022 );
xor mul_6_18_g1693( \3024 , \2862 , \2866 );
xor mul_6_18_g1694( \3025 , \3024 , \2871 );
and mul_6_18_g1695( \3026 , \3023 , \3025 );
xor mul_6_18_g1696( \3027 , \2878 , \2882 );
xor mul_6_18_g1697( \3028 , \3027 , \2887 );
and mul_6_18_g1698( \3029 , \3025 , \3028 );
and mul_6_18_g1699( \3030 , \3023 , \3028 );
or mul_6_18_g1700( \3031 , \3026 , \3029 , \3030 );
and mul_6_18_g1701( \3032 , \1368 , \1431 );
and mul_6_18_g1702( \3033 , \1470 , \1429 );
nor mul_6_18_g1703( \3034 , \3032 , \3033 );
xnor mul_6_18_g1704( \3035 , \3034 , \1438 );
and mul_6_18_g1705( \3036 , \1498 , \1395 );
not mul_6_18_g1706( \3037 , \3036 );
and mul_6_18_g1707( \3038 , \3037 , \1404 );
and mul_6_18_g1708( \3039 , \3035 , \3038 );
and mul_6_18_g1709( \3040 , \1526 , \1475 );
and mul_6_18_g1710( \3041 , \1622 , \1473 );
nor mul_6_18_g1711( \3042 , \3040 , \3041 );
xnor mul_6_18_g1712( \3043 , \3042 , \1482 );
and mul_6_18_g1713( \3044 , \3039 , \3043 );
xor mul_6_18_g1714( \3045 , \2947 , \2951 );
xor mul_6_18_g1715( \3046 , \3045 , \2809 );
and mul_6_18_g1716( \3047 , \3043 , \3046 );
and mul_6_18_g1717( \3048 , \3039 , \3046 );
or mul_6_18_g1718( \3049 , \3044 , \3047 , \3048 );
xor mul_6_18_g1719( \3050 , \2955 , \2971 );
xor mul_6_18_g1720( \3051 , \3050 , \2976 );
and mul_6_18_g1721( \3052 , \3049 , \3051 );
xor mul_6_18_g1722( \3053 , \2923 , \2927 );
xor mul_6_18_g1723( \3054 , \3053 , \2932 );
and mul_6_18_g1724( \3055 , \3051 , \3054 );
and mul_6_18_g1725( \3056 , \3049 , \3054 );
or mul_6_18_g1726( \3057 , \3052 , \3055 , \3056 );
and mul_6_18_g1727( \3058 , \3031 , \3057 );
xor mul_6_18_g1728( \3059 , \2935 , \2937 );
xor mul_6_18_g1729( \3060 , \3059 , \2940 );
and mul_6_18_g1730( \3061 , \3057 , \3060 );
and mul_6_18_g1731( \3062 , \3031 , \3060 );
or mul_6_18_g1732( \3063 , \3058 , \3061 , \3062 );
xor mul_6_18_g1733( \3064 , \2896 , \2898 );
xor mul_6_18_g1734( \3065 , \3064 , \2901 );
and mul_6_18_g1735( \3066 , \3063 , \3065 );
xor mul_6_18_g1736( \3067 , \2943 , \2987 );
xor mul_6_18_g1737( \3068 , \3067 , \2990 );
and mul_6_18_g1738( \3069 , \3065 , \3068 );
and mul_6_18_g1739( \3070 , \3063 , \3068 );
or mul_6_18_g1740( \3071 , \3066 , \3069 , \3070 );
and mul_6_18_g1741( \3072 , \3007 , \3071 );
xor mul_6_18_g1742( \3073 , \3007 , \3071 );
xor mul_6_18_g1743( \3074 , \3063 , \3065 );
xor mul_6_18_g1744( \3075 , \3074 , \3068 );
and mul_6_18_g1745( \3076 , \1477 , \1336 );
and mul_6_18_g1746( \3077 , \1454 , \1333 );
nor mul_6_18_g1747( \3078 , \3076 , \3077 );
xnor mul_6_18_g1748( \3079 , \3078 , \1332 );
and mul_6_18_g1749( \3080 , \1416 , \1382 );
and mul_6_18_g1750( \3081 , \1586 , \1380 );
nor mul_6_18_g1751( \3082 , \3080 , \3081 );
xnor mul_6_18_g1752( \3083 , \3082 , \1389 );
and mul_6_18_g1753( \3084 , \3079 , \3083 );
and mul_6_18_g1754( \3085 , \1498 , \1397 );
and mul_6_18_g1755( \3086 , \1553 , \1395 );
nor mul_6_18_g1756( \3087 , \3085 , \3086 );
xnor mul_6_18_g1757( \3088 , \3087 , \1404 );
and mul_6_18_g1758( \3089 , \3083 , \3088 );
and mul_6_18_g1759( \3090 , \3079 , \3088 );
or mul_6_18_g1760( \3091 , \3084 , \3089 , \3090 );
and mul_6_18_g1761( \3092 , \1399 , \1444 );
and mul_6_18_g1762( \3093 , \1359 , \1442 );
nor mul_6_18_g1763( \3094 , \3092 , \3093 );
xnor mul_6_18_g1764( \3095 , \3094 , \1451 );
and mul_6_18_g1765( \3096 , \1616 , \1349 );
and mul_6_18_g1766( \3097 , \1391 , \1347 );
nor mul_6_18_g1767( \3098 , \3096 , \3097 );
xnor mul_6_18_g1768( \3099 , \3098 , \1356 );
and mul_6_18_g1769( \3100 , \3095 , \3099 );
and mul_6_18_g1770( \3101 , \1533 , \1366 );
and mul_6_18_g1771( \3102 , \1540 , \1364 );
nor mul_6_18_g1772( \3103 , \3101 , \3102 );
xnor mul_6_18_g1773( \3104 , \3103 , \1373 );
and mul_6_18_g1774( \3105 , \3099 , \3104 );
and mul_6_18_g1775( \3106 , \3095 , \3104 );
or mul_6_18_g1776( \3107 , \3100 , \3105 , \3106 );
and mul_6_18_g1777( \3108 , \3091 , \3107 );
xor mul_6_18_g1778( \3109 , \3035 , \3038 );
and mul_6_18_g1779( \3110 , \1622 , \1460 );
and mul_6_18_g1780( \3111 , \1407 , \1458 );
nor mul_6_18_g1781( \3112 , \3110 , \3111 );
xnor mul_6_18_g1782( \3113 , \3112 , \1467 );
and mul_6_18_g1783( \3114 , \3109 , \3113 );
and mul_6_18_g1784( \3115 , \1517 , \1475 );
and mul_6_18_g1785( \3116 , \1526 , \1473 );
nor mul_6_18_g1786( \3117 , \3115 , \3116 );
xnor mul_6_18_g1787( \3118 , \3117 , \1482 );
and mul_6_18_g1788( \3119 , \3113 , \3118 );
and mul_6_18_g1789( \3120 , \3109 , \3118 );
or mul_6_18_g1790( \3121 , \3114 , \3119 , \3120 );
and mul_6_18_g1791( \3122 , \3107 , \3121 );
and mul_6_18_g1792( \3123 , \3091 , \3121 );
or mul_6_18_g1793( \3124 , \3108 , \3122 , \3123 );
and mul_6_18_g1794( \3125 , \1407 , \1382 );
and mul_6_18_g1795( \3126 , \1416 , \1380 );
nor mul_6_18_g1796( \3127 , \3125 , \3126 );
xnor mul_6_18_g1797( \3128 , \3127 , \1389 );
and mul_6_18_g1798( \3129 , \1526 , \1460 );
and mul_6_18_g1799( \3130 , \1622 , \1458 );
nor mul_6_18_g1800( \3131 , \3129 , \3130 );
xnor mul_6_18_g1801( \3132 , \3131 , \1467 );
and mul_6_18_g1802( \3133 , \3128 , \3132 );
and mul_6_18_g1803( \3134 , \1540 , \1475 );
and mul_6_18_g1804( \3135 , \1517 , \1473 );
nor mul_6_18_g1805( \3136 , \3134 , \3135 );
xnor mul_6_18_g1806( \3137 , \3136 , \1482 );
and mul_6_18_g1807( \3138 , \3132 , \3137 );
and mul_6_18_g1808( \3139 , \3128 , \3137 );
or mul_6_18_g1809( \3140 , \3133 , \3138 , \3139 );
and mul_6_18_g1810( \3141 , \1470 , \1336 );
and mul_6_18_g1811( \3142 , \1477 , \1333 );
nor mul_6_18_g1812( \3143 , \3141 , \3142 );
xnor mul_6_18_g1813( \3144 , \3143 , \1332 );
and mul_6_18_g1814( \3145 , \1586 , \1349 );
and mul_6_18_g1815( \3146 , \1616 , \1347 );
nor mul_6_18_g1816( \3147 , \3145 , \3146 );
xnor mul_6_18_g1817( \3148 , \3147 , \1356 );
and mul_6_18_g1818( \3149 , \3144 , \3148 );
and mul_6_18_g1819( \3150 , \1553 , \1366 );
and mul_6_18_g1820( \3151 , \1533 , \1364 );
nor mul_6_18_g1821( \3152 , \3150 , \3151 );
xnor mul_6_18_g1822( \3153 , \3152 , \1373 );
and mul_6_18_g1823( \3154 , \3148 , \3153 );
and mul_6_18_g1824( \3155 , \3144 , \3153 );
or mul_6_18_g1825( \3156 , \3149 , \3154 , \3155 );
and mul_6_18_g1826( \3157 , \3140 , \3156 );
and mul_6_18_g1827( \3158 , \1359 , \1431 );
and mul_6_18_g1828( \3159 , \1368 , \1429 );
nor mul_6_18_g1829( \3160 , \3158 , \3159 );
xnor mul_6_18_g1830( \3161 , \3160 , \1438 );
and mul_6_18_g1831( \3162 , \1391 , \1444 );
and mul_6_18_g1832( \3163 , \1399 , \1442 );
nor mul_6_18_g1833( \3164 , \3162 , \3163 );
xnor mul_6_18_g1834( \3165 , \3164 , \1451 );
and mul_6_18_g1835( \3166 , \3161 , \3165 );
and mul_6_18_g1836( \3167 , \3165 , \3036 );
and mul_6_18_g1837( \3168 , \3161 , \3036 );
or mul_6_18_g1838( \3169 , \3166 , \3167 , \3168 );
and mul_6_18_g1839( \3170 , \3156 , \3169 );
and mul_6_18_g1840( \3171 , \3140 , \3169 );
or mul_6_18_g1841( \3172 , \3157 , \3170 , \3171 );
xor mul_6_18_g1842( \3173 , \3011 , \3015 );
xor mul_6_18_g1843( \3174 , \3173 , \3020 );
and mul_6_18_g1844( \3175 , \3172 , \3174 );
xor mul_6_18_g1845( \3176 , \2959 , \2963 );
xor mul_6_18_g1846( \3177 , \3176 , \2968 );
and mul_6_18_g1847( \3178 , \3174 , \3177 );
and mul_6_18_g1848( \3179 , \3172 , \3177 );
or mul_6_18_g1849( \3180 , \3175 , \3178 , \3179 );
and mul_6_18_g1850( \3181 , \3124 , \3180 );
xor mul_6_18_g1851( \3182 , \3023 , \3025 );
xor mul_6_18_g1852( \3183 , \3182 , \3028 );
and mul_6_18_g1853( \3184 , \3180 , \3183 );
and mul_6_18_g1854( \3185 , \3124 , \3183 );
or mul_6_18_g1855( \3186 , \3181 , \3184 , \3185 );
xor mul_6_18_g1856( \3187 , \2979 , \2981 );
xor mul_6_18_g1857( \3188 , \3187 , \2984 );
and mul_6_18_g1858( \3189 , \3186 , \3188 );
xor mul_6_18_g1859( \3190 , \3031 , \3057 );
xor mul_6_18_g1860( \3191 , \3190 , \3060 );
and mul_6_18_g1861( \3192 , \3188 , \3191 );
and mul_6_18_g1862( \3193 , \3186 , \3191 );
or mul_6_18_g1863( \3194 , \3189 , \3192 , \3193 );
and mul_6_18_g1864( \3195 , \3075 , \3194 );
xor mul_6_18_g1865( \3196 , \3075 , \3194 );
xor mul_6_18_g1866( \3197 , \3186 , \3188 );
xor mul_6_18_g1867( \3198 , \3197 , \3191 );
xor mul_6_18_g1868( \3199 , \3079 , \3083 );
xor mul_6_18_g1869( \3200 , \3199 , \3088 );
xor mul_6_18_g1870( \3201 , \3095 , \3099 );
xor mul_6_18_g1871( \3202 , \3201 , \3104 );
and mul_6_18_g1872( \3203 , \3200 , \3202 );
xor mul_6_18_g1873( \3204 , \3109 , \3113 );
xor mul_6_18_g1874( \3205 , \3204 , \3118 );
and mul_6_18_g1875( \3206 , \3202 , \3205 );
and mul_6_18_g1876( \3207 , \3200 , \3205 );
or mul_6_18_g1877( \3208 , \3203 , \3206 , \3207 );
xor mul_6_18_g1878( \3209 , \3091 , \3107 );
xor mul_6_18_g1879( \3210 , \3209 , \3121 );
and mul_6_18_g1880( \3211 , \3208 , \3210 );
xor mul_6_18_g1881( \3212 , \3039 , \3043 );
xor mul_6_18_g1882( \3213 , \3212 , \3046 );
and mul_6_18_g1883( \3214 , \3210 , \3213 );
and mul_6_18_g1884( \3215 , \3208 , \3213 );
or mul_6_18_g1885( \3216 , \3211 , \3214 , \3215 );
xor mul_6_18_g1886( \3217 , \3049 , \3051 );
xor mul_6_18_g1887( \3218 , \3217 , \3054 );
and mul_6_18_g1888( \3219 , \3216 , \3218 );
xor mul_6_18_g1889( \3220 , \3124 , \3180 );
xor mul_6_18_g1890( \3221 , \3220 , \3183 );
and mul_6_18_g1891( \3222 , \3218 , \3221 );
and mul_6_18_g1892( \3223 , \3216 , \3221 );
or mul_6_18_g1893( \3224 , \3219 , \3222 , \3223 );
and mul_6_18_g1894( \3225 , \3198 , \3224 );
xor mul_6_18_g1895( \3226 , \3198 , \3224 );
xor mul_6_18_g1896( \3227 , \3216 , \3218 );
xor mul_6_18_g1897( \3228 , \3227 , \3221 );
and mul_6_18_g1898( \3229 , \1416 , \1349 );
and mul_6_18_g1899( \3230 , \1586 , \1347 );
nor mul_6_18_g1900( \3231 , \3229 , \3230 );
xnor mul_6_18_g1901( \3232 , \3231 , \1356 );
and mul_6_18_g1902( \3233 , \1622 , \1382 );
and mul_6_18_g1903( \3234 , \1407 , \1380 );
nor mul_6_18_g1904( \3235 , \3233 , \3234 );
xnor mul_6_18_g1905( \3236 , \3235 , \1389 );
and mul_6_18_g1906( \3237 , \3232 , \3236 );
and mul_6_18_g1907( \3238 , \1517 , \1460 );
and mul_6_18_g1908( \3239 , \1526 , \1458 );
nor mul_6_18_g1909( \3240 , \3238 , \3239 );
xnor mul_6_18_g1910( \3241 , \3240 , \1467 );
and mul_6_18_g1911( \3242 , \3236 , \3241 );
and mul_6_18_g1912( \3243 , \3232 , \3241 );
or mul_6_18_g1913( \3244 , \3237 , \3242 , \3243 );
xor mul_6_18_g1914( \3245 , \3128 , \3132 );
xor mul_6_18_g1915( \3246 , \3245 , \3137 );
and mul_6_18_g1916( \3247 , \3244 , \3246 );
xor mul_6_18_g1917( \3248 , \3144 , \3148 );
xor mul_6_18_g1918( \3249 , \3248 , \3153 );
and mul_6_18_g1919( \3250 , \3246 , \3249 );
and mul_6_18_g1920( \3251 , \3244 , \3249 );
or mul_6_18_g1921( \3252 , \3247 , \3250 , \3251 );
and mul_6_18_g1922( \3253 , \1368 , \1336 );
and mul_6_18_g1923( \3254 , \1470 , \1333 );
nor mul_6_18_g1924( \3255 , \3253 , \3254 );
xnor mul_6_18_g1925( \3256 , \3255 , \1332 );
and mul_6_18_g1926( \3257 , \1616 , \1444 );
and mul_6_18_g1927( \3258 , \1391 , \1442 );
nor mul_6_18_g1928( \3259 , \3257 , \3258 );
xnor mul_6_18_g1929( \3260 , \3259 , \1451 );
and mul_6_18_g1930( \3261 , \3256 , \3260 );
and mul_6_18_g1931( \3262 , \1498 , \1366 );
and mul_6_18_g1932( \3263 , \1553 , \1364 );
nor mul_6_18_g1933( \3264 , \3262 , \3263 );
xnor mul_6_18_g1934( \3265 , \3264 , \1373 );
and mul_6_18_g1935( \3266 , \3260 , \3265 );
and mul_6_18_g1936( \3267 , \3256 , \3265 );
or mul_6_18_g1937( \3268 , \3261 , \3266 , \3267 );
and mul_6_18_g1938( \3269 , \1399 , \1431 );
and mul_6_18_g1939( \3270 , \1359 , \1429 );
nor mul_6_18_g1940( \3271 , \3269 , \3270 );
xnor mul_6_18_g1941( \3272 , \3271 , \1438 );
and mul_6_18_g1942( \3273 , \1498 , \1364 );
not mul_6_18_g1943( \3274 , \3273 );
and mul_6_18_g1944( \3275 , \3274 , \1373 );
and mul_6_18_g1945( \3276 , \3272 , \3275 );
and mul_6_18_g1946( \3277 , \3268 , \3276 );
xor mul_6_18_g1947( \3278 , \3161 , \3165 );
xor mul_6_18_g1948( \3279 , \3278 , \3036 );
and mul_6_18_g1949( \3280 , \3276 , \3279 );
and mul_6_18_g1950( \3281 , \3268 , \3279 );
or mul_6_18_g1951( \3282 , \3277 , \3280 , \3281 );
and mul_6_18_g1952( \3283 , \3252 , \3282 );
xor mul_6_18_g1953( \3284 , \3140 , \3156 );
xor mul_6_18_g1954( \3285 , \3284 , \3169 );
and mul_6_18_g1955( \3286 , \3282 , \3285 );
and mul_6_18_g1956( \3287 , \3252 , \3285 );
or mul_6_18_g1957( \3288 , \3283 , \3286 , \3287 );
xor mul_6_18_g1958( \3289 , \3172 , \3174 );
xor mul_6_18_g1959( \3290 , \3289 , \3177 );
and mul_6_18_g1960( \3291 , \3288 , \3290 );
xor mul_6_18_g1961( \3292 , \3208 , \3210 );
xor mul_6_18_g1962( \3293 , \3292 , \3213 );
and mul_6_18_g1963( \3294 , \3290 , \3293 );
and mul_6_18_g1964( \3295 , \3288 , \3293 );
or mul_6_18_g1965( \3296 , \3291 , \3294 , \3295 );
and mul_6_18_g1966( \3297 , \3228 , \3296 );
xor mul_6_18_g1967( \3298 , \3228 , \3296 );
xor mul_6_18_g1968( \3299 , \3272 , \3275 );
and mul_6_18_g1969( \3300 , \1391 , \1431 );
and mul_6_18_g1970( \3301 , \1399 , \1429 );
nor mul_6_18_g1971( \3302 , \3300 , \3301 );
xnor mul_6_18_g1972( \3303 , \3302 , \1438 );
and mul_6_18_g1973( \3304 , \1586 , \1444 );
and mul_6_18_g1974( \3305 , \1616 , \1442 );
nor mul_6_18_g1975( \3306 , \3304 , \3305 );
xnor mul_6_18_g1976( \3307 , \3306 , \1451 );
and mul_6_18_g1977( \3308 , \3303 , \3307 );
and mul_6_18_g1978( \3309 , \3307 , \3273 );
and mul_6_18_g1979( \3310 , \3303 , \3273 );
or mul_6_18_g1980( \3311 , \3308 , \3309 , \3310 );
and mul_6_18_g1981( \3312 , \3299 , \3311 );
and mul_6_18_g1982( \3313 , \1533 , \1475 );
and mul_6_18_g1983( \3314 , \1540 , \1473 );
nor mul_6_18_g1984( \3315 , \3313 , \3314 );
xnor mul_6_18_g1985( \3316 , \3315 , \1482 );
and mul_6_18_g1986( \3317 , \3311 , \3316 );
and mul_6_18_g1987( \3318 , \3299 , \3316 );
or mul_6_18_g1988( \3319 , \3312 , \3317 , \3318 );
and mul_6_18_g1989( \3320 , \1359 , \1336 );
and mul_6_18_g1990( \3321 , \1368 , \1333 );
nor mul_6_18_g1991( \3322 , \3320 , \3321 );
xnor mul_6_18_g1992( \3323 , \3322 , \1332 );
and mul_6_18_g1993( \3324 , \1407 , \1349 );
and mul_6_18_g1994( \3325 , \1416 , \1347 );
nor mul_6_18_g1995( \3326 , \3324 , \3325 );
xnor mul_6_18_g1996( \3327 , \3326 , \1356 );
and mul_6_18_g1997( \3328 , \3323 , \3327 );
and mul_6_18_g1998( \3329 , \1526 , \1382 );
and mul_6_18_g1999( \3330 , \1622 , \1380 );
nor mul_6_18_g2000( \3331 , \3329 , \3330 );
xnor mul_6_18_g2001( \3332 , \3331 , \1389 );
and mul_6_18_g2002( \3333 , \3327 , \3332 );
and mul_6_18_g2003( \3334 , \3323 , \3332 );
or mul_6_18_g2004( \3335 , \3328 , \3333 , \3334 );
xor mul_6_18_g2005( \3336 , \3232 , \3236 );
xor mul_6_18_g2006( \3337 , \3336 , \3241 );
and mul_6_18_g2007( \3338 , \3335 , \3337 );
xor mul_6_18_g2008( \3339 , \3256 , \3260 );
xor mul_6_18_g2009( \3340 , \3339 , \3265 );
and mul_6_18_g2010( \3341 , \3337 , \3340 );
and mul_6_18_g2011( \3342 , \3335 , \3340 );
or mul_6_18_g2012( \3343 , \3338 , \3341 , \3342 );
and mul_6_18_g2013( \3344 , \3319 , \3343 );
xor mul_6_18_g2014( \3345 , \3268 , \3276 );
xor mul_6_18_g2015( \3346 , \3345 , \3279 );
and mul_6_18_g2016( \3347 , \3343 , \3346 );
and mul_6_18_g2017( \3348 , \3319 , \3346 );
or mul_6_18_g2018( \3349 , \3344 , \3347 , \3348 );
xor mul_6_18_g2019( \3350 , \3200 , \3202 );
xor mul_6_18_g2020( \3351 , \3350 , \3205 );
and mul_6_18_g2021( \3352 , \3349 , \3351 );
xor mul_6_18_g2022( \3353 , \3252 , \3282 );
xor mul_6_18_g2023( \3354 , \3353 , \3285 );
and mul_6_18_g2024( \3355 , \3351 , \3354 );
and mul_6_18_g2025( \3356 , \3349 , \3354 );
or mul_6_18_g2026( \3357 , \3352 , \3355 , \3356 );
xor mul_6_18_g2027( \3358 , \3288 , \3290 );
xor mul_6_18_g2028( \3359 , \3358 , \3293 );
and mul_6_18_g2029( \3360 , \3357 , \3359 );
xor mul_6_18_g2030( \3361 , \3357 , \3359 );
xor mul_6_18_g2031( \3362 , \3349 , \3351 );
xor mul_6_18_g2032( \3363 , \3362 , \3354 );
and mul_6_18_g2033( \3364 , \1616 , \1431 );
and mul_6_18_g2034( \3365 , \1391 , \1429 );
nor mul_6_18_g2035( \3366 , \3364 , \3365 );
xnor mul_6_18_g2036( \3367 , \3366 , \1438 );
and mul_6_18_g2037( \3368 , \1498 , \1473 );
not mul_6_18_g2038( \3369 , \3368 );
and mul_6_18_g2039( \3370 , \3369 , \1482 );
and mul_6_18_g2040( \3371 , \3367 , \3370 );
and mul_6_18_g2041( \3372 , \1540 , \1460 );
and mul_6_18_g2042( \3373 , \1517 , \1458 );
nor mul_6_18_g2043( \3374 , \3372 , \3373 );
xnor mul_6_18_g2044( \3375 , \3374 , \1467 );
and mul_6_18_g2045( \3376 , \3371 , \3375 );
and mul_6_18_g2046( \3377 , \1553 , \1475 );
and mul_6_18_g2047( \3378 , \1533 , \1473 );
nor mul_6_18_g2048( \3379 , \3377 , \3378 );
xnor mul_6_18_g2049( \3380 , \3379 , \1482 );
and mul_6_18_g2050( \3381 , \3375 , \3380 );
and mul_6_18_g2051( \3382 , \3371 , \3380 );
or mul_6_18_g2052( \3383 , \3376 , \3381 , \3382 );
and mul_6_18_g2053( \3384 , \1399 , \1336 );
and mul_6_18_g2054( \3385 , \1359 , \1333 );
nor mul_6_18_g2055( \3386 , \3384 , \3385 );
xnor mul_6_18_g2056( \3387 , \3386 , \1332 );
and mul_6_18_g2057( \3388 , \1416 , \1444 );
and mul_6_18_g2058( \3389 , \1586 , \1442 );
nor mul_6_18_g2059( \3390 , \3388 , \3389 );
xnor mul_6_18_g2060( \3391 , \3390 , \1451 );
and mul_6_18_g2061( \3392 , \3387 , \3391 );
and mul_6_18_g2062( \3393 , \1622 , \1349 );
and mul_6_18_g2063( \3394 , \1407 , \1347 );
nor mul_6_18_g2064( \3395 , \3393 , \3394 );
xnor mul_6_18_g2065( \3396 , \3395 , \1356 );
and mul_6_18_g2066( \3397 , \3391 , \3396 );
and mul_6_18_g2067( \3398 , \3387 , \3396 );
or mul_6_18_g2068( \3399 , \3392 , \3397 , \3398 );
and mul_6_18_g2069( \3400 , \1517 , \1382 );
and mul_6_18_g2070( \3401 , \1526 , \1380 );
nor mul_6_18_g2071( \3402 , \3400 , \3401 );
xnor mul_6_18_g2072( \3403 , \3402 , \1389 );
and mul_6_18_g2073( \3404 , \1533 , \1460 );
and mul_6_18_g2074( \3405 , \1540 , \1458 );
nor mul_6_18_g2075( \3406 , \3404 , \3405 );
xnor mul_6_18_g2076( \3407 , \3406 , \1467 );
and mul_6_18_g2077( \3408 , \3403 , \3407 );
and mul_6_18_g2078( \3409 , \1498 , \1475 );
and mul_6_18_g2079( \3410 , \1553 , \1473 );
nor mul_6_18_g2080( \3411 , \3409 , \3410 );
xnor mul_6_18_g2081( \3412 , \3411 , \1482 );
and mul_6_18_g2082( \3413 , \3407 , \3412 );
and mul_6_18_g2083( \3414 , \3403 , \3412 );
or mul_6_18_g2084( \3415 , \3408 , \3413 , \3414 );
and mul_6_18_g2085( \3416 , \3399 , \3415 );
xor mul_6_18_g2086( \3417 , \3303 , \3307 );
xor mul_6_18_g2087( \3418 , \3417 , \3273 );
and mul_6_18_g2088( \3419 , \3415 , \3418 );
and mul_6_18_g2089( \3420 , \3399 , \3418 );
or mul_6_18_g2090( \3421 , \3416 , \3419 , \3420 );
and mul_6_18_g2091( \3422 , \3383 , \3421 );
xor mul_6_18_g2092( \3423 , \3299 , \3311 );
xor mul_6_18_g2093( \3424 , \3423 , \3316 );
and mul_6_18_g2094( \3425 , \3421 , \3424 );
and mul_6_18_g2095( \3426 , \3383 , \3424 );
or mul_6_18_g2096( \3427 , \3422 , \3425 , \3426 );
xor mul_6_18_g2097( \3428 , \3244 , \3246 );
xor mul_6_18_g2098( \3429 , \3428 , \3249 );
and mul_6_18_g2099( \3430 , \3427 , \3429 );
xor mul_6_18_g2100( \3431 , \3319 , \3343 );
xor mul_6_18_g2101( \3432 , \3431 , \3346 );
and mul_6_18_g2102( \3433 , \3429 , \3432 );
and mul_6_18_g2103( \3434 , \3427 , \3432 );
or mul_6_18_g2104( \3435 , \3430 , \3433 , \3434 );
and mul_6_18_g2105( \3436 , \3363 , \3435 );
xor mul_6_18_g2106( \3437 , \3363 , \3435 );
xor mul_6_18_g2107( \3438 , \3427 , \3429 );
xor mul_6_18_g2108( \3439 , \3438 , \3432 );
xor mul_6_18_g2109( \3440 , \3367 , \3370 );
and mul_6_18_g2110( \3441 , \1586 , \1431 );
and mul_6_18_g2111( \3442 , \1616 , \1429 );
nor mul_6_18_g2112( \3443 , \3441 , \3442 );
xnor mul_6_18_g2113( \3444 , \3443 , \1438 );
and mul_6_18_g2114( \3445 , \1407 , \1444 );
and mul_6_18_g2115( \3446 , \1416 , \1442 );
nor mul_6_18_g2116( \3447 , \3445 , \3446 );
xnor mul_6_18_g2117( \3448 , \3447 , \1451 );
and mul_6_18_g2118( \3449 , \3444 , \3448 );
and mul_6_18_g2119( \3450 , \3448 , \3368 );
and mul_6_18_g2120( \3451 , \3444 , \3368 );
or mul_6_18_g2121( \3452 , \3449 , \3450 , \3451 );
and mul_6_18_g2122( \3453 , \3440 , \3452 );
and mul_6_18_g2123( \3454 , \1391 , \1336 );
and mul_6_18_g2124( \3455 , \1399 , \1333 );
nor mul_6_18_g2125( \3456 , \3454 , \3455 );
xnor mul_6_18_g2126( \3457 , \3456 , \1332 );
and mul_6_18_g2127( \3458 , \1526 , \1349 );
and mul_6_18_g2128( \3459 , \1622 , \1347 );
nor mul_6_18_g2129( \3460 , \3458 , \3459 );
xnor mul_6_18_g2130( \3461 , \3460 , \1356 );
and mul_6_18_g2131( \3462 , \3457 , \3461 );
and mul_6_18_g2132( \3463 , \1540 , \1382 );
and mul_6_18_g2133( \3464 , \1517 , \1380 );
nor mul_6_18_g2134( \3465 , \3463 , \3464 );
xnor mul_6_18_g2135( \3466 , \3465 , \1389 );
and mul_6_18_g2136( \3467 , \3461 , \3466 );
and mul_6_18_g2137( \3468 , \3457 , \3466 );
or mul_6_18_g2138( \3469 , \3462 , \3467 , \3468 );
and mul_6_18_g2139( \3470 , \3452 , \3469 );
and mul_6_18_g2140( \3471 , \3440 , \3469 );
or mul_6_18_g2141( \3472 , \3453 , \3470 , \3471 );
xor mul_6_18_g2142( \3473 , \3323 , \3327 );
xor mul_6_18_g2143( \3474 , \3473 , \3332 );
and mul_6_18_g2144( \3475 , \3472 , \3474 );
xor mul_6_18_g2145( \3476 , \3371 , \3375 );
xor mul_6_18_g2146( \3477 , \3476 , \3380 );
and mul_6_18_g2147( \3478 , \3474 , \3477 );
and mul_6_18_g2148( \3479 , \3472 , \3477 );
or mul_6_18_g2149( \3480 , \3475 , \3478 , \3479 );
xor mul_6_18_g2150( \3481 , \3335 , \3337 );
xor mul_6_18_g2151( \3482 , \3481 , \3340 );
and mul_6_18_g2152( \3483 , \3480 , \3482 );
xor mul_6_18_g2153( \3484 , \3383 , \3421 );
xor mul_6_18_g2154( \3485 , \3484 , \3424 );
and mul_6_18_g2155( \3486 , \3482 , \3485 );
and mul_6_18_g2156( \3487 , \3480 , \3485 );
or mul_6_18_g2157( \3488 , \3483 , \3486 , \3487 );
and mul_6_18_g2158( \3489 , \3439 , \3488 );
xor mul_6_18_g2159( \3490 , \3439 , \3488 );
xor mul_6_18_g2160( \3491 , \3480 , \3482 );
xor mul_6_18_g2161( \3492 , \3491 , \3485 );
and mul_6_18_g2162( \3493 , \1616 , \1336 );
and mul_6_18_g2163( \3494 , \1391 , \1333 );
nor mul_6_18_g2164( \3495 , \3493 , \3494 );
xnor mul_6_18_g2165( \3496 , \3495 , \1332 );
and mul_6_18_g2166( \3497 , \1622 , \1444 );
and mul_6_18_g2167( \3498 , \1407 , \1442 );
nor mul_6_18_g2168( \3499 , \3497 , \3498 );
xnor mul_6_18_g2169( \3500 , \3499 , \1451 );
and mul_6_18_g2170( \3501 , \3496 , \3500 );
and mul_6_18_g2171( \3502 , \1517 , \1349 );
and mul_6_18_g2172( \3503 , \1526 , \1347 );
nor mul_6_18_g2173( \3504 , \3502 , \3503 );
xnor mul_6_18_g2174( \3505 , \3504 , \1356 );
and mul_6_18_g2175( \3506 , \3500 , \3505 );
and mul_6_18_g2176( \3507 , \3496 , \3505 );
or mul_6_18_g2177( \3508 , \3501 , \3506 , \3507 );
and mul_6_18_g2178( \3509 , \1416 , \1431 );
and mul_6_18_g2179( \3510 , \1586 , \1429 );
nor mul_6_18_g2180( \3511 , \3509 , \3510 );
xnor mul_6_18_g2181( \3512 , \3511 , \1438 );
and mul_6_18_g2182( \3513 , \1498 , \1458 );
not mul_6_18_g2183( \3514 , \3513 );
and mul_6_18_g2184( \3515 , \3514 , \1467 );
and mul_6_18_g2185( \3516 , \3512 , \3515 );
and mul_6_18_g2186( \3517 , \3508 , \3516 );
and mul_6_18_g2187( \3518 , \1553 , \1460 );
and mul_6_18_g2188( \3519 , \1533 , \1458 );
nor mul_6_18_g2189( \3520 , \3518 , \3519 );
xnor mul_6_18_g2190( \3521 , \3520 , \1467 );
and mul_6_18_g2191( \3522 , \3516 , \3521 );
and mul_6_18_g2192( \3523 , \3508 , \3521 );
or mul_6_18_g2193( \3524 , \3517 , \3522 , \3523 );
xor mul_6_18_g2194( \3525 , \3387 , \3391 );
xor mul_6_18_g2195( \3526 , \3525 , \3396 );
and mul_6_18_g2196( \3527 , \3524 , \3526 );
xor mul_6_18_g2197( \3528 , \3403 , \3407 );
xor mul_6_18_g2198( \3529 , \3528 , \3412 );
and mul_6_18_g2199( \3530 , \3526 , \3529 );
and mul_6_18_g2200( \3531 , \3524 , \3529 );
or mul_6_18_g2201( \3532 , \3527 , \3530 , \3531 );
xor mul_6_18_g2202( \3533 , \3399 , \3415 );
xor mul_6_18_g2203( \3534 , \3533 , \3418 );
and mul_6_18_g2204( \3535 , \3532 , \3534 );
xor mul_6_18_g2205( \3536 , \3472 , \3474 );
xor mul_6_18_g2206( \3537 , \3536 , \3477 );
and mul_6_18_g2207( \3538 , \3534 , \3537 );
and mul_6_18_g2208( \3539 , \3532 , \3537 );
or mul_6_18_g2209( \3540 , \3535 , \3538 , \3539 );
and mul_6_18_g2210( \3541 , \3492 , \3540 );
xor mul_6_18_g2211( \3542 , \3492 , \3540 );
xor mul_6_18_g2212( \3543 , \3532 , \3534 );
xor mul_6_18_g2213( \3544 , \3543 , \3537 );
xor mul_6_18_g2214( \3545 , \3512 , \3515 );
and mul_6_18_g2215( \3546 , \1533 , \1382 );
and mul_6_18_g2216( \3547 , \1540 , \1380 );
nor mul_6_18_g2217( \3548 , \3546 , \3547 );
xnor mul_6_18_g2218( \3549 , \3548 , \1389 );
and mul_6_18_g2219( \3550 , \3545 , \3549 );
and mul_6_18_g2220( \3551 , \1498 , \1460 );
and mul_6_18_g2221( \3552 , \1553 , \1458 );
nor mul_6_18_g2222( \3553 , \3551 , \3552 );
xnor mul_6_18_g2223( \3554 , \3553 , \1467 );
and mul_6_18_g2224( \3555 , \3549 , \3554 );
and mul_6_18_g2225( \3556 , \3545 , \3554 );
or mul_6_18_g2226( \3557 , \3550 , \3555 , \3556 );
xor mul_6_18_g2227( \3558 , \3444 , \3448 );
xor mul_6_18_g2228( \3559 , \3558 , \3368 );
and mul_6_18_g2229( \3560 , \3557 , \3559 );
xor mul_6_18_g2230( \3561 , \3457 , \3461 );
xor mul_6_18_g2231( \3562 , \3561 , \3466 );
and mul_6_18_g2232( \3563 , \3559 , \3562 );
and mul_6_18_g2233( \3564 , \3557 , \3562 );
or mul_6_18_g2234( \3565 , \3560 , \3563 , \3564 );
xor mul_6_18_g2235( \3566 , \3440 , \3452 );
xor mul_6_18_g2236( \3567 , \3566 , \3469 );
and mul_6_18_g2237( \3568 , \3565 , \3567 );
xor mul_6_18_g2238( \3569 , \3524 , \3526 );
xor mul_6_18_g2239( \3570 , \3569 , \3529 );
and mul_6_18_g2240( \3571 , \3567 , \3570 );
and mul_6_18_g2241( \3572 , \3565 , \3570 );
or mul_6_18_g2242( \3573 , \3568 , \3571 , \3572 );
and mul_6_18_g2243( \3574 , \3544 , \3573 );
xor mul_6_18_g2244( \3575 , \3544 , \3573 );
xor mul_6_18_g2245( \3576 , \3565 , \3567 );
xor mul_6_18_g2246( \3577 , \3576 , \3570 );
and mul_6_18_g2247( \3578 , \1407 , \1431 );
and mul_6_18_g2248( \3579 , \1416 , \1429 );
nor mul_6_18_g2249( \3580 , \3578 , \3579 );
xnor mul_6_18_g2250( \3581 , \3580 , \1438 );
and mul_6_18_g2251( \3582 , \1526 , \1444 );
and mul_6_18_g2252( \3583 , \1622 , \1442 );
nor mul_6_18_g2253( \3584 , \3582 , \3583 );
xnor mul_6_18_g2254( \3585 , \3584 , \1451 );
and mul_6_18_g2255( \3586 , \3581 , \3585 );
and mul_6_18_g2256( \3587 , \3585 , \3513 );
and mul_6_18_g2257( \3588 , \3581 , \3513 );
or mul_6_18_g2258( \3589 , \3586 , \3587 , \3588 );
and mul_6_18_g2259( \3590 , \1586 , \1336 );
and mul_6_18_g2260( \3591 , \1616 , \1333 );
nor mul_6_18_g2261( \3592 , \3590 , \3591 );
xnor mul_6_18_g2262( \3593 , \3592 , \1332 );
and mul_6_18_g2263( \3594 , \1540 , \1349 );
and mul_6_18_g2264( \3595 , \1517 , \1347 );
nor mul_6_18_g2265( \3596 , \3594 , \3595 );
xnor mul_6_18_g2266( \3597 , \3596 , \1356 );
and mul_6_18_g2267( \3598 , \3593 , \3597 );
and mul_6_18_g2268( \3599 , \1553 , \1382 );
and mul_6_18_g2269( \3600 , \1533 , \1380 );
nor mul_6_18_g2270( \3601 , \3599 , \3600 );
xnor mul_6_18_g2271( \3602 , \3601 , \1389 );
and mul_6_18_g2272( \3603 , \3597 , \3602 );
and mul_6_18_g2273( \3604 , \3593 , \3602 );
or mul_6_18_g2274( \3605 , \3598 , \3603 , \3604 );
and mul_6_18_g2275( \3606 , \3589 , \3605 );
xor mul_6_18_g2276( \3607 , \3545 , \3549 );
xor mul_6_18_g2277( \3608 , \3607 , \3554 );
and mul_6_18_g2278( \3609 , \3605 , \3608 );
and mul_6_18_g2279( \3610 , \3589 , \3608 );
or mul_6_18_g2280( \3611 , \3606 , \3609 , \3610 );
xor mul_6_18_g2281( \3612 , \3508 , \3516 );
xor mul_6_18_g2282( \3613 , \3612 , \3521 );
and mul_6_18_g2283( \3614 , \3611 , \3613 );
xor mul_6_18_g2284( \3615 , \3557 , \3559 );
xor mul_6_18_g2285( \3616 , \3615 , \3562 );
and mul_6_18_g2286( \3617 , \3613 , \3616 );
and mul_6_18_g2287( \3618 , \3611 , \3616 );
or mul_6_18_g2288( \3619 , \3614 , \3617 , \3618 );
and mul_6_18_g2289( \3620 , \3577 , \3619 );
xor mul_6_18_g2290( \3621 , \3577 , \3619 );
xor mul_6_18_g2291( \3622 , \3611 , \3613 );
xor mul_6_18_g2292( \3623 , \3622 , \3616 );
and mul_6_18_g2293( \3624 , \1416 , \1336 );
and mul_6_18_g2294( \3625 , \1586 , \1333 );
nor mul_6_18_g2295( \3626 , \3624 , \3625 );
xnor mul_6_18_g2296( \3627 , \3626 , \1332 );
and mul_6_18_g2297( \3628 , \1517 , \1444 );
and mul_6_18_g2298( \3629 , \1526 , \1442 );
nor mul_6_18_g2299( \3630 , \3628 , \3629 );
xnor mul_6_18_g2300( \3631 , \3630 , \1451 );
and mul_6_18_g2301( \3632 , \3627 , \3631 );
and mul_6_18_g2302( \3633 , \1533 , \1349 );
and mul_6_18_g2303( \3634 , \1540 , \1347 );
nor mul_6_18_g2304( \3635 , \3633 , \3634 );
xnor mul_6_18_g2305( \3636 , \3635 , \1356 );
and mul_6_18_g2306( \3637 , \3631 , \3636 );
and mul_6_18_g2307( \3638 , \3627 , \3636 );
or mul_6_18_g2308( \3639 , \3632 , \3637 , \3638 );
and mul_6_18_g2309( \3640 , \1622 , \1431 );
and mul_6_18_g2310( \3641 , \1407 , \1429 );
nor mul_6_18_g2311( \3642 , \3640 , \3641 );
xnor mul_6_18_g2312( \3643 , \3642 , \1438 );
and mul_6_18_g2313( \3644 , \1498 , \1380 );
not mul_6_18_g2314( \3645 , \3644 );
and mul_6_18_g2315( \3646 , \3645 , \1389 );
and mul_6_18_g2316( \3647 , \3643 , \3646 );
and mul_6_18_g2317( \3648 , \3639 , \3647 );
xor mul_6_18_g2318( \3649 , \3581 , \3585 );
xor mul_6_18_g2319( \3650 , \3649 , \3513 );
and mul_6_18_g2320( \3651 , \3647 , \3650 );
and mul_6_18_g2321( \3652 , \3639 , \3650 );
or mul_6_18_g2322( \3653 , \3648 , \3651 , \3652 );
xor mul_6_18_g2323( \3654 , \3496 , \3500 );
xor mul_6_18_g2324( \3655 , \3654 , \3505 );
and mul_6_18_g2325( \3656 , \3653 , \3655 );
xor mul_6_18_g2326( \3657 , \3589 , \3605 );
xor mul_6_18_g2327( \3658 , \3657 , \3608 );
and mul_6_18_g2328( \3659 , \3655 , \3658 );
and mul_6_18_g2329( \3660 , \3653 , \3658 );
or mul_6_18_g2330( \3661 , \3656 , \3659 , \3660 );
and mul_6_18_g2331( \3662 , \3623 , \3661 );
xor mul_6_18_g2332( \3663 , \3623 , \3661 );
xor mul_6_18_g2333( \3664 , \3643 , \3646 );
and mul_6_18_g2334( \3665 , \1526 , \1431 );
and mul_6_18_g2335( \3666 , \1622 , \1429 );
nor mul_6_18_g2336( \3667 , \3665 , \3666 );
xnor mul_6_18_g2337( \3668 , \3667 , \1438 );
and mul_6_18_g2338( \3669 , \1540 , \1444 );
and mul_6_18_g2339( \3670 , \1517 , \1442 );
nor mul_6_18_g2340( \3671 , \3669 , \3670 );
xnor mul_6_18_g2341( \3672 , \3671 , \1451 );
and mul_6_18_g2342( \3673 , \3668 , \3672 );
and mul_6_18_g2343( \3674 , \3672 , \3644 );
and mul_6_18_g2344( \3675 , \3668 , \3644 );
or mul_6_18_g2345( \3676 , \3673 , \3674 , \3675 );
and mul_6_18_g2346( \3677 , \3664 , \3676 );
and mul_6_18_g2347( \3678 , \1498 , \1382 );
and mul_6_18_g2348( \3679 , \1553 , \1380 );
nor mul_6_18_g2349( \3680 , \3678 , \3679 );
xnor mul_6_18_g2350( \3681 , \3680 , \1389 );
and mul_6_18_g2351( \3682 , \3676 , \3681 );
and mul_6_18_g2352( \3683 , \3664 , \3681 );
or mul_6_18_g2353( \3684 , \3677 , \3682 , \3683 );
xor mul_6_18_g2354( \3685 , \3593 , \3597 );
xor mul_6_18_g2355( \3686 , \3685 , \3602 );
and mul_6_18_g2356( \3687 , \3684 , \3686 );
xor mul_6_18_g2357( \3688 , \3639 , \3647 );
xor mul_6_18_g2358( \3689 , \3688 , \3650 );
and mul_6_18_g2359( \3690 , \3686 , \3689 );
and mul_6_18_g2360( \3691 , \3684 , \3689 );
or mul_6_18_g2361( \3692 , \3687 , \3690 , \3691 );
xor mul_6_18_g2362( \3693 , \3653 , \3655 );
xor mul_6_18_g2363( \3694 , \3693 , \3658 );
and mul_6_18_g2364( \3695 , \3692 , \3694 );
xor mul_6_18_g2365( \3696 , \3692 , \3694 );
xor mul_6_18_g2366( \3697 , \3684 , \3686 );
xor mul_6_18_g2367( \3698 , \3697 , \3689 );
and mul_6_18_g2368( \3699 , \1517 , \1431 );
and mul_6_18_g2369( \3700 , \1526 , \1429 );
nor mul_6_18_g2370( \3701 , \3699 , \3700 );
xnor mul_6_18_g2371( \3702 , \3701 , \1438 );
and mul_6_18_g2372( \3703 , \1498 , \1347 );
not mul_6_18_g2373( \3704 , \3703 );
and mul_6_18_g2374( \3705 , \3704 , \1356 );
and mul_6_18_g2375( \3706 , \3702 , \3705 );
and mul_6_18_g2376( \3707 , \1407 , \1336 );
and mul_6_18_g2377( \3708 , \1416 , \1333 );
nor mul_6_18_g2378( \3709 , \3707 , \3708 );
xnor mul_6_18_g2379( \3710 , \3709 , \1332 );
and mul_6_18_g2380( \3711 , \3706 , \3710 );
and mul_6_18_g2381( \3712 , \1553 , \1349 );
and mul_6_18_g2382( \3713 , \1533 , \1347 );
nor mul_6_18_g2383( \3714 , \3712 , \3713 );
xnor mul_6_18_g2384( \3715 , \3714 , \1356 );
and mul_6_18_g2385( \3716 , \3710 , \3715 );
and mul_6_18_g2386( \3717 , \3706 , \3715 );
or mul_6_18_g2387( \3718 , \3711 , \3716 , \3717 );
xor mul_6_18_g2388( \3719 , \3627 , \3631 );
xor mul_6_18_g2389( \3720 , \3719 , \3636 );
and mul_6_18_g2390( \3721 , \3718 , \3720 );
xor mul_6_18_g2391( \3722 , \3664 , \3676 );
xor mul_6_18_g2392( \3723 , \3722 , \3681 );
and mul_6_18_g2393( \3724 , \3720 , \3723 );
and mul_6_18_g2394( \3725 , \3718 , \3723 );
or mul_6_18_g2395( \3726 , \3721 , \3724 , \3725 );
and mul_6_18_g2396( \3727 , \3698 , \3726 );
xor mul_6_18_g2397( \3728 , \3698 , \3726 );
xor mul_6_18_g2398( \3729 , \3718 , \3720 );
xor mul_6_18_g2399( \3730 , \3729 , \3723 );
and mul_6_18_g2400( \3731 , \1622 , \1336 );
and mul_6_18_g2401( \3732 , \1407 , \1333 );
nor mul_6_18_g2402( \3733 , \3731 , \3732 );
xnor mul_6_18_g2403( \3734 , \3733 , \1332 );
and mul_6_18_g2404( \3735 , \1533 , \1444 );
and mul_6_18_g2405( \3736 , \1540 , \1442 );
nor mul_6_18_g2406( \3737 , \3735 , \3736 );
xnor mul_6_18_g2407( \3738 , \3737 , \1451 );
and mul_6_18_g2408( \3739 , \3734 , \3738 );
and mul_6_18_g2409( \3740 , \1498 , \1349 );
and mul_6_18_g2410( \3741 , \1553 , \1347 );
nor mul_6_18_g2411( \3742 , \3740 , \3741 );
xnor mul_6_18_g2412( \3743 , \3742 , \1356 );
and mul_6_18_g2413( \3744 , \3738 , \3743 );
and mul_6_18_g2414( \3745 , \3734 , \3743 );
or mul_6_18_g2415( \3746 , \3739 , \3744 , \3745 );
xor mul_6_18_g2416( \3747 , \3668 , \3672 );
xor mul_6_18_g2417( \3748 , \3747 , \3644 );
and mul_6_18_g2418( \3749 , \3746 , \3748 );
xor mul_6_18_g2419( \3750 , \3706 , \3710 );
xor mul_6_18_g2420( \3751 , \3750 , \3715 );
and mul_6_18_g2421( \3752 , \3748 , \3751 );
and mul_6_18_g2422( \3753 , \3746 , \3751 );
or mul_6_18_g2423( \3754 , \3749 , \3752 , \3753 );
and mul_6_18_g2424( \3755 , \3730 , \3754 );
xor mul_6_18_g2425( \3756 , \3730 , \3754 );
xor mul_6_18_g2426( \3757 , \3702 , \3705 );
and mul_6_18_g2427( \3758 , \1540 , \1431 );
and mul_6_18_g2428( \3759 , \1517 , \1429 );
nor mul_6_18_g2429( \3760 , \3758 , \3759 );
xnor mul_6_18_g2430( \3761 , \3760 , \1438 );
and mul_6_18_g2431( \3762 , \1553 , \1444 );
and mul_6_18_g2432( \3763 , \1533 , \1442 );
nor mul_6_18_g2433( \3764 , \3762 , \3763 );
xnor mul_6_18_g2434( \3765 , \3764 , \1451 );
and mul_6_18_g2435( \3766 , \3761 , \3765 );
and mul_6_18_g2436( \3767 , \3765 , \3703 );
and mul_6_18_g2437( \3768 , \3761 , \3703 );
or mul_6_18_g2438( \3769 , \3766 , \3767 , \3768 );
and mul_6_18_g2439( \3770 , \3757 , \3769 );
xor mul_6_18_g2440( \3771 , \3734 , \3738 );
xor mul_6_18_g2441( \3772 , \3771 , \3743 );
and mul_6_18_g2442( \3773 , \3769 , \3772 );
and mul_6_18_g2443( \3774 , \3757 , \3772 );
or mul_6_18_g2444( \3775 , \3770 , \3773 , \3774 );
xor mul_6_18_g2445( \3776 , \3746 , \3748 );
xor mul_6_18_g2446( \3777 , \3776 , \3751 );
and mul_6_18_g2447( \3778 , \3775 , \3777 );
xor mul_6_18_g2448( \3779 , \3775 , \3777 );
xor mul_6_18_g2449( \3780 , \3757 , \3769 );
xor mul_6_18_g2450( \3781 , \3780 , \3772 );
and mul_6_18_g2451( \3782 , \1533 , \1431 );
and mul_6_18_g2452( \3783 , \1540 , \1429 );
nor mul_6_18_g2453( \3784 , \3782 , \3783 );
xnor mul_6_18_g2454( \3785 , \3784 , \1438 );
and mul_6_18_g2455( \3786 , \1498 , \1442 );
not mul_6_18_g2456( \3787 , \3786 );
and mul_6_18_g2457( \3788 , \3787 , \1451 );
and mul_6_18_g2458( \3789 , \3785 , \3788 );
and mul_6_18_g2459( \3790 , \1526 , \1336 );
and mul_6_18_g2460( \3791 , \1622 , \1333 );
nor mul_6_18_g2461( \3792 , \3790 , \3791 );
xnor mul_6_18_g2462( \3793 , \3792 , \1332 );
and mul_6_18_g2463( \3794 , \3789 , \3793 );
xor mul_6_18_g2464( \3795 , \3761 , \3765 );
xor mul_6_18_g2465( \3796 , \3795 , \3703 );
and mul_6_18_g2466( \3797 , \3793 , \3796 );
and mul_6_18_g2467( \3798 , \3789 , \3796 );
or mul_6_18_g2468( \3799 , \3794 , \3797 , \3798 );
and mul_6_18_g2469( \3800 , \3781 , \3799 );
xor mul_6_18_g2470( \3801 , \3781 , \3799 );
xor mul_6_18_g2471( \3802 , \3789 , \3793 );
xor mul_6_18_g2472( \3803 , \3802 , \3796 );
xor mul_6_18_g2473( \3804 , \3785 , \3788 );
and mul_6_18_g2474( \3805 , \1517 , \1336 );
and mul_6_18_g2475( \3806 , \1526 , \1333 );
nor mul_6_18_g2476( \3807 , \3805 , \3806 );
xnor mul_6_18_g2477( \3808 , \3807 , \1332 );
and mul_6_18_g2478( \3809 , \3804 , \3808 );
and mul_6_18_g2479( \3810 , \1498 , \1444 );
and mul_6_18_g2480( \3811 , \1553 , \1442 );
nor mul_6_18_g2481( \3812 , \3810 , \3811 );
xnor mul_6_18_g2482( \3813 , \3812 , \1451 );
and mul_6_18_g2483( \3814 , \3808 , \3813 );
and mul_6_18_g2484( \3815 , \3804 , \3813 );
or mul_6_18_g2485( \3816 , \3809 , \3814 , \3815 );
and mul_6_18_g2486( \3817 , \3803 , \3816 );
xor mul_6_18_g2487( \3818 , \3803 , \3816 );
and mul_6_18_g2488( \3819 , \1540 , \1336 );
and mul_6_18_g2489( \3820 , \1517 , \1333 );
nor mul_6_18_g2490( \3821 , \3819 , \3820 );
xnor mul_6_18_g2491( \3822 , \3821 , \1332 );
and mul_6_18_g2492( \3823 , \1553 , \1431 );
and mul_6_18_g2493( \3824 , \1533 , \1429 );
nor mul_6_18_g2494( \3825 , \3823 , \3824 );
xnor mul_6_18_g2495( \3826 , \3825 , \1438 );
and mul_6_18_g2496( \3827 , \3822 , \3826 );
and mul_6_18_g2497( \3828 , \3826 , \3786 );
and mul_6_18_g2498( \3829 , \3822 , \3786 );
or mul_6_18_g2499( \3830 , \3827 , \3828 , \3829 );
xor mul_6_18_g2500( \3831 , \3804 , \3808 );
xor mul_6_18_g2501( \3832 , \3831 , \3813 );
and mul_6_18_g2502( \3833 , \3830 , \3832 );
xor mul_6_18_g2503( \3834 , \3830 , \3832 );
xor mul_6_18_g2504( \3835 , \3822 , \3826 );
xor mul_6_18_g2505( \3836 , \3835 , \3786 );
and mul_6_18_g2506( \3837 , \1498 , \1429 );
not mul_6_18_g2507( \3838 , \3837 );
and mul_6_18_g2508( \3839 , \3838 , \1438 );
and mul_6_18_g2509( \3840 , \1498 , \1431 );
and mul_6_18_g2510( \3841 , \1553 , \1429 );
nor mul_6_18_g2511( \3842 , \3840 , \3841 );
xnor mul_6_18_g2512( \3843 , \3842 , \1438 );
and mul_6_18_g2513( \3844 , \3839 , \3843 );
and mul_6_18_g2514( \3845 , \3836 , \3844 );
xor mul_6_18_g2515( \3846 , \3836 , \3844 );
and mul_6_18_g2516( \3847 , \1533 , \1336 );
and mul_6_18_g2517( \3848 , \1540 , \1333 );
nor mul_6_18_g2518( \3849 , \3847 , \3848 );
xnor mul_6_18_g2519( \3850 , \3849 , \1332 );
xor mul_6_18_g2520( \3851 , \3839 , \3843 );
and mul_6_18_g2521( \3852 , \3850 , \3851 );
xor mul_6_18_g2522( \3853 , \3850 , \3851 );
and mul_6_18_g2523( \3854 , \1553 , \1336 );
and mul_6_18_g2524( \3855 , \1533 , \1333 );
nor mul_6_18_g2525( \3856 , \3854 , \3855 );
xnor mul_6_18_g2526( \3857 , \3856 , \1332 );
and mul_6_18_g2527( \3858 , \3857 , \3837 );
xor mul_6_18_g2528( \3859 , \3857 , \3837 );
and mul_6_18_g2529( \3860 , \1498 , \1336 );
and mul_6_18_g2530( \3861 , \1553 , \1333 );
nor mul_6_18_g2531( \3862 , \3860 , \3861 );
xnor mul_6_18_g2532( \3863 , \3862 , \1332 );
and mul_6_18_g2533( \3864 , \1498 , \1333 );
not mul_6_18_g2534( \3865 , \3864 );
and mul_6_18_g2535( \3866 , \3865 , \1332 );
and mul_6_18_g2536( \3867 , \3863 , \3866 );
and mul_6_18_g2537( \3868 , \3859 , \3867 );
or mul_6_18_g2538( \3869 , \3858 , \3868 );
and mul_6_18_g2539( \3870 , \3853 , \3869 );
or mul_6_18_g2540( \3871 , \3852 , \3870 );
and mul_6_18_g2541( \3872 , \3846 , \3871 );
or mul_6_18_g2542( \3873 , \3845 , \3872 );
and mul_6_18_g2543( \3874 , \3834 , \3873 );
or mul_6_18_g2544( \3875 , \3833 , \3874 );
and mul_6_18_g2545( \3876 , \3818 , \3875 );
or mul_6_18_g2546( \3877 , \3817 , \3876 );
and mul_6_18_g2547( \3878 , \3801 , \3877 );
or mul_6_18_g2548( \3879 , \3800 , \3878 );
and mul_6_18_g2549( \3880 , \3779 , \3879 );
or mul_6_18_g2550( \3881 , \3778 , \3880 );
and mul_6_18_g2551( \3882 , \3756 , \3881 );
or mul_6_18_g2552( \3883 , \3755 , \3882 );
and mul_6_18_g2553( \3884 , \3728 , \3883 );
or mul_6_18_g2554( \3885 , \3727 , \3884 );
and mul_6_18_g2555( \3886 , \3696 , \3885 );
or mul_6_18_g2556( \3887 , \3695 , \3886 );
and mul_6_18_g2557( \3888 , \3663 , \3887 );
or mul_6_18_g2558( \3889 , \3662 , \3888 );
and mul_6_18_g2559( \3890 , \3621 , \3889 );
or mul_6_18_g2560( \3891 , \3620 , \3890 );
and mul_6_18_g2561( \3892 , \3575 , \3891 );
or mul_6_18_g2562( \3893 , \3574 , \3892 );
and mul_6_18_g2563( \3894 , \3542 , \3893 );
or mul_6_18_g2564( \3895 , \3541 , \3894 );
and mul_6_18_g2565( \3896 , \3490 , \3895 );
or mul_6_18_g2566( \3897 , \3489 , \3896 );
and mul_6_18_g2567( \3898 , \3437 , \3897 );
or mul_6_18_g2568( \3899 , \3436 , \3898 );
and mul_6_18_g2569( \3900 , \3361 , \3899 );
or mul_6_18_g2570( \3901 , \3360 , \3900 );
and mul_6_18_g2571( \3902 , \3298 , \3901 );
or mul_6_18_g2572( \3903 , \3297 , \3902 );
and mul_6_18_g2573( \3904 , \3226 , \3903 );
or mul_6_18_g2574( \3905 , \3225 , \3904 );
and mul_6_18_g2575( \3906 , \3196 , \3905 );
or mul_6_18_g2576( \3907 , \3195 , \3906 );
and mul_6_18_g2577( \3908 , \3073 , \3907 );
or mul_6_18_g2578( \3909 , \3072 , \3908 );
and mul_6_18_g2579( \3910 , \3005 , \3909 );
or mul_6_18_g2580( \3911 , \3004 , \3910 );
and mul_6_18_g2581( \3912 , \2922 , \3911 );
or mul_6_18_g2582( \3913 , \2921 , \3912 );
and mul_6_18_g2583( \3914 , \2856 , \3913 );
or mul_6_18_g2584( \3915 , \2855 , \3914 );
and mul_6_18_g2585( \3916 , \2764 , \3915 );
or mul_6_18_g2586( \3917 , \2763 , \3916 );
and mul_6_18_g2587( \3918 , \2635 , \3917 );
or mul_6_18_g2588( \3919 , \2634 , \3918 );
and mul_6_18_g2589( \3920 , \2518 , \3919 );
or mul_6_18_g2590( \3921 , \2517 , \3920 );
and mul_6_18_g2591( \3922 , \2406 , \3921 );
or mul_6_18_g2592( \3923 , \2405 , \3922 );
and mul_6_18_g2593( \3924 , \2290 , \3923 );
or mul_6_18_g2594( \3925 , \2289 , \3924 );
xor mul_6_18_g2595( \3926 , \2252 , \3925 );
buf \mul_6_18/Z[31] ( \3927_Z[31] , \3926 );
xor mul_6_18_g2596( \3928 , \2290 , \3923 );
buf \mul_6_18/Z[30] ( \3929_Z[30] , \3928 );
xor mul_6_18_g2597( \3930 , \2406 , \3921 );
buf \mul_6_18/Z[29] ( \3931_Z[29] , \3930 );
xor mul_6_18_g2598( \3932 , \2518 , \3919 );
buf \mul_6_18/Z[28] ( \3933_Z[28] , \3932 );
xor mul_6_18_g2599( \3934 , \2635 , \3917 );
buf \mul_6_18/Z[27] ( \3935_Z[27] , \3934 );
xor mul_6_18_g2600( \3936 , \2764 , \3915 );
buf \mul_6_18/Z[26] ( \3937_Z[26] , \3936 );
xor mul_6_18_g2601( \3938 , \2856 , \3913 );
buf \mul_6_18/Z[25] ( \3939_Z[25] , \3938 );
xor mul_6_18_g2602( \3940 , \2922 , \3911 );
buf \mul_6_18/Z[24] ( \3941_Z[24] , \3940 );
xor mul_6_18_g2603( \3942 , \3005 , \3909 );
buf \mul_6_18/Z[23] ( \3943_Z[23] , \3942 );
xor mul_6_18_g2604( \3944 , \3073 , \3907 );
buf \mul_6_18/Z[22] ( \3945_Z[22] , \3944 );
xor mul_6_18_g2605( \3946 , \3196 , \3905 );
buf \mul_6_18/Z[21] ( \3947_Z[21] , \3946 );
xor mul_6_18_g2606( \3948 , \3226 , \3903 );
buf \mul_6_18/Z[20] ( \3949_Z[20] , \3948 );
xor mul_6_18_g2607( \3950 , \3298 , \3901 );
buf \mul_6_18/Z[19] ( \3951_Z[19] , \3950 );
xor mul_6_18_g2608( \3952 , \3361 , \3899 );
buf \mul_6_18/Z[18] ( \3953_Z[18] , \3952 );
xor mul_6_18_g2609( \3954 , \3437 , \3897 );
buf \mul_6_18/Z[17] ( \3955_Z[17] , \3954 );
xor mul_6_18_g2610( \3956 , \3490 , \3895 );
buf \mul_6_18/Z[16] ( \3957_Z[16] , \3956 );
xor mul_6_18_g2611( \3958 , \3542 , \3893 );
buf \mul_6_18/Z[15] ( \3959_Z[15] , \3958 );
xor mul_6_18_g2612( \3960 , \3575 , \3891 );
buf \mul_6_18/Z[14] ( \3961_Z[14] , \3960 );
xor mul_6_18_g2613( \3962 , \3621 , \3889 );
buf \mul_6_18/Z[13] ( \3963_Z[13] , \3962 );
xor mul_6_18_g2614( \3964 , \3663 , \3887 );
buf \mul_6_18/Z[12] ( \3965_Z[12] , \3964 );
xor mul_6_18_g2615( \3966 , \3696 , \3885 );
buf \mul_6_18/Z[11] ( \3967_Z[11] , \3966 );
xor mul_6_18_g2616( \3968 , \3728 , \3883 );
buf \mul_6_18/Z[10] ( \3969_Z[10] , \3968 );
xor mul_6_18_g2617( \3970 , \3756 , \3881 );
buf \mul_6_18/Z[9] ( \3971_Z[9] , \3970 );
xor mul_6_18_g2618( \3972 , \3779 , \3879 );
buf \mul_6_18/Z[8] ( \3973_Z[8] , \3972 );
xor mul_6_18_g2619( \3974 , \3801 , \3877 );
buf \mul_6_18/Z[7] ( \3975_Z[7] , \3974 );
xor mul_6_18_g2620( \3976 , \3818 , \3875 );
buf \mul_6_18/Z[6] ( \3977_Z[6] , \3976 );
xor mul_6_18_g2621( \3978 , \3834 , \3873 );
buf \mul_6_18/Z[5] ( \3979_Z[5] , \3978 );
xor mul_6_18_g2622( \3980 , \3846 , \3871 );
buf \mul_6_18/Z[4] ( \3981_Z[4] , \3980 );
xor mul_6_18_g2623( \3982 , \3853 , \3869 );
buf \mul_6_18/Z[3] ( \3983_Z[3] , \3982 );
xor mul_6_18_g2624( \3984 , \3859 , \3867 );
buf \mul_6_18/Z[2] ( \3985_Z[2] , \3984 );
xor mul_6_18_g2625( \3986 , \3863 , \3866 );
buf \mul_6_18/Z[1] ( \3987_Z[1] , \3986 );
buf mul_6_18_g2626( \3988 , \3864 );
buf \mul_6_18/Z[0] ( \3989_Z[0] , \3988 );
endmodule

