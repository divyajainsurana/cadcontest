//
// Conformal-LEC Version 20.10-d005 (29-Apr-2020)
//
module top(RI2b1c4342d4e0_65,RI2b1c4342c5e0_33,RI2b1c4342b6e0_1,RI2b1c4342d558_66,RI2b1c4342d5d0_67,RI2b1c4342d648_68,RI2b1c4342d6c0_69,RI2b1c4342d738_70,RI2b1c4342d7b0_71,
        RI2b1c4342d828_72,RI2b1c4342d8a0_73,RI2b1c4342d918_74,RI2b1c4342d990_75,RI2b1c4342da08_76,RI2b1c4342da80_77,RI2b1c4342daf8_78,RI2b1c4342db70_79,RI2b1c4342dbe8_80,RI2b1c4342dc60_81,
        RI2b1c4342dcd8_82,RI2b1c4342dd50_83,RI2b1c4342ddc8_84,RI2b1c4342de40_85,RI2b1c4342deb8_86,RI2b1c4342df30_87,RI2b1c4342dfa8_88,RI2b1c4342e020_89,RI2b1c4342e098_90,RI2b1c4342e110_91,
        RI2b1c4342e188_92,RI2b1c4342e200_93,RI2b1c4342e278_94,RI2b1c4342e2f0_95,RI2b1c4342e368_96,RI2b1c4342c658_34,RI2b1c4342b758_2,RI2b1c4342c6d0_35,RI2b1c4342b7d0_3,RI2b1c4342c748_36,
        RI2b1c4342b848_4,RI2b1c4342c7c0_37,RI2b1c4342b8c0_5,RI2b1c4342c838_38,RI2b1c4342b938_6,RI2b1c4342c8b0_39,RI2b1c4342b9b0_7,RI2b1c4342c928_40,RI2b1c4342ba28_8,RI2b1c4342c9a0_41,
        RI2b1c4342baa0_9,RI2b1c4342ca18_42,RI2b1c4342bb18_10,RI2b1c4342ca90_43,RI2b1c4342bb90_11,RI2b1c4342cb08_44,RI2b1c4342bc08_12,RI2b1c4342cb80_45,RI2b1c4342bc80_13,RI2b1c4342cbf8_46,
        RI2b1c4342bcf8_14,RI2b1c4342cc70_47,RI2b1c4342bd70_15,RI2b1c4342cce8_48,RI2b1c4342bde8_16,RI2b1c4342cd60_49,RI2b1c4342be60_17,RI2b1c4342cdd8_50,RI2b1c4342bed8_18,RI2b1c4342ce50_51,
        RI2b1c4342bf50_19,RI2b1c4342cec8_52,RI2b1c4342bfc8_20,RI2b1c4342cf40_53,RI2b1c4342c040_21,RI2b1c4342cfb8_54,RI2b1c4342c0b8_22,RI2b1c4342d030_55,RI2b1c4342c130_23,RI2b1c4342d0a8_56,
        RI2b1c4342c1a8_24,RI2b1c4342d120_57,RI2b1c4342c220_25,RI2b1c4342d198_58,RI2b1c4342c298_26,RI2b1c4342d210_59,RI2b1c4342c310_27,RI2b1c4342d288_60,RI2b1c4342c388_28,RI2b1c4342d300_61,
        RI2b1c4342c400_29,RI2b1c4342d378_62,RI2b1c4342c478_30,RI2b1c4342d3f0_63,RI2b1c4342c4f0_31,RI2b1c4342d468_64,RI2b1c4342c568_32,R_61_7d2b4e8,R_62_7d2b590,R_63_7d2b638,
        R_64_7d2b6e0,R_65_7d2b788,R_66_7d2b830,R_67_7d2b8d8,R_68_7d2b980,R_69_7d2ba28,R_6a_7d2bad0,R_6b_7d2bb78,R_6c_7d2bc20,R_6d_7d2bcc8,
        R_6e_7d2bd70,R_6f_7d2be18,R_70_7d2bec0,R_71_7d2bf68,R_72_7d2c010,R_73_7d2c0b8,R_74_7d2c160,R_75_7d2c208,R_76_7d2c2b0,R_77_7d2c358,
        R_78_7d2c400,R_79_7d2c4a8,R_7a_7d2c550,R_7b_7d2c5f8,R_7c_7d2c6a0,R_7d_7d2c748,R_7e_7d2c7f0,R_7f_7d2c898,R_80_7d2c940,R_81_7d2c9e8,
        R_82_7d2ca90,R_83_7d2cb38,R_84_7d2cbe0,R_85_7d2cc88,R_86_7d2cd30,R_87_7d2cdd8,R_88_7d2ce80,R_89_7d2cf28,R_8a_7d2cfd0,R_8b_7d2d078,
        R_8c_7d2d120,R_8d_7d2d1c8,R_8e_7d2d270,R_8f_7d2d318,R_90_7d2d3c0,R_91_7d2d468,R_92_7d2d510,R_93_7d2d5b8,R_94_7d2d660,R_95_7d2d708,
        R_96_7d2d7b0,R_97_7d2d858,R_98_7d2d900,R_99_7d2d9a8,R_9a_7d2da50,R_9b_7d2daf8);
input RI2b1c4342d4e0_65,RI2b1c4342c5e0_33,RI2b1c4342b6e0_1,RI2b1c4342d558_66,RI2b1c4342d5d0_67,RI2b1c4342d648_68,RI2b1c4342d6c0_69,RI2b1c4342d738_70,RI2b1c4342d7b0_71,
        RI2b1c4342d828_72,RI2b1c4342d8a0_73,RI2b1c4342d918_74,RI2b1c4342d990_75,RI2b1c4342da08_76,RI2b1c4342da80_77,RI2b1c4342daf8_78,RI2b1c4342db70_79,RI2b1c4342dbe8_80,RI2b1c4342dc60_81,
        RI2b1c4342dcd8_82,RI2b1c4342dd50_83,RI2b1c4342ddc8_84,RI2b1c4342de40_85,RI2b1c4342deb8_86,RI2b1c4342df30_87,RI2b1c4342dfa8_88,RI2b1c4342e020_89,RI2b1c4342e098_90,RI2b1c4342e110_91,
        RI2b1c4342e188_92,RI2b1c4342e200_93,RI2b1c4342e278_94,RI2b1c4342e2f0_95,RI2b1c4342e368_96,RI2b1c4342c658_34,RI2b1c4342b758_2,RI2b1c4342c6d0_35,RI2b1c4342b7d0_3,RI2b1c4342c748_36,
        RI2b1c4342b848_4,RI2b1c4342c7c0_37,RI2b1c4342b8c0_5,RI2b1c4342c838_38,RI2b1c4342b938_6,RI2b1c4342c8b0_39,RI2b1c4342b9b0_7,RI2b1c4342c928_40,RI2b1c4342ba28_8,RI2b1c4342c9a0_41,
        RI2b1c4342baa0_9,RI2b1c4342ca18_42,RI2b1c4342bb18_10,RI2b1c4342ca90_43,RI2b1c4342bb90_11,RI2b1c4342cb08_44,RI2b1c4342bc08_12,RI2b1c4342cb80_45,RI2b1c4342bc80_13,RI2b1c4342cbf8_46,
        RI2b1c4342bcf8_14,RI2b1c4342cc70_47,RI2b1c4342bd70_15,RI2b1c4342cce8_48,RI2b1c4342bde8_16,RI2b1c4342cd60_49,RI2b1c4342be60_17,RI2b1c4342cdd8_50,RI2b1c4342bed8_18,RI2b1c4342ce50_51,
        RI2b1c4342bf50_19,RI2b1c4342cec8_52,RI2b1c4342bfc8_20,RI2b1c4342cf40_53,RI2b1c4342c040_21,RI2b1c4342cfb8_54,RI2b1c4342c0b8_22,RI2b1c4342d030_55,RI2b1c4342c130_23,RI2b1c4342d0a8_56,
        RI2b1c4342c1a8_24,RI2b1c4342d120_57,RI2b1c4342c220_25,RI2b1c4342d198_58,RI2b1c4342c298_26,RI2b1c4342d210_59,RI2b1c4342c310_27,RI2b1c4342d288_60,RI2b1c4342c388_28,RI2b1c4342d300_61,
        RI2b1c4342c400_29,RI2b1c4342d378_62,RI2b1c4342c478_30,RI2b1c4342d3f0_63,RI2b1c4342c4f0_31,RI2b1c4342d468_64,RI2b1c4342c568_32;
output R_61_7d2b4e8,R_62_7d2b590,R_63_7d2b638,R_64_7d2b6e0,R_65_7d2b788,R_66_7d2b830,R_67_7d2b8d8,R_68_7d2b980,R_69_7d2ba28,
        R_6a_7d2bad0,R_6b_7d2bb78,R_6c_7d2bc20,R_6d_7d2bcc8,R_6e_7d2bd70,R_6f_7d2be18,R_70_7d2bec0,R_71_7d2bf68,R_72_7d2c010,R_73_7d2c0b8,
        R_74_7d2c160,R_75_7d2c208,R_76_7d2c2b0,R_77_7d2c358,R_78_7d2c400,R_79_7d2c4a8,R_7a_7d2c550,R_7b_7d2c5f8,R_7c_7d2c6a0,R_7d_7d2c748,
        R_7e_7d2c7f0,R_7f_7d2c898,R_80_7d2c940,R_81_7d2c9e8,R_82_7d2ca90,R_83_7d2cb38,R_84_7d2cbe0,R_85_7d2cc88,R_86_7d2cd30,R_87_7d2cdd8,
        R_88_7d2ce80,R_89_7d2cf28,R_8a_7d2cfd0,R_8b_7d2d078,R_8c_7d2d120,R_8d_7d2d1c8,R_8e_7d2d270,R_8f_7d2d318,R_90_7d2d3c0,R_91_7d2d468,
        R_92_7d2d510,R_93_7d2d5b8,R_94_7d2d660,R_95_7d2d708,R_96_7d2d7b0,R_97_7d2d858,R_98_7d2d900,R_99_7d2d9a8,R_9a_7d2da50,R_9b_7d2daf8;

wire \156 , \157 , \158 , \159 , \160 , \161 , \162 , \163 , \164 ,
         \165 , \166 , \167 , \168 , \169 , \170 , \171 , \172 , \173 , \174 ,
         \175 , \176 , \177 , \178 , \179 , \180 , \181 , \182 , \183 , \184 ,
         \185 , \186 , \187 , \188 , \189 , \190_N$1 , \191_N$2 , \192_N$3 , \193_N$4 , \194_N$5 ,
         \195_N$6 , \196_N$7 , \197_N$8 , \198_N$9 , \199_N$10 , \200_N$11 , \201_N$12 , \202_N$13 , \203_N$14 , \204_N$15 ,
         \205_N$16 , \206_N$17 , \207_N$18 , \208_N$19 , \209_N$20 , \210_N$21 , \211_N$22 , \212_N$23 , \213_N$24 , \214_N$25 ,
         \215_N$26 , \216_N$27 , \217_N$28 , \218_N$29 , \219_N$30 , \220_N$31 , \221_N$32 , \222_N$34 , \223_ZERO , \224 ,
         \225_N$33 , \226_ONE , \227 , \228_nG2cd , \229 , \230 , \231 , \232 , \233 , \234 ,
         \235 , \236 , \237 , \238 , \239 , \240 , \241 , \242 , \243 , \244 ,
         \245 , \246 , \247 , \248 , \249 , \250 , \251 , \252 , \253 , \254 ,
         \255 , \256 , \257 , \258 , \259 , \260 , \261_nG2cf , \262 , \263 , \264 ,
         \265_nG2bf , \266 , \267_nG2c1 , \268 , \269 , \270 , \271_nG2b1 , \272 , \273_nG2b3 , \274 ,
         \275 , \276 , \277_nG2a3 , \278 , \279_nG2a5 , \280 , \281 , \282 , \283_nG295 , \284 ,
         \285_nG297 , \286 , \287 , \288 , \289_nG287 , \290 , \291_nG289 , \292 , \293 , \294 ,
         \295_nG279 , \296 , \297_nG27b , \298 , \299 , \300 , \301_nG26b , \302 , \303_nG26d , \304 ,
         \305 , \306 , \307_nG25d , \308 , \309_nG25f , \310 , \311 , \312 , \313_nG24f , \314 ,
         \315_nG251 , \316 , \317 , \318 , \319_nG241 , \320 , \321_nG243 , \322 , \323 , \324 ,
         \325_nG233 , \326 , \327_nG235 , \328 , \329 , \330 , \331_nG225 , \332 , \333_nG227 , \334 ,
         \335 , \336 , \337_nG217 , \338 , \339_nG219 , \340 , \341 , \342 , \343_nG209 , \344 ,
         \345_nG20b , \346 , \347 , \348 , \349_nG1fb , \350 , \351_nG1fd , \352 , \353 , \354 ,
         \355_nG1ed , \356 , \357_nG1ef , \358 , \359 , \360 , \361_nG1df , \362 , \363_nG1e1 , \364 ,
         \365 , \366 , \367_nG1d1 , \368 , \369_nG1d3 , \370 , \371 , \372 , \373_nG1c3 , \374 ,
         \375_nG1c5 , \376 , \377 , \378 , \379_nG1b5 , \380 , \381_nG1b7 , \382 , \383 , \384 ,
         \385_nG1a7 , \386 , \387_nG1a9 , \388 , \389 , \390 , \391_nG199 , \392 , \393_nG19b , \394 ,
         \395 , \396 , \397_nG18b , \398 , \399_nG18d , \400 , \401 , \402 , \403_nG17d , \404 ,
         \405_nG17f , \406 , \407 , \408 , \409_nG16f , \410 , \411_nG171 , \412 , \413 , \414 ,
         \415_nG161 , \416 , \417_nG163 , \418 , \419 , \420 , \421_nG153 , \422 , \423_nG155 , \424 ,
         \425 , \426 , \427_nG145 , \428 , \429_nG147 , \430 , \431 , \432 , \433_nG137 , \434 ,
         \435_nG139 , \436 , \437 , \438 , \439_nG12c , \440 , \441_nG12e , \442 , \443 , \444 ,
         \445_nG104 , \446 , \447_nG106 , \448 , \449 , \450 , \451 , \452 , \453 , \454 ,
         \455 , \456 , \457 , \458 , \459 , \460 , \461 , \462 , \463 , \464 ,
         \465 , \466 , \467 , \468 , \469 , \470 , \471 , \472 , \473 , \474 ,
         \475 , \476 , \477 , \478 , \479 , \480 , \481 , \482 , \483 , \484 ,
         \485 , \486 , \487 , \488 , \489 , \490 , \491 , \492 , \493 , \494 ,
         \495 , \496 , \497 , \498 , \499 , \500 , \501 , \502 , \503 , \504 ,
         \505 , \506 , \507 , \508 , \509 , \510 , \511 , \512 , \513 , \514 ,
         \515 , \516 , \517 , \518 , \519 , \520 , \521 , \522 , \523 , \524 ,
         \525 , \526 , \527 , \528 , \529 , \530 , \531 , \532 , \533 , \534 ,
         \535 , \536 , \537 , \538 , \539 , \540 , \541 , \542 , \543 , \544_nG2da ,
         \545 , \546 , \547 , \548 , \549 , \550_nG2cc , \551 , \552 , \553 , \554 ,
         \555 , \556 , \557_nG2be , \558 , \559 , \560 , \561 , \562 , \563 , \564 ,
         \565 , \566 , \567 , \568 , \569 , \570 , \571 , \572 , \573 , \574 ,
         \575 , \576 , \577 , \578 , \579 , \580 , \581 , \582 , \583 , \584_nG2b0 ,
         \585 , \586 , \587 , \588 , \589 , \590_nG2a2 , \591 , \592 , \593 , \594 ,
         \595 , \596 , \597 , \598 , \599 , \600 , \601 , \602 , \603 , \604 ,
         \605 , \606 , \607 , \608 , \609 , \610 , \611 , \612 , \613 , \614 ,
         \615 , \616 , \617 , \618_nG294 , \619 , \620 , \621 , \622 , \623 , \624_nG286 ,
         \625 , \626 , \627 , \628 , \629 , \630 , \631 , \632 , \633 , \634_nG136 ,
         \635 , \636 , \637 , \638 , \639 , \640 , \641 , \642 , \643 , \644 ,
         \645 , \646 , \647 , \648 , \649 , \650 , \651 , \652 , \653 , \654 ,
         \655 , \656 , \657 , \658 , \659 , \660 , \661 , \662 , \663 , \664 ,
         \665 , \666 , \667 , \668 , \669 , \670_nG12b , \671 , \672 , \673 , \674 ,
         \675 , \676 , \677 , \678 , \679 , \680 , \681 , \682 , \683 , \684 ,
         \685 , \686_nG152 , \687 , \688 , \689 , \690 , \691 , \692_nG144 , \693 , \694 ,
         \695 , \696 , \697 , \698 , \699 , \700 , \701 , \702 , \703 , \704 ,
         \705 , \706 , \707 , \708 , \709 , \710 , \711 , \712 , \713 , \714_nG16e ,
         \715 , \716 , \717 , \718 , \719 , \720_nG160 , \721 , \722 , \723 , \724 ,
         \725 , \726 , \727 , \728 , \729 , \730 , \731 , \732 , \733 , \734 ,
         \735 , \736 , \737 , \738 , \739_nG18a , \740 , \741 , \742 , \743 , \744 ,
         \745_nG17c , \746 , \747 , \748 , \749 , \750 , \751 , \752 , \753 , \754 ,
         \755 , \756 , \757 , \758 , \759 , \760 , \761 , \762 , \763 , \764 ,
         \765_nG1a6 , \766 , \767 , \768 , \769 , \770 , \771_nG198 , \772 , \773 , \774 ,
         \775 , \776 , \777 , \778 , \779 , \780 , \781 , \782 , \783 , \784 ,
         \785 , \786 , \787 , \788 , \789 , \790 , \791 , \792 , \793 , \794_nG1c2 ,
         \795 , \796 , \797 , \798 , \799 , \800_nG1b4 , \801 , \802 , \803 , \804 ,
         \805 , \806 , \807 , \808 , \809 , \810 , \811 , \812 , \813 , \814 ,
         \815 , \816 , \817 , \818 , \819_nG1de , \820 , \821 , \822 , \823 , \824 ,
         \825_nG1d0 , \826 , \827 , \828 , \829 , \830 , \831 , \832 , \833 , \834 ,
         \835 , \836 , \837 , \838 , \839 , \840 , \841 , \842 , \843 , \844 ,
         \845_nG1fa , \846 , \847 , \848 , \849 , \850 , \851_nG1ec , \852 , \853 , \854 ,
         \855 , \856 , \857 , \858 , \859 , \860 , \861 , \862 , \863 , \864 ,
         \865 , \866 , \867 , \868 , \869 , \870 , \871 , \872 , \873 , \874 ,
         \875 , \876_nG216 , \877 , \878 , \879 , \880 , \881 , \882_nG208 , \883 , \884 ,
         \885 , \886 , \887 , \888 , \889 , \890 , \891 , \892 , \893 , \894 ,
         \895 , \896 , \897 , \898 , \899 , \900 , \901_nG232 , \902 , \903 , \904 ,
         \905 , \906 , \907_nG224 , \908 , \909 , \910 , \911 , \912 , \913 , \914 ,
         \915 , \916 , \917 , \918 , \919 , \920 , \921 , \922 , \923 , \924 ,
         \925 , \926 , \927_nG24e , \928 , \929 , \930 , \931 , \932 , \933_nG240 , \934 ,
         \935 , \936 , \937 , \938 , \939 , \940 , \941 , \942 , \943 , \944 ,
         \945 , \946 , \947 , \948 , \949 , \950 , \951 , \952 , \953 , \954 ,
         \955_nG26a , \956 , \957 , \958 , \959 , \960 , \961_nG25c , \962 , \963 , \964 ,
         \965 , \966 , \967 , \968 , \969 , \970 , \971 , \972 , \973 , \974 ,
         \975 , \976 , \977 , \978 , \979 , \980_nG278 , \981 , \982 , \983 , \984 ,
         \985 , \986 , \987 , \988 , \989 , \990 , \991 , \992 , \993 , \994 ,
         \995 , \996 , \997 , \998 , \999 , \1000 , \1001 , \1002 , \1003 , \1004 ,
         \1005 , \1006 , \1007 , \1008 , \1009 , \1010 , \1011 , \1012 , \1013 , \1014 ,
         \1015 , \1016 , \1017 , \1018 , \1019 , \1020 , \1021 , \1022 , \1023 , \1024 ,
         \1025 , \1026 , \1027 , \1028 , \1029 , \1030 , \1031 , \1032 , \1033 , \1034 ,
         \1035 , \1036 , \1037 , \1038 , \1039 , \1040 , \1041 , \1042 , \1043 , \1044 ,
         \1045 , \1046 , \1047 , \1048 , \1049 , \1050 , \1051 , \1052 , \1053 , \1054 ,
         \1055 , \1056 , \1057 , \1058 , \1059 , \1060 , \1061 , \1062 , \1063 , \1064 ,
         \1065 , \1066 , \1067 , \1068 , \1069 , \1070 , \1071 , \1072 , \1073 , \1074 ,
         \1075 , \1076 , \1077 , \1078 , \1079 , \1080 , \1081 , \1082 , \1083 , \1084 ,
         \1085 , \1086 , \1087 , \1088 , \1089 , \1090 , \1091 , \1092 , \1093 , \1094 ,
         \1095 , \1096 , \1097 , \1098 , \1099 , \1100 , \1101 , \1102 , \1103 , \1104 ,
         \1105 , \1106 , \1107 , \1108 , \1109 , \1110 , \1111 , \1112 , \1113 , \1114 ,
         \1115 , \1116 , \1117 , \1118 , \1119 , \1120 , \1121 , \1122 , \1123 , \1124 ,
         \1125 , \1126 , \1127 , \1128 , \1129 , \1130 , \1131 , \1132 , \1133 , \1134 ,
         \1135 , \1136 , \1137 , \1138 , \1139 , \1140 , \1141 , \1142 , \1143 , \1144 ,
         \1145 , \1146 , \1147 , \1148 , \1149 , \1150 , \1151 , \1152 , \1153 , \1154 ,
         \1155 , \1156 , \1157 , \1158 , \1159 , \1160 , \1161 , \1162 , \1163 , \1164 ,
         \1165 , \1166 , \1167 , \1168 , \1169 , \1170 , \1171 , \1172 , \1173 , \1174 ,
         \1175 , \1176 , \1177 , \1178 , \1179 , \1180 , \1181 , \1182 , \1183 , \1184 ,
         \1185 , \1186 , \1187 , \1188 , \1189 , \1190 , \1191 , \1192 , \1193 , \1194 ,
         \1195 , \1196 , \1197 , \1198 , \1199 , \1200 , \1201 , \1202 , \1203 , \1204 ,
         \1205 , \1206 , \1207 , \1208 , \1209 , \1210 , \1211 , \1212 , \1213 , \1214 ,
         \1215 , \1216 , \1217 , \1218 , \1219 , \1220 , \1221 , \1222 , \1223 , \1224 ,
         \1225 , \1226 , \1227 , \1228 , \1229 , \1230 , \1231 , \1232 , \1233 , \1234 ,
         \1235 , \1236 , \1237 , \1238 , \1239 , \1240 , \1241 , \1242 , \1243 , \1244 ,
         \1245 , \1246 , \1247 , \1248 , \1249 , \1250 , \1251 , \1252 , \1253 , \1254 ,
         \1255 , \1256 , \1257 , \1258 , \1259 , \1260 , \1261 , \1262 , \1263 , \1264 ,
         \1265 , \1266 , \1267 , \1268 , \1269 , \1270 , \1271 , \1272 , \1273 , \1274 ,
         \1275 , \1276 , \1277 , \1278 , \1279 , \1280 , \1281 , \1282 , \1283 , \1284 ,
         \1285 , \1286 , \1287 , \1288 , \1289 , \1290 , \1291 , \1292 , \1293 , \1294 ,
         \1295 , \1296 , \1297 , \1298 , \1299 , \1300 , \1301 , \1302 , \1303 , \1304 ,
         \1305 , \1306 , \1307 , \1308 , \1309 , \1310 , \1311 , \1312 , \1313 , \1314 ,
         \1315 , \1316 , \1317 , \1318 , \1319 , \1320 , \1321 , \1322 , \1323 , \1324 ,
         \1325 , \1326 , \1327 , \1328 , \1329 , \1330 , \1331 , \1332 , \1333 , \1334 ,
         \1335 , \1336 , \1337 , \1338 , \1339 , \1340 , \1341 , \1342 , \1343 , \1344 ,
         \1345 , \1346 , \1347 , \1348 , \1349 , \1350 , \1351 , \1352 , \1353 , \1354 ,
         \1355 , \1356 , \1357 , \1358 , \1359 , \1360 , \1361 , \1362 , \1363 , \1364 ,
         \1365 , \1366 , \1367 , \1368 , \1369 , \1370 , \1371 , \1372 , \1373 , \1374 ,
         \1375 , \1376 , \1377 , \1378 , \1379 , \1380 , \1381 , \1382 , \1383 , \1384 ,
         \1385 , \1386 , \1387 , \1388 , \1389 , \1390 , \1391 , \1392 , \1393 , \1394 ,
         \1395 , \1396 , \1397 , \1398 , \1399 , \1400 , \1401 , \1402 , \1403 , \1404 ,
         \1405 , \1406 , \1407 , \1408 , \1409 , \1410 , \1411 , \1412 , \1413 , \1414 ,
         \1415 , \1416 , \1417 , \1418 , \1419 , \1420 , \1421 , \1422 , \1423 , \1424 ,
         \1425 , \1426 , \1427 , \1428 , \1429 , \1430 , \1431 , \1432 , \1433 , \1434 ,
         \1435 , \1436 , \1437 , \1438 , \1439 , \1440 , \1441 , \1442 , \1443 , \1444 ,
         \1445 , \1446 , \1447 , \1448 , \1449 , \1450 , \1451 , \1452 , \1453 , \1454 ,
         \1455 , \1456 , \1457 , \1458 , \1459 , \1460 , \1461 , \1462 , \1463 , \1464 ,
         \1465 , \1466 , \1467 , \1468 , \1469 , \1470 , \1471 , \1472 , \1473 , \1474 ,
         \1475 , \1476 , \1477 , \1478 , \1479 , \1480 , \1481 , \1482 , \1483 , \1484 ,
         \1485 , \1486 , \1487 , \1488 , \1489 , \1490 , \1491 , \1492 , \1493 , \1494 ,
         \1495 , \1496 , \1497 , \1498 , \1499 , \1500 , \1501 , \1502 , \1503 , \1504 ,
         \1505 , \1506 , \1507 , \1508 , \1509 , \1510 , \1511 , \1512 , \1513 , \1514 ,
         \1515 , \1516 , \1517 , \1518 , \1519 , \1520 , \1521 , \1522 , \1523 , \1524 ,
         \1525 , \1526 , \1527 , \1528 , \1529 , \1530 , \1531 , \1532 , \1533 , \1534 ,
         \1535 , \1536 , \1537 , \1538 , \1539 , \1540 , \1541 , \1542 , \1543 , \1544 ,
         \1545 , \1546 , \1547 , \1548 , \1549 , \1550 , \1551 , \1552 , \1553 , \1554 ,
         \1555 , \1556 , \1557 , \1558 , \1559 , \1560 , \1561 , \1562 , \1563 , \1564 ,
         \1565 , \1566 , \1567 , \1568 , \1569 , \1570 , \1571 , \1572 , \1573 , \1574 ,
         \1575 , \1576 , \1577 , \1578 , \1579 , \1580 , \1581 , \1582 , \1583 , \1584 ,
         \1585 , \1586 , \1587 , \1588 , \1589 , \1590 , \1591 , \1592 , \1593 , \1594 ,
         \1595 , \1596 , \1597 , \1598 , \1599 , \1600 , \1601 , \1602 , \1603 , \1604 ,
         \1605 , \1606 , \1607 , \1608 , \1609 , \1610 , \1611 , \1612 , \1613 , \1614 ,
         \1615 , \1616 , \1617 , \1618 , \1619 , \1620 , \1621 , \1622 , \1623 , \1624 ,
         \1625 , \1626 , \1627 , \1628 , \1629 , \1630 , \1631 , \1632 , \1633 , \1634 ,
         \1635 , \1636 , \1637 , \1638 , \1639 , \1640 , \1641 , \1642 , \1643 , \1644 ,
         \1645 , \1646 , \1647 , \1648 , \1649 , \1650 , \1651 , \1652 , \1653 , \1654 ,
         \1655 , \1656 , \1657 , \1658 , \1659 , \1660 , \1661 , \1662 , \1663 , \1664 ,
         \1665 , \1666 , \1667 , \1668 , \1669 , \1670 , \1671 , \1672 , \1673 , \1674 ,
         \1675 , \1676 , \1677 , \1678 , \1679 , \1680 , \1681 , \1682 , \1683 , \1684 ,
         \1685 , \1686 , \1687 , \1688 , \1689 , \1690 , \1691 , \1692 , \1693 , \1694 ,
         \1695 , \1696 , \1697 , \1698 , \1699 , \1700 , \1701 , \1702 , \1703 , \1704 ,
         \1705 , \1706 , \1707 , \1708 , \1709 , \1710 , \1711 , \1712 , \1713 , \1714 ,
         \1715 , \1716 , \1717 , \1718 , \1719 , \1720 , \1721 , \1722 , \1723 , \1724 ,
         \1725 , \1726 , \1727 , \1728 , \1729 , \1730 , \1731 , \1732 , \1733 , \1734 ,
         \1735 , \1736 , \1737 , \1738 , \1739 , \1740 , \1741 , \1742 , \1743 , \1744 ,
         \1745 , \1746 , \1747 , \1748 , \1749 , \1750 , \1751 , \1752 , \1753 , \1754 ,
         \1755 , \1756 , \1757 , \1758 , \1759 , \1760 , \1761 , \1762 , \1763 , \1764 ,
         \1765 , \1766 , \1767 , \1768 , \1769 , \1770 , \1771 , \1772 , \1773 , \1774 ,
         \1775 , \1776 , \1777 , \1778 , \1779 , \1780 , \1781 , \1782 , \1783 , \1784 ,
         \1785 , \1786 , \1787 , \1788 , \1789 , \1790 , \1791 , \1792 , \1793 , \1794 ,
         \1795 , \1796 , \1797 , \1798 , \1799 , \1800 , \1801 , \1802 , \1803 , \1804 ,
         \1805 , \1806 , \1807 , \1808 , \1809 , \1810 , \1811 , \1812 , \1813 , \1814 ,
         \1815 , \1816 , \1817 , \1818 , \1819 , \1820 , \1821 , \1822 , \1823 , \1824 ,
         \1825 , \1826 , \1827 , \1828 , \1829 , \1830 , \1831 , \1832 , \1833 , \1834 ,
         \1835 , \1836 , \1837 , \1838 , \1839 , \1840 , \1841 , \1842 , \1843 , \1844 ,
         \1845 , \1846 , \1847 , \1848 , \1849 , \1850 , \1851 , \1852 , \1853 , \1854 ,
         \1855 , \1856 , \1857 , \1858 , \1859 , \1860 , \1861 , \1862 , \1863 , \1864 ,
         \1865 , \1866 , \1867 , \1868 , \1869 , \1870 , \1871 , \1872 , \1873 , \1874 ,
         \1875 , \1876 , \1877 , \1878 , \1879 , \1880 , \1881 , \1882 , \1883 , \1884 ,
         \1885 , \1886 , \1887 , \1888 , \1889 , \1890 , \1891 , \1892 , \1893 , \1894 ,
         \1895 , \1896 , \1897 , \1898 , \1899 , \1900 , \1901 , \1902 , \1903 , \1904 ,
         \1905 , \1906 , \1907 , \1908 , \1909 , \1910 , \1911 , \1912 , \1913 , \1914 ,
         \1915 , \1916 , \1917 , \1918 , \1919 , \1920 , \1921 , \1922 , \1923 , \1924 ,
         \1925 , \1926 , \1927 , \1928 , \1929 , \1930 , \1931 , \1932 , \1933 , \1934 ,
         \1935 , \1936 , \1937 , \1938 , \1939 , \1940 , \1941 , \1942 , \1943 , \1944 ,
         \1945 , \1946 , \1947 , \1948 , \1949 , \1950 , \1951 , \1952 , \1953 , \1954 ,
         \1955 , \1956 , \1957 , \1958 , \1959 , \1960 , \1961 , \1962 , \1963 , \1964 ,
         \1965 , \1966 , \1967 , \1968 , \1969 , \1970 , \1971 , \1972 , \1973 , \1974 ,
         \1975 , \1976 , \1977 , \1978 , \1979 , \1980 , \1981 , \1982 , \1983 , \1984 ,
         \1985 , \1986 , \1987 , \1988 , \1989 , \1990 , \1991 , \1992 , \1993 , \1994 ,
         \1995 , \1996 , \1997 , \1998 , \1999 , \2000 , \2001 , \2002 , \2003 , \2004 ,
         \2005 , \2006 , \2007 , \2008 , \2009 , \2010 , \2011 , \2012 , \2013 , \2014 ,
         \2015 , \2016 , \2017 , \2018 , \2019 , \2020 , \2021 , \2022 , \2023 , \2024 ,
         \2025 , \2026 , \2027 , \2028 , \2029 , \2030 , \2031 , \2032 , \2033 , \2034 ,
         \2035 , \2036 , \2037 , \2038 , \2039 , \2040 , \2041 , \2042 , \2043 , \2044 ,
         \2045 , \2046 , \2047 , \2048 , \2049 , \2050 , \2051 , \2052 , \2053 , \2054 ,
         \2055 , \2056 , \2057 , \2058 , \2059 , \2060 , \2061 , \2062 , \2063 , \2064 ,
         \2065 , \2066 , \2067 , \2068 , \2069 , \2070 , \2071 , \2072 , \2073 , \2074 ,
         \2075 , \2076 , \2077 , \2078 , \2079 , \2080 , \2081 , \2082 , \2083 , \2084 ,
         \2085 , \2086 , \2087 , \2088 , \2089 , \2090 , \2091 , \2092 , \2093 , \2094 ,
         \2095 , \2096 , \2097 , \2098 , \2099 , \2100 , \2101 , \2102 , \2103 , \2104 ,
         \2105 , \2106 , \2107 , \2108 , \2109 , \2110 , \2111 , \2112 , \2113 , \2114 ,
         \2115 , \2116 , \2117 , \2118 , \2119 , \2120 , \2121 , \2122 , \2123 , \2124 ,
         \2125 , \2126 , \2127 , \2128 , \2129 , \2130 , \2131 , \2132 , \2133 , \2134 ,
         \2135 , \2136 , \2137 , \2138 , \2139 , \2140 , \2141 , \2142 , \2143 , \2144 ,
         \2145 , \2146 , \2147 , \2148 , \2149 , \2150 , \2151 , \2152 , \2153 , \2154 ,
         \2155 , \2156 , \2157 , \2158 , \2159 , \2160 , \2161 , \2162 , \2163 , \2164 ,
         \2165 , \2166 , \2167 , \2168 , \2169 , \2170 , \2171 , \2172 , \2173 , \2174 ,
         \2175 , \2176 , \2177 , \2178 , \2179 , \2180 , \2181 , \2182 , \2183 , \2184 ,
         \2185 , \2186 , \2187 , \2188 , \2189 , \2190 , \2191 , \2192 , \2193 , \2194 ,
         \2195 , \2196 , \2197 , \2198 , \2199 , \2200 , \2201 , \2202 , \2203 , \2204 ,
         \2205 , \2206 , \2207 , \2208 , \2209 , \2210 , \2211 , \2212 , \2213 , \2214 ,
         \2215 , \2216 , \2217 , \2218 , \2219 , \2220 , \2221 , \2222 , \2223 , \2224 ,
         \2225 , \2226 , \2227 , \2228 , \2229 , \2230 , \2231 , \2232 , \2233 , \2234 ,
         \2235 , \2236 , \2237 , \2238 , \2239 , \2240 , \2241 , \2242 , \2243 , \2244 ,
         \2245 , \2246 , \2247 , \2248 , \2249 , \2250 , \2251 , \2252 , \2253 , \2254 ,
         \2255 , \2256 , \2257 , \2258 , \2259 , \2260 , \2261 , \2262 , \2263 , \2264 ,
         \2265 , \2266 , \2267 , \2268 , \2269 , \2270 , \2271 , \2272 , \2273 , \2274 ,
         \2275 , \2276 , \2277 , \2278 , \2279 , \2280 , \2281 , \2282 , \2283 , \2284 ,
         \2285 , \2286 , \2287 , \2288 , \2289 , \2290 , \2291 , \2292 , \2293 , \2294 ,
         \2295 , \2296 , \2297 , \2298 , \2299 , \2300 , \2301 , \2302 , \2303 , \2304 ,
         \2305 , \2306 , \2307 , \2308 , \2309 , \2310 , \2311 , \2312 , \2313 , \2314 ,
         \2315 , \2316 , \2317 , \2318 , \2319 , \2320 , \2321 , \2322 , \2323 , \2324 ,
         \2325 , \2326 , \2327 , \2328 , \2329 , \2330 , \2331 , \2332 , \2333 , \2334 ,
         \2335 , \2336 , \2337 , \2338 , \2339 , \2340 , \2341 , \2342 , \2343 , \2344 ,
         \2345 , \2346 , \2347 , \2348 , \2349 , \2350 , \2351 , \2352 , \2353 , \2354 ,
         \2355 , \2356 , \2357 , \2358 , \2359 , \2360 , \2361 , \2362 , \2363 , \2364 ,
         \2365 , \2366 , \2367 , \2368 , \2369 , \2370 , \2371 , \2372 , \2373 , \2374 ,
         \2375 , \2376 , \2377 , \2378 , \2379 , \2380 , \2381 , \2382 , \2383 , \2384 ,
         \2385 , \2386 , \2387 , \2388 , \2389 , \2390 , \2391 , \2392 , \2393 , \2394 ,
         \2395 , \2396 , \2397 , \2398 , \2399 , \2400 , \2401 , \2402 , \2403 , \2404 ,
         \2405 , \2406 , \2407 , \2408 , \2409 , \2410 , \2411 , \2412 , \2413 , \2414 ,
         \2415 , \2416 , \2417 , \2418 , \2419 , \2420 , \2421 , \2422 , \2423 , \2424 ,
         \2425 , \2426 , \2427 , \2428 , \2429 , \2430 , \2431 , \2432 , \2433 , \2434 ,
         \2435 , \2436 , \2437 , \2438 , \2439 , \2440 , \2441 , \2442 , \2443 , \2444 ,
         \2445 , \2446 , \2447 , \2448 , \2449 , \2450 , \2451 , \2452 , \2453 , \2454 ,
         \2455 , \2456 , \2457 , \2458 , \2459 , \2460 , \2461 , \2462 , \2463 , \2464 ,
         \2465 , \2466 , \2467 , \2468 , \2469 , \2470 , \2471 , \2472 , \2473 , \2474 ,
         \2475 , \2476 , \2477 , \2478 , \2479 , \2480 , \2481 , \2482 , \2483 , \2484 ,
         \2485 , \2486 , \2487 , \2488 , \2489 , \2490 , \2491 , \2492 , \2493 , \2494 ,
         \2495 , \2496 , \2497 , \2498 , \2499 , \2500 , \2501 , \2502 , \2503 , \2504 ,
         \2505 , \2506 , \2507 , \2508 , \2509 , \2510 , \2511 , \2512 , \2513 , \2514 ,
         \2515 , \2516 , \2517 , \2518 , \2519 , \2520 , \2521 , \2522 , \2523 , \2524 ,
         \2525 , \2526 , \2527 , \2528 , \2529 , \2530 , \2531 , \2532 , \2533 , \2534 ,
         \2535 , \2536 , \2537 , \2538 , \2539 , \2540 , \2541 , \2542 , \2543 , \2544 ,
         \2545 , \2546 , \2547 , \2548 , \2549 , \2550 , \2551 , \2552 , \2553 , \2554 ,
         \2555 , \2556 , \2557 , \2558 , \2559 , \2560 , \2561 , \2562 , \2563 , \2564 ,
         \2565 , \2566 , \2567 , \2568 , \2569 , \2570 , \2571 , \2572 , \2573 , \2574 ,
         \2575 , \2576 , \2577 , \2578 , \2579 , \2580 , \2581 , \2582 , \2583 , \2584 ,
         \2585 , \2586 , \2587 , \2588 , \2589 , \2590 , \2591 , \2592 , \2593 , \2594 ,
         \2595 , \2596 , \2597 , \2598 , \2599 , \2600 , \2601 , \2602 , \2603 , \2604 ,
         \2605 , \2606 , \2607 , \2608 , \2609 , \2610 , \2611 , \2612 , \2613 , \2614 ,
         \2615 , \2616 , \2617 , \2618 , \2619 , \2620 , \2621 , \2622 , \2623 , \2624 ,
         \2625 , \2626 , \2627 , \2628 , \2629 , \2630 , \2631 , \2632 , \2633 , \2634 ,
         \2635 , \2636 , \2637 , \2638 , \2639 , \2640 , \2641 , \2642 , \2643 , \2644 ,
         \2645 , \2646 , \2647 , \2648 , \2649 , \2650 , \2651 , \2652 , \2653 , \2654 ,
         \2655 , \2656 , \2657 , \2658 , \2659 , \2660 , \2661 , \2662 , \2663 , \2664 ,
         \2665 , \2666 , \2667 , \2668 , \2669 , \2670 , \2671 , \2672 , \2673 , \2674 ,
         \2675 , \2676 , \2677 , \2678 , \2679 , \2680 , \2681 , \2682 , \2683 , \2684 ,
         \2685 , \2686 , \2687 , \2688 , \2689 , \2690 , \2691 , \2692 , \2693 , \2694 ,
         \2695 , \2696 , \2697 , \2698 , \2699 , \2700 , \2701 , \2702 , \2703 , \2704 ,
         \2705 , \2706 , \2707 , \2708 , \2709 , \2710 , \2711 , \2712 , \2713 , \2714 ,
         \2715 , \2716 , \2717 , \2718 , \2719 , \2720 , \2721 , \2722 , \2723 , \2724 ,
         \2725 , \2726 , \2727 , \2728 , \2729 , \2730 , \2731 , \2732 , \2733 , \2734 ,
         \2735 , \2736 , \2737 , \2738 , \2739 , \2740 , \2741 , \2742 , \2743 , \2744 ,
         \2745 , \2746 , \2747 , \2748 , \2749 , \2750 , \2751 , \2752 , \2753 , \2754 ,
         \2755 , \2756 , \2757 , \2758 , \2759 , \2760 , \2761 , \2762 , \2763 , \2764 ,
         \2765 , \2766 , \2767 , \2768 , \2769 , \2770 , \2771 , \2772 , \2773 , \2774 ,
         \2775 , \2776 , \2777 , \2778 , \2779 , \2780 , \2781 , \2782 , \2783 , \2784 ,
         \2785 , \2786 , \2787 , \2788 , \2789 , \2790 , \2791 , \2792 , \2793 , \2794 ,
         \2795 , \2796 , \2797 , \2798 , \2799 , \2800 , \2801 , \2802 , \2803 , \2804 ,
         \2805 , \2806 , \2807 , \2808 , \2809 , \2810 , \2811 , \2812 , \2813 , \2814 ,
         \2815 , \2816 , \2817 , \2818 , \2819 , \2820 , \2821 , \2822 , \2823 , \2824 ,
         \2825 , \2826 , \2827 , \2828 , \2829 , \2830 , \2831 , \2832 , \2833 , \2834 ,
         \2835 , \2836 , \2837 , \2838 , \2839 , \2840 , \2841 , \2842 , \2843 , \2844 ,
         \2845 , \2846 , \2847 , \2848 , \2849 , \2850 , \2851 , \2852 , \2853 , \2854 ,
         \2855 , \2856 , \2857 , \2858 , \2859 , \2860 , \2861 , \2862 , \2863 , \2864 ,
         \2865 , \2866 , \2867 , \2868 , \2869 , \2870 , \2871 , \2872 , \2873 , \2874 ,
         \2875 , \2876 , \2877 , \2878 , \2879 , \2880 , \2881 , \2882 , \2883 , \2884 ,
         \2885 , \2886 , \2887 , \2888 , \2889 , \2890 , \2891 , \2892 , \2893 , \2894 ,
         \2895 , \2896 , \2897 , \2898 , \2899 , \2900 , \2901 , \2902 , \2903 , \2904 ,
         \2905 , \2906 , \2907 , \2908 , \2909 , \2910 , \2911 , \2912 , \2913 , \2914 ,
         \2915 , \2916 , \2917 , \2918 , \2919 , \2920 , \2921 , \2922 , \2923 , \2924 ,
         \2925 , \2926 , \2927 , \2928 , \2929 , \2930 , \2931 , \2932 , \2933 , \2934 ,
         \2935 , \2936 , \2937 , \2938 , \2939 , \2940 , \2941 , \2942 , \2943 , \2944 ,
         \2945 , \2946 , \2947 , \2948 , \2949 , \2950 , \2951 , \2952 , \2953 , \2954 ,
         \2955 , \2956 , \2957 , \2958 , \2959 , \2960 , \2961 , \2962 , \2963 , \2964 ,
         \2965 , \2966 , \2967 , \2968 , \2969 , \2970 , \2971 , \2972 , \2973 , \2974 ,
         \2975 , \2976 , \2977 , \2978 , \2979 , \2980 , \2981 , \2982 , \2983 , \2984 ,
         \2985 , \2986 , \2987 , \2988 , \2989 , \2990 , \2991 , \2992 , \2993 , \2994 ,
         \2995 , \2996 , \2997 , \2998 , \2999 , \3000 , \3001 , \3002 , \3003 , \3004 ,
         \3005 , \3006 , \3007 , \3008 , \3009 , \3010 , \3011 , \3012 , \3013 , \3014 ,
         \3015 , \3016 , \3017 , \3018 , \3019 , \3020 , \3021 , \3022 , \3023 , \3024 ,
         \3025 , \3026 , \3027 , \3028 , \3029 , \3030 , \3031 , \3032 , \3033 , \3034 ,
         \3035 , \3036 , \3037 , \3038 , \3039 , \3040 , \3041 , \3042 , \3043 , \3044 ,
         \3045 , \3046 , \3047 , \3048 , \3049 , \3050 , \3051 , \3052 , \3053 , \3054 ,
         \3055 , \3056 , \3057 , \3058 , \3059 , \3060 , \3061 , \3062 , \3063 , \3064 ,
         \3065 , \3066 , \3067 , \3068 , \3069 , \3070 , \3071 , \3072 , \3073 , \3074 ,
         \3075 , \3076 , \3077 , \3078 , \3079 , \3080 , \3081 , \3082 , \3083 , \3084 ,
         \3085 , \3086 , \3087 , \3088 , \3089 , \3090 , \3091 , \3092 , \3093 , \3094 ,
         \3095 , \3096 , \3097 , \3098 , \3099 , \3100 , \3101 , \3102 , \3103 , \3104 ,
         \3105 , \3106 , \3107 , \3108 , \3109 , \3110 , \3111 , \3112 , \3113 , \3114 ,
         \3115 , \3116 , \3117 , \3118 , \3119 , \3120 , \3121 , \3122 , \3123 , \3124 ,
         \3125 , \3126 , \3127 , \3128 , \3129 , \3130 , \3131 , \3132 , \3133 , \3134 ,
         \3135 , \3136 , \3137 , \3138 , \3139 , \3140 , \3141 , \3142 , \3143 , \3144 ,
         \3145 , \3146 , \3147 , \3148 , \3149 , \3150 , \3151 , \3152 , \3153 , \3154 ,
         \3155 , \3156 , \3157 , \3158 , \3159 , \3160 , \3161 , \3162 , \3163 , \3164 ,
         \3165 , \3166 , \3167 , \3168 , \3169 , \3170 , \3171 , \3172 , \3173 , \3174 ,
         \3175 , \3176 , \3177 , \3178 , \3179 , \3180 , \3181 , \3182 , \3183 , \3184 ,
         \3185 , \3186 , \3187 , \3188 , \3189 , \3190 , \3191 , \3192 , \3193 , \3194 ,
         \3195 , \3196 , \3197 , \3198 , \3199 , \3200 , \3201 , \3202 , \3203 , \3204 ,
         \3205 , \3206 , \3207 , \3208 , \3209 , \3210 , \3211 , \3212 , \3213 , \3214 ,
         \3215 , \3216 , \3217 , \3218 , \3219 , \3220 , \3221 , \3222 , \3223 , \3224 ,
         \3225 , \3226 , \3227 , \3228 , \3229 , \3230 , \3231 , \3232 , \3233 , \3234 ,
         \3235 , \3236 , \3237 , \3238 , \3239 , \3240 , \3241 , \3242 , \3243 , \3244 ,
         \3245 , \3246 , \3247 , \3248 , \3249 , \3250 , \3251 , \3252 , \3253 , \3254 ,
         \3255 , \3256 , \3257 , \3258 , \3259 , \3260 , \3261 , \3262 , \3263 , \3264 ,
         \3265 , \3266 , \3267 , \3268 , \3269 , \3270 , \3271 , \3272 , \3273 , \3274 ,
         \3275 , \3276 , \3277 , \3278 , \3279 , \3280 , \3281 , \3282 , \3283 , \3284 ,
         \3285 , \3286 , \3287 , \3288 , \3289 , \3290 , \3291 , \3292 , \3293 , \3294 ,
         \3295 , \3296 , \3297 , \3298 , \3299 , \3300 , \3301 , \3302 , \3303 , \3304 ,
         \3305 , \3306 , \3307 , \3308 , \3309 , \3310 , \3311 , \3312 , \3313 , \3314 ,
         \3315 , \3316 , \3317 , \3318 , \3319 , \3320 , \3321 , \3322 , \3323 , \3324 ,
         \3325 , \3326 , \3327 , \3328 , \3329 , \3330 , \3331 , \3332 , \3333 , \3334 ,
         \3335 , \3336 , \3337 , \3338 , \3339 , \3340 , \3341 , \3342 , \3343 , \3344 ,
         \3345 , \3346 , \3347 , \3348 , \3349 , \3350 , \3351 , \3352 , \3353 , \3354 ,
         \3355 , \3356 , \3357 , \3358 , \3359 , \3360 , \3361 , \3362 , \3363 , \3364 ,
         \3365 , \3366 , \3367 , \3368 , \3369 , \3370 , \3371 , \3372 , \3373 , \3374 ,
         \3375 , \3376 , \3377 , \3378 , \3379 , \3380 , \3381 , \3382 , \3383 , \3384 ,
         \3385 , \3386 , \3387 , \3388 , \3389 , \3390 , \3391 , \3392 , \3393 , \3394 ,
         \3395 , \3396 , \3397 , \3398 , \3399 , \3400 , \3401 , \3402 , \3403 , \3404 ,
         \3405 , \3406 , \3407 , \3408 , \3409 , \3410 , \3411 , \3412 , \3413 , \3414 ,
         \3415 , \3416 , \3417 , \3418 , \3419 , \3420 , \3421 , \3422 , \3423 , \3424 ,
         \3425 , \3426 , \3427 , \3428 , \3429 , \3430 , \3431 , \3432 , \3433 , \3434 ,
         \3435 , \3436 , \3437 , \3438 , \3439 , \3440 , \3441 , \3442 , \3443 , \3444 ,
         \3445 , \3446 , \3447 , \3448 , \3449 , \3450 , \3451 , \3452 , \3453 , \3454 ,
         \3455 , \3456 , \3457 , \3458 , \3459 , \3460 , \3461 , \3462 , \3463 , \3464 ,
         \3465 , \3466 , \3467 , \3468 , \3469 , \3470 , \3471 , \3472 , \3473 , \3474 ,
         \3475 , \3476 , \3477 , \3478 , \3479 , \3480 , \3481 , \3482 , \3483 , \3484 ,
         \3485 , \3486 , \3487 , \3488 , \3489 , \3490 , \3491 , \3492 , \3493 , \3494 ,
         \3495 , \3496 , \3497 , \3498 , \3499 , \3500 , \3501 , \3502 , \3503 , \3504 ,
         \3505 , \3506 , \3507 , \3508 , \3509 , \3510 , \3511 , \3512 , \3513 , \3514 ,
         \3515 , \3516 , \3517 , \3518 , \3519 , \3520 , \3521 , \3522 , \3523 , \3524 ,
         \3525 , \3526 , \3527 , \3528 , \3529 , \3530 , \3531 , \3532 , \3533 , \3534 ,
         \3535 , \3536 , \3537 , \3538 , \3539 , \3540 , \3541 , \3542 , \3543 , \3544 ,
         \3545 , \3546 , \3547 , \3548 , \3549 , \3550 , \3551 , \3552 , \3553 , \3554 ,
         \3555 , \3556 , \3557 , \3558 , \3559 , \3560 , \3561 , \3562 , \3563 , \3564 ,
         \3565 , \3566 , \3567 , \3568 , \3569 , \3570 , \3571 , \3572 , \3573 , \3574 ,
         \3575 , \3576 , \3577 , \3578 , \3579 , \3580 , \3581 , \3582 , \3583 , \3584 ,
         \3585 , \3586 , \3587 , \3588 , \3589 , \3590 , \3591 , \3592 , \3593 , \3594 ,
         \3595 , \3596 , \3597 , \3598 , \3599 , \3600 , \3601 , \3602 , \3603 , \3604 ,
         \3605 , \3606 , \3607 , \3608 , \3609 , \3610 , \3611 , \3612 , \3613 , \3614 ,
         \3615 , \3616 , \3617 , \3618 , \3619 , \3620 , \3621 , \3622 , \3623 , \3624 ,
         \3625 , \3626 , \3627 , \3628 , \3629 , \3630 , \3631 , \3632 , \3633 , \3634 ,
         \3635 , \3636 , \3637 , \3638 , \3639 , \3640 , \3641 , \3642 , \3643 , \3644 ,
         \3645 , \3646 , \3647 , \3648 , \3649 , \3650 , \3651 , \3652 , \3653 , \3654 ,
         \3655 , \3656 , \3657 , \3658 , \3659 , \3660 , \3661 , \3662 , \3663 , \3664 ,
         \3665 , \3666 , \3667 , \3668 , \3669 , \3670 , \3671 , \3672 , \3673 , \3674 ,
         \3675 , \3676 , \3677 , \3678 , \3679 , \3680 , \3681 , \3682 , \3683 , \3684 ,
         \3685 , \3686 , \3687 , \3688 , \3689 , \3690 , \3691 , \3692 , \3693 , \3694 ,
         \3695 , \3696 , \3697 , \3698 , \3699 , \3700 , \3701 , \3702 , \3703 , \3704 ,
         \3705 , \3706 , \3707 , \3708 , \3709 , \3710 , \3711 , \3712 , \3713 , \3714 ,
         \3715 , \3716 , \3717 , \3718 , \3719 , \3720 , \3721 , \3722 , \3723 , \3724 ,
         \3725 , \3726 , \3727 , \3728 , \3729 , \3730 , \3731 , \3732 , \3733 , \3734 ,
         \3735 , \3736 , \3737 , \3738 , \3739 , \3740 , \3741 , \3742 , \3743 , \3744 ,
         \3745 , \3746 , \3747 , \3748 , \3749 , \3750 , \3751 , \3752 , \3753 , \3754 ,
         \3755 , \3756 , \3757 , \3758 , \3759 , \3760 , \3761 , \3762 , \3763 , \3764 ,
         \3765 , \3766 , \3767 , \3768 , \3769 , \3770 , \3771 , \3772 , \3773 , \3774 ,
         \3775 , \3776 , \3777 , \3778 , \3779 , \3780 , \3781 , \3782 , \3783 , \3784 ,
         \3785 , \3786 , \3787 , \3788 , \3789 , \3790 , \3791 , \3792 , \3793 , \3794 ,
         \3795 , \3796 , \3797 , \3798 , \3799 , \3800 , \3801 , \3802 , \3803 , \3804 ,
         \3805 , \3806 , \3807 , \3808 , \3809 , \3810 , \3811 , \3812 , \3813 , \3814 ,
         \3815 , \3816 , \3817 , \3818 , \3819 , \3820 , \3821 , \3822 , \3823 , \3824 ,
         \3825 , \3826 , \3827 , \3828 , \3829 , \3830 , \3831 , \3832 , \3833 , \3834 ,
         \3835 , \3836 , \3837 , \3838 , \3839 , \3840 , \3841 , \3842 , \3843 , \3844 ,
         \3845 , \3846 , \3847 , \3848 , \3849 , \3850 , \3851 , \3852 , \3853 , \3854 ,
         \3855 , \3856 , \3857 , \3858 , \3859 , \3860 , \3861 , \3862 , \3863 , \3864 ,
         \3865 , \3866 , \3867 , \3868 , \3869 , \3870 , \3871 , \3872 , \3873 , \3874 ,
         \3875 , \3876 , \3877 , \3878 , \3879 , \3880 , \3881 , \3882 , \3883 , \3884 ,
         \3885 , \3886 , \3887 , \3888 , \3889 , \3890 , \3891 , \3892 , \3893 , \3894 ,
         \3895 , \3896 , \3897 , \3898 , \3899 , \3900 , \3901 , \3902 , \3903 , \3904 ,
         \3905 , \3906 , \3907 , \3908 , \3909 , \3910 , \3911 , \3912 , \3913 , \3914 ,
         \3915 , \3916 , \3917 , \3918 , \3919 , \3920 , \3921 , \3922 , \3923 , \3924 ,
         \3925 , \3926 , \3927 , \3928 , \3929 , \3930 , \3931 , \3932 , \3933 , \3934 ,
         \3935 , \3936 , \3937 , \3938 , \3939 , \3940 , \3941 , \3942 , \3943 , \3944 ,
         \3945 , \3946 , \3947 , \3948 , \3949 , \3950 , \3951 , \3952 , \3953 , \3954 ,
         \3955 , \3956 , \3957 , \3958 , \3959 , \3960 , \3961 , \3962 , \3963 , \3964 ,
         \3965 , \3966 , \3967 , \3968 , \3969 , \3970 , \3971 , \3972 , \3973 , \3974 ,
         \3975 , \3976 , \3977 , \3978 , \3979 , \3980 , \3981 , \3982 , \3983 , \3984 ,
         \3985 , \3986 , \3987 , \3988 , \3989 , \3990 , \3991 , \3992 , \3993 , \3994 ,
         \3995 , \3996 , \3997 , \3998 , \3999 , \4000 , \4001 , \4002 , \4003 , \4004 ,
         \4005 , \4006 , \4007 , \4008 , \4009 , \4010 , \4011 , \4012 , \4013 , \4014 ,
         \4015 , \4016 , \4017 , \4018 , \4019 , \4020 , \4021 , \4022 , \4023 , \4024 ,
         \4025 , \4026 , \4027 , \4028 , \4029 , \4030 , \4031 , \4032 , \4033 , \4034 ,
         \4035 , \4036 , \4037 , \4038 , \4039 , \4040 , \4041 , \4042 , \4043 , \4044 ,
         \4045 , \4046 , \4047 , \4048 , \4049 , \4050 , \4051 , \4052 , \4053 , \4054 ,
         \4055 , \4056 , \4057 , \4058 , \4059 , \4060 , \4061 , \4062 , \4063 , \4064 ,
         \4065 , \4066 , \4067 , \4068 , \4069 , \4070 , \4071 , \4072 , \4073 , \4074 ,
         \4075 , \4076 , \4077 , \4078 , \4079 , \4080 , \4081 , \4082 , \4083 , \4084 ,
         \4085 , \4086 , \4087 , \4088 , \4089 , \4090 , \4091 , \4092 , \4093 , \4094 ,
         \4095 , \4096 , \4097 , \4098 , \4099 , \4100 , \4101 , \4102 , \4103 , \4104 ,
         \4105 , \4106 , \4107 , \4108 , \4109 , \4110 , \4111 , \4112 , \4113 , \4114 ,
         \4115 , \4116 , \4117 , \4118 , \4119 , \4120 , \4121 , \4122 , \4123 , \4124 ,
         \4125 , \4126 , \4127 , \4128 , \4129 , \4130 , \4131 , \4132 , \4133 , \4134 ,
         \4135 , \4136 , \4137 , \4138 , \4139 , \4140 , \4141 , \4142 , \4143 , \4144 ,
         \4145 , \4146 , \4147 , \4148 , \4149 , \4150 , \4151 , \4152 , \4153 , \4154 ,
         \4155 , \4156 , \4157 , \4158 , \4159 , \4160 , \4161 , \4162 , \4163 , \4164 ,
         \4165 , \4166 , \4167 , \4168 , \4169 , \4170 , \4171 , \4172 , \4173 , \4174 ,
         \4175 , \4176 , \4177 , \4178 , \4179 , \4180 , \4181 , \4182 , \4183 , \4184 ,
         \4185 , \4186 , \4187 , \4188 , \4189 , \4190 , \4191 , \4192 , \4193 , \4194 ,
         \4195 , \4196 , \4197 , \4198 , \4199 , \4200 , \4201 , \4202 , \4203 , \4204 ,
         \4205 , \4206 , \4207 , \4208 , \4209 , \4210 , \4211 , \4212 , \4213 , \4214 ,
         \4215 , \4216 , \4217 , \4218 , \4219 , \4220 , \4221 , \4222 , \4223 , \4224 ,
         \4225 , \4226 , \4227 , \4228 , \4229 , \4230 , \4231 , \4232 , \4233 , \4234 ,
         \4235 , \4236 , \4237 , \4238 , \4239 , \4240 , \4241 , \4242 , \4243 , \4244 ,
         \4245 , \4246 , \4247 , \4248 , \4249 , \4250 , \4251 , \4252 , \4253 , \4254 ,
         \4255 , \4256 , \4257 , \4258 , \4259 , \4260 , \4261 , \4262 , \4263 , \4264 ,
         \4265 , \4266 , \4267 , \4268 , \4269 , \4270 , \4271 , \4272 , \4273 , \4274 ,
         \4275 , \4276 , \4277 , \4278 , \4279 , \4280 , \4281 , \4282 , \4283 , \4284 ,
         \4285 , \4286 , \4287 , \4288 , \4289 , \4290 , \4291 , \4292 , \4293 , \4294 ,
         \4295 , \4296 , \4297 , \4298 , \4299 , \4300 , \4301 , \4302 , \4303 , \4304 ,
         \4305 , \4306 , \4307 , \4308 , \4309 , \4310 , \4311 , \4312 , \4313 , \4314 ,
         \4315 , \4316 , \4317 , \4318 , \4319 , \4320 , \4321 , \4322 , \4323 , \4324 ,
         \4325 , \4326 , \4327 , \4328 , \4329 , \4330 , \4331 , \4332 , \4333 , \4334 ,
         \4335 , \4336 , \4337 , \4338 , \4339 , \4340 , \4341 , \4342 , \4343 , \4344 ,
         \4345 , \4346 , \4347 , \4348 , \4349 , \4350 , \4351 , \4352 , \4353 , \4354 ,
         \4355 , \4356 , \4357 , \4358 , \4359 , \4360 , \4361 , \4362 , \4363 , \4364 ,
         \4365 , \4366 , \4367 , \4368 , \4369 , \4370 , \4371 , \4372 , \4373 , \4374 ,
         \4375 , \4376 , \4377 , \4378 , \4379 , \4380 , \4381 , \4382 , \4383 , \4384 ,
         \4385 , \4386 , \4387 , \4388 , \4389 , \4390 , \4391 , \4392 , \4393 , \4394 ,
         \4395 , \4396 , \4397 , \4398 , \4399 , \4400 , \4401 , \4402 , \4403 , \4404 ,
         \4405 , \4406 , \4407 , \4408 , \4409 , \4410 , \4411 , \4412 , \4413 , \4414 ,
         \4415 , \4416 , \4417 , \4418 , \4419 , \4420 , \4421 , \4422 , \4423 , \4424 ,
         \4425 , \4426 , \4427 , \4428 , \4429 , \4430 , \4431 , \4432 , \4433 , \4434 ,
         \4435 , \4436 , \4437 , \4438 , \4439 , \4440 , \4441 , \4442 , \4443 , \4444 ,
         \4445 , \4446 , \4447 , \4448 , \4449 , \4450 , \4451 , \4452 , \4453 , \4454 ,
         \4455 , \4456 , \4457 , \4458 , \4459 , \4460 , \4461 , \4462 , \4463 , \4464 ,
         \4465 , \4466 , \4467 , \4468 , \4469 , \4470 , \4471 , \4472 , \4473 , \4474 ,
         \4475 , \4476 , \4477 , \4478 , \4479 , \4480 , \4481 , \4482 , \4483 , \4484 ,
         \4485 , \4486 , \4487 , \4488 , \4489 , \4490 , \4491 , \4492 , \4493 , \4494 ,
         \4495 , \4496 , \4497 , \4498 , \4499 , \4500 , \4501 , \4502 , \4503 , \4504 ,
         \4505 , \4506 , \4507 , \4508 , \4509 , \4510 , \4511 , \4512 , \4513 , \4514 ,
         \4515 , \4516 , \4517 , \4518 , \4519 , \4520 , \4521 , \4522 , \4523 , \4524 ,
         \4525 , \4526 , \4527 , \4528 , \4529 , \4530 , \4531 , \4532 , \4533 , \4534 ,
         \4535 , \4536 , \4537 , \4538 , \4539 , \4540 , \4541 , \4542 , \4543 , \4544 ,
         \4545 , \4546 , \4547 , \4548 , \4549 , \4550 , \4551 , \4552 , \4553 , \4554 ,
         \4555 , \4556 , \4557 , \4558 , \4559 , \4560 , \4561 , \4562 , \4563 , \4564 ,
         \4565 , \4566 , \4567 , \4568 , \4569 , \4570 , \4571 , \4572 , \4573 , \4574 ,
         \4575 , \4576 , \4577 , \4578 , \4579 , \4580 , \4581 , \4582 , \4583 , \4584 ,
         \4585 , \4586 , \4587 , \4588 , \4589 , \4590 , \4591 , \4592 , \4593 , \4594 ,
         \4595 , \4596 , \4597 , \4598 , \4599 , \4600 , \4601 , \4602 , \4603 , \4604 ,
         \4605 , \4606 , \4607 , \4608 , \4609 , \4610 , \4611 , \4612 , \4613 , \4614 ,
         \4615 , \4616 , \4617 , \4618 , \4619 , \4620 , \4621 , \4622 , \4623 , \4624 ,
         \4625 , \4626 , \4627 , \4628 , \4629 , \4630 , \4631 , \4632 , \4633 , \4634 ,
         \4635 , \4636 , \4637 , \4638 , \4639 , \4640 , \4641 , \4642 , \4643 , \4644 ,
         \4645 , \4646 , \4647 , \4648 , \4649 , \4650 , \4651 , \4652 , \4653 , \4654 ,
         \4655 , \4656 , \4657 , \4658 , \4659 , \4660 , \4661 , \4662 , \4663 , \4664 ,
         \4665 , \4666 , \4667 , \4668 , \4669 , \4670 , \4671 , \4672 , \4673 , \4674 ,
         \4675 , \4676 , \4677 , \4678 , \4679 , \4680 , \4681 , \4682 , \4683 , \4684 ,
         \4685 , \4686 , \4687 , \4688 , \4689 , \4690 , \4691 , \4692 , \4693 , \4694 ,
         \4695 , \4696 , \4697 , \4698 , \4699 , \4700 , \4701 , \4702 , \4703 , \4704 ,
         \4705 , \4706 , \4707 , \4708 , \4709 , \4710 , \4711 , \4712 , \4713 , \4714 ,
         \4715 , \4716 , \4717 , \4718 , \4719 , \4720 , \4721 , \4722 , \4723 , \4724 ,
         \4725 , \4726 , \4727 , \4728 , \4729 , \4730 , \4731 , \4732 , \4733 , \4734 ,
         \4735 , \4736 , \4737 , \4738 , \4739 , \4740 , \4741 , \4742 , \4743 , \4744 ,
         \4745 , \4746 , \4747 , \4748 , \4749 , \4750 , \4751 , \4752 , \4753 , \4754 ,
         \4755 , \4756 , \4757 , \4758 , \4759 , \4760 , \4761 , \4762 , \4763 , \4764 ,
         \4765 , \4766 , \4767 , \4768 , \4769 , \4770 , \4771 , \4772 , \4773 , \4774 ,
         \4775 , \4776 , \4777 , \4778 , \4779 , \4780 , \4781 , \4782 , \4783 , \4784 ,
         \4785 , \4786 , \4787 , \4788 , \4789 , \4790 , \4791 , \4792 , \4793 , \4794 ,
         \4795 , \4796 , \4797 , \4798 , \4799 , \4800 , \4801 , \4802 , \4803 , \4804 ,
         \4805 , \4806 , \4807 , \4808 , \4809 , \4810 , \4811 , \4812 , \4813 , \4814 ,
         \4815 , \4816 , \4817 , \4818 , \4819 , \4820 , \4821 , \4822 , \4823 , \4824 ,
         \4825 , \4826 , \4827 , \4828 , \4829 , \4830 , \4831 , \4832 , \4833 , \4834 ,
         \4835 , \4836 , \4837 , \4838 , \4839 , \4840 , \4841 , \4842 , \4843 , \4844 ,
         \4845 , \4846 , \4847 , \4848 , \4849 , \4850 , \4851 , \4852 , \4853 , \4854 ,
         \4855 , \4856 , \4857 , \4858 , \4859 , \4860 , \4861 , \4862 , \4863 , \4864 ,
         \4865 , \4866 , \4867 , \4868 , \4869 , \4870 , \4871 , \4872 , \4873 , \4874 ,
         \4875 , \4876 , \4877 , \4878 , \4879 , \4880 , \4881 , \4882 , \4883 , \4884 ,
         \4885 , \4886 , \4887 , \4888 , \4889 , \4890 , \4891 , \4892 , \4893 , \4894 ,
         \4895 , \4896 , \4897 , \4898 , \4899 , \4900 , \4901 , \4902 , \4903 , \4904 ,
         \4905 , \4906 , \4907 , \4908 , \4909 , \4910 , \4911 , \4912 , \4913 , \4914 ,
         \4915 , \4916 , \4917 , \4918 , \4919 , \4920 , \4921 , \4922 , \4923 , \4924 ,
         \4925 , \4926 , \4927 , \4928 , \4929 , \4930 , \4931 , \4932 , \4933 , \4934 ,
         \4935 , \4936 , \4937 , \4938 , \4939 , \4940 , \4941 , \4942 , \4943 , \4944 ,
         \4945 , \4946 , \4947 , \4948 , \4949 , \4950 , \4951 , \4952 , \4953 , \4954 ,
         \4955 , \4956 , \4957 , \4958 , \4959 , \4960 , \4961 , \4962 , \4963 , \4964 ,
         \4965 , \4966 , \4967 , \4968 , \4969 , \4970 , \4971 , \4972 , \4973 , \4974 ,
         \4975 , \4976 , \4977 , \4978 , \4979 , \4980 , \4981 , \4982 , \4983 , \4984 ,
         \4985 , \4986 , \4987 , \4988 , \4989 , \4990 , \4991 , \4992 , \4993 , \4994 ,
         \4995 , \4996 , \4997 , \4998 , \4999 , \5000 , \5001 , \5002 , \5003 , \5004 ,
         \5005 , \5006 , \5007 , \5008 , \5009 , \5010 , \5011 , \5012 , \5013 , \5014 ,
         \5015 , \5016 , \5017 , \5018 , \5019 , \5020 , \5021 , \5022 , \5023 , \5024 ,
         \5025 , \5026 , \5027 , \5028 , \5029 , \5030 , \5031 , \5032 , \5033 , \5034 ,
         \5035 , \5036 , \5037 , \5038 , \5039 , \5040 , \5041 , \5042 , \5043 , \5044 ,
         \5045 , \5046 , \5047 , \5048 , \5049 , \5050 , \5051 , \5052 , \5053 , \5054 ,
         \5055 , \5056 , \5057 , \5058 , \5059 , \5060 , \5061 , \5062 , \5063 , \5064 ,
         \5065 , \5066 , \5067 , \5068 , \5069 , \5070 , \5071 , \5072 , \5073 , \5074 ,
         \5075 , \5076 , \5077 , \5078 , \5079 , \5080 , \5081 , \5082 , \5083 , \5084 ,
         \5085 , \5086 , \5087 , \5088 , \5089 , \5090 , \5091 , \5092 , \5093 , \5094 ,
         \5095 , \5096 , \5097 , \5098 , \5099 , \5100 , \5101 , \5102 , \5103 , \5104 ,
         \5105 , \5106 , \5107 , \5108 , \5109 , \5110 , \5111 , \5112 , \5113 , \5114 ,
         \5115 , \5116 , \5117 , \5118 , \5119 , \5120 , \5121 , \5122 , \5123 , \5124 ,
         \5125 , \5126 , \5127 , \5128 , \5129 , \5130 , \5131 , \5132 , \5133 , \5134 ,
         \5135 , \5136 , \5137 , \5138 , \5139 , \5140 , \5141 , \5142 , \5143 , \5144 ,
         \5145 , \5146 , \5147 , \5148 , \5149 , \5150 , \5151 , \5152 , \5153 , \5154 ,
         \5155 , \5156 , \5157 , \5158 , \5159 , \5160 , \5161 , \5162 , \5163 , \5164 ,
         \5165 , \5166 , \5167 , \5168 , \5169 , \5170 , \5171 , \5172 , \5173 , \5174 ,
         \5175 , \5176 , \5177 , \5178 , \5179 , \5180 , \5181 , \5182 , \5183 , \5184 ,
         \5185 , \5186 , \5187 , \5188 , \5189 , \5190 , \5191 , \5192 , \5193 , \5194 ,
         \5195 , \5196 , \5197 , \5198 , \5199 , \5200 , \5201 , \5202 , \5203 , \5204 ,
         \5205 , \5206 , \5207 , \5208 , \5209 , \5210 , \5211 , \5212 , \5213 , \5214 ,
         \5215 , \5216 , \5217 , \5218 , \5219 , \5220 , \5221 , \5222 , \5223 , \5224 ,
         \5225 , \5226 , \5227 , \5228 , \5229 , \5230 , \5231 , \5232 , \5233 , \5234 ,
         \5235 , \5236 , \5237 , \5238 , \5239 , \5240 , \5241 , \5242 , \5243 , \5244 ,
         \5245 , \5246 , \5247 , \5248 , \5249 , \5250 , \5251 , \5252 , \5253 , \5254 ,
         \5255 , \5256 , \5257 , \5258 , \5259 , \5260 , \5261 , \5262 , \5263 , \5264 ,
         \5265 , \5266 , \5267 , \5268 , \5269 , \5270 , \5271 , \5272 , \5273 , \5274 ,
         \5275 , \5276 , \5277 , \5278 , \5279 , \5280 , \5281 , \5282 , \5283 , \5284 ,
         \5285 , \5286 , \5287 , \5288 , \5289 , \5290 , \5291 , \5292 , \5293 , \5294 ,
         \5295 , \5296 , \5297 , \5298 , \5299 , \5300 , \5301 , \5302 , \5303 , \5304 ,
         \5305 , \5306 , \5307 , \5308 , \5309 , \5310 , \5311 , \5312 , \5313 , \5314 ,
         \5315 , \5316 , \5317 , \5318 , \5319 , \5320 , \5321 , \5322 , \5323 , \5324 ,
         \5325 , \5326 , \5327 , \5328 , \5329 , \5330 , \5331 , \5332 , \5333 , \5334 ,
         \5335 , \5336 , \5337 , \5338 , \5339 , \5340 , \5341 , \5342 , \5343 , \5344 ,
         \5345 , \5346 , \5347 , \5348 , \5349 , \5350 , \5351 , \5352 , \5353 , \5354 ,
         \5355 , \5356 , \5357 , \5358 , \5359 , \5360 , \5361 , \5362 , \5363 , \5364 ,
         \5365 , \5366 , \5367 , \5368 , \5369 , \5370 , \5371 , \5372 , \5373 , \5374 ,
         \5375 , \5376 , \5377 , \5378 , \5379 , \5380 , \5381 , \5382 , \5383 , \5384 ,
         \5385 , \5386 , \5387 , \5388 , \5389 , \5390 , \5391 , \5392 , \5393 , \5394 ,
         \5395 , \5396 , \5397 , \5398 , \5399 , \5400 , \5401 , \5402 , \5403 , \5404 ,
         \5405 , \5406 , \5407 , \5408 , \5409 , \5410 , \5411 , \5412 , \5413 , \5414 ,
         \5415 , \5416 , \5417 , \5418 , \5419 , \5420 , \5421 , \5422 , \5423 , \5424 ,
         \5425 , \5426 , \5427 , \5428 , \5429 , \5430 , \5431 , \5432 , \5433 , \5434 ,
         \5435 , \5436 , \5437 , \5438 , \5439 , \5440 , \5441 , \5442 , \5443 , \5444 ,
         \5445 , \5446 , \5447 , \5448 , \5449 , \5450 , \5451 , \5452 , \5453 , \5454 ,
         \5455 , \5456 , \5457 , \5458 , \5459 , \5460 , \5461 , \5462 , \5463 , \5464 ,
         \5465 , \5466 , \5467 , \5468 , \5469 , \5470 , \5471 , \5472 , \5473 , \5474 ,
         \5475 , \5476 , \5477 , \5478 , \5479 , \5480 , \5481 , \5482 , \5483 , \5484 ,
         \5485 , \5486 , \5487 , \5488 , \5489 , \5490 , \5491 , \5492 , \5493 , \5494 ,
         \5495 , \5496 , \5497 , \5498 , \5499 , \5500 , \5501 , \5502 , \5503 , \5504 ,
         \5505 , \5506 , \5507 , \5508 , \5509 , \5510 , \5511 , \5512 , \5513 , \5514 ,
         \5515 , \5516 , \5517 , \5518 , \5519 , \5520 , \5521 , \5522 , \5523 , \5524 ,
         \5525 , \5526 , \5527 , \5528 , \5529 , \5530 , \5531 , \5532 , \5533 , \5534 ,
         \5535 , \5536 , \5537 , \5538 , \5539 , \5540 , \5541 , \5542 , \5543 , \5544 ,
         \5545 , \5546 , \5547 , \5548 , \5549 , \5550 , \5551 , \5552 , \5553 , \5554 ,
         \5555 , \5556 , \5557 , \5558 , \5559 , \5560 , \5561 , \5562 , \5563 , \5564 ,
         \5565 , \5566 , \5567 , \5568 , \5569 , \5570 , \5571 , \5572 , \5573 , \5574 ,
         \5575 , \5576 , \5577 , \5578 , \5579 , \5580 , \5581 , \5582 , \5583 , \5584 ,
         \5585 , \5586 , \5587 , \5588 , \5589 , \5590 , \5591 , \5592 , \5593 , \5594 ,
         \5595 , \5596 , \5597 , \5598 , \5599 , \5600 , \5601 , \5602 , \5603 , \5604 ,
         \5605 , \5606 , \5607 , \5608 , \5609 , \5610 , \5611 , \5612 , \5613 , \5614 ,
         \5615 , \5616 , \5617 , \5618 , \5619 , \5620 , \5621 , \5622 , \5623 , \5624 ,
         \5625 , \5626 , \5627 , \5628 , \5629 , \5630 , \5631 , \5632 , \5633 , \5634 ,
         \5635 , \5636 , \5637 , \5638 , \5639 , \5640 , \5641 , \5642 , \5643 , \5644 ,
         \5645 , \5646 , \5647 , \5648 , \5649 , \5650 , \5651 , \5652 , \5653 , \5654 ,
         \5655 , \5656 , \5657 , \5658 , \5659 , \5660 , \5661 , \5662 , \5663 , \5664 ,
         \5665 , \5666 , \5667 , \5668 , \5669 , \5670 , \5671 , \5672 , \5673 , \5674 ,
         \5675 , \5676 , \5677 , \5678 , \5679 , \5680 , \5681 , \5682 , \5683 , \5684 ,
         \5685 , \5686 , \5687 , \5688 , \5689 , \5690 , \5691 , \5692 , \5693 , \5694 ,
         \5695 , \5696 , \5697 , \5698 , \5699 , \5700 , \5701 , \5702 , \5703 , \5704 ,
         \5705 , \5706 , \5707 , \5708 , \5709 , \5710 , \5711 , \5712 , \5713 , \5714 ,
         \5715 , \5716 , \5717 , \5718 , \5719 , \5720 , \5721 , \5722 , \5723 , \5724 ,
         \5725 , \5726 , \5727 , \5728 , \5729 , \5730 , \5731 , \5732 , \5733 , \5734 ,
         \5735 , \5736 , \5737 , \5738 , \5739 , \5740 , \5741 , \5742 , \5743 , \5744 ,
         \5745 , \5746 , \5747 , \5748 , \5749 , \5750 , \5751 , \5752 , \5753 , \5754 ,
         \5755 , \5756 , \5757 , \5758 , \5759 , \5760 , \5761 , \5762 , \5763 , \5764 ,
         \5765 , \5766 , \5767 , \5768 , \5769 , \5770 , \5771 , \5772 , \5773 , \5774 ,
         \5775 , \5776 , \5777 , \5778 , \5779 , \5780 , \5781 , \5782 , \5783 , \5784 ,
         \5785 , \5786 , \5787 , \5788 , \5789 , \5790 , \5791 , \5792 , \5793 , \5794 ,
         \5795 , \5796 , \5797 , \5798 , \5799 , \5800 , \5801 , \5802 , \5803 , \5804 ,
         \5805 , \5806 , \5807 , \5808 , \5809 , \5810 , \5811 , \5812 , \5813 , \5814 ,
         \5815 , \5816 , \5817 , \5818 , \5819 , \5820 , \5821 , \5822 , \5823 , \5824 ,
         \5825 , \5826 , \5827 , \5828 , \5829 , \5830 , \5831 , \5832 , \5833 , \5834 ,
         \5835 , \5836 , \5837 , \5838 , \5839 , \5840 , \5841 , \5842 , \5843 , \5844 ,
         \5845 , \5846 , \5847 , \5848 , \5849 , \5850 , \5851 , \5852 , \5853 , \5854 ,
         \5855 , \5856 , \5857 , \5858 , \5859 , \5860 , \5861 , \5862 , \5863 , \5864 ,
         \5865 , \5866 , \5867 , \5868 , \5869 , \5870 , \5871 , \5872 , \5873 , \5874 ,
         \5875 , \5876 , \5877 , \5878 , \5879 , \5880 , \5881 , \5882 , \5883 , \5884 ,
         \5885 , \5886 , \5887 , \5888 , \5889 , \5890 , \5891 , \5892 , \5893 , \5894 ,
         \5895 , \5896 , \5897 , \5898 , \5899 , \5900 , \5901 , \5902 , \5903 , \5904 ,
         \5905 , \5906 , \5907 , \5908 , \5909 , \5910 , \5911 , \5912 , \5913 , \5914 ,
         \5915 , \5916 , \5917 , \5918 , \5919 , \5920 , \5921 , \5922 , \5923 , \5924 ,
         \5925 , \5926 , \5927 , \5928 , \5929 , \5930 , \5931 , \5932 , \5933 , \5934 ,
         \5935 , \5936 , \5937 , \5938 , \5939 , \5940 , \5941 , \5942 , \5943 , \5944 ,
         \5945 , \5946 , \5947 , \5948 , \5949 , \5950 , \5951 , \5952 , \5953 , \5954 ,
         \5955 , \5956 , \5957 , \5958 , \5959 , \5960 , \5961 , \5962 , \5963 , \5964 ,
         \5965 , \5966 , \5967 , \5968 , \5969 , \5970 , \5971 , \5972 , \5973 , \5974 ,
         \5975 , \5976 , \5977 , \5978 , \5979 , \5980 , \5981 , \5982 , \5983 , \5984 ,
         \5985 , \5986 , \5987 , \5988 , \5989 , \5990 , \5991 , \5992 , \5993 , \5994 ,
         \5995 , \5996 , \5997 , \5998 , \5999 , \6000 , \6001 , \6002 , \6003 , \6004 ,
         \6005 , \6006 , \6007 , \6008 , \6009 , \6010 , \6011 , \6012 , \6013 , \6014 ,
         \6015 , \6016 , \6017 , \6018 , \6019 , \6020 , \6021 , \6022 , \6023 , \6024 ,
         \6025 , \6026 , \6027 , \6028 , \6029 , \6030 , \6031 , \6032 , \6033 , \6034 ,
         \6035 , \6036 , \6037 , \6038 , \6039 , \6040 , \6041 , \6042 , \6043 , \6044 ,
         \6045 , \6046 , \6047 , \6048 , \6049 , \6050 , \6051 , \6052 , \6053 , \6054 ,
         \6055 , \6056 , \6057 , \6058 , \6059 , \6060 , \6061 , \6062 , \6063 , \6064 ,
         \6065 , \6066 , \6067 , \6068 , \6069 , \6070 , \6071 , \6072 , \6073 , \6074 ,
         \6075 , \6076 , \6077 , \6078 , \6079 , \6080 , \6081 , \6082 , \6083 , \6084 ,
         \6085 , \6086 , \6087 , \6088 , \6089 , \6090 , \6091 , \6092 , \6093 , \6094 ,
         \6095 , \6096 , \6097 , \6098 , \6099 , \6100 , \6101 , \6102 , \6103 , \6104 ,
         \6105 , \6106 , \6107 , \6108 , \6109 , \6110 , \6111 , \6112 , \6113 , \6114 ,
         \6115 , \6116 , \6117 , \6118 , \6119 , \6120 , \6121 , \6122 , \6123 , \6124 ,
         \6125 , \6126 , \6127 , \6128 , \6129 , \6130 , \6131 , \6132 , \6133 , \6134 ,
         \6135 , \6136 , \6137 , \6138 , \6139 , \6140 , \6141 , \6142 , \6143 , \6144 ,
         \6145 , \6146 , \6147 , \6148 , \6149 , \6150 , \6151 , \6152 , \6153 , \6154 ,
         \6155 , \6156 , \6157 , \6158 , \6159 , \6160 , \6161 , \6162 , \6163 , \6164 ,
         \6165 , \6166 , \6167 , \6168 , \6169 , \6170 , \6171 , \6172 , \6173 , \6174 ,
         \6175 , \6176 , \6177 , \6178 , \6179 , \6180 , \6181 , \6182 , \6183 , \6184 ,
         \6185 , \6186 , \6187 , \6188 , \6189 , \6190 , \6191 , \6192 , \6193 , \6194 ,
         \6195 , \6196 , \6197 , \6198 , \6199 , \6200 , \6201 , \6202 , \6203 , \6204 ,
         \6205 , \6206 , \6207 , \6208 , \6209 , \6210 , \6211 , \6212 , \6213 , \6214 ,
         \6215 , \6216 , \6217 , \6218 , \6219 , \6220 , \6221 , \6222 , \6223 , \6224 ,
         \6225 , \6226 , \6227 , \6228 , \6229 , \6230 , \6231 , \6232 , \6233 , \6234 ,
         \6235 , \6236 , \6237 , \6238 , \6239 , \6240 , \6241 , \6242 , \6243 , \6244 ,
         \6245 , \6246 , \6247 , \6248 , \6249 , \6250 , \6251 , \6252 , \6253 , \6254 ,
         \6255 , \6256 , \6257 , \6258 , \6259 , \6260 , \6261 , \6262 , \6263 , \6264 ,
         \6265 , \6266 , \6267 , \6268 , \6269 , \6270 , \6271 , \6272 , \6273 , \6274 ,
         \6275 , \6276 , \6277 , \6278 , \6279 , \6280 , \6281 , \6282 , \6283 , \6284 ,
         \6285 , \6286 , \6287 , \6288 , \6289 , \6290 , \6291 , \6292 , \6293 , \6294 ,
         \6295 , \6296 , \6297 , \6298 , \6299 , \6300 , \6301 , \6302 , \6303 , \6304 ,
         \6305 , \6306 , \6307 , \6308 , \6309 , \6310 , \6311 , \6312 , \6313 , \6314 ,
         \6315 , \6316 , \6317 , \6318 , \6319 , \6320 , \6321 , \6322 , \6323 , \6324 ,
         \6325 , \6326 , \6327 , \6328 , \6329 , \6330 , \6331 , \6332_nG18bf , \6333 , \6334 ,
         \6335 , \6336 , \6337 , \6338 , \6339 , \6340 , \6341 , \6342 , \6343 , \6344 ,
         \6345 , \6346 , \6347 , \6348 , \6349 , \6350 , \6351 , \6352 , \6353 , \6354 ,
         \6355 , \6356 , \6357 , \6358 , \6359 , \6360 , \6361 , \6362 , \6363 , \6364 ,
         \6365 , \6366 , \6367 , \6368 , \6369 , \6370 , \6371 , \6372 , \6373 , \6374 ,
         \6375 , \6376 , \6377 , \6378 , \6379 , \6380 , \6381 , \6382 , \6383 , \6384 ,
         \6385 , \6386 , \6387 , \6388 , \6389 , \6390 , \6391 , \6392 , \6393 , \6394 ,
         \6395 , \6396 , \6397 , \6398 , \6399 , \6400 , \6401 , \6402 , \6403 , \6404 ,
         \6405 , \6406 , \6407 , \6408 , \6409 , \6410 , \6411 , \6412 , \6413 , \6414 ,
         \6415 , \6416 , \6417 , \6418 , \6419 , \6420 , \6421 , \6422 , \6423 , \6424 ,
         \6425 , \6426 , \6427 , \6428 , \6429 , \6430 , \6431 , \6432 , \6433 , \6434 ,
         \6435 , \6436 , \6437 , \6438 , \6439 , \6440 , \6441 , \6442 , \6443 , \6444 ,
         \6445 , \6446 , \6447 , \6448 , \6449 , \6450 , \6451 , \6452 , \6453 , \6454 ,
         \6455 , \6456 , \6457 , \6458 , \6459 , \6460 , \6461 , \6462 , \6463 , \6464 ,
         \6465 , \6466 , \6467 , \6468 , \6469 , \6470 , \6471 , \6472 , \6473 , \6474 ,
         \6475 , \6476 , \6477 , \6478 , \6479 , \6480 , \6481 , \6482 , \6483 , \6484 ,
         \6485 , \6486 , \6487 , \6488 , \6489 , \6490 , \6491 , \6492 , \6493 , \6494 ,
         \6495 , \6496 , \6497 , \6498 , \6499 , \6500 , \6501 , \6502 , \6503 , \6504 ,
         \6505 , \6506 , \6507 , \6508 , \6509 , \6510 , \6511 , \6512 , \6513 , \6514_nG1974 ,
         \6515 , \6516 , \6517 , \6518 , \6519 , \6520 , \6521 , \6522 , \6523 , \6524 ,
         \6525 , \6526 , \6527 , \6528 , \6529 , \6530 , \6531 , \6532 , \6533 , \6534 ,
         \6535 , \6536 , \6537 , \6538 , \6539 , \6540 , \6541 , \6542 , \6543 , \6544 ,
         \6545 , \6546 , \6547 , \6548 , \6549 , \6550 , \6551 , \6552 , \6553 , \6554 ,
         \6555 , \6556 , \6557 , \6558 , \6559 , \6560 , \6561 , \6562 , \6563 , \6564 ,
         \6565 , \6566 , \6567 , \6568 , \6569 , \6570 , \6571 , \6572 , \6573 , \6574 ,
         \6575 , \6576 , \6577 , \6578 , \6579 , \6580 , \6581 , \6582 , \6583 , \6584 ,
         \6585 , \6586 , \6587 , \6588 , \6589 , \6590 , \6591 , \6592 , \6593 , \6594 ,
         \6595 , \6596 , \6597 , \6598 , \6599 , \6600 , \6601 , \6602 , \6603 , \6604_nG19cd ,
         \6605 , \6606 , \6607 , \6608 , \6609 , \6610 , \6611 , \6612 , \6613 , \6614 ,
         \6615 , \6616 , \6617 , \6618 , \6619 , \6620 , \6621 , \6622 , \6623 , \6624 ,
         \6625 , \6626 , \6627 , \6628 , \6629 , \6630 , \6631 , \6632 , \6633 , \6634 ,
         \6635 , \6636 , \6637 , \6638 , \6639 , \6640 , \6641 , \6642 , \6643 , \6644 ,
         \6645 , \6646 , \6647 , \6648 , \6649 , \6650 , \6651 , \6652 , \6653 , \6654 ,
         \6655 , \6656 , \6657 , \6658 , \6659 , \6660 , \6661 , \6662 , \6663 , \6664 ,
         \6665 , \6666 , \6667 , \6668 , \6669 , \6670 , \6671 , \6672 , \6673 , \6674 ,
         \6675 , \6676 , \6677 , \6678 , \6679 , \6680 , \6681 , \6682 , \6683 , \6684 ,
         \6685 , \6686 , \6687 , \6688 , \6689 , \6690 , \6691 , \6692 , \6693 , \6694 ,
         \6695_nG1a27 , \6696 , \6697 , \6698 , \6699 , \6700 , \6701 , \6702 , \6703 , \6704 ,
         \6705 , \6706 , \6707 , \6708 , \6709 , \6710 , \6711 , \6712 , \6713 , \6714 ,
         \6715 , \6716 , \6717 , \6718 , \6719 , \6720 , \6721 , \6722 , \6723 , \6724 ,
         \6725 , \6726 , \6727 , \6728 , \6729 , \6730 , \6731 , \6732 , \6733 , \6734 ,
         \6735 , \6736 , \6737 , \6738 , \6739 , \6740_nG1a53 , \6741 , \6742 , \6743 , \6744 ,
         \6745 , \6746 , \6747 , \6748 , \6749 , \6750 , \6751 , \6752 , \6753 , \6754 ,
         \6755 , \6756 , \6757 , \6758 , \6759 , \6760 , \6761 , \6762 , \6763 , \6764 ,
         \6765 , \6766 , \6767 , \6768 , \6769 , \6770 , \6771 , \6772 , \6773 , \6774 ,
         \6775 , \6776 , \6777 , \6778 , \6779 , \6780 , \6781 , \6782 , \6783 , \6784 ,
         \6785_nG1a7f , \6786 , \6787 , \6788 , \6789 , \6790 , \6791 , \6792 , \6793 , \6794 ,
         \6795 , \6796 , \6797 , \6798 , \6799 , \6800 , \6801 , \6802 , \6803 , \6804 ,
         \6805 , \6806 , \6807 , \6808 , \6809 , \6810 , \6811 , \6812 , \6813 , \6814 ,
         \6815 , \6816 , \6817 , \6818 , \6819 , \6820 , \6821 , \6822 , \6823 , \6824 ,
         \6825 , \6826 , \6827 , \6828_nG1aa9 , \6829 , \6830 , \6831 , \6832 , \6833 , \6834 ,
         \6835 , \6836 , \6837 , \6838 , \6839 , \6840 , \6841 , \6842 , \6843 , \6844 ,
         \6845 , \6846 , \6847 , \6848 , \6849 , \6850 , \6851 , \6852 , \6853 , \6854 ,
         \6855 , \6856 , \6857 , \6858 , \6859 , \6860 , \6861 , \6862 , \6863 , \6864 ,
         \6865 , \6866 , \6867 , \6868 , \6869 , \6870 , \6871_nG1ad3 , \6872 , \6873 , \6874 ,
         \6875 , \6876 , \6877 , \6878 , \6879 , \6880 , \6881 , \6882 , \6883 , \6884 ,
         \6885 , \6886 , \6887 , \6888 , \6889 , \6890 , \6891 , \6892 , \6893 , \6894_nG1ae9 ,
         \6895 , \6896 , \6897 , \6898 , \6899 , \6900 , \6901 , \6902 , \6903 , \6904 ,
         \6905 , \6906 , \6907 , \6908 , \6909 , \6910 , \6911 , \6912 , \6913 , \6914 ,
         \6915 , \6916 , \6917_nG1aff , \6918 , \6919 , \6920 , \6921 , \6922 , \6923 , \6924 ,
         \6925 , \6926 , \6927 , \6928 , \6929 , \6930 , \6931 , \6932 , \6933 , \6934 ,
         \6935 , \6936 , \6937 , \6938 , \6939_nG1b14 , \6940 , \6941 , \6942 , \6943 , \6944 ,
         \6945 , \6946 , \6947 , \6948 , \6949 , \6950 , \6951 , \6952 , \6953 , \6954 ,
         \6955 , \6956 , \6957 , \6958 , \6959 , \6960 , \6961_nG1b29 , \6962 , \6963 , \6964 ,
         \6965 , \6966 , \6967 , \6968 , \6969 , \6970 , \6971 , \6972 , \6973 , \6974 ,
         \6975 , \6976 , \6977 , \6978 , \6979 , \6980 , \6981 , \6982 , \6983_nG1b3e , \6984 ,
         \6985 , \6986 , \6987 , \6988 , \6989 , \6990 , \6991 , \6992 , \6993 , \6994 ,
         \6995 , \6996 , \6997 , \6998 , \6999 , \7000 , \7001 , \7002 , \7003 , \7004 ,
         \7005_nG1b53 , \7006 , \7007 , \7008 , \7009 , \7010 , \7011 , \7012 , \7013 , \7014 ,
         \7015 , \7016 , \7017 , \7018 , \7019 , \7020 , \7021 , \7022 , \7023 , \7024 ,
         \7025_nG1b66 , \7026 , \7027 , \7028 , \7029 , \7030 , \7031 , \7032 , \7033 , \7034 ,
         \7035 , \7036 , \7037 , \7038 , \7039 , \7040 , \7041 , \7042 , \7043 , \7044 ,
         \7045_nG1b79 , \7046 , \7047 , \7048 , \7049 , \7050 , \7051 , \7052 , \7053 , \7054 ,
         \7055 , \7056 , \7057_nG1b84 , \7058 , \7059 , \7060 , \7061 , \7062 , \7063 , \7064 ,
         \7065 , \7066 , \7067 , \7068 , \7069_nG1b8f , \7070 , \7071 , \7072 , \7073 , \7074 ,
         \7075 , \7076 , \7077 , \7078 , \7079 , \7080 , \7081_nG1b9a , \7082 , \7083 , \7084 ,
         \7085 , \7086 , \7087 , \7088 , \7089 , \7090 , \7091 , \7092 , \7093_nG1ba5 , \7094 ,
         \7095 , \7096 , \7097 , \7098 , \7099 , \7100 , \7101 , \7102 , \7103 , \7104 ,
         \7105_nG1bb0 , \7106 , \7107 , \7108 , \7109 , \7110 , \7111 , \7112 , \7113 , \7114 ,
         \7115 , \7116 , \7117_nG1bbb , \7118 , \7119 , \7120 , \7121 , \7122 , \7123 , \7124 ,
         \7125 , \7126 , \7127 , \7128_nG1bc5 , \7129 , \7130 , \7131 , \7132 , \7133 , \7134 ,
         \7135 , \7136 , \7137 , \7138 , \7139_nG1bcf , \7140 , \7141 , \7142 , \7143 , \7144 ,
         \7145 , \7146 , \7147 , \7148 , \7149 , \7150_nG1bd9 , \7151 , \7152 , \7153 , \7154 ,
         \7155 , \7156 , \7157 , \7158 , \7159 , \7160 , \7161_nG1be3 , \7162 , \7163 , \7164 ,
         \7165 , \7166 , \7167 , \7168 , \7169 , \7170 , \7171 , \7172_nG1bed , \7173 , \7174 ,
         \7175 , \7176 , \7177 , \7178 , \7179 , \7180 , \7181 , \7182 , \7183_nG1bf7 , \7184 ,
         \7185 , \7186 , \7187 , \7188 , \7189 , \7190 , \7191 , \7192 , \7193 , \7194_nG1c01 ,
         \7195 , \7196 , \7197 , \7198 , \7199 , \7200 , \7201 , \7202 , \7203 , \7204 ,
         \7205_nG1c0b , \7206 , \7207 , \7208 , \7209 , \7210 , \7211 , \7212_nG1c11 , \7213 , \7214 ,
         \7215 , \7216 , \7217 , \7218 , \7219_nG1c17 , \7220 , \7221 , \7222 , \7223 , \7224_nG1c1b ,
         \7225 , \7226 , \7227 , \7228 , \7229_nG1c1f , \7230 , \7231 , \7232 , \7233 , \7234_nG1c23 ,
         \7235 , \7236 , \7237 , \7238 , \7239_nG1c27 , \7240 , \7241 , \7242 , \7243 , \7244_nG1c2b ,
         \7245 , \7246 , \7247 , \7248 , \7249_nG1c2f , \7250 , \7251 , \7252 , \7253 , \7254_nG1c33 ,
         \7255 , \7256 , \7257 , \7258 , \7259_nG1c37 , \7260 , \7261 , \7262 , \7263 , \7264_nG1c3b ,
         \7265 , \7266 , \7267 , \7268 , \7269_nG1c3f , \7270 , \7271 , \7272 , \7273 , \7274_nG1c43 ,
         \7275 , \7276 , \7277 , \7278 , \7279_nG1c47 , \7280 , \7281 , \7282 , \7283 , \7284_nG1c4b ,
         \7285 , \7286 , \7287 , \7288 , \7289_nG1c4f , \7290 , \7291 , \7292 , \7293 , \7294_nG1c53 ,
         \7295 , \7296 , \7297 , \7298 , \7299_nG1c57 , \7300 , \7301 , \7302 , \7303 , \7304_nG1c5b ,
         \7305 , \7306 , \7307 , \7308 , \7309_nG1c5f , \7310 , \7311 , \7312 , \7313 , \7314_nG1c63 ,
         \7315 , \7316 , \7317 , \7318 , \7319_nG1c67 , \7320 , \7321 , \7322 , \7323 , \7324_nG1c6b ,
         \7325 , \7326 , \7327 , \7328 , \7329_nG1c6f , \7330 , \7331 , \7332 , \7333 , \7334_nG1c73 ,
         \7335 , \7336 , \7337 , \7338 , \7339_nG1c77 , \7340 , \7341 , \7342 , \7343 , \7344_nG1c7b ,
         \7345 , \7346 , \7347 , \7348 , \7349_nG1c7f , \7350 , \7351 , \7352 , \7353 , \7354_nG1c83 ,
         \7355 ;
buf \U$labaj758 ( R_61_7d2b4e8, \6333 );
buf \U$labaj759 ( R_62_7d2b590, \6515 );
buf \U$labaj760 ( R_63_7d2b638, \6605 );
buf \U$labaj761 ( R_64_7d2b6e0, \6696 );
buf \U$labaj762 ( R_65_7d2b788, \6741 );
buf \U$labaj763 ( R_66_7d2b830, \6786 );
buf \U$labaj764 ( R_67_7d2b8d8, \6829 );
buf \U$labaj765 ( R_68_7d2b980, \6872 );
buf \U$labaj766 ( R_69_7d2ba28, \6895 );
buf \U$labaj767 ( R_6a_7d2bad0, \6918 );
buf \U$labaj768 ( R_6b_7d2bb78, \6940 );
buf \U$labaj769 ( R_6c_7d2bc20, \6962 );
buf \U$labaj770 ( R_6d_7d2bcc8, \6984 );
buf \U$labaj771 ( R_6e_7d2bd70, \7006 );
buf \U$labaj772 ( R_6f_7d2be18, \7026 );
buf \U$labaj773 ( R_70_7d2bec0, \7046 );
buf \U$labaj774 ( R_71_7d2bf68, \7058 );
buf \U$labaj775 ( R_72_7d2c010, \7070 );
buf \U$labaj776 ( R_73_7d2c0b8, \7082 );
buf \U$labaj777 ( R_74_7d2c160, \7094 );
buf \U$labaj778 ( R_75_7d2c208, \7106 );
buf \U$labaj779 ( R_76_7d2c2b0, \7118 );
buf \U$labaj780 ( R_77_7d2c358, \7129 );
buf \U$labaj781 ( R_78_7d2c400, \7140 );
buf \U$labaj782 ( R_79_7d2c4a8, \7151 );
buf \U$labaj783 ( R_7a_7d2c550, \7162 );
buf \U$labaj784 ( R_7b_7d2c5f8, \7173 );
buf \U$labaj785 ( R_7c_7d2c6a0, \7184 );
buf \U$labaj786 ( R_7d_7d2c748, \7195 );
buf \U$labaj787 ( R_7e_7d2c7f0, \7206 );
buf \U$labaj788 ( R_7f_7d2c898, \7213 );
buf \U$labaj789 ( R_80_7d2c940, \7220 );
buf \U$labaj790 ( R_81_7d2c9e8, \7225 );
buf \U$labaj791 ( R_82_7d2ca90, \7230 );
buf \U$labaj792 ( R_83_7d2cb38, \7235 );
buf \U$labaj793 ( R_84_7d2cbe0, \7240 );
buf \U$labaj794 ( R_85_7d2cc88, \7245 );
buf \U$labaj795 ( R_86_7d2cd30, \7250 );
buf \U$labaj796 ( R_87_7d2cdd8, \7255 );
buf \U$labaj797 ( R_88_7d2ce80, \7260 );
buf \U$labaj798 ( R_89_7d2cf28, \7265 );
buf \U$labaj799 ( R_8a_7d2cfd0, \7270 );
buf \U$labaj800 ( R_8b_7d2d078, \7275 );
buf \U$labaj801 ( R_8c_7d2d120, \7280 );
buf \U$labaj802 ( R_8d_7d2d1c8, \7285 );
buf \U$labaj803 ( R_8e_7d2d270, \7290 );
buf \U$labaj804 ( R_8f_7d2d318, \7295 );
buf \U$labaj805 ( R_90_7d2d3c0, \7300 );
buf \U$labaj806 ( R_91_7d2d468, \7305 );
buf \U$labaj807 ( R_92_7d2d510, \7310 );
buf \U$labaj808 ( R_93_7d2d5b8, \7315 );
buf \U$labaj809 ( R_94_7d2d660, \7320 );
buf \U$labaj810 ( R_95_7d2d708, \7325 );
buf \U$labaj811 ( R_96_7d2d7b0, \7330 );
buf \U$labaj812 ( R_97_7d2d858, \7335 );
buf \U$labaj813 ( R_98_7d2d900, \7340 );
buf \U$labaj814 ( R_99_7d2d9a8, \7345 );
buf \U$labaj815 ( R_9a_7d2da50, \7350 );
buf \U$labaj816 ( R_9b_7d2daf8, \7355 );
buf \U$1 ( \227 , RI2b1c4342d4e0_65);
_DC g2cd ( \228_nG2cd , 1'b0 , 1'b1 );
and \U$4 ( \229 , RI2b1c4342c5e0_33, \228_nG2cd );
xor \U$5 ( \230 , RI2b1c4342d4e0_65, RI2b1c4342d558_66);
xor \U$6 ( \231 , RI2b1c4342d5d0_67, RI2b1c4342d648_68);
xor \U$7 ( \232 , \230 , \231 );
xor \U$8 ( \233 , RI2b1c4342d6c0_69, RI2b1c4342d738_70);
xor \U$9 ( \234 , RI2b1c4342d7b0_71, RI2b1c4342d828_72);
xor \U$10 ( \235 , \233 , \234 );
xor \U$11 ( \236 , \232 , \235 );
xor \U$12 ( \237 , RI2b1c4342d8a0_73, RI2b1c4342d918_74);
xor \U$13 ( \238 , RI2b1c4342d990_75, RI2b1c4342da08_76);
xor \U$14 ( \239 , \237 , \238 );
xor \U$15 ( \240 , RI2b1c4342da80_77, RI2b1c4342daf8_78);
xor \U$16 ( \241 , RI2b1c4342db70_79, RI2b1c4342dbe8_80);
xor \U$17 ( \242 , \240 , \241 );
xor \U$18 ( \243 , \239 , \242 );
xor \U$19 ( \244 , \236 , \243 );
xor \U$20 ( \245 , RI2b1c4342dc60_81, RI2b1c4342dcd8_82);
xor \U$21 ( \246 , RI2b1c4342dd50_83, RI2b1c4342ddc8_84);
xor \U$22 ( \247 , \245 , \246 );
xor \U$23 ( \248 , RI2b1c4342de40_85, RI2b1c4342deb8_86);
xor \U$24 ( \249 , RI2b1c4342df30_87, RI2b1c4342dfa8_88);
xor \U$25 ( \250 , \248 , \249 );
xor \U$26 ( \251 , \247 , \250 );
xor \U$27 ( \252 , RI2b1c4342e020_89, RI2b1c4342e098_90);
xor \U$28 ( \253 , RI2b1c4342e110_91, RI2b1c4342e188_92);
xor \U$29 ( \254 , \252 , \253 );
xor \U$30 ( \255 , RI2b1c4342e200_93, RI2b1c4342e278_94);
xor \U$31 ( \256 , RI2b1c4342e2f0_95, RI2b1c4342e368_96);
xor \U$32 ( \257 , \255 , \256 );
xor \U$33 ( \258 , \254 , \257 );
xor \U$34 ( \259 , \251 , \258 );
xor \U$35 ( \260 , \244 , \259 );
_HMUX g2cf ( \261_nG2cf , \229 , RI2b1c4342b6e0_1 , \260 );
buf \U$36 ( \262 , \261_nG2cf );
buf \U$37 ( \263 , RI2b1c4342c5e0_33);
xor \U$38 ( \264 , \262 , \263 );
_DC g2bf ( \265_nG2bf , 1'b0 , 1'b1 );
and \U$39 ( \266 , RI2b1c4342c658_34, \265_nG2bf );
_HMUX g2c1 ( \267_nG2c1 , \266 , RI2b1c4342b758_2 , \260 );
buf \U$40 ( \268 , \267_nG2c1 );
buf \U$41 ( \269 , RI2b1c4342c658_34);
and \U$42 ( \270 , \268 , \269 );
_DC g2b1 ( \271_nG2b1 , 1'b0 , 1'b1 );
and \U$43 ( \272 , RI2b1c4342c6d0_35, \271_nG2b1 );
_HMUX g2b3 ( \273_nG2b3 , \272 , RI2b1c4342b7d0_3 , \260 );
buf \U$44 ( \274 , \273_nG2b3 );
buf \U$45 ( \275 , RI2b1c4342c6d0_35);
and \U$46 ( \276 , \274 , \275 );
_DC g2a3 ( \277_nG2a3 , 1'b0 , 1'b1 );
and \U$47 ( \278 , RI2b1c4342c748_36, \277_nG2a3 );
_HMUX g2a5 ( \279_nG2a5 , \278 , RI2b1c4342b848_4 , \260 );
buf \U$48 ( \280 , \279_nG2a5 );
buf \U$49 ( \281 , RI2b1c4342c748_36);
and \U$50 ( \282 , \280 , \281 );
_DC g295 ( \283_nG295 , 1'b0 , 1'b1 );
and \U$51 ( \284 , RI2b1c4342c7c0_37, \283_nG295 );
_HMUX g297 ( \285_nG297 , \284 , RI2b1c4342b8c0_5 , \260 );
buf \U$52 ( \286 , \285_nG297 );
buf \U$53 ( \287 , RI2b1c4342c7c0_37);
and \U$54 ( \288 , \286 , \287 );
_DC g287 ( \289_nG287 , 1'b0 , 1'b1 );
and \U$55 ( \290 , RI2b1c4342c838_38, \289_nG287 );
_HMUX g289 ( \291_nG289 , \290 , RI2b1c4342b938_6 , \260 );
buf \U$56 ( \292 , \291_nG289 );
buf \U$57 ( \293 , RI2b1c4342c838_38);
and \U$58 ( \294 , \292 , \293 );
_DC g279 ( \295_nG279 , 1'b0 , 1'b1 );
and \U$59 ( \296 , RI2b1c4342c8b0_39, \295_nG279 );
_HMUX g27b ( \297_nG27b , \296 , RI2b1c4342b9b0_7 , \260 );
buf \U$60 ( \298 , \297_nG27b );
buf \U$61 ( \299 , RI2b1c4342c8b0_39);
and \U$62 ( \300 , \298 , \299 );
_DC g26b ( \301_nG26b , 1'b0 , 1'b1 );
and \U$63 ( \302 , RI2b1c4342c928_40, \301_nG26b );
_HMUX g26d ( \303_nG26d , \302 , RI2b1c4342ba28_8 , \260 );
buf \U$64 ( \304 , \303_nG26d );
buf \U$65 ( \305 , RI2b1c4342c928_40);
and \U$66 ( \306 , \304 , \305 );
_DC g25d ( \307_nG25d , 1'b0 , 1'b1 );
and \U$67 ( \308 , RI2b1c4342c9a0_41, \307_nG25d );
_HMUX g25f ( \309_nG25f , \308 , RI2b1c4342baa0_9 , \260 );
buf \U$68 ( \310 , \309_nG25f );
buf \U$69 ( \311 , RI2b1c4342c9a0_41);
and \U$70 ( \312 , \310 , \311 );
_DC g24f ( \313_nG24f , 1'b0 , 1'b1 );
and \U$71 ( \314 , RI2b1c4342ca18_42, \313_nG24f );
_HMUX g251 ( \315_nG251 , \314 , RI2b1c4342bb18_10 , \260 );
buf \U$72 ( \316 , \315_nG251 );
buf \U$73 ( \317 , RI2b1c4342ca18_42);
and \U$74 ( \318 , \316 , \317 );
_DC g241 ( \319_nG241 , 1'b0 , 1'b1 );
and \U$75 ( \320 , RI2b1c4342ca90_43, \319_nG241 );
_HMUX g243 ( \321_nG243 , \320 , RI2b1c4342bb90_11 , \260 );
buf \U$76 ( \322 , \321_nG243 );
buf \U$77 ( \323 , RI2b1c4342ca90_43);
and \U$78 ( \324 , \322 , \323 );
_DC g233 ( \325_nG233 , 1'b0 , 1'b1 );
and \U$79 ( \326 , RI2b1c4342cb08_44, \325_nG233 );
_HMUX g235 ( \327_nG235 , \326 , RI2b1c4342bc08_12 , \260 );
buf \U$80 ( \328 , \327_nG235 );
buf \U$81 ( \329 , RI2b1c4342cb08_44);
and \U$82 ( \330 , \328 , \329 );
_DC g225 ( \331_nG225 , 1'b0 , 1'b1 );
and \U$83 ( \332 , RI2b1c4342cb80_45, \331_nG225 );
_HMUX g227 ( \333_nG227 , \332 , RI2b1c4342bc80_13 , \260 );
buf \U$84 ( \334 , \333_nG227 );
buf \U$85 ( \335 , RI2b1c4342cb80_45);
and \U$86 ( \336 , \334 , \335 );
_DC g217 ( \337_nG217 , 1'b0 , 1'b1 );
and \U$87 ( \338 , RI2b1c4342cbf8_46, \337_nG217 );
_HMUX g219 ( \339_nG219 , \338 , RI2b1c4342bcf8_14 , \260 );
buf \U$88 ( \340 , \339_nG219 );
buf \U$89 ( \341 , RI2b1c4342cbf8_46);
and \U$90 ( \342 , \340 , \341 );
_DC g209 ( \343_nG209 , 1'b0 , 1'b1 );
and \U$91 ( \344 , RI2b1c4342cc70_47, \343_nG209 );
_HMUX g20b ( \345_nG20b , \344 , RI2b1c4342bd70_15 , \260 );
buf \U$92 ( \346 , \345_nG20b );
buf \U$93 ( \347 , RI2b1c4342cc70_47);
and \U$94 ( \348 , \346 , \347 );
_DC g1fb ( \349_nG1fb , 1'b0 , 1'b1 );
and \U$95 ( \350 , RI2b1c4342cce8_48, \349_nG1fb );
_HMUX g1fd ( \351_nG1fd , \350 , RI2b1c4342bde8_16 , \260 );
buf \U$96 ( \352 , \351_nG1fd );
buf \U$97 ( \353 , RI2b1c4342cce8_48);
and \U$98 ( \354 , \352 , \353 );
_DC g1ed ( \355_nG1ed , 1'b0 , 1'b1 );
and \U$99 ( \356 , RI2b1c4342cd60_49, \355_nG1ed );
_HMUX g1ef ( \357_nG1ef , \356 , RI2b1c4342be60_17 , \260 );
buf \U$100 ( \358 , \357_nG1ef );
buf \U$101 ( \359 , RI2b1c4342cd60_49);
and \U$102 ( \360 , \358 , \359 );
_DC g1df ( \361_nG1df , 1'b0 , 1'b1 );
and \U$103 ( \362 , RI2b1c4342cdd8_50, \361_nG1df );
_HMUX g1e1 ( \363_nG1e1 , \362 , RI2b1c4342bed8_18 , \260 );
buf \U$104 ( \364 , \363_nG1e1 );
buf \U$105 ( \365 , RI2b1c4342cdd8_50);
and \U$106 ( \366 , \364 , \365 );
_DC g1d1 ( \367_nG1d1 , 1'b0 , 1'b1 );
and \U$107 ( \368 , RI2b1c4342ce50_51, \367_nG1d1 );
_HMUX g1d3 ( \369_nG1d3 , \368 , RI2b1c4342bf50_19 , \260 );
buf \U$108 ( \370 , \369_nG1d3 );
buf \U$109 ( \371 , RI2b1c4342ce50_51);
and \U$110 ( \372 , \370 , \371 );
_DC g1c3 ( \373_nG1c3 , 1'b0 , 1'b1 );
and \U$111 ( \374 , RI2b1c4342cec8_52, \373_nG1c3 );
_HMUX g1c5 ( \375_nG1c5 , \374 , RI2b1c4342bfc8_20 , \260 );
buf \U$112 ( \376 , \375_nG1c5 );
buf \U$113 ( \377 , RI2b1c4342cec8_52);
and \U$114 ( \378 , \376 , \377 );
_DC g1b5 ( \379_nG1b5 , 1'b0 , 1'b1 );
and \U$115 ( \380 , RI2b1c4342cf40_53, \379_nG1b5 );
_HMUX g1b7 ( \381_nG1b7 , \380 , RI2b1c4342c040_21 , \260 );
buf \U$116 ( \382 , \381_nG1b7 );
buf \U$117 ( \383 , RI2b1c4342cf40_53);
and \U$118 ( \384 , \382 , \383 );
_DC g1a7 ( \385_nG1a7 , 1'b0 , 1'b1 );
and \U$119 ( \386 , RI2b1c4342cfb8_54, \385_nG1a7 );
_HMUX g1a9 ( \387_nG1a9 , \386 , RI2b1c4342c0b8_22 , \260 );
buf \U$120 ( \388 , \387_nG1a9 );
buf \U$121 ( \389 , RI2b1c4342cfb8_54);
and \U$122 ( \390 , \388 , \389 );
_DC g199 ( \391_nG199 , 1'b0 , 1'b1 );
and \U$123 ( \392 , RI2b1c4342d030_55, \391_nG199 );
_HMUX g19b ( \393_nG19b , \392 , RI2b1c4342c130_23 , \260 );
buf \U$124 ( \394 , \393_nG19b );
buf \U$125 ( \395 , RI2b1c4342d030_55);
and \U$126 ( \396 , \394 , \395 );
_DC g18b ( \397_nG18b , 1'b0 , 1'b1 );
and \U$127 ( \398 , RI2b1c4342d0a8_56, \397_nG18b );
_HMUX g18d ( \399_nG18d , \398 , RI2b1c4342c1a8_24 , \260 );
buf \U$128 ( \400 , \399_nG18d );
buf \U$129 ( \401 , RI2b1c4342d0a8_56);
and \U$130 ( \402 , \400 , \401 );
_DC g17d ( \403_nG17d , 1'b0 , 1'b1 );
and \U$131 ( \404 , RI2b1c4342d120_57, \403_nG17d );
_HMUX g17f ( \405_nG17f , \404 , RI2b1c4342c220_25 , \260 );
buf \U$132 ( \406 , \405_nG17f );
buf \U$133 ( \407 , RI2b1c4342d120_57);
and \U$134 ( \408 , \406 , \407 );
_DC g16f ( \409_nG16f , 1'b0 , 1'b1 );
and \U$135 ( \410 , RI2b1c4342d198_58, \409_nG16f );
_HMUX g171 ( \411_nG171 , \410 , RI2b1c4342c298_26 , \260 );
buf \U$136 ( \412 , \411_nG171 );
buf \U$137 ( \413 , RI2b1c4342d198_58);
and \U$138 ( \414 , \412 , \413 );
_DC g161 ( \415_nG161 , 1'b0 , 1'b1 );
and \U$139 ( \416 , RI2b1c4342d210_59, \415_nG161 );
_HMUX g163 ( \417_nG163 , \416 , RI2b1c4342c310_27 , \260 );
buf \U$140 ( \418 , \417_nG163 );
buf \U$141 ( \419 , RI2b1c4342d210_59);
and \U$142 ( \420 , \418 , \419 );
_DC g153 ( \421_nG153 , 1'b0 , 1'b1 );
and \U$143 ( \422 , RI2b1c4342d288_60, \421_nG153 );
_HMUX g155 ( \423_nG155 , \422 , RI2b1c4342c388_28 , \260 );
buf \U$144 ( \424 , \423_nG155 );
buf \U$145 ( \425 , RI2b1c4342d288_60);
and \U$146 ( \426 , \424 , \425 );
_DC g145 ( \427_nG145 , 1'b0 , 1'b1 );
and \U$147 ( \428 , RI2b1c4342d300_61, \427_nG145 );
_HMUX g147 ( \429_nG147 , \428 , RI2b1c4342c400_29 , \260 );
buf \U$148 ( \430 , \429_nG147 );
buf \U$149 ( \431 , RI2b1c4342d300_61);
and \U$150 ( \432 , \430 , \431 );
_DC g137 ( \433_nG137 , 1'b0 , 1'b1 );
and \U$151 ( \434 , RI2b1c4342d378_62, \433_nG137 );
_HMUX g139 ( \435_nG139 , \434 , RI2b1c4342c478_30 , \260 );
buf \U$152 ( \436 , \435_nG139 );
buf \U$153 ( \437 , RI2b1c4342d378_62);
and \U$154 ( \438 , \436 , \437 );
_DC g12c ( \439_nG12c , 1'b0 , 1'b1 );
and \U$155 ( \440 , RI2b1c4342d3f0_63, \439_nG12c );
_HMUX g12e ( \441_nG12e , \440 , RI2b1c4342c4f0_31 , \260 );
buf \U$156 ( \442 , \441_nG12e );
buf \U$157 ( \443 , RI2b1c4342d3f0_63);
and \U$158 ( \444 , \442 , \443 );
_DC g104 ( \445_nG104 , 1'b0 , 1'b1 );
and \U$159 ( \446 , RI2b1c4342d468_64, \445_nG104 );
_HMUX g106 ( \447_nG106 , \446 , RI2b1c4342c568_32 , \260 );
buf \U$160 ( \448 , \447_nG106 );
buf \U$161 ( \449 , RI2b1c4342d468_64);
and \U$162 ( \450 , \448 , \449 );
and \U$163 ( \451 , \443 , \450 );
and \U$164 ( \452 , \442 , \450 );
or \U$165 ( \453 , \444 , \451 , \452 );
and \U$166 ( \454 , \437 , \453 );
and \U$167 ( \455 , \436 , \453 );
or \U$168 ( \456 , \438 , \454 , \455 );
and \U$169 ( \457 , \431 , \456 );
and \U$170 ( \458 , \430 , \456 );
or \U$171 ( \459 , \432 , \457 , \458 );
and \U$172 ( \460 , \425 , \459 );
and \U$173 ( \461 , \424 , \459 );
or \U$174 ( \462 , \426 , \460 , \461 );
and \U$175 ( \463 , \419 , \462 );
and \U$176 ( \464 , \418 , \462 );
or \U$177 ( \465 , \420 , \463 , \464 );
and \U$178 ( \466 , \413 , \465 );
and \U$179 ( \467 , \412 , \465 );
or \U$180 ( \468 , \414 , \466 , \467 );
and \U$181 ( \469 , \407 , \468 );
and \U$182 ( \470 , \406 , \468 );
or \U$183 ( \471 , \408 , \469 , \470 );
and \U$184 ( \472 , \401 , \471 );
and \U$185 ( \473 , \400 , \471 );
or \U$186 ( \474 , \402 , \472 , \473 );
and \U$187 ( \475 , \395 , \474 );
and \U$188 ( \476 , \394 , \474 );
or \U$189 ( \477 , \396 , \475 , \476 );
and \U$190 ( \478 , \389 , \477 );
and \U$191 ( \479 , \388 , \477 );
or \U$192 ( \480 , \390 , \478 , \479 );
and \U$193 ( \481 , \383 , \480 );
and \U$194 ( \482 , \382 , \480 );
or \U$195 ( \483 , \384 , \481 , \482 );
and \U$196 ( \484 , \377 , \483 );
and \U$197 ( \485 , \376 , \483 );
or \U$198 ( \486 , \378 , \484 , \485 );
and \U$199 ( \487 , \371 , \486 );
and \U$200 ( \488 , \370 , \486 );
or \U$201 ( \489 , \372 , \487 , \488 );
and \U$202 ( \490 , \365 , \489 );
and \U$203 ( \491 , \364 , \489 );
or \U$204 ( \492 , \366 , \490 , \491 );
and \U$205 ( \493 , \359 , \492 );
and \U$206 ( \494 , \358 , \492 );
or \U$207 ( \495 , \360 , \493 , \494 );
and \U$208 ( \496 , \353 , \495 );
and \U$209 ( \497 , \352 , \495 );
or \U$210 ( \498 , \354 , \496 , \497 );
and \U$211 ( \499 , \347 , \498 );
and \U$212 ( \500 , \346 , \498 );
or \U$213 ( \501 , \348 , \499 , \500 );
and \U$214 ( \502 , \341 , \501 );
and \U$215 ( \503 , \340 , \501 );
or \U$216 ( \504 , \342 , \502 , \503 );
and \U$217 ( \505 , \335 , \504 );
and \U$218 ( \506 , \334 , \504 );
or \U$219 ( \507 , \336 , \505 , \506 );
and \U$220 ( \508 , \329 , \507 );
and \U$221 ( \509 , \328 , \507 );
or \U$222 ( \510 , \330 , \508 , \509 );
and \U$223 ( \511 , \323 , \510 );
and \U$224 ( \512 , \322 , \510 );
or \U$225 ( \513 , \324 , \511 , \512 );
and \U$226 ( \514 , \317 , \513 );
and \U$227 ( \515 , \316 , \513 );
or \U$228 ( \516 , \318 , \514 , \515 );
and \U$229 ( \517 , \311 , \516 );
and \U$230 ( \518 , \310 , \516 );
or \U$231 ( \519 , \312 , \517 , \518 );
and \U$232 ( \520 , \305 , \519 );
and \U$233 ( \521 , \304 , \519 );
or \U$234 ( \522 , \306 , \520 , \521 );
and \U$235 ( \523 , \299 , \522 );
and \U$236 ( \524 , \298 , \522 );
or \U$237 ( \525 , \300 , \523 , \524 );
and \U$238 ( \526 , \293 , \525 );
and \U$239 ( \527 , \292 , \525 );
or \U$240 ( \528 , \294 , \526 , \527 );
and \U$241 ( \529 , \287 , \528 );
and \U$242 ( \530 , \286 , \528 );
or \U$243 ( \531 , \288 , \529 , \530 );
and \U$244 ( \532 , \281 , \531 );
and \U$245 ( \533 , \280 , \531 );
or \U$246 ( \534 , \282 , \532 , \533 );
and \U$247 ( \535 , \275 , \534 );
and \U$248 ( \536 , \274 , \534 );
or \U$249 ( \537 , \276 , \535 , \536 );
and \U$250 ( \538 , \269 , \537 );
and \U$251 ( \539 , \268 , \537 );
or \U$252 ( \540 , \270 , \538 , \539 );
xor \U$253 ( \541 , \264 , \540 );
buf \U$254 ( \542 , \541 );
buf \U$255 ( \543 , RI2b1c4342b6e0_1);
and g2da ( \544_nG2da , \542 , \543 );
buf \U$256 ( \545 , \544_nG2da );
xor \U$257 ( \546 , \268 , \269 );
xor \U$258 ( \547 , \546 , \537 );
buf \U$259 ( \548 , \547 );
buf \U$260 ( \549 , RI2b1c4342b758_2);
and g2cc ( \550_nG2cc , \548 , \549 );
buf \U$261 ( \551 , \550_nG2cc );
xor \U$262 ( \552 , \545 , \551 );
xor \U$263 ( \553 , \274 , \275 );
xor \U$264 ( \554 , \553 , \534 );
buf \U$265 ( \555 , \554 );
buf \U$266 ( \556 , RI2b1c4342b7d0_3);
and g2be ( \557_nG2be , \555 , \556 );
buf \U$267 ( \558 , \557_nG2be );
xor \U$268 ( \559 , \551 , \558 );
not \U$269 ( \560 , \559 );
and \U$270 ( \561 , \552 , \560 );
and \U$271 ( \562 , \227 , \561 );
not \U$272 ( \563 , \562 );
and \U$273 ( \564 , \551 , \558 );
not \U$274 ( \565 , \564 );
and \U$275 ( \566 , \545 , \565 );
xnor \U$276 ( \567 , \563 , \566 );
buf \U$278 ( \568 , RI2b1c4342d558_66);
xor \U$281 ( \569 , 1'b0 , \545 );
and \U$282 ( \570 , \568 , \569 );
nor \U$283 ( \571 , 1'b0 , \570 );
not \U$284 ( \572 , \571 );
or \U$285 ( \573 , \567 , \572 );
not \U$286 ( \574 , \566 );
xor \U$287 ( \575 , \573 , \574 );
and \U$289 ( \576 , \227 , \569 );
nor \U$290 ( \577 , 1'b0 , \576 );
not \U$291 ( \578 , \577 );
xor \U$292 ( \579 , \575 , \578 );
xor \U$293 ( \580 , \280 , \281 );
xor \U$294 ( \581 , \580 , \531 );
buf \U$295 ( \582 , \581 );
buf \U$296 ( \583 , RI2b1c4342b848_4);
and g2b0 ( \584_nG2b0 , \582 , \583 );
buf \U$297 ( \585 , \584_nG2b0 );
xor \U$298 ( \586 , \286 , \287 );
xor \U$299 ( \587 , \586 , \528 );
buf \U$300 ( \588 , \587 );
buf \U$301 ( \589 , RI2b1c4342b8c0_5);
and g2a2 ( \590_nG2a2 , \588 , \589 );
buf \U$302 ( \591 , \590_nG2a2 );
and \U$303 ( \592 , \585 , \591 );
not \U$304 ( \593 , \592 );
and \U$305 ( \594 , \558 , \593 );
not \U$306 ( \595 , \594 );
and \U$307 ( \596 , \568 , \561 );
and \U$308 ( \597 , \227 , \559 );
nor \U$309 ( \598 , \596 , \597 );
xnor \U$310 ( \599 , \598 , \566 );
and \U$311 ( \600 , \595 , \599 );
buf \U$313 ( \601 , RI2b1c4342d5d0_67);
and \U$314 ( \602 , \601 , \569 );
nor \U$315 ( \603 , 1'b0 , \602 );
not \U$316 ( \604 , \603 );
and \U$317 ( \605 , \599 , \604 );
and \U$318 ( \606 , \595 , \604 );
or \U$319 ( \607 , \600 , \605 , \606 );
xnor \U$320 ( \608 , \567 , \572 );
and \U$321 ( \609 , \607 , \608 );
nand \U$322 ( \610 , \579 , \609 );
nor \U$323 ( \611 , \579 , \609 );
not \U$324 ( \612 , \611 );
nand \U$325 ( \613 , \610 , \612 );
xor \U$326 ( \614 , \292 , \293 );
xor \U$327 ( \615 , \614 , \525 );
buf \U$328 ( \616 , \615 );
buf \U$329 ( \617 , RI2b1c4342b938_6);
and g294 ( \618_nG294 , \616 , \617 );
buf \U$330 ( \619 , \618_nG294 );
xor \U$331 ( \620 , \298 , \299 );
xor \U$332 ( \621 , \620 , \522 );
buf \U$333 ( \622 , \621 );
buf \U$334 ( \623 , RI2b1c4342b9b0_7);
and g286 ( \624_nG286 , \622 , \623 );
buf \U$335 ( \625 , \624_nG286 );
and \U$336 ( \626 , \619 , \625 );
not \U$337 ( \627 , \626 );
and \U$338 ( \628 , \591 , \627 );
buf \U$339 ( \629 , RI2b1c4342d7b0_71);
xor \U$340 ( \630 , \442 , \443 );
xor \U$341 ( \631 , \630 , \450 );
buf \U$342 ( \632 , \631 );
buf \U$343 ( \633 , RI2b1c4342c4f0_31);
and g136 ( \634_nG136 , \632 , \633 );
buf \U$344 ( \635 , \634_nG136 );
xor \U$345 ( \636 , \448 , \449 );
buf \U$346 ( \637 , \636 );
xor \U$347 ( \638 , RI2b1c4342c5e0_33, RI2b1c4342c658_34);
xor \U$348 ( \639 , RI2b1c4342c6d0_35, RI2b1c4342c748_36);
xor \U$349 ( \640 , \638 , \639 );
xor \U$350 ( \641 , RI2b1c4342c7c0_37, RI2b1c4342c838_38);
xor \U$351 ( \642 , RI2b1c4342c8b0_39, RI2b1c4342c928_40);
xor \U$352 ( \643 , \641 , \642 );
xor \U$353 ( \644 , \640 , \643 );
xor \U$354 ( \645 , RI2b1c4342c9a0_41, RI2b1c4342ca18_42);
xor \U$355 ( \646 , RI2b1c4342ca90_43, RI2b1c4342cb08_44);
xor \U$356 ( \647 , \645 , \646 );
xor \U$357 ( \648 , RI2b1c4342cb80_45, RI2b1c4342cbf8_46);
xor \U$358 ( \649 , RI2b1c4342cc70_47, RI2b1c4342cce8_48);
xor \U$359 ( \650 , \648 , \649 );
xor \U$360 ( \651 , \647 , \650 );
xor \U$361 ( \652 , \644 , \651 );
xor \U$362 ( \653 , RI2b1c4342cd60_49, RI2b1c4342cdd8_50);
xor \U$363 ( \654 , RI2b1c4342ce50_51, RI2b1c4342cec8_52);
xor \U$364 ( \655 , \653 , \654 );
xor \U$365 ( \656 , RI2b1c4342cf40_53, RI2b1c4342cfb8_54);
xor \U$366 ( \657 , RI2b1c4342d030_55, RI2b1c4342d0a8_56);
xor \U$367 ( \658 , \656 , \657 );
xor \U$368 ( \659 , \655 , \658 );
xor \U$369 ( \660 , RI2b1c4342d120_57, RI2b1c4342d198_58);
xor \U$370 ( \661 , RI2b1c4342d210_59, RI2b1c4342d288_60);
xor \U$371 ( \662 , \660 , \661 );
xor \U$372 ( \663 , RI2b1c4342d300_61, RI2b1c4342d378_62);
xor \U$373 ( \664 , RI2b1c4342d3f0_63, RI2b1c4342d468_64);
xor \U$374 ( \665 , \663 , \664 );
xor \U$375 ( \666 , \662 , \665 );
xor \U$376 ( \667 , \659 , \666 );
xor \U$377 ( \668 , \652 , \667 );
xor \U$378 ( \669 , \668 , RI2b1c4342c568_32);
and g12b ( \670_nG12b , \637 , \669 );
buf \U$379 ( \671 , \670_nG12b );
xor \U$380 ( \672 , \635 , \671 );
not \U$381 ( \673 , \671 );
and \U$382 ( \674 , \672 , \673 );
and \U$383 ( \675 , \629 , \674 );
buf \U$384 ( \676 , RI2b1c4342d738_70);
and \U$385 ( \677 , \676 , \671 );
nor \U$386 ( \678 , \675 , \677 );
xnor \U$387 ( \679 , \678 , \635 );
and \U$388 ( \680 , \628 , \679 );
buf \U$389 ( \681 , RI2b1c4342d8a0_73);
xor \U$390 ( \682 , \430 , \431 );
xor \U$391 ( \683 , \682 , \456 );
buf \U$392 ( \684 , \683 );
buf \U$393 ( \685 , RI2b1c4342c400_29);
and g152 ( \686_nG152 , \684 , \685 );
buf \U$394 ( \687 , \686_nG152 );
xor \U$395 ( \688 , \436 , \437 );
xor \U$396 ( \689 , \688 , \453 );
buf \U$397 ( \690 , \689 );
buf \U$398 ( \691 , RI2b1c4342c478_30);
and g144 ( \692_nG144 , \690 , \691 );
buf \U$399 ( \693 , \692_nG144 );
xor \U$400 ( \694 , \687 , \693 );
xor \U$401 ( \695 , \693 , \635 );
not \U$402 ( \696 , \695 );
and \U$403 ( \697 , \694 , \696 );
and \U$404 ( \698 , \681 , \697 );
buf \U$405 ( \699 , RI2b1c4342d828_72);
and \U$406 ( \700 , \699 , \695 );
nor \U$407 ( \701 , \698 , \700 );
and \U$408 ( \702 , \693 , \635 );
not \U$409 ( \703 , \702 );
and \U$410 ( \704 , \687 , \703 );
xnor \U$411 ( \705 , \701 , \704 );
and \U$412 ( \706 , \679 , \705 );
and \U$413 ( \707 , \628 , \705 );
or \U$414 ( \708 , \680 , \706 , \707 );
buf \U$415 ( \709 , RI2b1c4342d990_75);
xor \U$416 ( \710 , \418 , \419 );
xor \U$417 ( \711 , \710 , \462 );
buf \U$418 ( \712 , \711 );
buf \U$419 ( \713 , RI2b1c4342c310_27);
and g16e ( \714_nG16e , \712 , \713 );
buf \U$420 ( \715 , \714_nG16e );
xor \U$421 ( \716 , \424 , \425 );
xor \U$422 ( \717 , \716 , \459 );
buf \U$423 ( \718 , \717 );
buf \U$424 ( \719 , RI2b1c4342c388_28);
and g160 ( \720_nG160 , \718 , \719 );
buf \U$425 ( \721 , \720_nG160 );
xor \U$426 ( \722 , \715 , \721 );
xor \U$427 ( \723 , \721 , \687 );
not \U$428 ( \724 , \723 );
and \U$429 ( \725 , \722 , \724 );
and \U$430 ( \726 , \709 , \725 );
buf \U$431 ( \727 , RI2b1c4342d918_74);
and \U$432 ( \728 , \727 , \723 );
nor \U$433 ( \729 , \726 , \728 );
and \U$434 ( \730 , \721 , \687 );
not \U$435 ( \731 , \730 );
and \U$436 ( \732 , \715 , \731 );
xnor \U$437 ( \733 , \729 , \732 );
buf \U$438 ( \734 , RI2b1c4342da80_77);
xor \U$439 ( \735 , \406 , \407 );
xor \U$440 ( \736 , \735 , \468 );
buf \U$441 ( \737 , \736 );
buf \U$442 ( \738 , RI2b1c4342c220_25);
and g18a ( \739_nG18a , \737 , \738 );
buf \U$443 ( \740 , \739_nG18a );
xor \U$444 ( \741 , \412 , \413 );
xor \U$445 ( \742 , \741 , \465 );
buf \U$446 ( \743 , \742 );
buf \U$447 ( \744 , RI2b1c4342c298_26);
and g17c ( \745_nG17c , \743 , \744 );
buf \U$448 ( \746 , \745_nG17c );
xor \U$449 ( \747 , \740 , \746 );
xor \U$450 ( \748 , \746 , \715 );
not \U$451 ( \749 , \748 );
and \U$452 ( \750 , \747 , \749 );
and \U$453 ( \751 , \734 , \750 );
buf \U$454 ( \752 , RI2b1c4342da08_76);
and \U$455 ( \753 , \752 , \748 );
nor \U$456 ( \754 , \751 , \753 );
and \U$457 ( \755 , \746 , \715 );
not \U$458 ( \756 , \755 );
and \U$459 ( \757 , \740 , \756 );
xnor \U$460 ( \758 , \754 , \757 );
and \U$461 ( \759 , \733 , \758 );
buf \U$462 ( \760 , RI2b1c4342db70_79);
xor \U$463 ( \761 , \394 , \395 );
xor \U$464 ( \762 , \761 , \474 );
buf \U$465 ( \763 , \762 );
buf \U$466 ( \764 , RI2b1c4342c130_23);
and g1a6 ( \765_nG1a6 , \763 , \764 );
buf \U$467 ( \766 , \765_nG1a6 );
xor \U$468 ( \767 , \400 , \401 );
xor \U$469 ( \768 , \767 , \471 );
buf \U$470 ( \769 , \768 );
buf \U$471 ( \770 , RI2b1c4342c1a8_24);
and g198 ( \771_nG198 , \769 , \770 );
buf \U$472 ( \772 , \771_nG198 );
xor \U$473 ( \773 , \766 , \772 );
xor \U$474 ( \774 , \772 , \740 );
not \U$475 ( \775 , \774 );
and \U$476 ( \776 , \773 , \775 );
and \U$477 ( \777 , \760 , \776 );
buf \U$478 ( \778 , RI2b1c4342daf8_78);
and \U$479 ( \779 , \778 , \774 );
nor \U$480 ( \780 , \777 , \779 );
and \U$481 ( \781 , \772 , \740 );
not \U$482 ( \782 , \781 );
and \U$483 ( \783 , \766 , \782 );
xnor \U$484 ( \784 , \780 , \783 );
and \U$485 ( \785 , \758 , \784 );
and \U$486 ( \786 , \733 , \784 );
or \U$487 ( \787 , \759 , \785 , \786 );
and \U$488 ( \788 , \708 , \787 );
buf \U$489 ( \789 , RI2b1c4342dc60_81);
xor \U$490 ( \790 , \382 , \383 );
xor \U$491 ( \791 , \790 , \480 );
buf \U$492 ( \792 , \791 );
buf \U$493 ( \793 , RI2b1c4342c040_21);
and g1c2 ( \794_nG1c2 , \792 , \793 );
buf \U$494 ( \795 , \794_nG1c2 );
xor \U$495 ( \796 , \388 , \389 );
xor \U$496 ( \797 , \796 , \477 );
buf \U$497 ( \798 , \797 );
buf \U$498 ( \799 , RI2b1c4342c0b8_22);
and g1b4 ( \800_nG1b4 , \798 , \799 );
buf \U$499 ( \801 , \800_nG1b4 );
xor \U$500 ( \802 , \795 , \801 );
xor \U$501 ( \803 , \801 , \766 );
not \U$502 ( \804 , \803 );
and \U$503 ( \805 , \802 , \804 );
and \U$504 ( \806 , \789 , \805 );
buf \U$505 ( \807 , RI2b1c4342dbe8_80);
and \U$506 ( \808 , \807 , \803 );
nor \U$507 ( \809 , \806 , \808 );
and \U$508 ( \810 , \801 , \766 );
not \U$509 ( \811 , \810 );
and \U$510 ( \812 , \795 , \811 );
xnor \U$511 ( \813 , \809 , \812 );
buf \U$512 ( \814 , RI2b1c4342dd50_83);
xor \U$513 ( \815 , \370 , \371 );
xor \U$514 ( \816 , \815 , \486 );
buf \U$515 ( \817 , \816 );
buf \U$516 ( \818 , RI2b1c4342bf50_19);
and g1de ( \819_nG1de , \817 , \818 );
buf \U$517 ( \820 , \819_nG1de );
xor \U$518 ( \821 , \376 , \377 );
xor \U$519 ( \822 , \821 , \483 );
buf \U$520 ( \823 , \822 );
buf \U$521 ( \824 , RI2b1c4342bfc8_20);
and g1d0 ( \825_nG1d0 , \823 , \824 );
buf \U$522 ( \826 , \825_nG1d0 );
xor \U$523 ( \827 , \820 , \826 );
xor \U$524 ( \828 , \826 , \795 );
not \U$525 ( \829 , \828 );
and \U$526 ( \830 , \827 , \829 );
and \U$527 ( \831 , \814 , \830 );
buf \U$528 ( \832 , RI2b1c4342dcd8_82);
and \U$529 ( \833 , \832 , \828 );
nor \U$530 ( \834 , \831 , \833 );
and \U$531 ( \835 , \826 , \795 );
not \U$532 ( \836 , \835 );
and \U$533 ( \837 , \820 , \836 );
xnor \U$534 ( \838 , \834 , \837 );
and \U$535 ( \839 , \813 , \838 );
buf \U$536 ( \840 , RI2b1c4342de40_85);
xor \U$537 ( \841 , \358 , \359 );
xor \U$538 ( \842 , \841 , \492 );
buf \U$539 ( \843 , \842 );
buf \U$540 ( \844 , RI2b1c4342be60_17);
and g1fa ( \845_nG1fa , \843 , \844 );
buf \U$541 ( \846 , \845_nG1fa );
xor \U$542 ( \847 , \364 , \365 );
xor \U$543 ( \848 , \847 , \489 );
buf \U$544 ( \849 , \848 );
buf \U$545 ( \850 , RI2b1c4342bed8_18);
and g1ec ( \851_nG1ec , \849 , \850 );
buf \U$546 ( \852 , \851_nG1ec );
xor \U$547 ( \853 , \846 , \852 );
xor \U$548 ( \854 , \852 , \820 );
not \U$549 ( \855 , \854 );
and \U$550 ( \856 , \853 , \855 );
and \U$551 ( \857 , \840 , \856 );
buf \U$552 ( \858 , RI2b1c4342ddc8_84);
and \U$553 ( \859 , \858 , \854 );
nor \U$554 ( \860 , \857 , \859 );
and \U$555 ( \861 , \852 , \820 );
not \U$556 ( \862 , \861 );
and \U$557 ( \863 , \846 , \862 );
xnor \U$558 ( \864 , \860 , \863 );
and \U$559 ( \865 , \838 , \864 );
and \U$560 ( \866 , \813 , \864 );
or \U$561 ( \867 , \839 , \865 , \866 );
and \U$562 ( \868 , \787 , \867 );
and \U$563 ( \869 , \708 , \867 );
or \U$564 ( \870 , \788 , \868 , \869 );
buf \U$565 ( \871 , RI2b1c4342df30_87);
xor \U$566 ( \872 , \346 , \347 );
xor \U$567 ( \873 , \872 , \498 );
buf \U$568 ( \874 , \873 );
buf \U$569 ( \875 , RI2b1c4342bd70_15);
and g216 ( \876_nG216 , \874 , \875 );
buf \U$570 ( \877 , \876_nG216 );
xor \U$571 ( \878 , \352 , \353 );
xor \U$572 ( \879 , \878 , \495 );
buf \U$573 ( \880 , \879 );
buf \U$574 ( \881 , RI2b1c4342bde8_16);
and g208 ( \882_nG208 , \880 , \881 );
buf \U$575 ( \883 , \882_nG208 );
xor \U$576 ( \884 , \877 , \883 );
xor \U$577 ( \885 , \883 , \846 );
not \U$578 ( \886 , \885 );
and \U$579 ( \887 , \884 , \886 );
and \U$580 ( \888 , \871 , \887 );
buf \U$581 ( \889 , RI2b1c4342deb8_86);
and \U$582 ( \890 , \889 , \885 );
nor \U$583 ( \891 , \888 , \890 );
and \U$584 ( \892 , \883 , \846 );
not \U$585 ( \893 , \892 );
and \U$586 ( \894 , \877 , \893 );
xnor \U$587 ( \895 , \891 , \894 );
buf \U$588 ( \896 , RI2b1c4342e020_89);
xor \U$589 ( \897 , \334 , \335 );
xor \U$590 ( \898 , \897 , \504 );
buf \U$591 ( \899 , \898 );
buf \U$592 ( \900 , RI2b1c4342bc80_13);
and g232 ( \901_nG232 , \899 , \900 );
buf \U$593 ( \902 , \901_nG232 );
xor \U$594 ( \903 , \340 , \341 );
xor \U$595 ( \904 , \903 , \501 );
buf \U$596 ( \905 , \904 );
buf \U$597 ( \906 , RI2b1c4342bcf8_14);
and g224 ( \907_nG224 , \905 , \906 );
buf \U$598 ( \908 , \907_nG224 );
xor \U$599 ( \909 , \902 , \908 );
xor \U$600 ( \910 , \908 , \877 );
not \U$601 ( \911 , \910 );
and \U$602 ( \912 , \909 , \911 );
and \U$603 ( \913 , \896 , \912 );
buf \U$604 ( \914 , RI2b1c4342dfa8_88);
and \U$605 ( \915 , \914 , \910 );
nor \U$606 ( \916 , \913 , \915 );
and \U$607 ( \917 , \908 , \877 );
not \U$608 ( \918 , \917 );
and \U$609 ( \919 , \902 , \918 );
xnor \U$610 ( \920 , \916 , \919 );
and \U$611 ( \921 , \895 , \920 );
buf \U$612 ( \922 , RI2b1c4342e110_91);
xor \U$613 ( \923 , \322 , \323 );
xor \U$614 ( \924 , \923 , \510 );
buf \U$615 ( \925 , \924 );
buf \U$616 ( \926 , RI2b1c4342bb90_11);
and g24e ( \927_nG24e , \925 , \926 );
buf \U$617 ( \928 , \927_nG24e );
xor \U$618 ( \929 , \328 , \329 );
xor \U$619 ( \930 , \929 , \507 );
buf \U$620 ( \931 , \930 );
buf \U$621 ( \932 , RI2b1c4342bc08_12);
and g240 ( \933_nG240 , \931 , \932 );
buf \U$622 ( \934 , \933_nG240 );
xor \U$623 ( \935 , \928 , \934 );
xor \U$624 ( \936 , \934 , \902 );
not \U$625 ( \937 , \936 );
and \U$626 ( \938 , \935 , \937 );
and \U$627 ( \939 , \922 , \938 );
buf \U$628 ( \940 , RI2b1c4342e098_90);
and \U$629 ( \941 , \940 , \936 );
nor \U$630 ( \942 , \939 , \941 );
and \U$631 ( \943 , \934 , \902 );
not \U$632 ( \944 , \943 );
and \U$633 ( \945 , \928 , \944 );
xnor \U$634 ( \946 , \942 , \945 );
and \U$635 ( \947 , \920 , \946 );
and \U$636 ( \948 , \895 , \946 );
or \U$637 ( \949 , \921 , \947 , \948 );
buf \U$638 ( \950 , RI2b1c4342e200_93);
xor \U$639 ( \951 , \310 , \311 );
xor \U$640 ( \952 , \951 , \516 );
buf \U$641 ( \953 , \952 );
buf \U$642 ( \954 , RI2b1c4342baa0_9);
and g26a ( \955_nG26a , \953 , \954 );
buf \U$643 ( \956 , \955_nG26a );
xor \U$644 ( \957 , \316 , \317 );
xor \U$645 ( \958 , \957 , \513 );
buf \U$646 ( \959 , \958 );
buf \U$647 ( \960 , RI2b1c4342bb18_10);
and g25c ( \961_nG25c , \959 , \960 );
buf \U$648 ( \962 , \961_nG25c );
xor \U$649 ( \963 , \956 , \962 );
xor \U$650 ( \964 , \962 , \928 );
not \U$651 ( \965 , \964 );
and \U$652 ( \966 , \963 , \965 );
and \U$653 ( \967 , \950 , \966 );
buf \U$654 ( \968 , RI2b1c4342e188_92);
and \U$655 ( \969 , \968 , \964 );
nor \U$656 ( \970 , \967 , \969 );
and \U$657 ( \971 , \962 , \928 );
not \U$658 ( \972 , \971 );
and \U$659 ( \973 , \956 , \972 );
xnor \U$660 ( \974 , \970 , \973 );
buf \U$661 ( \975 , RI2b1c4342e2f0_95);
xor \U$662 ( \976 , \304 , \305 );
xor \U$663 ( \977 , \976 , \519 );
buf \U$664 ( \978 , \977 );
buf \U$665 ( \979 , RI2b1c4342ba28_8);
and g278 ( \980_nG278 , \978 , \979 );
buf \U$666 ( \981 , \980_nG278 );
xor \U$667 ( \982 , \625 , \981 );
xor \U$668 ( \983 , \981 , \956 );
not \U$669 ( \984 , \983 );
and \U$670 ( \985 , \982 , \984 );
and \U$671 ( \986 , \975 , \985 );
buf \U$672 ( \987 , RI2b1c4342e278_94);
and \U$673 ( \988 , \987 , \983 );
nor \U$674 ( \989 , \986 , \988 );
and \U$675 ( \990 , \981 , \956 );
not \U$676 ( \991 , \990 );
and \U$677 ( \992 , \625 , \991 );
xnor \U$678 ( \993 , \989 , \992 );
and \U$679 ( \994 , \974 , \993 );
buf \U$680 ( \995 , RI2b1c4342e368_96);
xor \U$681 ( \996 , \619 , \625 );
nand \U$682 ( \997 , \995 , \996 );
xnor \U$683 ( \998 , \997 , \628 );
and \U$684 ( \999 , \993 , \998 );
and \U$685 ( \1000 , \974 , \998 );
or \U$686 ( \1001 , \994 , \999 , \1000 );
and \U$687 ( \1002 , \949 , \1001 );
and \U$688 ( \1003 , \987 , \985 );
and \U$689 ( \1004 , \950 , \983 );
nor \U$690 ( \1005 , \1003 , \1004 );
xnor \U$691 ( \1006 , \1005 , \992 );
and \U$692 ( \1007 , \1001 , \1006 );
and \U$693 ( \1008 , \949 , \1006 );
or \U$694 ( \1009 , \1002 , \1007 , \1008 );
and \U$695 ( \1010 , \870 , \1009 );
xor \U$696 ( \1011 , \591 , \619 );
not \U$697 ( \1012 , \996 );
and \U$698 ( \1013 , \1011 , \1012 );
and \U$699 ( \1014 , \995 , \1013 );
and \U$700 ( \1015 , \975 , \996 );
nor \U$701 ( \1016 , \1014 , \1015 );
xnor \U$702 ( \1017 , \1016 , \628 );
and \U$703 ( \1018 , \914 , \912 );
and \U$704 ( \1019 , \871 , \910 );
nor \U$705 ( \1020 , \1018 , \1019 );
xnor \U$706 ( \1021 , \1020 , \919 );
and \U$707 ( \1022 , \940 , \938 );
and \U$708 ( \1023 , \896 , \936 );
nor \U$709 ( \1024 , \1022 , \1023 );
xnor \U$710 ( \1025 , \1024 , \945 );
xor \U$711 ( \1026 , \1021 , \1025 );
and \U$712 ( \1027 , \968 , \966 );
and \U$713 ( \1028 , \922 , \964 );
nor \U$714 ( \1029 , \1027 , \1028 );
xnor \U$715 ( \1030 , \1029 , \973 );
xor \U$716 ( \1031 , \1026 , \1030 );
and \U$717 ( \1032 , \1017 , \1031 );
and \U$718 ( \1033 , \832 , \830 );
and \U$719 ( \1034 , \789 , \828 );
nor \U$720 ( \1035 , \1033 , \1034 );
xnor \U$721 ( \1036 , \1035 , \837 );
and \U$722 ( \1037 , \858 , \856 );
and \U$723 ( \1038 , \814 , \854 );
nor \U$724 ( \1039 , \1037 , \1038 );
xnor \U$725 ( \1040 , \1039 , \863 );
xor \U$726 ( \1041 , \1036 , \1040 );
and \U$727 ( \1042 , \889 , \887 );
and \U$728 ( \1043 , \840 , \885 );
nor \U$729 ( \1044 , \1042 , \1043 );
xnor \U$730 ( \1045 , \1044 , \894 );
xor \U$731 ( \1046 , \1041 , \1045 );
and \U$732 ( \1047 , \1031 , \1046 );
and \U$733 ( \1048 , \1017 , \1046 );
or \U$734 ( \1049 , \1032 , \1047 , \1048 );
and \U$735 ( \1050 , \1009 , \1049 );
and \U$736 ( \1051 , \870 , \1049 );
or \U$737 ( \1052 , \1010 , \1050 , \1051 );
buf \U$738 ( \1053 , RI2b1c4342d6c0_69);
and \U$739 ( \1054 , \1053 , \674 );
buf \U$740 ( \1055 , RI2b1c4342d648_68);
and \U$741 ( \1056 , \1055 , \671 );
nor \U$742 ( \1057 , \1054 , \1056 );
xnor \U$743 ( \1058 , \1057 , \635 );
xor \U$744 ( \1059 , \594 , \1058 );
and \U$745 ( \1060 , \629 , \697 );
and \U$746 ( \1061 , \676 , \695 );
nor \U$747 ( \1062 , \1060 , \1061 );
xnor \U$748 ( \1063 , \1062 , \704 );
xor \U$749 ( \1064 , \1059 , \1063 );
and \U$750 ( \1065 , \840 , \887 );
and \U$751 ( \1066 , \858 , \885 );
nor \U$752 ( \1067 , \1065 , \1066 );
xnor \U$753 ( \1068 , \1067 , \894 );
and \U$754 ( \1069 , \871 , \912 );
and \U$755 ( \1070 , \889 , \910 );
nor \U$756 ( \1071 , \1069 , \1070 );
xnor \U$757 ( \1072 , \1071 , \919 );
xor \U$758 ( \1073 , \1068 , \1072 );
and \U$759 ( \1074 , \896 , \938 );
and \U$760 ( \1075 , \914 , \936 );
nor \U$761 ( \1076 , \1074 , \1075 );
xnor \U$762 ( \1077 , \1076 , \945 );
xor \U$763 ( \1078 , \1073 , \1077 );
and \U$764 ( \1079 , \760 , \805 );
and \U$765 ( \1080 , \778 , \803 );
nor \U$766 ( \1081 , \1079 , \1080 );
xnor \U$767 ( \1082 , \1081 , \812 );
and \U$768 ( \1083 , \789 , \830 );
and \U$769 ( \1084 , \807 , \828 );
nor \U$770 ( \1085 , \1083 , \1084 );
xnor \U$771 ( \1086 , \1085 , \837 );
xor \U$772 ( \1087 , \1082 , \1086 );
and \U$773 ( \1088 , \814 , \856 );
and \U$774 ( \1089 , \832 , \854 );
nor \U$775 ( \1090 , \1088 , \1089 );
xnor \U$776 ( \1091 , \1090 , \863 );
xor \U$777 ( \1092 , \1087 , \1091 );
xor \U$778 ( \1093 , \1078 , \1092 );
and \U$779 ( \1094 , \681 , \725 );
and \U$780 ( \1095 , \699 , \723 );
nor \U$781 ( \1096 , \1094 , \1095 );
xnor \U$782 ( \1097 , \1096 , \732 );
and \U$783 ( \1098 , \709 , \750 );
and \U$784 ( \1099 , \727 , \748 );
nor \U$785 ( \1100 , \1098 , \1099 );
xnor \U$786 ( \1101 , \1100 , \757 );
xor \U$787 ( \1102 , \1097 , \1101 );
and \U$788 ( \1103 , \734 , \776 );
and \U$789 ( \1104 , \752 , \774 );
nor \U$790 ( \1105 , \1103 , \1104 );
xnor \U$791 ( \1106 , \1105 , \783 );
xor \U$792 ( \1107 , \1102 , \1106 );
xor \U$793 ( \1108 , \1093 , \1107 );
and \U$794 ( \1109 , \1064 , \1108 );
and \U$795 ( \1110 , \1021 , \1025 );
and \U$796 ( \1111 , \1025 , \1030 );
and \U$797 ( \1112 , \1021 , \1030 );
or \U$798 ( \1113 , \1110 , \1111 , \1112 );
xor \U$799 ( \1114 , \585 , \591 );
nand \U$800 ( \1115 , \995 , \1114 );
xnor \U$801 ( \1116 , \1115 , \594 );
xor \U$802 ( \1117 , \1113 , \1116 );
and \U$803 ( \1118 , \922 , \966 );
and \U$804 ( \1119 , \940 , \964 );
nor \U$805 ( \1120 , \1118 , \1119 );
xnor \U$806 ( \1121 , \1120 , \973 );
and \U$807 ( \1122 , \950 , \985 );
and \U$808 ( \1123 , \968 , \983 );
nor \U$809 ( \1124 , \1122 , \1123 );
xnor \U$810 ( \1125 , \1124 , \992 );
xor \U$811 ( \1126 , \1121 , \1125 );
and \U$812 ( \1127 , \975 , \1013 );
and \U$813 ( \1128 , \987 , \996 );
nor \U$814 ( \1129 , \1127 , \1128 );
xnor \U$815 ( \1130 , \1129 , \628 );
xor \U$816 ( \1131 , \1126 , \1130 );
xor \U$817 ( \1132 , \1117 , \1131 );
and \U$818 ( \1133 , \1108 , \1132 );
and \U$819 ( \1134 , \1064 , \1132 );
or \U$820 ( \1135 , \1109 , \1133 , \1134 );
and \U$821 ( \1136 , \1052 , \1135 );
and \U$822 ( \1137 , \594 , \1058 );
and \U$823 ( \1138 , \1058 , \1063 );
and \U$824 ( \1139 , \594 , \1063 );
or \U$825 ( \1140 , \1137 , \1138 , \1139 );
and \U$826 ( \1141 , \1097 , \1101 );
and \U$827 ( \1142 , \1101 , \1106 );
and \U$828 ( \1143 , \1097 , \1106 );
or \U$829 ( \1144 , \1141 , \1142 , \1143 );
xor \U$830 ( \1145 , \1140 , \1144 );
and \U$831 ( \1146 , \1082 , \1086 );
and \U$832 ( \1147 , \1086 , \1091 );
and \U$833 ( \1148 , \1082 , \1091 );
or \U$834 ( \1149 , \1146 , \1147 , \1148 );
xor \U$835 ( \1150 , \1145 , \1149 );
and \U$836 ( \1151 , \1135 , \1150 );
and \U$837 ( \1152 , \1052 , \1150 );
or \U$838 ( \1153 , \1136 , \1151 , \1152 );
and \U$839 ( \1154 , \1055 , \674 );
and \U$840 ( \1155 , \601 , \671 );
nor \U$841 ( \1156 , \1154 , \1155 );
xnor \U$842 ( \1157 , \1156 , \635 );
and \U$843 ( \1158 , \676 , \697 );
and \U$844 ( \1159 , \1053 , \695 );
nor \U$845 ( \1160 , \1158 , \1159 );
xnor \U$846 ( \1161 , \1160 , \704 );
xor \U$847 ( \1162 , \1157 , \1161 );
and \U$848 ( \1163 , \699 , \725 );
and \U$849 ( \1164 , \629 , \723 );
nor \U$850 ( \1165 , \1163 , \1164 );
xnor \U$851 ( \1166 , \1165 , \732 );
xor \U$852 ( \1167 , \1162 , \1166 );
and \U$853 ( \1168 , \889 , \912 );
and \U$854 ( \1169 , \840 , \910 );
nor \U$855 ( \1170 , \1168 , \1169 );
xnor \U$856 ( \1171 , \1170 , \919 );
and \U$857 ( \1172 , \914 , \938 );
and \U$858 ( \1173 , \871 , \936 );
nor \U$859 ( \1174 , \1172 , \1173 );
xnor \U$860 ( \1175 , \1174 , \945 );
xor \U$861 ( \1176 , \1171 , \1175 );
and \U$862 ( \1177 , \940 , \966 );
and \U$863 ( \1178 , \896 , \964 );
nor \U$864 ( \1179 , \1177 , \1178 );
xnor \U$865 ( \1180 , \1179 , \973 );
xor \U$866 ( \1181 , \1176 , \1180 );
and \U$867 ( \1182 , \807 , \830 );
and \U$868 ( \1183 , \760 , \828 );
nor \U$869 ( \1184 , \1182 , \1183 );
xnor \U$870 ( \1185 , \1184 , \837 );
and \U$871 ( \1186 , \832 , \856 );
and \U$872 ( \1187 , \789 , \854 );
nor \U$873 ( \1188 , \1186 , \1187 );
xnor \U$874 ( \1189 , \1188 , \863 );
xor \U$875 ( \1190 , \1185 , \1189 );
and \U$876 ( \1191 , \858 , \887 );
and \U$877 ( \1192 , \814 , \885 );
nor \U$878 ( \1193 , \1191 , \1192 );
xnor \U$879 ( \1194 , \1193 , \894 );
xor \U$880 ( \1195 , \1190 , \1194 );
xor \U$881 ( \1196 , \1181 , \1195 );
and \U$882 ( \1197 , \727 , \750 );
and \U$883 ( \1198 , \681 , \748 );
nor \U$884 ( \1199 , \1197 , \1198 );
xnor \U$885 ( \1200 , \1199 , \757 );
and \U$886 ( \1201 , \752 , \776 );
and \U$887 ( \1202 , \709 , \774 );
nor \U$888 ( \1203 , \1201 , \1202 );
xnor \U$889 ( \1204 , \1203 , \783 );
xor \U$890 ( \1205 , \1200 , \1204 );
and \U$891 ( \1206 , \778 , \805 );
and \U$892 ( \1207 , \734 , \803 );
nor \U$893 ( \1208 , \1206 , \1207 );
xnor \U$894 ( \1209 , \1208 , \812 );
xor \U$895 ( \1210 , \1205 , \1209 );
xor \U$896 ( \1211 , \1196 , \1210 );
xor \U$897 ( \1212 , \1167 , \1211 );
and \U$898 ( \1213 , \1068 , \1072 );
and \U$899 ( \1214 , \1072 , \1077 );
and \U$900 ( \1215 , \1068 , \1077 );
or \U$901 ( \1216 , \1213 , \1214 , \1215 );
and \U$902 ( \1217 , \1121 , \1125 );
and \U$903 ( \1218 , \1125 , \1130 );
and \U$904 ( \1219 , \1121 , \1130 );
or \U$905 ( \1220 , \1217 , \1218 , \1219 );
xor \U$906 ( \1221 , \1216 , \1220 );
and \U$907 ( \1222 , \968 , \985 );
and \U$908 ( \1223 , \922 , \983 );
nor \U$909 ( \1224 , \1222 , \1223 );
xnor \U$910 ( \1225 , \1224 , \992 );
and \U$911 ( \1226 , \987 , \1013 );
and \U$912 ( \1227 , \950 , \996 );
nor \U$913 ( \1228 , \1226 , \1227 );
xnor \U$914 ( \1229 , \1228 , \628 );
xor \U$915 ( \1230 , \1225 , \1229 );
xor \U$916 ( \1231 , \558 , \585 );
not \U$917 ( \1232 , \1114 );
and \U$918 ( \1233 , \1231 , \1232 );
and \U$919 ( \1234 , \995 , \1233 );
and \U$920 ( \1235 , \975 , \1114 );
nor \U$921 ( \1236 , \1234 , \1235 );
xnor \U$922 ( \1237 , \1236 , \594 );
xor \U$923 ( \1238 , \1230 , \1237 );
xor \U$924 ( \1239 , \1221 , \1238 );
xor \U$925 ( \1240 , \1212 , \1239 );
and \U$926 ( \1241 , \676 , \674 );
and \U$927 ( \1242 , \1053 , \671 );
nor \U$928 ( \1243 , \1241 , \1242 );
xnor \U$929 ( \1244 , \1243 , \635 );
and \U$930 ( \1245 , \699 , \697 );
and \U$931 ( \1246 , \629 , \695 );
nor \U$932 ( \1247 , \1245 , \1246 );
xnor \U$933 ( \1248 , \1247 , \704 );
and \U$934 ( \1249 , \1244 , \1248 );
and \U$935 ( \1250 , \727 , \725 );
and \U$936 ( \1251 , \681 , \723 );
nor \U$937 ( \1252 , \1250 , \1251 );
xnor \U$938 ( \1253 , \1252 , \732 );
and \U$939 ( \1254 , \1248 , \1253 );
and \U$940 ( \1255 , \1244 , \1253 );
or \U$941 ( \1256 , \1249 , \1254 , \1255 );
and \U$942 ( \1257 , \752 , \750 );
and \U$943 ( \1258 , \709 , \748 );
nor \U$944 ( \1259 , \1257 , \1258 );
xnor \U$945 ( \1260 , \1259 , \757 );
and \U$946 ( \1261 , \778 , \776 );
and \U$947 ( \1262 , \734 , \774 );
nor \U$948 ( \1263 , \1261 , \1262 );
xnor \U$949 ( \1264 , \1263 , \783 );
and \U$950 ( \1265 , \1260 , \1264 );
and \U$951 ( \1266 , \807 , \805 );
and \U$952 ( \1267 , \760 , \803 );
nor \U$953 ( \1268 , \1266 , \1267 );
xnor \U$954 ( \1269 , \1268 , \812 );
and \U$955 ( \1270 , \1264 , \1269 );
and \U$956 ( \1271 , \1260 , \1269 );
or \U$957 ( \1272 , \1265 , \1270 , \1271 );
and \U$958 ( \1273 , \1256 , \1272 );
and \U$959 ( \1274 , \1036 , \1040 );
and \U$960 ( \1275 , \1040 , \1045 );
and \U$961 ( \1276 , \1036 , \1045 );
or \U$962 ( \1277 , \1274 , \1275 , \1276 );
and \U$963 ( \1278 , \1272 , \1277 );
and \U$964 ( \1279 , \1256 , \1277 );
or \U$965 ( \1280 , \1273 , \1278 , \1279 );
and \U$966 ( \1281 , \1113 , \1116 );
and \U$967 ( \1282 , \1116 , \1131 );
and \U$968 ( \1283 , \1113 , \1131 );
or \U$969 ( \1284 , \1281 , \1282 , \1283 );
xor \U$970 ( \1285 , \1280 , \1284 );
and \U$971 ( \1286 , \1078 , \1092 );
and \U$972 ( \1287 , \1092 , \1107 );
and \U$973 ( \1288 , \1078 , \1107 );
or \U$974 ( \1289 , \1286 , \1287 , \1288 );
xor \U$975 ( \1290 , \1285 , \1289 );
and \U$976 ( \1291 , \1240 , \1290 );
and \U$977 ( \1292 , \1153 , \1291 );
and \U$978 ( \1293 , \734 , \805 );
and \U$979 ( \1294 , \752 , \803 );
nor \U$980 ( \1295 , \1293 , \1294 );
xnor \U$981 ( \1296 , \1295 , \812 );
and \U$982 ( \1297 , \760 , \830 );
and \U$983 ( \1298 , \778 , \828 );
nor \U$984 ( \1299 , \1297 , \1298 );
xnor \U$985 ( \1300 , \1299 , \837 );
xor \U$986 ( \1301 , \1296 , \1300 );
and \U$987 ( \1302 , \789 , \856 );
and \U$988 ( \1303 , \807 , \854 );
nor \U$989 ( \1304 , \1302 , \1303 );
xnor \U$990 ( \1305 , \1304 , \863 );
xor \U$991 ( \1306 , \1301 , \1305 );
and \U$992 ( \1307 , \629 , \725 );
and \U$993 ( \1308 , \676 , \723 );
nor \U$994 ( \1309 , \1307 , \1308 );
xnor \U$995 ( \1310 , \1309 , \732 );
and \U$996 ( \1311 , \681 , \750 );
and \U$997 ( \1312 , \699 , \748 );
nor \U$998 ( \1313 , \1311 , \1312 );
xnor \U$999 ( \1314 , \1313 , \757 );
xor \U$1000 ( \1315 , \1310 , \1314 );
and \U$1001 ( \1316 , \709 , \776 );
and \U$1002 ( \1317 , \727 , \774 );
nor \U$1003 ( \1318 , \1316 , \1317 );
xnor \U$1004 ( \1319 , \1318 , \783 );
xor \U$1005 ( \1320 , \1315 , \1319 );
xor \U$1006 ( \1321 , \1306 , \1320 );
and \U$1007 ( \1322 , \601 , \674 );
and \U$1008 ( \1323 , \568 , \671 );
nor \U$1009 ( \1324 , \1322 , \1323 );
xnor \U$1010 ( \1325 , \1324 , \635 );
xor \U$1011 ( \1326 , \566 , \1325 );
and \U$1012 ( \1327 , \1053 , \697 );
and \U$1013 ( \1328 , \1055 , \695 );
nor \U$1014 ( \1329 , \1327 , \1328 );
xnor \U$1015 ( \1330 , \1329 , \704 );
xor \U$1016 ( \1331 , \1326 , \1330 );
xor \U$1017 ( \1332 , \1321 , \1331 );
nand \U$1018 ( \1333 , \995 , \559 );
xnor \U$1019 ( \1334 , \1333 , \566 );
and \U$1020 ( \1335 , \896 , \966 );
and \U$1021 ( \1336 , \914 , \964 );
nor \U$1022 ( \1337 , \1335 , \1336 );
xnor \U$1023 ( \1338 , \1337 , \973 );
and \U$1024 ( \1339 , \922 , \985 );
and \U$1025 ( \1340 , \940 , \983 );
nor \U$1026 ( \1341 , \1339 , \1340 );
xnor \U$1027 ( \1342 , \1341 , \992 );
xor \U$1028 ( \1343 , \1338 , \1342 );
and \U$1029 ( \1344 , \950 , \1013 );
and \U$1030 ( \1345 , \968 , \996 );
nor \U$1031 ( \1346 , \1344 , \1345 );
xnor \U$1032 ( \1347 , \1346 , \628 );
xor \U$1033 ( \1348 , \1343 , \1347 );
xor \U$1034 ( \1349 , \1334 , \1348 );
and \U$1035 ( \1350 , \814 , \887 );
and \U$1036 ( \1351 , \832 , \885 );
nor \U$1037 ( \1352 , \1350 , \1351 );
xnor \U$1038 ( \1353 , \1352 , \894 );
and \U$1039 ( \1354 , \840 , \912 );
and \U$1040 ( \1355 , \858 , \910 );
nor \U$1041 ( \1356 , \1354 , \1355 );
xnor \U$1042 ( \1357 , \1356 , \919 );
xor \U$1043 ( \1358 , \1353 , \1357 );
and \U$1044 ( \1359 , \871 , \938 );
and \U$1045 ( \1360 , \889 , \936 );
nor \U$1046 ( \1361 , \1359 , \1360 );
xnor \U$1047 ( \1362 , \1361 , \945 );
xor \U$1048 ( \1363 , \1358 , \1362 );
xor \U$1049 ( \1364 , \1349 , \1363 );
xor \U$1050 ( \1365 , \1332 , \1364 );
and \U$1051 ( \1366 , \1171 , \1175 );
and \U$1052 ( \1367 , \1175 , \1180 );
and \U$1053 ( \1368 , \1171 , \1180 );
or \U$1054 ( \1369 , \1366 , \1367 , \1368 );
and \U$1055 ( \1370 , \1225 , \1229 );
and \U$1056 ( \1371 , \1229 , \1237 );
and \U$1057 ( \1372 , \1225 , \1237 );
or \U$1058 ( \1373 , \1370 , \1371 , \1372 );
xor \U$1059 ( \1374 , \1369 , \1373 );
and \U$1060 ( \1375 , \975 , \1233 );
and \U$1061 ( \1376 , \987 , \1114 );
nor \U$1062 ( \1377 , \1375 , \1376 );
xnor \U$1063 ( \1378 , \1377 , \594 );
xor \U$1064 ( \1379 , \1374 , \1378 );
xor \U$1065 ( \1380 , \1365 , \1379 );
and \U$1066 ( \1381 , \1291 , \1380 );
and \U$1067 ( \1382 , \1153 , \1380 );
or \U$1068 ( \1383 , \1292 , \1381 , \1382 );
and \U$1069 ( \1384 , \1140 , \1144 );
and \U$1070 ( \1385 , \1144 , \1149 );
and \U$1071 ( \1386 , \1140 , \1149 );
or \U$1072 ( \1387 , \1384 , \1385 , \1386 );
and \U$1073 ( \1388 , \1216 , \1220 );
and \U$1074 ( \1389 , \1220 , \1238 );
and \U$1075 ( \1390 , \1216 , \1238 );
or \U$1076 ( \1391 , \1388 , \1389 , \1390 );
xor \U$1077 ( \1392 , \1387 , \1391 );
and \U$1078 ( \1393 , \1181 , \1195 );
and \U$1079 ( \1394 , \1195 , \1210 );
and \U$1080 ( \1395 , \1181 , \1210 );
or \U$1081 ( \1396 , \1393 , \1394 , \1395 );
xor \U$1082 ( \1397 , \1392 , \1396 );
and \U$1083 ( \1398 , \1280 , \1284 );
and \U$1084 ( \1399 , \1284 , \1289 );
and \U$1085 ( \1400 , \1280 , \1289 );
or \U$1086 ( \1401 , \1398 , \1399 , \1400 );
and \U$1087 ( \1402 , \1167 , \1211 );
and \U$1088 ( \1403 , \1211 , \1239 );
and \U$1089 ( \1404 , \1167 , \1239 );
or \U$1090 ( \1405 , \1402 , \1403 , \1404 );
xor \U$1091 ( \1406 , \1401 , \1405 );
and \U$1092 ( \1407 , \1157 , \1161 );
and \U$1093 ( \1408 , \1161 , \1166 );
and \U$1094 ( \1409 , \1157 , \1166 );
or \U$1095 ( \1410 , \1407 , \1408 , \1409 );
and \U$1096 ( \1411 , \1200 , \1204 );
and \U$1097 ( \1412 , \1204 , \1209 );
and \U$1098 ( \1413 , \1200 , \1209 );
or \U$1099 ( \1414 , \1411 , \1412 , \1413 );
xor \U$1100 ( \1415 , \1410 , \1414 );
and \U$1101 ( \1416 , \1185 , \1189 );
and \U$1102 ( \1417 , \1189 , \1194 );
and \U$1103 ( \1418 , \1185 , \1194 );
or \U$1104 ( \1419 , \1416 , \1417 , \1418 );
xor \U$1105 ( \1420 , \1415 , \1419 );
xor \U$1106 ( \1421 , \1406 , \1420 );
and \U$1107 ( \1422 , \1397 , \1421 );
xor \U$1108 ( \1423 , \1383 , \1422 );
and \U$1109 ( \1424 , \1401 , \1405 );
and \U$1110 ( \1425 , \1405 , \1420 );
and \U$1111 ( \1426 , \1401 , \1420 );
or \U$1112 ( \1427 , \1424 , \1425 , \1426 );
and \U$1113 ( \1428 , \1306 , \1320 );
and \U$1114 ( \1429 , \1320 , \1331 );
and \U$1115 ( \1430 , \1306 , \1331 );
or \U$1116 ( \1431 , \1428 , \1429 , \1430 );
and \U$1117 ( \1432 , \699 , \750 );
and \U$1118 ( \1433 , \629 , \748 );
nor \U$1119 ( \1434 , \1432 , \1433 );
xnor \U$1120 ( \1435 , \1434 , \757 );
and \U$1121 ( \1436 , \727 , \776 );
and \U$1122 ( \1437 , \681 , \774 );
nor \U$1123 ( \1438 , \1436 , \1437 );
xnor \U$1124 ( \1439 , \1438 , \783 );
xor \U$1125 ( \1440 , \1435 , \1439 );
and \U$1126 ( \1441 , \752 , \805 );
and \U$1127 ( \1442 , \709 , \803 );
nor \U$1128 ( \1443 , \1441 , \1442 );
xnor \U$1129 ( \1444 , \1443 , \812 );
xor \U$1130 ( \1445 , \1440 , \1444 );
xor \U$1131 ( \1446 , \1431 , \1445 );
and \U$1132 ( \1447 , \568 , \674 );
and \U$1133 ( \1448 , \227 , \671 );
nor \U$1134 ( \1449 , \1447 , \1448 );
xnor \U$1135 ( \1450 , \1449 , \635 );
and \U$1136 ( \1451 , \1055 , \697 );
and \U$1137 ( \1452 , \601 , \695 );
nor \U$1138 ( \1453 , \1451 , \1452 );
xnor \U$1139 ( \1454 , \1453 , \704 );
xor \U$1140 ( \1455 , \1450 , \1454 );
and \U$1141 ( \1456 , \676 , \725 );
and \U$1142 ( \1457 , \1053 , \723 );
nor \U$1143 ( \1458 , \1456 , \1457 );
xnor \U$1144 ( \1459 , \1458 , \732 );
xor \U$1145 ( \1460 , \1455 , \1459 );
xor \U$1146 ( \1461 , \1446 , \1460 );
and \U$1147 ( \1462 , \1410 , \1414 );
and \U$1148 ( \1463 , \1414 , \1419 );
and \U$1149 ( \1464 , \1410 , \1419 );
or \U$1150 ( \1465 , \1462 , \1463 , \1464 );
and \U$1151 ( \1466 , \1369 , \1373 );
and \U$1152 ( \1467 , \1373 , \1378 );
and \U$1153 ( \1468 , \1369 , \1378 );
or \U$1154 ( \1469 , \1466 , \1467 , \1468 );
xor \U$1155 ( \1470 , \1465 , \1469 );
and \U$1156 ( \1471 , \1334 , \1348 );
and \U$1157 ( \1472 , \1348 , \1363 );
and \U$1158 ( \1473 , \1334 , \1363 );
or \U$1159 ( \1474 , \1471 , \1472 , \1473 );
xor \U$1160 ( \1475 , \1470 , \1474 );
xor \U$1161 ( \1476 , \1461 , \1475 );
xor \U$1162 ( \1477 , \1427 , \1476 );
and \U$1163 ( \1478 , \1387 , \1391 );
and \U$1164 ( \1479 , \1391 , \1396 );
and \U$1165 ( \1480 , \1387 , \1396 );
or \U$1166 ( \1481 , \1478 , \1479 , \1480 );
and \U$1167 ( \1482 , \1332 , \1364 );
and \U$1168 ( \1483 , \1364 , \1379 );
and \U$1169 ( \1484 , \1332 , \1379 );
or \U$1170 ( \1485 , \1482 , \1483 , \1484 );
xor \U$1171 ( \1486 , \1481 , \1485 );
and \U$1172 ( \1487 , \940 , \985 );
and \U$1173 ( \1488 , \896 , \983 );
nor \U$1174 ( \1489 , \1487 , \1488 );
xnor \U$1175 ( \1490 , \1489 , \992 );
and \U$1176 ( \1491 , \968 , \1013 );
and \U$1177 ( \1492 , \922 , \996 );
nor \U$1178 ( \1493 , \1491 , \1492 );
xnor \U$1179 ( \1494 , \1493 , \628 );
xor \U$1180 ( \1495 , \1490 , \1494 );
and \U$1181 ( \1496 , \987 , \1233 );
and \U$1182 ( \1497 , \950 , \1114 );
nor \U$1183 ( \1498 , \1496 , \1497 );
xnor \U$1184 ( \1499 , \1498 , \594 );
xor \U$1185 ( \1500 , \1495 , \1499 );
and \U$1186 ( \1501 , \858 , \912 );
and \U$1187 ( \1502 , \814 , \910 );
nor \U$1188 ( \1503 , \1501 , \1502 );
xnor \U$1189 ( \1504 , \1503 , \919 );
and \U$1190 ( \1505 , \889 , \938 );
and \U$1191 ( \1506 , \840 , \936 );
nor \U$1192 ( \1507 , \1505 , \1506 );
xnor \U$1193 ( \1508 , \1507 , \945 );
xor \U$1194 ( \1509 , \1504 , \1508 );
and \U$1195 ( \1510 , \914 , \966 );
and \U$1196 ( \1511 , \871 , \964 );
nor \U$1197 ( \1512 , \1510 , \1511 );
xnor \U$1198 ( \1513 , \1512 , \973 );
xor \U$1199 ( \1514 , \1509 , \1513 );
xor \U$1200 ( \1515 , \1500 , \1514 );
and \U$1201 ( \1516 , \778 , \830 );
and \U$1202 ( \1517 , \734 , \828 );
nor \U$1203 ( \1518 , \1516 , \1517 );
xnor \U$1204 ( \1519 , \1518 , \837 );
and \U$1205 ( \1520 , \807 , \856 );
and \U$1206 ( \1521 , \760 , \854 );
nor \U$1207 ( \1522 , \1520 , \1521 );
xnor \U$1208 ( \1523 , \1522 , \863 );
xor \U$1209 ( \1524 , \1519 , \1523 );
and \U$1210 ( \1525 , \832 , \887 );
and \U$1211 ( \1526 , \789 , \885 );
nor \U$1212 ( \1527 , \1525 , \1526 );
xnor \U$1213 ( \1528 , \1527 , \894 );
xor \U$1214 ( \1529 , \1524 , \1528 );
xor \U$1215 ( \1530 , \1515 , \1529 );
and \U$1216 ( \1531 , \1353 , \1357 );
and \U$1217 ( \1532 , \1357 , \1362 );
and \U$1218 ( \1533 , \1353 , \1362 );
or \U$1219 ( \1534 , \1531 , \1532 , \1533 );
and \U$1220 ( \1535 , \1338 , \1342 );
and \U$1221 ( \1536 , \1342 , \1347 );
and \U$1222 ( \1537 , \1338 , \1347 );
or \U$1223 ( \1538 , \1535 , \1536 , \1537 );
xor \U$1224 ( \1539 , \1534 , \1538 );
and \U$1225 ( \1540 , \995 , \561 );
and \U$1226 ( \1541 , \975 , \559 );
nor \U$1227 ( \1542 , \1540 , \1541 );
xnor \U$1228 ( \1543 , \1542 , \566 );
xor \U$1229 ( \1544 , \1539 , \1543 );
xor \U$1230 ( \1545 , \1530 , \1544 );
and \U$1231 ( \1546 , \566 , \1325 );
and \U$1232 ( \1547 , \1325 , \1330 );
and \U$1233 ( \1548 , \566 , \1330 );
or \U$1234 ( \1549 , \1546 , \1547 , \1548 );
and \U$1235 ( \1550 , \1310 , \1314 );
and \U$1236 ( \1551 , \1314 , \1319 );
and \U$1237 ( \1552 , \1310 , \1319 );
or \U$1238 ( \1553 , \1550 , \1551 , \1552 );
xor \U$1239 ( \1554 , \1549 , \1553 );
and \U$1240 ( \1555 , \1296 , \1300 );
and \U$1241 ( \1556 , \1300 , \1305 );
and \U$1242 ( \1557 , \1296 , \1305 );
or \U$1243 ( \1558 , \1555 , \1556 , \1557 );
xor \U$1244 ( \1559 , \1554 , \1558 );
xor \U$1245 ( \1560 , \1545 , \1559 );
xor \U$1246 ( \1561 , \1486 , \1560 );
xor \U$1247 ( \1562 , \1477 , \1561 );
xor \U$1248 ( \1563 , \1423 , \1562 );
and \U$1249 ( \1564 , \699 , \674 );
and \U$1250 ( \1565 , \629 , \671 );
nor \U$1251 ( \1566 , \1564 , \1565 );
xnor \U$1252 ( \1567 , \1566 , \635 );
and \U$1253 ( \1568 , \727 , \697 );
and \U$1254 ( \1569 , \681 , \695 );
nor \U$1255 ( \1570 , \1568 , \1569 );
xnor \U$1256 ( \1571 , \1570 , \704 );
and \U$1257 ( \1572 , \1567 , \1571 );
and \U$1258 ( \1573 , \752 , \725 );
and \U$1259 ( \1574 , \709 , \723 );
nor \U$1260 ( \1575 , \1573 , \1574 );
xnor \U$1261 ( \1576 , \1575 , \732 );
and \U$1262 ( \1577 , \1571 , \1576 );
and \U$1263 ( \1578 , \1567 , \1576 );
or \U$1264 ( \1579 , \1572 , \1577 , \1578 );
and \U$1265 ( \1580 , \778 , \750 );
and \U$1266 ( \1581 , \734 , \748 );
nor \U$1267 ( \1582 , \1580 , \1581 );
xnor \U$1268 ( \1583 , \1582 , \757 );
and \U$1269 ( \1584 , \807 , \776 );
and \U$1270 ( \1585 , \760 , \774 );
nor \U$1271 ( \1586 , \1584 , \1585 );
xnor \U$1272 ( \1587 , \1586 , \783 );
and \U$1273 ( \1588 , \1583 , \1587 );
and \U$1274 ( \1589 , \832 , \805 );
and \U$1275 ( \1590 , \789 , \803 );
nor \U$1276 ( \1591 , \1589 , \1590 );
xnor \U$1277 ( \1592 , \1591 , \812 );
and \U$1278 ( \1593 , \1587 , \1592 );
and \U$1279 ( \1594 , \1583 , \1592 );
or \U$1280 ( \1595 , \1588 , \1593 , \1594 );
and \U$1281 ( \1596 , \1579 , \1595 );
and \U$1282 ( \1597 , \858 , \830 );
and \U$1283 ( \1598 , \814 , \828 );
nor \U$1284 ( \1599 , \1597 , \1598 );
xnor \U$1285 ( \1600 , \1599 , \837 );
and \U$1286 ( \1601 , \889 , \856 );
and \U$1287 ( \1602 , \840 , \854 );
nor \U$1288 ( \1603 , \1601 , \1602 );
xnor \U$1289 ( \1604 , \1603 , \863 );
and \U$1290 ( \1605 , \1600 , \1604 );
and \U$1291 ( \1606 , \914 , \887 );
and \U$1292 ( \1607 , \871 , \885 );
nor \U$1293 ( \1608 , \1606 , \1607 );
xnor \U$1294 ( \1609 , \1608 , \894 );
and \U$1295 ( \1610 , \1604 , \1609 );
and \U$1296 ( \1611 , \1600 , \1609 );
or \U$1297 ( \1612 , \1605 , \1610 , \1611 );
and \U$1298 ( \1613 , \1595 , \1612 );
and \U$1299 ( \1614 , \1579 , \1612 );
or \U$1300 ( \1615 , \1596 , \1613 , \1614 );
and \U$1301 ( \1616 , \940 , \912 );
and \U$1302 ( \1617 , \896 , \910 );
nor \U$1303 ( \1618 , \1616 , \1617 );
xnor \U$1304 ( \1619 , \1618 , \919 );
and \U$1305 ( \1620 , \968 , \938 );
and \U$1306 ( \1621 , \922 , \936 );
nor \U$1307 ( \1622 , \1620 , \1621 );
xnor \U$1308 ( \1623 , \1622 , \945 );
and \U$1309 ( \1624 , \1619 , \1623 );
and \U$1310 ( \1625 , \987 , \966 );
and \U$1311 ( \1626 , \950 , \964 );
nor \U$1312 ( \1627 , \1625 , \1626 );
xnor \U$1313 ( \1628 , \1627 , \973 );
and \U$1314 ( \1629 , \1623 , \1628 );
and \U$1315 ( \1630 , \1619 , \1628 );
or \U$1316 ( \1631 , \1624 , \1629 , \1630 );
xor \U$1317 ( \1632 , \974 , \993 );
xor \U$1318 ( \1633 , \1632 , \998 );
and \U$1319 ( \1634 , \1631 , \1633 );
xor \U$1320 ( \1635 , \895 , \920 );
xor \U$1321 ( \1636 , \1635 , \946 );
and \U$1322 ( \1637 , \1633 , \1636 );
and \U$1323 ( \1638 , \1631 , \1636 );
or \U$1324 ( \1639 , \1634 , \1637 , \1638 );
and \U$1325 ( \1640 , \1615 , \1639 );
xor \U$1326 ( \1641 , \813 , \838 );
xor \U$1327 ( \1642 , \1641 , \864 );
xor \U$1328 ( \1643 , \733 , \758 );
xor \U$1329 ( \1644 , \1643 , \784 );
and \U$1330 ( \1645 , \1642 , \1644 );
xor \U$1331 ( \1646 , \628 , \679 );
xor \U$1332 ( \1647 , \1646 , \705 );
and \U$1333 ( \1648 , \1644 , \1647 );
and \U$1334 ( \1649 , \1642 , \1647 );
or \U$1335 ( \1650 , \1645 , \1648 , \1649 );
and \U$1336 ( \1651 , \1639 , \1650 );
and \U$1337 ( \1652 , \1615 , \1650 );
or \U$1338 ( \1653 , \1640 , \1651 , \1652 );
xor \U$1339 ( \1654 , \1260 , \1264 );
xor \U$1340 ( \1655 , \1654 , \1269 );
xor \U$1341 ( \1656 , \1244 , \1248 );
xor \U$1342 ( \1657 , \1656 , \1253 );
and \U$1343 ( \1658 , \1655 , \1657 );
xor \U$1344 ( \1659 , \1017 , \1031 );
xor \U$1345 ( \1660 , \1659 , \1046 );
and \U$1346 ( \1661 , \1657 , \1660 );
and \U$1347 ( \1662 , \1655 , \1660 );
or \U$1348 ( \1663 , \1658 , \1661 , \1662 );
and \U$1349 ( \1664 , \1653 , \1663 );
xor \U$1350 ( \1665 , \1256 , \1272 );
xor \U$1351 ( \1666 , \1665 , \1277 );
and \U$1352 ( \1667 , \1663 , \1666 );
and \U$1353 ( \1668 , \1653 , \1666 );
or \U$1354 ( \1669 , \1664 , \1667 , \1668 );
xor \U$1355 ( \1670 , \1240 , \1290 );
and \U$1356 ( \1671 , \1669 , \1670 );
xor \U$1357 ( \1672 , \1052 , \1135 );
xor \U$1358 ( \1673 , \1672 , \1150 );
and \U$1359 ( \1674 , \1670 , \1673 );
and \U$1360 ( \1675 , \1669 , \1673 );
or \U$1361 ( \1676 , \1671 , \1674 , \1675 );
xor \U$1362 ( \1677 , \1397 , \1421 );
and \U$1363 ( \1678 , \1676 , \1677 );
xor \U$1364 ( \1679 , \1153 , \1291 );
xor \U$1365 ( \1680 , \1679 , \1380 );
and \U$1366 ( \1681 , \1677 , \1680 );
and \U$1367 ( \1682 , \1676 , \1680 );
or \U$1368 ( \1683 , \1678 , \1681 , \1682 );
nor \U$1369 ( \1684 , \1563 , \1683 );
and \U$1370 ( \1685 , \1427 , \1476 );
and \U$1371 ( \1686 , \1476 , \1561 );
and \U$1372 ( \1687 , \1427 , \1561 );
or \U$1373 ( \1688 , \1685 , \1686 , \1687 );
and \U$1374 ( \1689 , \1465 , \1469 );
and \U$1375 ( \1690 , \1469 , \1474 );
and \U$1376 ( \1691 , \1465 , \1474 );
or \U$1377 ( \1692 , \1689 , \1690 , \1691 );
and \U$1378 ( \1693 , \1431 , \1445 );
and \U$1379 ( \1694 , \1445 , \1460 );
and \U$1380 ( \1695 , \1431 , \1460 );
or \U$1381 ( \1696 , \1693 , \1694 , \1695 );
xor \U$1382 ( \1697 , \1692 , \1696 );
and \U$1383 ( \1698 , \1530 , \1544 );
and \U$1384 ( \1699 , \1544 , \1559 );
and \U$1385 ( \1700 , \1530 , \1559 );
or \U$1386 ( \1701 , \1698 , \1699 , \1700 );
xor \U$1387 ( \1702 , \1697 , \1701 );
xor \U$1388 ( \1703 , \1688 , \1702 );
and \U$1389 ( \1704 , \1481 , \1485 );
and \U$1390 ( \1705 , \1485 , \1560 );
and \U$1391 ( \1706 , \1481 , \1560 );
or \U$1392 ( \1707 , \1704 , \1705 , \1706 );
and \U$1393 ( \1708 , \1461 , \1475 );
xor \U$1394 ( \1709 , \1707 , \1708 );
and \U$1395 ( \1710 , \1504 , \1508 );
and \U$1396 ( \1711 , \1508 , \1513 );
and \U$1397 ( \1712 , \1504 , \1513 );
or \U$1398 ( \1713 , \1710 , \1711 , \1712 );
and \U$1399 ( \1714 , \1490 , \1494 );
and \U$1400 ( \1715 , \1494 , \1499 );
and \U$1401 ( \1716 , \1490 , \1499 );
or \U$1402 ( \1717 , \1714 , \1715 , \1716 );
xor \U$1403 ( \1718 , \1713 , \1717 );
and \U$1404 ( \1719 , \950 , \1233 );
and \U$1405 ( \1720 , \968 , \1114 );
nor \U$1406 ( \1721 , \1719 , \1720 );
xnor \U$1407 ( \1722 , \1721 , \594 );
and \U$1408 ( \1723 , \975 , \561 );
and \U$1409 ( \1724 , \987 , \559 );
nor \U$1410 ( \1725 , \1723 , \1724 );
xnor \U$1411 ( \1726 , \1725 , \566 );
xor \U$1412 ( \1727 , \1722 , \1726 );
nand \U$1413 ( \1728 , \995 , \569 );
not \U$1414 ( \1729 , \1728 );
xor \U$1415 ( \1730 , \1727 , \1729 );
xor \U$1416 ( \1731 , \1718 , \1730 );
and \U$1417 ( \1732 , \1450 , \1454 );
and \U$1418 ( \1733 , \1454 , \1459 );
and \U$1419 ( \1734 , \1450 , \1459 );
or \U$1420 ( \1735 , \1732 , \1733 , \1734 );
and \U$1421 ( \1736 , \1435 , \1439 );
and \U$1422 ( \1737 , \1439 , \1444 );
and \U$1423 ( \1738 , \1435 , \1444 );
or \U$1424 ( \1739 , \1736 , \1737 , \1738 );
xor \U$1425 ( \1740 , \1735 , \1739 );
and \U$1426 ( \1741 , \1519 , \1523 );
and \U$1427 ( \1742 , \1523 , \1528 );
and \U$1428 ( \1743 , \1519 , \1528 );
or \U$1429 ( \1744 , \1741 , \1742 , \1743 );
xor \U$1430 ( \1745 , \1740 , \1744 );
xor \U$1431 ( \1746 , \1731 , \1745 );
and \U$1432 ( \1747 , \1053 , \725 );
and \U$1433 ( \1748 , \1055 , \723 );
nor \U$1434 ( \1749 , \1747 , \1748 );
xnor \U$1435 ( \1750 , \1749 , \732 );
and \U$1436 ( \1751 , \629 , \750 );
and \U$1437 ( \1752 , \676 , \748 );
nor \U$1438 ( \1753 , \1751 , \1752 );
xnor \U$1439 ( \1754 , \1753 , \757 );
xor \U$1440 ( \1755 , \1750 , \1754 );
and \U$1441 ( \1756 , \681 , \776 );
and \U$1442 ( \1757 , \699 , \774 );
nor \U$1443 ( \1758 , \1756 , \1757 );
xnor \U$1444 ( \1759 , \1758 , \783 );
xor \U$1445 ( \1760 , \1755 , \1759 );
and \U$1446 ( \1761 , \227 , \674 );
not \U$1447 ( \1762 , \1761 );
xnor \U$1448 ( \1763 , \1762 , \635 );
and \U$1449 ( \1764 , \601 , \697 );
and \U$1450 ( \1765 , \568 , \695 );
nor \U$1451 ( \1766 , \1764 , \1765 );
xnor \U$1452 ( \1767 , \1766 , \704 );
xor \U$1453 ( \1768 , \1763 , \1767 );
xor \U$1454 ( \1769 , \1760 , \1768 );
and \U$1455 ( \1770 , \871 , \966 );
and \U$1456 ( \1771 , \889 , \964 );
nor \U$1457 ( \1772 , \1770 , \1771 );
xnor \U$1458 ( \1773 , \1772 , \973 );
and \U$1459 ( \1774 , \896 , \985 );
and \U$1460 ( \1775 , \914 , \983 );
nor \U$1461 ( \1776 , \1774 , \1775 );
xnor \U$1462 ( \1777 , \1776 , \992 );
xor \U$1463 ( \1778 , \1773 , \1777 );
and \U$1464 ( \1779 , \922 , \1013 );
and \U$1465 ( \1780 , \940 , \996 );
nor \U$1466 ( \1781 , \1779 , \1780 );
xnor \U$1467 ( \1782 , \1781 , \628 );
xor \U$1468 ( \1783 , \1778 , \1782 );
and \U$1469 ( \1784 , \789 , \887 );
and \U$1470 ( \1785 , \807 , \885 );
nor \U$1471 ( \1786 , \1784 , \1785 );
xnor \U$1472 ( \1787 , \1786 , \894 );
and \U$1473 ( \1788 , \814 , \912 );
and \U$1474 ( \1789 , \832 , \910 );
nor \U$1475 ( \1790 , \1788 , \1789 );
xnor \U$1476 ( \1791 , \1790 , \919 );
xor \U$1477 ( \1792 , \1787 , \1791 );
and \U$1478 ( \1793 , \840 , \938 );
and \U$1479 ( \1794 , \858 , \936 );
nor \U$1480 ( \1795 , \1793 , \1794 );
xnor \U$1481 ( \1796 , \1795 , \945 );
xor \U$1482 ( \1797 , \1792 , \1796 );
xor \U$1483 ( \1798 , \1783 , \1797 );
and \U$1484 ( \1799 , \709 , \805 );
and \U$1485 ( \1800 , \727 , \803 );
nor \U$1486 ( \1801 , \1799 , \1800 );
xnor \U$1487 ( \1802 , \1801 , \812 );
and \U$1488 ( \1803 , \734 , \830 );
and \U$1489 ( \1804 , \752 , \828 );
nor \U$1490 ( \1805 , \1803 , \1804 );
xnor \U$1491 ( \1806 , \1805 , \837 );
xor \U$1492 ( \1807 , \1802 , \1806 );
and \U$1493 ( \1808 , \760 , \856 );
and \U$1494 ( \1809 , \778 , \854 );
nor \U$1495 ( \1810 , \1808 , \1809 );
xnor \U$1496 ( \1811 , \1810 , \863 );
xor \U$1497 ( \1812 , \1807 , \1811 );
xor \U$1498 ( \1813 , \1798 , \1812 );
xor \U$1499 ( \1814 , \1769 , \1813 );
xor \U$1500 ( \1815 , \1746 , \1814 );
and \U$1501 ( \1816 , \1549 , \1553 );
and \U$1502 ( \1817 , \1553 , \1558 );
and \U$1503 ( \1818 , \1549 , \1558 );
or \U$1504 ( \1819 , \1816 , \1817 , \1818 );
and \U$1505 ( \1820 , \1534 , \1538 );
and \U$1506 ( \1821 , \1538 , \1543 );
and \U$1507 ( \1822 , \1534 , \1543 );
or \U$1508 ( \1823 , \1820 , \1821 , \1822 );
xor \U$1509 ( \1824 , \1819 , \1823 );
and \U$1510 ( \1825 , \1500 , \1514 );
and \U$1511 ( \1826 , \1514 , \1529 );
and \U$1512 ( \1827 , \1500 , \1529 );
or \U$1513 ( \1828 , \1825 , \1826 , \1827 );
xor \U$1514 ( \1829 , \1824 , \1828 );
xor \U$1515 ( \1830 , \1815 , \1829 );
xor \U$1516 ( \1831 , \1709 , \1830 );
xor \U$1517 ( \1832 , \1703 , \1831 );
and \U$1518 ( \1833 , \1383 , \1422 );
and \U$1519 ( \1834 , \1422 , \1562 );
and \U$1520 ( \1835 , \1383 , \1562 );
or \U$1521 ( \1836 , \1833 , \1834 , \1835 );
nor \U$1522 ( \1837 , \1832 , \1836 );
nor \U$1523 ( \1838 , \1684 , \1837 );
and \U$1524 ( \1839 , \1707 , \1708 );
and \U$1525 ( \1840 , \1708 , \1830 );
and \U$1526 ( \1841 , \1707 , \1830 );
or \U$1527 ( \1842 , \1839 , \1840 , \1841 );
and \U$1528 ( \1843 , \1819 , \1823 );
and \U$1529 ( \1844 , \1823 , \1828 );
and \U$1530 ( \1845 , \1819 , \1828 );
or \U$1531 ( \1846 , \1843 , \1844 , \1845 );
and \U$1532 ( \1847 , \1760 , \1768 );
and \U$1533 ( \1848 , \1768 , \1813 );
and \U$1534 ( \1849 , \1760 , \1813 );
or \U$1535 ( \1850 , \1847 , \1848 , \1849 );
xor \U$1536 ( \1851 , \1846 , \1850 );
and \U$1537 ( \1852 , \1731 , \1745 );
xor \U$1538 ( \1853 , \1851 , \1852 );
xor \U$1539 ( \1854 , \1842 , \1853 );
and \U$1540 ( \1855 , \1692 , \1696 );
and \U$1541 ( \1856 , \1696 , \1701 );
and \U$1542 ( \1857 , \1692 , \1701 );
or \U$1543 ( \1858 , \1855 , \1856 , \1857 );
and \U$1544 ( \1859 , \1746 , \1814 );
and \U$1545 ( \1860 , \1814 , \1829 );
and \U$1546 ( \1861 , \1746 , \1829 );
or \U$1547 ( \1862 , \1859 , \1860 , \1861 );
xor \U$1548 ( \1863 , \1858 , \1862 );
and \U$1549 ( \1864 , \1763 , \1767 );
and \U$1550 ( \1865 , \1750 , \1754 );
and \U$1551 ( \1866 , \1754 , \1759 );
and \U$1552 ( \1867 , \1750 , \1759 );
or \U$1553 ( \1868 , \1865 , \1866 , \1867 );
xor \U$1554 ( \1869 , \1864 , \1868 );
and \U$1555 ( \1870 , \1802 , \1806 );
and \U$1556 ( \1871 , \1806 , \1811 );
and \U$1557 ( \1872 , \1802 , \1811 );
or \U$1558 ( \1873 , \1870 , \1871 , \1872 );
xor \U$1559 ( \1874 , \1869 , \1873 );
and \U$1560 ( \1875 , \752 , \830 );
and \U$1561 ( \1876 , \709 , \828 );
nor \U$1562 ( \1877 , \1875 , \1876 );
xnor \U$1563 ( \1878 , \1877 , \837 );
and \U$1564 ( \1879 , \778 , \856 );
and \U$1565 ( \1880 , \734 , \854 );
nor \U$1566 ( \1881 , \1879 , \1880 );
xnor \U$1567 ( \1882 , \1881 , \863 );
xor \U$1568 ( \1883 , \1878 , \1882 );
and \U$1569 ( \1884 , \807 , \887 );
and \U$1570 ( \1885 , \760 , \885 );
nor \U$1571 ( \1886 , \1884 , \1885 );
xnor \U$1572 ( \1887 , \1886 , \894 );
xor \U$1573 ( \1888 , \1883 , \1887 );
and \U$1574 ( \1889 , \676 , \750 );
and \U$1575 ( \1890 , \1053 , \748 );
nor \U$1576 ( \1891 , \1889 , \1890 );
xnor \U$1577 ( \1892 , \1891 , \757 );
and \U$1578 ( \1893 , \699 , \776 );
and \U$1579 ( \1894 , \629 , \774 );
nor \U$1580 ( \1895 , \1893 , \1894 );
xnor \U$1581 ( \1896 , \1895 , \783 );
xor \U$1582 ( \1897 , \1892 , \1896 );
and \U$1583 ( \1898 , \727 , \805 );
and \U$1584 ( \1899 , \681 , \803 );
nor \U$1585 ( \1900 , \1898 , \1899 );
xnor \U$1586 ( \1901 , \1900 , \812 );
xor \U$1587 ( \1902 , \1897 , \1901 );
xor \U$1588 ( \1903 , \1888 , \1902 );
not \U$1589 ( \1904 , \635 );
and \U$1590 ( \1905 , \568 , \697 );
and \U$1591 ( \1906 , \227 , \695 );
nor \U$1592 ( \1907 , \1905 , \1906 );
xnor \U$1593 ( \1908 , \1907 , \704 );
xor \U$1594 ( \1909 , \1904 , \1908 );
and \U$1595 ( \1910 , \1055 , \725 );
and \U$1596 ( \1911 , \601 , \723 );
nor \U$1597 ( \1912 , \1910 , \1911 );
xnor \U$1598 ( \1913 , \1912 , \732 );
xor \U$1599 ( \1914 , \1909 , \1913 );
xor \U$1600 ( \1915 , \1903 , \1914 );
and \U$1601 ( \1916 , \987 , \561 );
and \U$1602 ( \1917 , \950 , \559 );
nor \U$1603 ( \1918 , \1916 , \1917 );
xnor \U$1604 ( \1919 , \1918 , \566 );
and \U$1606 ( \1920 , \975 , \569 );
nor \U$1607 ( \1921 , 1'b0 , \1920 );
not \U$1608 ( \1922 , \1921 );
xnor \U$1609 ( \1923 , \1919 , \1922 );
and \U$1610 ( \1924 , \914 , \985 );
and \U$1611 ( \1925 , \871 , \983 );
nor \U$1612 ( \1926 , \1924 , \1925 );
xnor \U$1613 ( \1927 , \1926 , \992 );
and \U$1614 ( \1928 , \940 , \1013 );
and \U$1615 ( \1929 , \896 , \996 );
nor \U$1616 ( \1930 , \1928 , \1929 );
xnor \U$1617 ( \1931 , \1930 , \628 );
xor \U$1618 ( \1932 , \1927 , \1931 );
and \U$1619 ( \1933 , \968 , \1233 );
and \U$1620 ( \1934 , \922 , \1114 );
nor \U$1621 ( \1935 , \1933 , \1934 );
xnor \U$1622 ( \1936 , \1935 , \594 );
xor \U$1623 ( \1937 , \1932 , \1936 );
xor \U$1624 ( \1938 , \1923 , \1937 );
and \U$1625 ( \1939 , \832 , \912 );
and \U$1626 ( \1940 , \789 , \910 );
nor \U$1627 ( \1941 , \1939 , \1940 );
xnor \U$1628 ( \1942 , \1941 , \919 );
and \U$1629 ( \1943 , \858 , \938 );
and \U$1630 ( \1944 , \814 , \936 );
nor \U$1631 ( \1945 , \1943 , \1944 );
xnor \U$1632 ( \1946 , \1945 , \945 );
xor \U$1633 ( \1947 , \1942 , \1946 );
and \U$1634 ( \1948 , \889 , \966 );
and \U$1635 ( \1949 , \840 , \964 );
nor \U$1636 ( \1950 , \1948 , \1949 );
xnor \U$1637 ( \1951 , \1950 , \973 );
xor \U$1638 ( \1952 , \1947 , \1951 );
xor \U$1639 ( \1953 , \1938 , \1952 );
xor \U$1640 ( \1954 , \1915 , \1953 );
and \U$1641 ( \1955 , \1787 , \1791 );
and \U$1642 ( \1956 , \1791 , \1796 );
and \U$1643 ( \1957 , \1787 , \1796 );
or \U$1644 ( \1958 , \1955 , \1956 , \1957 );
and \U$1645 ( \1959 , \1773 , \1777 );
and \U$1646 ( \1960 , \1777 , \1782 );
and \U$1647 ( \1961 , \1773 , \1782 );
or \U$1648 ( \1962 , \1959 , \1960 , \1961 );
xor \U$1649 ( \1963 , \1958 , \1962 );
and \U$1650 ( \1964 , \1722 , \1726 );
and \U$1651 ( \1965 , \1726 , \1729 );
and \U$1652 ( \1966 , \1722 , \1729 );
or \U$1653 ( \1967 , \1964 , \1965 , \1966 );
xor \U$1654 ( \1968 , \1963 , \1967 );
xor \U$1655 ( \1969 , \1954 , \1968 );
xor \U$1656 ( \1970 , \1874 , \1969 );
and \U$1657 ( \1971 , \1735 , \1739 );
and \U$1658 ( \1972 , \1739 , \1744 );
and \U$1659 ( \1973 , \1735 , \1744 );
or \U$1660 ( \1974 , \1971 , \1972 , \1973 );
and \U$1661 ( \1975 , \1713 , \1717 );
and \U$1662 ( \1976 , \1717 , \1730 );
and \U$1663 ( \1977 , \1713 , \1730 );
or \U$1664 ( \1978 , \1975 , \1976 , \1977 );
xor \U$1665 ( \1979 , \1974 , \1978 );
and \U$1666 ( \1980 , \1783 , \1797 );
and \U$1667 ( \1981 , \1797 , \1812 );
and \U$1668 ( \1982 , \1783 , \1812 );
or \U$1669 ( \1983 , \1980 , \1981 , \1982 );
xor \U$1670 ( \1984 , \1979 , \1983 );
xor \U$1671 ( \1985 , \1970 , \1984 );
xor \U$1672 ( \1986 , \1863 , \1985 );
xor \U$1673 ( \1987 , \1854 , \1986 );
and \U$1674 ( \1988 , \1688 , \1702 );
and \U$1675 ( \1989 , \1702 , \1831 );
and \U$1676 ( \1990 , \1688 , \1831 );
or \U$1677 ( \1991 , \1988 , \1989 , \1990 );
nor \U$1678 ( \1992 , \1987 , \1991 );
and \U$1679 ( \1993 , \1858 , \1862 );
and \U$1680 ( \1994 , \1862 , \1985 );
and \U$1681 ( \1995 , \1858 , \1985 );
or \U$1682 ( \1996 , \1993 , \1994 , \1995 );
and \U$1683 ( \1997 , \1974 , \1978 );
and \U$1684 ( \1998 , \1978 , \1983 );
and \U$1685 ( \1999 , \1974 , \1983 );
or \U$1686 ( \2000 , \1997 , \1998 , \1999 );
and \U$1687 ( \2001 , \1915 , \1953 );
and \U$1688 ( \2002 , \1953 , \1968 );
and \U$1689 ( \2003 , \1915 , \1968 );
or \U$1690 ( \2004 , \2001 , \2002 , \2003 );
xor \U$1691 ( \2005 , \2000 , \2004 );
and \U$1692 ( \2006 , \1942 , \1946 );
and \U$1693 ( \2007 , \1946 , \1951 );
and \U$1694 ( \2008 , \1942 , \1951 );
or \U$1695 ( \2009 , \2006 , \2007 , \2008 );
and \U$1696 ( \2010 , \1927 , \1931 );
and \U$1697 ( \2011 , \1931 , \1936 );
and \U$1698 ( \2012 , \1927 , \1936 );
or \U$1699 ( \2013 , \2010 , \2011 , \2012 );
xor \U$1700 ( \2014 , \2009 , \2013 );
or \U$1701 ( \2015 , \1919 , \1922 );
xor \U$1702 ( \2016 , \2014 , \2015 );
xor \U$1703 ( \2017 , \2005 , \2016 );
xor \U$1704 ( \2018 , \1996 , \2017 );
and \U$1705 ( \2019 , \1846 , \1850 );
and \U$1706 ( \2020 , \1850 , \1852 );
and \U$1707 ( \2021 , \1846 , \1852 );
or \U$1708 ( \2022 , \2019 , \2020 , \2021 );
and \U$1709 ( \2023 , \1874 , \1969 );
and \U$1710 ( \2024 , \1969 , \1984 );
and \U$1711 ( \2025 , \1874 , \1984 );
or \U$1712 ( \2026 , \2023 , \2024 , \2025 );
xor \U$1713 ( \2027 , \2022 , \2026 );
and \U$1714 ( \2028 , \1904 , \1908 );
and \U$1715 ( \2029 , \1908 , \1913 );
and \U$1716 ( \2030 , \1904 , \1913 );
or \U$1717 ( \2031 , \2028 , \2029 , \2030 );
and \U$1718 ( \2032 , \1892 , \1896 );
and \U$1719 ( \2033 , \1896 , \1901 );
and \U$1720 ( \2034 , \1892 , \1901 );
or \U$1721 ( \2035 , \2032 , \2033 , \2034 );
xor \U$1722 ( \2036 , \2031 , \2035 );
and \U$1723 ( \2037 , \1878 , \1882 );
and \U$1724 ( \2038 , \1882 , \1887 );
and \U$1725 ( \2039 , \1878 , \1887 );
or \U$1726 ( \2040 , \2037 , \2038 , \2039 );
xor \U$1727 ( \2041 , \2036 , \2040 );
and \U$1728 ( \2042 , \1888 , \1902 );
and \U$1729 ( \2043 , \1902 , \1914 );
and \U$1730 ( \2044 , \1888 , \1914 );
or \U$1731 ( \2045 , \2042 , \2043 , \2044 );
and \U$1732 ( \2046 , \734 , \856 );
and \U$1733 ( \2047 , \752 , \854 );
nor \U$1734 ( \2048 , \2046 , \2047 );
xnor \U$1735 ( \2049 , \2048 , \863 );
and \U$1736 ( \2050 , \760 , \887 );
and \U$1737 ( \2051 , \778 , \885 );
nor \U$1738 ( \2052 , \2050 , \2051 );
xnor \U$1739 ( \2053 , \2052 , \894 );
xor \U$1740 ( \2054 , \2049 , \2053 );
and \U$1741 ( \2055 , \789 , \912 );
and \U$1742 ( \2056 , \807 , \910 );
nor \U$1743 ( \2057 , \2055 , \2056 );
xnor \U$1744 ( \2058 , \2057 , \919 );
xor \U$1745 ( \2059 , \2054 , \2058 );
and \U$1746 ( \2060 , \629 , \776 );
and \U$1747 ( \2061 , \676 , \774 );
nor \U$1748 ( \2062 , \2060 , \2061 );
xnor \U$1749 ( \2063 , \2062 , \783 );
and \U$1750 ( \2064 , \681 , \805 );
and \U$1751 ( \2065 , \699 , \803 );
nor \U$1752 ( \2066 , \2064 , \2065 );
xnor \U$1753 ( \2067 , \2066 , \812 );
xor \U$1754 ( \2068 , \2063 , \2067 );
and \U$1755 ( \2069 , \709 , \830 );
and \U$1756 ( \2070 , \727 , \828 );
nor \U$1757 ( \2071 , \2069 , \2070 );
xnor \U$1758 ( \2072 , \2071 , \837 );
xor \U$1759 ( \2073 , \2068 , \2072 );
xor \U$1760 ( \2074 , \2059 , \2073 );
and \U$1761 ( \2075 , \227 , \697 );
not \U$1762 ( \2076 , \2075 );
xnor \U$1763 ( \2077 , \2076 , \704 );
and \U$1764 ( \2078 , \601 , \725 );
and \U$1765 ( \2079 , \568 , \723 );
nor \U$1766 ( \2080 , \2078 , \2079 );
xnor \U$1767 ( \2081 , \2080 , \732 );
xor \U$1768 ( \2082 , \2077 , \2081 );
and \U$1769 ( \2083 , \1053 , \750 );
and \U$1770 ( \2084 , \1055 , \748 );
nor \U$1771 ( \2085 , \2083 , \2084 );
xnor \U$1772 ( \2086 , \2085 , \757 );
xor \U$1773 ( \2087 , \2082 , \2086 );
xor \U$1774 ( \2088 , \2074 , \2087 );
xor \U$1775 ( \2089 , \2045 , \2088 );
and \U$1777 ( \2090 , \987 , \569 );
nor \U$1778 ( \2091 , 1'b0 , \2090 );
and \U$1779 ( \2092 , \896 , \1013 );
and \U$1780 ( \2093 , \914 , \996 );
nor \U$1781 ( \2094 , \2092 , \2093 );
xnor \U$1782 ( \2095 , \2094 , \628 );
and \U$1783 ( \2096 , \922 , \1233 );
and \U$1784 ( \2097 , \940 , \1114 );
nor \U$1785 ( \2098 , \2096 , \2097 );
xnor \U$1786 ( \2099 , \2098 , \594 );
xor \U$1787 ( \2100 , \2095 , \2099 );
and \U$1788 ( \2101 , \950 , \561 );
and \U$1789 ( \2102 , \968 , \559 );
nor \U$1790 ( \2103 , \2101 , \2102 );
xnor \U$1791 ( \2104 , \2103 , \566 );
xor \U$1792 ( \2105 , \2100 , \2104 );
xor \U$1793 ( \2106 , \2091 , \2105 );
and \U$1794 ( \2107 , \814 , \938 );
and \U$1795 ( \2108 , \832 , \936 );
nor \U$1796 ( \2109 , \2107 , \2108 );
xnor \U$1797 ( \2110 , \2109 , \945 );
and \U$1798 ( \2111 , \840 , \966 );
and \U$1799 ( \2112 , \858 , \964 );
nor \U$1800 ( \2113 , \2111 , \2112 );
xnor \U$1801 ( \2114 , \2113 , \973 );
xor \U$1802 ( \2115 , \2110 , \2114 );
and \U$1803 ( \2116 , \871 , \985 );
and \U$1804 ( \2117 , \889 , \983 );
nor \U$1805 ( \2118 , \2116 , \2117 );
xnor \U$1806 ( \2119 , \2118 , \992 );
xor \U$1807 ( \2120 , \2115 , \2119 );
xor \U$1808 ( \2121 , \2106 , \2120 );
xor \U$1809 ( \2122 , \2089 , \2121 );
xor \U$1810 ( \2123 , \2041 , \2122 );
and \U$1811 ( \2124 , \1864 , \1868 );
and \U$1812 ( \2125 , \1868 , \1873 );
and \U$1813 ( \2126 , \1864 , \1873 );
or \U$1814 ( \2127 , \2124 , \2125 , \2126 );
and \U$1815 ( \2128 , \1958 , \1962 );
and \U$1816 ( \2129 , \1962 , \1967 );
and \U$1817 ( \2130 , \1958 , \1967 );
or \U$1818 ( \2131 , \2128 , \2129 , \2130 );
xor \U$1819 ( \2132 , \2127 , \2131 );
and \U$1820 ( \2133 , \1923 , \1937 );
and \U$1821 ( \2134 , \1937 , \1952 );
and \U$1822 ( \2135 , \1923 , \1952 );
or \U$1823 ( \2136 , \2133 , \2134 , \2135 );
xor \U$1824 ( \2137 , \2132 , \2136 );
xor \U$1825 ( \2138 , \2123 , \2137 );
xor \U$1826 ( \2139 , \2027 , \2138 );
xor \U$1827 ( \2140 , \2018 , \2139 );
and \U$1828 ( \2141 , \1842 , \1853 );
and \U$1829 ( \2142 , \1853 , \1986 );
and \U$1830 ( \2143 , \1842 , \1986 );
or \U$1831 ( \2144 , \2141 , \2142 , \2143 );
nor \U$1832 ( \2145 , \2140 , \2144 );
nor \U$1833 ( \2146 , \1992 , \2145 );
nand \U$1834 ( \2147 , \1838 , \2146 );
and \U$1835 ( \2148 , \2022 , \2026 );
and \U$1836 ( \2149 , \2026 , \2138 );
and \U$1837 ( \2150 , \2022 , \2138 );
or \U$1838 ( \2151 , \2148 , \2149 , \2150 );
and \U$1839 ( \2152 , \2127 , \2131 );
and \U$1840 ( \2153 , \2131 , \2136 );
and \U$1841 ( \2154 , \2127 , \2136 );
or \U$1842 ( \2155 , \2152 , \2153 , \2154 );
and \U$1843 ( \2156 , \2045 , \2088 );
and \U$1844 ( \2157 , \2088 , \2121 );
and \U$1845 ( \2158 , \2045 , \2121 );
or \U$1846 ( \2159 , \2156 , \2157 , \2158 );
xor \U$1847 ( \2160 , \2155 , \2159 );
and \U$1848 ( \2161 , \2110 , \2114 );
and \U$1849 ( \2162 , \2114 , \2119 );
and \U$1850 ( \2163 , \2110 , \2119 );
or \U$1851 ( \2164 , \2161 , \2162 , \2163 );
and \U$1852 ( \2165 , \2095 , \2099 );
and \U$1853 ( \2166 , \2099 , \2104 );
and \U$1854 ( \2167 , \2095 , \2104 );
or \U$1855 ( \2168 , \2165 , \2166 , \2167 );
xor \U$1856 ( \2169 , \2164 , \2168 );
not \U$1857 ( \2170 , \2091 );
xor \U$1858 ( \2171 , \2169 , \2170 );
xor \U$1859 ( \2172 , \2160 , \2171 );
xor \U$1860 ( \2173 , \2151 , \2172 );
and \U$1861 ( \2174 , \2000 , \2004 );
and \U$1862 ( \2175 , \2004 , \2016 );
and \U$1863 ( \2176 , \2000 , \2016 );
or \U$1864 ( \2177 , \2174 , \2175 , \2176 );
and \U$1865 ( \2178 , \2041 , \2122 );
and \U$1866 ( \2179 , \2122 , \2137 );
and \U$1867 ( \2180 , \2041 , \2137 );
or \U$1868 ( \2181 , \2178 , \2179 , \2180 );
xor \U$1869 ( \2182 , \2177 , \2181 );
and \U$1870 ( \2183 , \2077 , \2081 );
and \U$1871 ( \2184 , \2081 , \2086 );
and \U$1872 ( \2185 , \2077 , \2086 );
or \U$1873 ( \2186 , \2183 , \2184 , \2185 );
and \U$1874 ( \2187 , \2063 , \2067 );
and \U$1875 ( \2188 , \2067 , \2072 );
and \U$1876 ( \2189 , \2063 , \2072 );
or \U$1877 ( \2190 , \2187 , \2188 , \2189 );
xor \U$1878 ( \2191 , \2186 , \2190 );
and \U$1879 ( \2192 , \2049 , \2053 );
and \U$1880 ( \2193 , \2053 , \2058 );
and \U$1881 ( \2194 , \2049 , \2058 );
or \U$1882 ( \2195 , \2192 , \2193 , \2194 );
xor \U$1883 ( \2196 , \2191 , \2195 );
and \U$1884 ( \2197 , \2059 , \2073 );
and \U$1885 ( \2198 , \2073 , \2087 );
and \U$1886 ( \2199 , \2059 , \2087 );
or \U$1887 ( \2200 , \2197 , \2198 , \2199 );
and \U$1888 ( \2201 , \752 , \856 );
and \U$1889 ( \2202 , \709 , \854 );
nor \U$1890 ( \2203 , \2201 , \2202 );
xnor \U$1891 ( \2204 , \2203 , \863 );
and \U$1892 ( \2205 , \778 , \887 );
and \U$1893 ( \2206 , \734 , \885 );
nor \U$1894 ( \2207 , \2205 , \2206 );
xnor \U$1895 ( \2208 , \2207 , \894 );
xor \U$1896 ( \2209 , \2204 , \2208 );
and \U$1897 ( \2210 , \807 , \912 );
and \U$1898 ( \2211 , \760 , \910 );
nor \U$1899 ( \2212 , \2210 , \2211 );
xnor \U$1900 ( \2213 , \2212 , \919 );
xor \U$1901 ( \2214 , \2209 , \2213 );
and \U$1902 ( \2215 , \676 , \776 );
and \U$1903 ( \2216 , \1053 , \774 );
nor \U$1904 ( \2217 , \2215 , \2216 );
xnor \U$1905 ( \2218 , \2217 , \783 );
and \U$1906 ( \2219 , \699 , \805 );
and \U$1907 ( \2220 , \629 , \803 );
nor \U$1908 ( \2221 , \2219 , \2220 );
xnor \U$1909 ( \2222 , \2221 , \812 );
xor \U$1910 ( \2223 , \2218 , \2222 );
and \U$1911 ( \2224 , \727 , \830 );
and \U$1912 ( \2225 , \681 , \828 );
nor \U$1913 ( \2226 , \2224 , \2225 );
xnor \U$1914 ( \2227 , \2226 , \837 );
xor \U$1915 ( \2228 , \2223 , \2227 );
xor \U$1916 ( \2229 , \2214 , \2228 );
not \U$1917 ( \2230 , \704 );
and \U$1918 ( \2231 , \568 , \725 );
and \U$1919 ( \2232 , \227 , \723 );
nor \U$1920 ( \2233 , \2231 , \2232 );
xnor \U$1921 ( \2234 , \2233 , \732 );
xor \U$1922 ( \2235 , \2230 , \2234 );
and \U$1923 ( \2236 , \1055 , \750 );
and \U$1924 ( \2237 , \601 , \748 );
nor \U$1925 ( \2238 , \2236 , \2237 );
xnor \U$1926 ( \2239 , \2238 , \757 );
xor \U$1927 ( \2240 , \2235 , \2239 );
xor \U$1928 ( \2241 , \2229 , \2240 );
xor \U$1929 ( \2242 , \2200 , \2241 );
and \U$1931 ( \2243 , \950 , \569 );
nor \U$1932 ( \2244 , 1'b0 , \2243 );
not \U$1933 ( \2245 , \2244 );
and \U$1934 ( \2246 , \914 , \1013 );
and \U$1935 ( \2247 , \871 , \996 );
nor \U$1936 ( \2248 , \2246 , \2247 );
xnor \U$1937 ( \2249 , \2248 , \628 );
and \U$1938 ( \2250 , \940 , \1233 );
and \U$1939 ( \2251 , \896 , \1114 );
nor \U$1940 ( \2252 , \2250 , \2251 );
xnor \U$1941 ( \2253 , \2252 , \594 );
xor \U$1942 ( \2254 , \2249 , \2253 );
and \U$1943 ( \2255 , \968 , \561 );
and \U$1944 ( \2256 , \922 , \559 );
nor \U$1945 ( \2257 , \2255 , \2256 );
xnor \U$1946 ( \2258 , \2257 , \566 );
xor \U$1947 ( \2259 , \2254 , \2258 );
xor \U$1948 ( \2260 , \2245 , \2259 );
and \U$1949 ( \2261 , \832 , \938 );
and \U$1950 ( \2262 , \789 , \936 );
nor \U$1951 ( \2263 , \2261 , \2262 );
xnor \U$1952 ( \2264 , \2263 , \945 );
and \U$1953 ( \2265 , \858 , \966 );
and \U$1954 ( \2266 , \814 , \964 );
nor \U$1955 ( \2267 , \2265 , \2266 );
xnor \U$1956 ( \2268 , \2267 , \973 );
xor \U$1957 ( \2269 , \2264 , \2268 );
and \U$1958 ( \2270 , \889 , \985 );
and \U$1959 ( \2271 , \840 , \983 );
nor \U$1960 ( \2272 , \2270 , \2271 );
xnor \U$1961 ( \2273 , \2272 , \992 );
xor \U$1962 ( \2274 , \2269 , \2273 );
xor \U$1963 ( \2275 , \2260 , \2274 );
xor \U$1964 ( \2276 , \2242 , \2275 );
xor \U$1965 ( \2277 , \2196 , \2276 );
and \U$1966 ( \2278 , \2031 , \2035 );
and \U$1967 ( \2279 , \2035 , \2040 );
and \U$1968 ( \2280 , \2031 , \2040 );
or \U$1969 ( \2281 , \2278 , \2279 , \2280 );
and \U$1970 ( \2282 , \2009 , \2013 );
and \U$1971 ( \2283 , \2013 , \2015 );
and \U$1972 ( \2284 , \2009 , \2015 );
or \U$1973 ( \2285 , \2282 , \2283 , \2284 );
xor \U$1974 ( \2286 , \2281 , \2285 );
and \U$1975 ( \2287 , \2091 , \2105 );
and \U$1976 ( \2288 , \2105 , \2120 );
and \U$1977 ( \2289 , \2091 , \2120 );
or \U$1978 ( \2290 , \2287 , \2288 , \2289 );
xor \U$1979 ( \2291 , \2286 , \2290 );
xor \U$1980 ( \2292 , \2277 , \2291 );
xor \U$1981 ( \2293 , \2182 , \2292 );
xor \U$1982 ( \2294 , \2173 , \2293 );
and \U$1983 ( \2295 , \1996 , \2017 );
and \U$1984 ( \2296 , \2017 , \2139 );
and \U$1985 ( \2297 , \1996 , \2139 );
or \U$1986 ( \2298 , \2295 , \2296 , \2297 );
nor \U$1987 ( \2299 , \2294 , \2298 );
and \U$1988 ( \2300 , \2177 , \2181 );
and \U$1989 ( \2301 , \2181 , \2292 );
and \U$1990 ( \2302 , \2177 , \2292 );
or \U$1991 ( \2303 , \2300 , \2301 , \2302 );
and \U$1992 ( \2304 , \2186 , \2190 );
and \U$1993 ( \2305 , \2190 , \2195 );
and \U$1994 ( \2306 , \2186 , \2195 );
or \U$1995 ( \2307 , \2304 , \2305 , \2306 );
and \U$1996 ( \2308 , \2164 , \2168 );
and \U$1997 ( \2309 , \2168 , \2170 );
and \U$1998 ( \2310 , \2164 , \2170 );
or \U$1999 ( \2311 , \2308 , \2309 , \2310 );
xor \U$2000 ( \2312 , \2307 , \2311 );
and \U$2001 ( \2313 , \2245 , \2259 );
and \U$2002 ( \2314 , \2259 , \2274 );
and \U$2003 ( \2315 , \2245 , \2274 );
or \U$2004 ( \2316 , \2313 , \2314 , \2315 );
xor \U$2005 ( \2317 , \2312 , \2316 );
and \U$2006 ( \2318 , \2281 , \2285 );
and \U$2007 ( \2319 , \2285 , \2290 );
and \U$2008 ( \2320 , \2281 , \2290 );
or \U$2009 ( \2321 , \2318 , \2319 , \2320 );
and \U$2010 ( \2322 , \2200 , \2241 );
and \U$2011 ( \2323 , \2241 , \2275 );
and \U$2012 ( \2324 , \2200 , \2275 );
or \U$2013 ( \2325 , \2322 , \2323 , \2324 );
xor \U$2014 ( \2326 , \2321 , \2325 );
and \U$2015 ( \2327 , \896 , \1233 );
and \U$2016 ( \2328 , \914 , \1114 );
nor \U$2017 ( \2329 , \2327 , \2328 );
xnor \U$2018 ( \2330 , \2329 , \594 );
and \U$2019 ( \2331 , \922 , \561 );
and \U$2020 ( \2332 , \940 , \559 );
nor \U$2021 ( \2333 , \2331 , \2332 );
xnor \U$2022 ( \2334 , \2333 , \566 );
xor \U$2023 ( \2335 , \2330 , \2334 );
and \U$2025 ( \2336 , \968 , \569 );
nor \U$2026 ( \2337 , 1'b0 , \2336 );
not \U$2027 ( \2338 , \2337 );
xor \U$2028 ( \2339 , \2335 , \2338 );
and \U$2029 ( \2340 , \814 , \966 );
and \U$2030 ( \2341 , \832 , \964 );
nor \U$2031 ( \2342 , \2340 , \2341 );
xnor \U$2032 ( \2343 , \2342 , \973 );
and \U$2033 ( \2344 , \840 , \985 );
and \U$2034 ( \2345 , \858 , \983 );
nor \U$2035 ( \2346 , \2344 , \2345 );
xnor \U$2036 ( \2347 , \2346 , \992 );
xor \U$2037 ( \2348 , \2343 , \2347 );
and \U$2038 ( \2349 , \871 , \1013 );
and \U$2039 ( \2350 , \889 , \996 );
nor \U$2040 ( \2351 , \2349 , \2350 );
xnor \U$2041 ( \2352 , \2351 , \628 );
xor \U$2042 ( \2353 , \2348 , \2352 );
xor \U$2043 ( \2354 , \2339 , \2353 );
and \U$2044 ( \2355 , \734 , \887 );
and \U$2045 ( \2356 , \752 , \885 );
nor \U$2046 ( \2357 , \2355 , \2356 );
xnor \U$2047 ( \2358 , \2357 , \894 );
and \U$2048 ( \2359 , \760 , \912 );
and \U$2049 ( \2360 , \778 , \910 );
nor \U$2050 ( \2361 , \2359 , \2360 );
xnor \U$2051 ( \2362 , \2361 , \919 );
xor \U$2052 ( \2363 , \2358 , \2362 );
and \U$2053 ( \2364 , \789 , \938 );
and \U$2054 ( \2365 , \807 , \936 );
nor \U$2055 ( \2366 , \2364 , \2365 );
xnor \U$2056 ( \2367 , \2366 , \945 );
xor \U$2057 ( \2368 , \2363 , \2367 );
xor \U$2058 ( \2369 , \2354 , \2368 );
and \U$2059 ( \2370 , \2264 , \2268 );
and \U$2060 ( \2371 , \2268 , \2273 );
and \U$2061 ( \2372 , \2264 , \2273 );
or \U$2062 ( \2373 , \2370 , \2371 , \2372 );
and \U$2063 ( \2374 , \2249 , \2253 );
and \U$2064 ( \2375 , \2253 , \2258 );
and \U$2065 ( \2376 , \2249 , \2258 );
or \U$2066 ( \2377 , \2374 , \2375 , \2376 );
xnor \U$2067 ( \2378 , \2373 , \2377 );
xor \U$2068 ( \2379 , \2369 , \2378 );
and \U$2069 ( \2380 , \2230 , \2234 );
and \U$2070 ( \2381 , \2234 , \2239 );
and \U$2071 ( \2382 , \2230 , \2239 );
or \U$2072 ( \2383 , \2380 , \2381 , \2382 );
and \U$2073 ( \2384 , \2218 , \2222 );
and \U$2074 ( \2385 , \2222 , \2227 );
and \U$2075 ( \2386 , \2218 , \2227 );
or \U$2076 ( \2387 , \2384 , \2385 , \2386 );
xor \U$2077 ( \2388 , \2383 , \2387 );
and \U$2078 ( \2389 , \2204 , \2208 );
and \U$2079 ( \2390 , \2208 , \2213 );
and \U$2080 ( \2391 , \2204 , \2213 );
or \U$2081 ( \2392 , \2389 , \2390 , \2391 );
xor \U$2082 ( \2393 , \2388 , \2392 );
xor \U$2083 ( \2394 , \2379 , \2393 );
xor \U$2084 ( \2395 , \2326 , \2394 );
xor \U$2085 ( \2396 , \2317 , \2395 );
xor \U$2086 ( \2397 , \2303 , \2396 );
and \U$2087 ( \2398 , \2155 , \2159 );
and \U$2088 ( \2399 , \2159 , \2171 );
and \U$2089 ( \2400 , \2155 , \2171 );
or \U$2090 ( \2401 , \2398 , \2399 , \2400 );
and \U$2091 ( \2402 , \2196 , \2276 );
and \U$2092 ( \2403 , \2276 , \2291 );
and \U$2093 ( \2404 , \2196 , \2291 );
or \U$2094 ( \2405 , \2402 , \2403 , \2404 );
xor \U$2095 ( \2406 , \2401 , \2405 );
and \U$2096 ( \2407 , \2214 , \2228 );
and \U$2097 ( \2408 , \2228 , \2240 );
and \U$2098 ( \2409 , \2214 , \2240 );
or \U$2099 ( \2410 , \2407 , \2408 , \2409 );
and \U$2100 ( \2411 , \629 , \805 );
and \U$2101 ( \2412 , \676 , \803 );
nor \U$2102 ( \2413 , \2411 , \2412 );
xnor \U$2103 ( \2414 , \2413 , \812 );
and \U$2104 ( \2415 , \681 , \830 );
and \U$2105 ( \2416 , \699 , \828 );
nor \U$2106 ( \2417 , \2415 , \2416 );
xnor \U$2107 ( \2418 , \2417 , \837 );
xor \U$2108 ( \2419 , \2414 , \2418 );
and \U$2109 ( \2420 , \709 , \856 );
and \U$2110 ( \2421 , \727 , \854 );
nor \U$2111 ( \2422 , \2420 , \2421 );
xnor \U$2112 ( \2423 , \2422 , \863 );
xor \U$2113 ( \2424 , \2419 , \2423 );
xor \U$2114 ( \2425 , \2410 , \2424 );
and \U$2115 ( \2426 , \227 , \725 );
not \U$2116 ( \2427 , \2426 );
xnor \U$2117 ( \2428 , \2427 , \732 );
and \U$2118 ( \2429 , \601 , \750 );
and \U$2119 ( \2430 , \568 , \748 );
nor \U$2120 ( \2431 , \2429 , \2430 );
xnor \U$2121 ( \2432 , \2431 , \757 );
xor \U$2122 ( \2433 , \2428 , \2432 );
and \U$2123 ( \2434 , \1053 , \776 );
and \U$2124 ( \2435 , \1055 , \774 );
nor \U$2125 ( \2436 , \2434 , \2435 );
xnor \U$2126 ( \2437 , \2436 , \783 );
xor \U$2127 ( \2438 , \2433 , \2437 );
xor \U$2128 ( \2439 , \2425 , \2438 );
xor \U$2129 ( \2440 , \2406 , \2439 );
xor \U$2130 ( \2441 , \2397 , \2440 );
and \U$2131 ( \2442 , \2151 , \2172 );
and \U$2132 ( \2443 , \2172 , \2293 );
and \U$2133 ( \2444 , \2151 , \2293 );
or \U$2134 ( \2445 , \2442 , \2443 , \2444 );
nor \U$2135 ( \2446 , \2441 , \2445 );
nor \U$2136 ( \2447 , \2299 , \2446 );
and \U$2137 ( \2448 , \2401 , \2405 );
and \U$2138 ( \2449 , \2405 , \2439 );
and \U$2139 ( \2450 , \2401 , \2439 );
or \U$2140 ( \2451 , \2448 , \2449 , \2450 );
and \U$2141 ( \2452 , \2317 , \2395 );
xor \U$2142 ( \2453 , \2451 , \2452 );
and \U$2143 ( \2454 , \2321 , \2325 );
and \U$2144 ( \2455 , \2325 , \2394 );
and \U$2145 ( \2456 , \2321 , \2394 );
or \U$2146 ( \2457 , \2454 , \2455 , \2456 );
and \U$2147 ( \2458 , \2428 , \2432 );
and \U$2148 ( \2459 , \2432 , \2437 );
and \U$2149 ( \2460 , \2428 , \2437 );
or \U$2150 ( \2461 , \2458 , \2459 , \2460 );
and \U$2151 ( \2462 , \2414 , \2418 );
and \U$2152 ( \2463 , \2418 , \2423 );
and \U$2153 ( \2464 , \2414 , \2423 );
or \U$2154 ( \2465 , \2462 , \2463 , \2464 );
xor \U$2155 ( \2466 , \2461 , \2465 );
and \U$2156 ( \2467 , \2358 , \2362 );
and \U$2157 ( \2468 , \2362 , \2367 );
and \U$2158 ( \2469 , \2358 , \2367 );
or \U$2159 ( \2470 , \2467 , \2468 , \2469 );
xor \U$2160 ( \2471 , \2466 , \2470 );
not \U$2161 ( \2472 , \732 );
and \U$2162 ( \2473 , \568 , \750 );
and \U$2163 ( \2474 , \227 , \748 );
nor \U$2164 ( \2475 , \2473 , \2474 );
xnor \U$2165 ( \2476 , \2475 , \757 );
xor \U$2166 ( \2477 , \2472 , \2476 );
and \U$2167 ( \2478 , \1055 , \776 );
and \U$2168 ( \2479 , \601 , \774 );
nor \U$2169 ( \2480 , \2478 , \2479 );
xnor \U$2170 ( \2481 , \2480 , \783 );
xor \U$2171 ( \2482 , \2477 , \2481 );
and \U$2172 ( \2483 , \832 , \966 );
and \U$2173 ( \2484 , \789 , \964 );
nor \U$2174 ( \2485 , \2483 , \2484 );
xnor \U$2175 ( \2486 , \2485 , \973 );
and \U$2176 ( \2487 , \858 , \985 );
and \U$2177 ( \2488 , \814 , \983 );
nor \U$2178 ( \2489 , \2487 , \2488 );
xnor \U$2179 ( \2490 , \2489 , \992 );
xor \U$2180 ( \2491 , \2486 , \2490 );
and \U$2181 ( \2492 , \889 , \1013 );
and \U$2182 ( \2493 , \840 , \996 );
nor \U$2183 ( \2494 , \2492 , \2493 );
xnor \U$2184 ( \2495 , \2494 , \628 );
xor \U$2185 ( \2496 , \2491 , \2495 );
and \U$2186 ( \2497 , \752 , \887 );
and \U$2187 ( \2498 , \709 , \885 );
nor \U$2188 ( \2499 , \2497 , \2498 );
xnor \U$2189 ( \2500 , \2499 , \894 );
and \U$2190 ( \2501 , \778 , \912 );
and \U$2191 ( \2502 , \734 , \910 );
nor \U$2192 ( \2503 , \2501 , \2502 );
xnor \U$2193 ( \2504 , \2503 , \919 );
xor \U$2194 ( \2505 , \2500 , \2504 );
and \U$2195 ( \2506 , \807 , \938 );
and \U$2196 ( \2507 , \760 , \936 );
nor \U$2197 ( \2508 , \2506 , \2507 );
xnor \U$2198 ( \2509 , \2508 , \945 );
xor \U$2199 ( \2510 , \2505 , \2509 );
xor \U$2200 ( \2511 , \2496 , \2510 );
and \U$2201 ( \2512 , \676 , \805 );
and \U$2202 ( \2513 , \1053 , \803 );
nor \U$2203 ( \2514 , \2512 , \2513 );
xnor \U$2204 ( \2515 , \2514 , \812 );
and \U$2205 ( \2516 , \699 , \830 );
and \U$2206 ( \2517 , \629 , \828 );
nor \U$2207 ( \2518 , \2516 , \2517 );
xnor \U$2208 ( \2519 , \2518 , \837 );
xor \U$2209 ( \2520 , \2515 , \2519 );
and \U$2210 ( \2521 , \727 , \856 );
and \U$2211 ( \2522 , \681 , \854 );
nor \U$2212 ( \2523 , \2521 , \2522 );
xnor \U$2213 ( \2524 , \2523 , \863 );
xor \U$2214 ( \2525 , \2520 , \2524 );
xor \U$2215 ( \2526 , \2511 , \2525 );
xor \U$2216 ( \2527 , \2482 , \2526 );
and \U$2217 ( \2528 , \2343 , \2347 );
and \U$2218 ( \2529 , \2347 , \2352 );
and \U$2219 ( \2530 , \2343 , \2352 );
or \U$2220 ( \2531 , \2528 , \2529 , \2530 );
and \U$2221 ( \2532 , \2330 , \2334 );
and \U$2222 ( \2533 , \2334 , \2338 );
and \U$2223 ( \2534 , \2330 , \2338 );
or \U$2224 ( \2535 , \2532 , \2533 , \2534 );
xor \U$2225 ( \2536 , \2531 , \2535 );
and \U$2226 ( \2537 , \914 , \1233 );
and \U$2227 ( \2538 , \871 , \1114 );
nor \U$2228 ( \2539 , \2537 , \2538 );
xnor \U$2229 ( \2540 , \2539 , \594 );
and \U$2230 ( \2541 , \940 , \561 );
and \U$2231 ( \2542 , \896 , \559 );
nor \U$2232 ( \2543 , \2541 , \2542 );
xnor \U$2233 ( \2544 , \2543 , \566 );
xor \U$2234 ( \2545 , \2540 , \2544 );
and \U$2236 ( \2546 , \922 , \569 );
nor \U$2237 ( \2547 , 1'b0 , \2546 );
not \U$2238 ( \2548 , \2547 );
xor \U$2239 ( \2549 , \2545 , \2548 );
xor \U$2240 ( \2550 , \2536 , \2549 );
xor \U$2241 ( \2551 , \2527 , \2550 );
xor \U$2242 ( \2552 , \2471 , \2551 );
and \U$2243 ( \2553 , \2383 , \2387 );
and \U$2244 ( \2554 , \2387 , \2392 );
and \U$2245 ( \2555 , \2383 , \2392 );
or \U$2246 ( \2556 , \2553 , \2554 , \2555 );
or \U$2247 ( \2557 , \2373 , \2377 );
xor \U$2248 ( \2558 , \2556 , \2557 );
and \U$2249 ( \2559 , \2339 , \2353 );
and \U$2250 ( \2560 , \2353 , \2368 );
and \U$2251 ( \2561 , \2339 , \2368 );
or \U$2252 ( \2562 , \2559 , \2560 , \2561 );
xor \U$2253 ( \2563 , \2558 , \2562 );
xor \U$2254 ( \2564 , \2552 , \2563 );
xor \U$2255 ( \2565 , \2457 , \2564 );
and \U$2256 ( \2566 , \2307 , \2311 );
and \U$2257 ( \2567 , \2311 , \2316 );
and \U$2258 ( \2568 , \2307 , \2316 );
or \U$2259 ( \2569 , \2566 , \2567 , \2568 );
and \U$2260 ( \2570 , \2410 , \2424 );
and \U$2261 ( \2571 , \2424 , \2438 );
and \U$2262 ( \2572 , \2410 , \2438 );
or \U$2263 ( \2573 , \2570 , \2571 , \2572 );
xor \U$2264 ( \2574 , \2569 , \2573 );
and \U$2265 ( \2575 , \2369 , \2378 );
and \U$2266 ( \2576 , \2378 , \2393 );
and \U$2267 ( \2577 , \2369 , \2393 );
or \U$2268 ( \2578 , \2575 , \2576 , \2577 );
xor \U$2269 ( \2579 , \2574 , \2578 );
xor \U$2270 ( \2580 , \2565 , \2579 );
xor \U$2271 ( \2581 , \2453 , \2580 );
and \U$2272 ( \2582 , \2303 , \2396 );
and \U$2273 ( \2583 , \2396 , \2440 );
and \U$2274 ( \2584 , \2303 , \2440 );
or \U$2275 ( \2585 , \2582 , \2583 , \2584 );
nor \U$2276 ( \2586 , \2581 , \2585 );
and \U$2277 ( \2587 , \2457 , \2564 );
and \U$2278 ( \2588 , \2564 , \2579 );
and \U$2279 ( \2589 , \2457 , \2579 );
or \U$2280 ( \2590 , \2587 , \2588 , \2589 );
and \U$2281 ( \2591 , \2461 , \2465 );
and \U$2282 ( \2592 , \2465 , \2470 );
and \U$2283 ( \2593 , \2461 , \2470 );
or \U$2284 ( \2594 , \2591 , \2592 , \2593 );
and \U$2285 ( \2595 , \2531 , \2535 );
and \U$2286 ( \2596 , \2535 , \2549 );
and \U$2287 ( \2597 , \2531 , \2549 );
or \U$2288 ( \2598 , \2595 , \2596 , \2597 );
xor \U$2289 ( \2599 , \2594 , \2598 );
and \U$2290 ( \2600 , \2496 , \2510 );
and \U$2291 ( \2601 , \2510 , \2525 );
and \U$2292 ( \2602 , \2496 , \2525 );
or \U$2293 ( \2603 , \2600 , \2601 , \2602 );
xor \U$2294 ( \2604 , \2599 , \2603 );
and \U$2295 ( \2605 , \2556 , \2557 );
and \U$2296 ( \2606 , \2557 , \2562 );
and \U$2297 ( \2607 , \2556 , \2562 );
or \U$2298 ( \2608 , \2605 , \2606 , \2607 );
and \U$2299 ( \2609 , \2482 , \2526 );
and \U$2300 ( \2610 , \2526 , \2550 );
and \U$2301 ( \2611 , \2482 , \2550 );
or \U$2302 ( \2612 , \2609 , \2610 , \2611 );
xor \U$2303 ( \2613 , \2608 , \2612 );
and \U$2304 ( \2614 , \2472 , \2476 );
and \U$2305 ( \2615 , \2476 , \2481 );
and \U$2306 ( \2616 , \2472 , \2481 );
or \U$2307 ( \2617 , \2614 , \2615 , \2616 );
and \U$2308 ( \2618 , \2515 , \2519 );
and \U$2309 ( \2619 , \2519 , \2524 );
and \U$2310 ( \2620 , \2515 , \2524 );
or \U$2311 ( \2621 , \2618 , \2619 , \2620 );
xor \U$2312 ( \2622 , \2617 , \2621 );
and \U$2313 ( \2623 , \2500 , \2504 );
and \U$2314 ( \2624 , \2504 , \2509 );
and \U$2315 ( \2625 , \2500 , \2509 );
or \U$2316 ( \2626 , \2623 , \2624 , \2625 );
xor \U$2317 ( \2627 , \2622 , \2626 );
xor \U$2318 ( \2628 , \2613 , \2627 );
xor \U$2319 ( \2629 , \2604 , \2628 );
xor \U$2320 ( \2630 , \2590 , \2629 );
and \U$2321 ( \2631 , \2569 , \2573 );
and \U$2322 ( \2632 , \2573 , \2578 );
and \U$2323 ( \2633 , \2569 , \2578 );
or \U$2324 ( \2634 , \2631 , \2632 , \2633 );
and \U$2325 ( \2635 , \2471 , \2551 );
and \U$2326 ( \2636 , \2551 , \2563 );
and \U$2327 ( \2637 , \2471 , \2563 );
or \U$2328 ( \2638 , \2635 , \2636 , \2637 );
xor \U$2329 ( \2639 , \2634 , \2638 );
and \U$2330 ( \2640 , \227 , \750 );
not \U$2331 ( \2641 , \2640 );
xnor \U$2332 ( \2642 , \2641 , \757 );
and \U$2333 ( \2643 , \601 , \776 );
and \U$2334 ( \2644 , \568 , \774 );
nor \U$2335 ( \2645 , \2643 , \2644 );
xnor \U$2336 ( \2646 , \2645 , \783 );
xor \U$2337 ( \2647 , \2642 , \2646 );
and \U$2338 ( \2648 , \1053 , \805 );
and \U$2339 ( \2649 , \1055 , \803 );
nor \U$2340 ( \2650 , \2648 , \2649 );
xnor \U$2341 ( \2651 , \2650 , \812 );
xor \U$2342 ( \2652 , \2647 , \2651 );
and \U$2343 ( \2653 , \814 , \985 );
and \U$2344 ( \2654 , \832 , \983 );
nor \U$2345 ( \2655 , \2653 , \2654 );
xnor \U$2346 ( \2656 , \2655 , \992 );
and \U$2347 ( \2657 , \840 , \1013 );
and \U$2348 ( \2658 , \858 , \996 );
nor \U$2349 ( \2659 , \2657 , \2658 );
xnor \U$2350 ( \2660 , \2659 , \628 );
xor \U$2351 ( \2661 , \2656 , \2660 );
and \U$2352 ( \2662 , \871 , \1233 );
and \U$2353 ( \2663 , \889 , \1114 );
nor \U$2354 ( \2664 , \2662 , \2663 );
xnor \U$2355 ( \2665 , \2664 , \594 );
xor \U$2356 ( \2666 , \2661 , \2665 );
and \U$2357 ( \2667 , \734 , \912 );
and \U$2358 ( \2668 , \752 , \910 );
nor \U$2359 ( \2669 , \2667 , \2668 );
xnor \U$2360 ( \2670 , \2669 , \919 );
and \U$2361 ( \2671 , \760 , \938 );
and \U$2362 ( \2672 , \778 , \936 );
nor \U$2363 ( \2673 , \2671 , \2672 );
xnor \U$2364 ( \2674 , \2673 , \945 );
xor \U$2365 ( \2675 , \2670 , \2674 );
and \U$2366 ( \2676 , \789 , \966 );
and \U$2367 ( \2677 , \807 , \964 );
nor \U$2368 ( \2678 , \2676 , \2677 );
xnor \U$2369 ( \2679 , \2678 , \973 );
xor \U$2370 ( \2680 , \2675 , \2679 );
xor \U$2371 ( \2681 , \2666 , \2680 );
and \U$2372 ( \2682 , \629 , \830 );
and \U$2373 ( \2683 , \676 , \828 );
nor \U$2374 ( \2684 , \2682 , \2683 );
xnor \U$2375 ( \2685 , \2684 , \837 );
and \U$2376 ( \2686 , \681 , \856 );
and \U$2377 ( \2687 , \699 , \854 );
nor \U$2378 ( \2688 , \2686 , \2687 );
xnor \U$2379 ( \2689 , \2688 , \863 );
xor \U$2380 ( \2690 , \2685 , \2689 );
and \U$2381 ( \2691 , \709 , \887 );
and \U$2382 ( \2692 , \727 , \885 );
nor \U$2383 ( \2693 , \2691 , \2692 );
xnor \U$2384 ( \2694 , \2693 , \894 );
xor \U$2385 ( \2695 , \2690 , \2694 );
xor \U$2386 ( \2696 , \2681 , \2695 );
xor \U$2387 ( \2697 , \2652 , \2696 );
and \U$2388 ( \2698 , \2486 , \2490 );
and \U$2389 ( \2699 , \2490 , \2495 );
and \U$2390 ( \2700 , \2486 , \2495 );
or \U$2391 ( \2701 , \2698 , \2699 , \2700 );
and \U$2392 ( \2702 , \2540 , \2544 );
and \U$2393 ( \2703 , \2544 , \2548 );
and \U$2394 ( \2704 , \2540 , \2548 );
or \U$2395 ( \2705 , \2702 , \2703 , \2704 );
xor \U$2396 ( \2706 , \2701 , \2705 );
and \U$2397 ( \2707 , \896 , \561 );
and \U$2398 ( \2708 , \914 , \559 );
nor \U$2399 ( \2709 , \2707 , \2708 );
xnor \U$2400 ( \2710 , \2709 , \566 );
and \U$2402 ( \2711 , \940 , \569 );
nor \U$2403 ( \2712 , 1'b0 , \2711 );
not \U$2404 ( \2713 , \2712 );
xnor \U$2405 ( \2714 , \2710 , \2713 );
xor \U$2406 ( \2715 , \2706 , \2714 );
xor \U$2407 ( \2716 , \2697 , \2715 );
xor \U$2408 ( \2717 , \2639 , \2716 );
xor \U$2409 ( \2718 , \2630 , \2717 );
and \U$2410 ( \2719 , \2451 , \2452 );
and \U$2411 ( \2720 , \2452 , \2580 );
and \U$2412 ( \2721 , \2451 , \2580 );
or \U$2413 ( \2722 , \2719 , \2720 , \2721 );
nor \U$2414 ( \2723 , \2718 , \2722 );
nor \U$2415 ( \2724 , \2586 , \2723 );
nand \U$2416 ( \2725 , \2447 , \2724 );
nor \U$2417 ( \2726 , \2147 , \2725 );
and \U$2418 ( \2727 , \2634 , \2638 );
and \U$2419 ( \2728 , \2638 , \2716 );
and \U$2420 ( \2729 , \2634 , \2716 );
or \U$2421 ( \2730 , \2727 , \2728 , \2729 );
and \U$2422 ( \2731 , \2604 , \2628 );
xor \U$2423 ( \2732 , \2730 , \2731 );
and \U$2424 ( \2733 , \2608 , \2612 );
and \U$2425 ( \2734 , \2612 , \2627 );
and \U$2426 ( \2735 , \2608 , \2627 );
or \U$2427 ( \2736 , \2733 , \2734 , \2735 );
and \U$2428 ( \2737 , \2642 , \2646 );
and \U$2429 ( \2738 , \2646 , \2651 );
and \U$2430 ( \2739 , \2642 , \2651 );
or \U$2431 ( \2740 , \2737 , \2738 , \2739 );
and \U$2432 ( \2741 , \2685 , \2689 );
and \U$2433 ( \2742 , \2689 , \2694 );
and \U$2434 ( \2743 , \2685 , \2694 );
or \U$2435 ( \2744 , \2741 , \2742 , \2743 );
xor \U$2436 ( \2745 , \2740 , \2744 );
and \U$2437 ( \2746 , \2670 , \2674 );
and \U$2438 ( \2747 , \2674 , \2679 );
and \U$2439 ( \2748 , \2670 , \2679 );
or \U$2440 ( \2749 , \2746 , \2747 , \2748 );
xor \U$2441 ( \2750 , \2745 , \2749 );
and \U$2442 ( \2751 , \676 , \830 );
and \U$2443 ( \2752 , \1053 , \828 );
nor \U$2444 ( \2753 , \2751 , \2752 );
xnor \U$2445 ( \2754 , \2753 , \837 );
and \U$2446 ( \2755 , \699 , \856 );
and \U$2447 ( \2756 , \629 , \854 );
nor \U$2448 ( \2757 , \2755 , \2756 );
xnor \U$2449 ( \2758 , \2757 , \863 );
xor \U$2450 ( \2759 , \2754 , \2758 );
and \U$2451 ( \2760 , \727 , \887 );
and \U$2452 ( \2761 , \681 , \885 );
nor \U$2453 ( \2762 , \2760 , \2761 );
xnor \U$2454 ( \2763 , \2762 , \894 );
xor \U$2455 ( \2764 , \2759 , \2763 );
not \U$2456 ( \2765 , \757 );
and \U$2457 ( \2766 , \568 , \776 );
and \U$2458 ( \2767 , \227 , \774 );
nor \U$2459 ( \2768 , \2766 , \2767 );
xnor \U$2460 ( \2769 , \2768 , \783 );
xor \U$2461 ( \2770 , \2765 , \2769 );
and \U$2462 ( \2771 , \1055 , \805 );
and \U$2463 ( \2772 , \601 , \803 );
nor \U$2464 ( \2773 , \2771 , \2772 );
xnor \U$2465 ( \2774 , \2773 , \812 );
xor \U$2466 ( \2775 , \2770 , \2774 );
xor \U$2467 ( \2776 , \2764 , \2775 );
and \U$2469 ( \2777 , \896 , \569 );
nor \U$2470 ( \2778 , 1'b0 , \2777 );
not \U$2471 ( \2779 , \2778 );
and \U$2472 ( \2780 , \832 , \985 );
and \U$2473 ( \2781 , \789 , \983 );
nor \U$2474 ( \2782 , \2780 , \2781 );
xnor \U$2475 ( \2783 , \2782 , \992 );
and \U$2476 ( \2784 , \858 , \1013 );
and \U$2477 ( \2785 , \814 , \996 );
nor \U$2478 ( \2786 , \2784 , \2785 );
xnor \U$2479 ( \2787 , \2786 , \628 );
xor \U$2480 ( \2788 , \2783 , \2787 );
and \U$2481 ( \2789 , \889 , \1233 );
and \U$2482 ( \2790 , \840 , \1114 );
nor \U$2483 ( \2791 , \2789 , \2790 );
xnor \U$2484 ( \2792 , \2791 , \594 );
xor \U$2485 ( \2793 , \2788 , \2792 );
xor \U$2486 ( \2794 , \2779 , \2793 );
and \U$2487 ( \2795 , \752 , \912 );
and \U$2488 ( \2796 , \709 , \910 );
nor \U$2489 ( \2797 , \2795 , \2796 );
xnor \U$2490 ( \2798 , \2797 , \919 );
and \U$2491 ( \2799 , \778 , \938 );
and \U$2492 ( \2800 , \734 , \936 );
nor \U$2493 ( \2801 , \2799 , \2800 );
xnor \U$2494 ( \2802 , \2801 , \945 );
xor \U$2495 ( \2803 , \2798 , \2802 );
and \U$2496 ( \2804 , \807 , \966 );
and \U$2497 ( \2805 , \760 , \964 );
nor \U$2498 ( \2806 , \2804 , \2805 );
xnor \U$2499 ( \2807 , \2806 , \973 );
xor \U$2500 ( \2808 , \2803 , \2807 );
xor \U$2501 ( \2809 , \2794 , \2808 );
xor \U$2502 ( \2810 , \2776 , \2809 );
xor \U$2503 ( \2811 , \2750 , \2810 );
and \U$2504 ( \2812 , \2617 , \2621 );
and \U$2505 ( \2813 , \2621 , \2626 );
and \U$2506 ( \2814 , \2617 , \2626 );
or \U$2507 ( \2815 , \2812 , \2813 , \2814 );
and \U$2508 ( \2816 , \2701 , \2705 );
and \U$2509 ( \2817 , \2705 , \2714 );
and \U$2510 ( \2818 , \2701 , \2714 );
or \U$2511 ( \2819 , \2816 , \2817 , \2818 );
xor \U$2512 ( \2820 , \2815 , \2819 );
and \U$2513 ( \2821 , \2666 , \2680 );
and \U$2514 ( \2822 , \2680 , \2695 );
and \U$2515 ( \2823 , \2666 , \2695 );
or \U$2516 ( \2824 , \2821 , \2822 , \2823 );
xor \U$2517 ( \2825 , \2820 , \2824 );
xor \U$2518 ( \2826 , \2811 , \2825 );
xor \U$2519 ( \2827 , \2736 , \2826 );
and \U$2520 ( \2828 , \2594 , \2598 );
and \U$2521 ( \2829 , \2598 , \2603 );
and \U$2522 ( \2830 , \2594 , \2603 );
or \U$2523 ( \2831 , \2828 , \2829 , \2830 );
and \U$2524 ( \2832 , \2652 , \2696 );
and \U$2525 ( \2833 , \2696 , \2715 );
and \U$2526 ( \2834 , \2652 , \2715 );
or \U$2527 ( \2835 , \2832 , \2833 , \2834 );
xor \U$2528 ( \2836 , \2831 , \2835 );
and \U$2529 ( \2837 , \2656 , \2660 );
and \U$2530 ( \2838 , \2660 , \2665 );
and \U$2531 ( \2839 , \2656 , \2665 );
or \U$2532 ( \2840 , \2837 , \2838 , \2839 );
or \U$2533 ( \2841 , \2710 , \2713 );
xor \U$2534 ( \2842 , \2840 , \2841 );
and \U$2535 ( \2843 , \914 , \561 );
and \U$2536 ( \2844 , \871 , \559 );
nor \U$2537 ( \2845 , \2843 , \2844 );
xnor \U$2538 ( \2846 , \2845 , \566 );
xor \U$2539 ( \2847 , \2842 , \2846 );
xor \U$2540 ( \2848 , \2836 , \2847 );
xor \U$2541 ( \2849 , \2827 , \2848 );
xor \U$2542 ( \2850 , \2732 , \2849 );
and \U$2543 ( \2851 , \2590 , \2629 );
and \U$2544 ( \2852 , \2629 , \2717 );
and \U$2545 ( \2853 , \2590 , \2717 );
or \U$2546 ( \2854 , \2851 , \2852 , \2853 );
nor \U$2547 ( \2855 , \2850 , \2854 );
and \U$2548 ( \2856 , \2736 , \2826 );
and \U$2549 ( \2857 , \2826 , \2848 );
and \U$2550 ( \2858 , \2736 , \2848 );
or \U$2551 ( \2859 , \2856 , \2857 , \2858 );
and \U$2552 ( \2860 , \2815 , \2819 );
and \U$2553 ( \2861 , \2819 , \2824 );
and \U$2554 ( \2862 , \2815 , \2824 );
or \U$2555 ( \2863 , \2860 , \2861 , \2862 );
and \U$2556 ( \2864 , \2764 , \2775 );
and \U$2557 ( \2865 , \2775 , \2809 );
and \U$2558 ( \2866 , \2764 , \2809 );
or \U$2559 ( \2867 , \2864 , \2865 , \2866 );
xor \U$2560 ( \2868 , \2863 , \2867 );
and \U$2561 ( \2869 , \734 , \938 );
and \U$2562 ( \2870 , \752 , \936 );
nor \U$2563 ( \2871 , \2869 , \2870 );
xnor \U$2564 ( \2872 , \2871 , \945 );
and \U$2565 ( \2873 , \760 , \966 );
and \U$2566 ( \2874 , \778 , \964 );
nor \U$2567 ( \2875 , \2873 , \2874 );
xnor \U$2568 ( \2876 , \2875 , \973 );
xor \U$2569 ( \2877 , \2872 , \2876 );
and \U$2570 ( \2878 , \789 , \985 );
and \U$2571 ( \2879 , \807 , \983 );
nor \U$2572 ( \2880 , \2878 , \2879 );
xnor \U$2573 ( \2881 , \2880 , \992 );
xor \U$2574 ( \2882 , \2877 , \2881 );
and \U$2575 ( \2883 , \629 , \856 );
and \U$2576 ( \2884 , \676 , \854 );
nor \U$2577 ( \2885 , \2883 , \2884 );
xnor \U$2578 ( \2886 , \2885 , \863 );
and \U$2579 ( \2887 , \681 , \887 );
and \U$2580 ( \2888 , \699 , \885 );
nor \U$2581 ( \2889 , \2887 , \2888 );
xnor \U$2582 ( \2890 , \2889 , \894 );
xor \U$2583 ( \2891 , \2886 , \2890 );
and \U$2584 ( \2892 , \709 , \912 );
and \U$2585 ( \2893 , \727 , \910 );
nor \U$2586 ( \2894 , \2892 , \2893 );
xnor \U$2587 ( \2895 , \2894 , \919 );
xor \U$2588 ( \2896 , \2891 , \2895 );
xor \U$2589 ( \2897 , \2882 , \2896 );
and \U$2590 ( \2898 , \227 , \776 );
not \U$2591 ( \2899 , \2898 );
xnor \U$2592 ( \2900 , \2899 , \783 );
and \U$2593 ( \2901 , \601 , \805 );
and \U$2594 ( \2902 , \568 , \803 );
nor \U$2595 ( \2903 , \2901 , \2902 );
xnor \U$2596 ( \2904 , \2903 , \812 );
xor \U$2597 ( \2905 , \2900 , \2904 );
and \U$2598 ( \2906 , \1053 , \830 );
and \U$2599 ( \2907 , \1055 , \828 );
nor \U$2600 ( \2908 , \2906 , \2907 );
xnor \U$2601 ( \2909 , \2908 , \837 );
xor \U$2602 ( \2910 , \2905 , \2909 );
xor \U$2603 ( \2911 , \2897 , \2910 );
and \U$2604 ( \2912 , \2783 , \2787 );
and \U$2605 ( \2913 , \2787 , \2792 );
and \U$2606 ( \2914 , \2783 , \2792 );
or \U$2607 ( \2915 , \2912 , \2913 , \2914 );
and \U$2609 ( \2916 , \914 , \569 );
nor \U$2610 ( \2917 , 1'b0 , \2916 );
xor \U$2611 ( \2918 , \2915 , \2917 );
and \U$2612 ( \2919 , \814 , \1013 );
and \U$2613 ( \2920 , \832 , \996 );
nor \U$2614 ( \2921 , \2919 , \2920 );
xnor \U$2615 ( \2922 , \2921 , \628 );
and \U$2616 ( \2923 , \840 , \1233 );
and \U$2617 ( \2924 , \858 , \1114 );
nor \U$2618 ( \2925 , \2923 , \2924 );
xnor \U$2619 ( \2926 , \2925 , \594 );
xor \U$2620 ( \2927 , \2922 , \2926 );
and \U$2621 ( \2928 , \871 , \561 );
and \U$2622 ( \2929 , \889 , \559 );
nor \U$2623 ( \2930 , \2928 , \2929 );
xnor \U$2624 ( \2931 , \2930 , \566 );
xor \U$2625 ( \2932 , \2927 , \2931 );
xor \U$2626 ( \2933 , \2918 , \2932 );
xor \U$2627 ( \2934 , \2911 , \2933 );
and \U$2628 ( \2935 , \2765 , \2769 );
and \U$2629 ( \2936 , \2769 , \2774 );
and \U$2630 ( \2937 , \2765 , \2774 );
or \U$2631 ( \2938 , \2935 , \2936 , \2937 );
and \U$2632 ( \2939 , \2754 , \2758 );
and \U$2633 ( \2940 , \2758 , \2763 );
and \U$2634 ( \2941 , \2754 , \2763 );
or \U$2635 ( \2942 , \2939 , \2940 , \2941 );
xor \U$2636 ( \2943 , \2938 , \2942 );
and \U$2637 ( \2944 , \2798 , \2802 );
and \U$2638 ( \2945 , \2802 , \2807 );
and \U$2639 ( \2946 , \2798 , \2807 );
or \U$2640 ( \2947 , \2944 , \2945 , \2946 );
xor \U$2641 ( \2948 , \2943 , \2947 );
xor \U$2642 ( \2949 , \2934 , \2948 );
xor \U$2643 ( \2950 , \2868 , \2949 );
xor \U$2644 ( \2951 , \2859 , \2950 );
and \U$2645 ( \2952 , \2831 , \2835 );
and \U$2646 ( \2953 , \2835 , \2847 );
and \U$2647 ( \2954 , \2831 , \2847 );
or \U$2648 ( \2955 , \2952 , \2953 , \2954 );
and \U$2649 ( \2956 , \2750 , \2810 );
and \U$2650 ( \2957 , \2810 , \2825 );
and \U$2651 ( \2958 , \2750 , \2825 );
or \U$2652 ( \2959 , \2956 , \2957 , \2958 );
xor \U$2653 ( \2960 , \2955 , \2959 );
and \U$2654 ( \2961 , \2740 , \2744 );
and \U$2655 ( \2962 , \2744 , \2749 );
and \U$2656 ( \2963 , \2740 , \2749 );
or \U$2657 ( \2964 , \2961 , \2962 , \2963 );
and \U$2658 ( \2965 , \2840 , \2841 );
and \U$2659 ( \2966 , \2841 , \2846 );
and \U$2660 ( \2967 , \2840 , \2846 );
or \U$2661 ( \2968 , \2965 , \2966 , \2967 );
xor \U$2662 ( \2969 , \2964 , \2968 );
and \U$2663 ( \2970 , \2779 , \2793 );
and \U$2664 ( \2971 , \2793 , \2808 );
and \U$2665 ( \2972 , \2779 , \2808 );
or \U$2666 ( \2973 , \2970 , \2971 , \2972 );
xor \U$2667 ( \2974 , \2969 , \2973 );
xor \U$2668 ( \2975 , \2960 , \2974 );
xor \U$2669 ( \2976 , \2951 , \2975 );
and \U$2670 ( \2977 , \2730 , \2731 );
and \U$2671 ( \2978 , \2731 , \2849 );
and \U$2672 ( \2979 , \2730 , \2849 );
or \U$2673 ( \2980 , \2977 , \2978 , \2979 );
nor \U$2674 ( \2981 , \2976 , \2980 );
nor \U$2675 ( \2982 , \2855 , \2981 );
and \U$2676 ( \2983 , \2955 , \2959 );
and \U$2677 ( \2984 , \2959 , \2974 );
and \U$2678 ( \2985 , \2955 , \2974 );
or \U$2679 ( \2986 , \2983 , \2984 , \2985 );
and \U$2680 ( \2987 , \2863 , \2867 );
and \U$2681 ( \2988 , \2867 , \2949 );
and \U$2682 ( \2989 , \2863 , \2949 );
or \U$2683 ( \2990 , \2987 , \2988 , \2989 );
not \U$2684 ( \2991 , \783 );
and \U$2685 ( \2992 , \568 , \805 );
and \U$2686 ( \2993 , \227 , \803 );
nor \U$2687 ( \2994 , \2992 , \2993 );
xnor \U$2688 ( \2995 , \2994 , \812 );
xor \U$2689 ( \2996 , \2991 , \2995 );
and \U$2690 ( \2997 , \1055 , \830 );
and \U$2691 ( \2998 , \601 , \828 );
nor \U$2692 ( \2999 , \2997 , \2998 );
xnor \U$2693 ( \3000 , \2999 , \837 );
xor \U$2694 ( \3001 , \2996 , \3000 );
and \U$2695 ( \3002 , \832 , \1013 );
and \U$2696 ( \3003 , \789 , \996 );
nor \U$2697 ( \3004 , \3002 , \3003 );
xnor \U$2698 ( \3005 , \3004 , \628 );
and \U$2699 ( \3006 , \858 , \1233 );
and \U$2700 ( \3007 , \814 , \1114 );
nor \U$2701 ( \3008 , \3006 , \3007 );
xnor \U$2702 ( \3009 , \3008 , \594 );
xor \U$2703 ( \3010 , \3005 , \3009 );
and \U$2704 ( \3011 , \889 , \561 );
and \U$2705 ( \3012 , \840 , \559 );
nor \U$2706 ( \3013 , \3011 , \3012 );
xnor \U$2707 ( \3014 , \3013 , \566 );
xor \U$2708 ( \3015 , \3010 , \3014 );
and \U$2709 ( \3016 , \752 , \938 );
and \U$2710 ( \3017 , \709 , \936 );
nor \U$2711 ( \3018 , \3016 , \3017 );
xnor \U$2712 ( \3019 , \3018 , \945 );
and \U$2713 ( \3020 , \778 , \966 );
and \U$2714 ( \3021 , \734 , \964 );
nor \U$2715 ( \3022 , \3020 , \3021 );
xnor \U$2716 ( \3023 , \3022 , \973 );
xor \U$2717 ( \3024 , \3019 , \3023 );
and \U$2718 ( \3025 , \807 , \985 );
and \U$2719 ( \3026 , \760 , \983 );
nor \U$2720 ( \3027 , \3025 , \3026 );
xnor \U$2721 ( \3028 , \3027 , \992 );
xor \U$2722 ( \3029 , \3024 , \3028 );
xor \U$2723 ( \3030 , \3015 , \3029 );
and \U$2724 ( \3031 , \676 , \856 );
and \U$2725 ( \3032 , \1053 , \854 );
nor \U$2726 ( \3033 , \3031 , \3032 );
xnor \U$2727 ( \3034 , \3033 , \863 );
and \U$2728 ( \3035 , \699 , \887 );
and \U$2729 ( \3036 , \629 , \885 );
nor \U$2730 ( \3037 , \3035 , \3036 );
xnor \U$2731 ( \3038 , \3037 , \894 );
xor \U$2732 ( \3039 , \3034 , \3038 );
and \U$2733 ( \3040 , \727 , \912 );
and \U$2734 ( \3041 , \681 , \910 );
nor \U$2735 ( \3042 , \3040 , \3041 );
xnor \U$2736 ( \3043 , \3042 , \919 );
xor \U$2737 ( \3044 , \3039 , \3043 );
xor \U$2738 ( \3045 , \3030 , \3044 );
xor \U$2739 ( \3046 , \3001 , \3045 );
and \U$2740 ( \3047 , \2922 , \2926 );
and \U$2741 ( \3048 , \2926 , \2931 );
and \U$2742 ( \3049 , \2922 , \2931 );
or \U$2743 ( \3050 , \3047 , \3048 , \3049 );
not \U$2744 ( \3051 , \2917 );
xor \U$2745 ( \3052 , \3050 , \3051 );
and \U$2747 ( \3053 , \871 , \569 );
nor \U$2748 ( \3054 , 1'b0 , \3053 );
not \U$2749 ( \3055 , \3054 );
xor \U$2750 ( \3056 , \3052 , \3055 );
xor \U$2751 ( \3057 , \3046 , \3056 );
and \U$2752 ( \3058 , \2938 , \2942 );
and \U$2753 ( \3059 , \2942 , \2947 );
and \U$2754 ( \3060 , \2938 , \2947 );
or \U$2755 ( \3061 , \3058 , \3059 , \3060 );
and \U$2756 ( \3062 , \2915 , \2917 );
and \U$2757 ( \3063 , \2917 , \2932 );
and \U$2758 ( \3064 , \2915 , \2932 );
or \U$2759 ( \3065 , \3062 , \3063 , \3064 );
xor \U$2760 ( \3066 , \3061 , \3065 );
and \U$2761 ( \3067 , \2882 , \2896 );
and \U$2762 ( \3068 , \2896 , \2910 );
and \U$2763 ( \3069 , \2882 , \2910 );
or \U$2764 ( \3070 , \3067 , \3068 , \3069 );
xor \U$2765 ( \3071 , \3066 , \3070 );
xor \U$2766 ( \3072 , \3057 , \3071 );
xor \U$2767 ( \3073 , \2990 , \3072 );
and \U$2768 ( \3074 , \2964 , \2968 );
and \U$2769 ( \3075 , \2968 , \2973 );
and \U$2770 ( \3076 , \2964 , \2973 );
or \U$2771 ( \3077 , \3074 , \3075 , \3076 );
and \U$2772 ( \3078 , \2911 , \2933 );
and \U$2773 ( \3079 , \2933 , \2948 );
and \U$2774 ( \3080 , \2911 , \2948 );
or \U$2775 ( \3081 , \3078 , \3079 , \3080 );
xor \U$2776 ( \3082 , \3077 , \3081 );
and \U$2777 ( \3083 , \2900 , \2904 );
and \U$2778 ( \3084 , \2904 , \2909 );
and \U$2779 ( \3085 , \2900 , \2909 );
or \U$2780 ( \3086 , \3083 , \3084 , \3085 );
and \U$2781 ( \3087 , \2886 , \2890 );
and \U$2782 ( \3088 , \2890 , \2895 );
and \U$2783 ( \3089 , \2886 , \2895 );
or \U$2784 ( \3090 , \3087 , \3088 , \3089 );
xor \U$2785 ( \3091 , \3086 , \3090 );
and \U$2786 ( \3092 , \2872 , \2876 );
and \U$2787 ( \3093 , \2876 , \2881 );
and \U$2788 ( \3094 , \2872 , \2881 );
or \U$2789 ( \3095 , \3092 , \3093 , \3094 );
xor \U$2790 ( \3096 , \3091 , \3095 );
xor \U$2791 ( \3097 , \3082 , \3096 );
xor \U$2792 ( \3098 , \3073 , \3097 );
xor \U$2793 ( \3099 , \2986 , \3098 );
and \U$2794 ( \3100 , \2859 , \2950 );
and \U$2795 ( \3101 , \2950 , \2975 );
and \U$2796 ( \3102 , \2859 , \2975 );
or \U$2797 ( \3103 , \3100 , \3101 , \3102 );
nor \U$2798 ( \3104 , \3099 , \3103 );
and \U$2799 ( \3105 , \2990 , \3072 );
and \U$2800 ( \3106 , \3072 , \3097 );
and \U$2801 ( \3107 , \2990 , \3097 );
or \U$2802 ( \3108 , \3105 , \3106 , \3107 );
and \U$2803 ( \3109 , \3061 , \3065 );
and \U$2804 ( \3110 , \3065 , \3070 );
and \U$2805 ( \3111 , \3061 , \3070 );
or \U$2806 ( \3112 , \3109 , \3110 , \3111 );
and \U$2807 ( \3113 , \3001 , \3045 );
and \U$2808 ( \3114 , \3045 , \3056 );
and \U$2809 ( \3115 , \3001 , \3056 );
or \U$2810 ( \3116 , \3113 , \3114 , \3115 );
xor \U$2811 ( \3117 , \3112 , \3116 );
and \U$2812 ( \3118 , \734 , \966 );
and \U$2813 ( \3119 , \752 , \964 );
nor \U$2814 ( \3120 , \3118 , \3119 );
xnor \U$2815 ( \3121 , \3120 , \973 );
and \U$2816 ( \3122 , \760 , \985 );
and \U$2817 ( \3123 , \778 , \983 );
nor \U$2818 ( \3124 , \3122 , \3123 );
xnor \U$2819 ( \3125 , \3124 , \992 );
xor \U$2820 ( \3126 , \3121 , \3125 );
and \U$2821 ( \3127 , \789 , \1013 );
and \U$2822 ( \3128 , \807 , \996 );
nor \U$2823 ( \3129 , \3127 , \3128 );
xnor \U$2824 ( \3130 , \3129 , \628 );
xor \U$2825 ( \3131 , \3126 , \3130 );
and \U$2826 ( \3132 , \629 , \887 );
and \U$2827 ( \3133 , \676 , \885 );
nor \U$2828 ( \3134 , \3132 , \3133 );
xnor \U$2829 ( \3135 , \3134 , \894 );
and \U$2830 ( \3136 , \681 , \912 );
and \U$2831 ( \3137 , \699 , \910 );
nor \U$2832 ( \3138 , \3136 , \3137 );
xnor \U$2833 ( \3139 , \3138 , \919 );
xor \U$2834 ( \3140 , \3135 , \3139 );
and \U$2835 ( \3141 , \709 , \938 );
and \U$2836 ( \3142 , \727 , \936 );
nor \U$2837 ( \3143 , \3141 , \3142 );
xnor \U$2838 ( \3144 , \3143 , \945 );
xor \U$2839 ( \3145 , \3140 , \3144 );
xor \U$2840 ( \3146 , \3131 , \3145 );
and \U$2841 ( \3147 , \227 , \805 );
not \U$2842 ( \3148 , \3147 );
xnor \U$2843 ( \3149 , \3148 , \812 );
and \U$2844 ( \3150 , \601 , \830 );
and \U$2845 ( \3151 , \568 , \828 );
nor \U$2846 ( \3152 , \3150 , \3151 );
xnor \U$2847 ( \3153 , \3152 , \837 );
xor \U$2848 ( \3154 , \3149 , \3153 );
and \U$2849 ( \3155 , \1053 , \856 );
and \U$2850 ( \3156 , \1055 , \854 );
nor \U$2851 ( \3157 , \3155 , \3156 );
xnor \U$2852 ( \3158 , \3157 , \863 );
xor \U$2853 ( \3159 , \3154 , \3158 );
xor \U$2854 ( \3160 , \3146 , \3159 );
and \U$2855 ( \3161 , \3005 , \3009 );
and \U$2856 ( \3162 , \3009 , \3014 );
and \U$2857 ( \3163 , \3005 , \3014 );
or \U$2858 ( \3164 , \3161 , \3162 , \3163 );
and \U$2859 ( \3165 , \814 , \1233 );
and \U$2860 ( \3166 , \832 , \1114 );
nor \U$2861 ( \3167 , \3165 , \3166 );
xnor \U$2862 ( \3168 , \3167 , \594 );
and \U$2863 ( \3169 , \840 , \561 );
and \U$2864 ( \3170 , \858 , \559 );
nor \U$2865 ( \3171 , \3169 , \3170 );
xnor \U$2866 ( \3172 , \3171 , \566 );
xor \U$2867 ( \3173 , \3168 , \3172 );
and \U$2869 ( \3174 , \889 , \569 );
nor \U$2870 ( \3175 , 1'b0 , \3174 );
not \U$2871 ( \3176 , \3175 );
xor \U$2872 ( \3177 , \3173 , \3176 );
xnor \U$2873 ( \3178 , \3164 , \3177 );
xor \U$2874 ( \3179 , \3160 , \3178 );
and \U$2875 ( \3180 , \2991 , \2995 );
and \U$2876 ( \3181 , \2995 , \3000 );
and \U$2877 ( \3182 , \2991 , \3000 );
or \U$2878 ( \3183 , \3180 , \3181 , \3182 );
and \U$2879 ( \3184 , \3034 , \3038 );
and \U$2880 ( \3185 , \3038 , \3043 );
and \U$2881 ( \3186 , \3034 , \3043 );
or \U$2882 ( \3187 , \3184 , \3185 , \3186 );
xor \U$2883 ( \3188 , \3183 , \3187 );
and \U$2884 ( \3189 , \3019 , \3023 );
and \U$2885 ( \3190 , \3023 , \3028 );
and \U$2886 ( \3191 , \3019 , \3028 );
or \U$2887 ( \3192 , \3189 , \3190 , \3191 );
xor \U$2888 ( \3193 , \3188 , \3192 );
xor \U$2889 ( \3194 , \3179 , \3193 );
xor \U$2890 ( \3195 , \3117 , \3194 );
xor \U$2891 ( \3196 , \3108 , \3195 );
and \U$2892 ( \3197 , \3077 , \3081 );
and \U$2893 ( \3198 , \3081 , \3096 );
and \U$2894 ( \3199 , \3077 , \3096 );
or \U$2895 ( \3200 , \3197 , \3198 , \3199 );
and \U$2896 ( \3201 , \3057 , \3071 );
xor \U$2897 ( \3202 , \3200 , \3201 );
and \U$2898 ( \3203 , \3086 , \3090 );
and \U$2899 ( \3204 , \3090 , \3095 );
and \U$2900 ( \3205 , \3086 , \3095 );
or \U$2901 ( \3206 , \3203 , \3204 , \3205 );
and \U$2902 ( \3207 , \3050 , \3051 );
and \U$2903 ( \3208 , \3051 , \3055 );
and \U$2904 ( \3209 , \3050 , \3055 );
or \U$2905 ( \3210 , \3207 , \3208 , \3209 );
xor \U$2906 ( \3211 , \3206 , \3210 );
and \U$2907 ( \3212 , \3015 , \3029 );
and \U$2908 ( \3213 , \3029 , \3044 );
and \U$2909 ( \3214 , \3015 , \3044 );
or \U$2910 ( \3215 , \3212 , \3213 , \3214 );
xor \U$2911 ( \3216 , \3211 , \3215 );
xor \U$2912 ( \3217 , \3202 , \3216 );
xor \U$2913 ( \3218 , \3196 , \3217 );
and \U$2914 ( \3219 , \2986 , \3098 );
nor \U$2915 ( \3220 , \3218 , \3219 );
nor \U$2916 ( \3221 , \3104 , \3220 );
nand \U$2917 ( \3222 , \2982 , \3221 );
and \U$2918 ( \3223 , \3200 , \3201 );
and \U$2919 ( \3224 , \3201 , \3216 );
and \U$2920 ( \3225 , \3200 , \3216 );
or \U$2921 ( \3226 , \3223 , \3224 , \3225 );
and \U$2922 ( \3227 , \3112 , \3116 );
and \U$2923 ( \3228 , \3116 , \3194 );
and \U$2924 ( \3229 , \3112 , \3194 );
or \U$2925 ( \3230 , \3227 , \3228 , \3229 );
and \U$2926 ( \3231 , \3183 , \3187 );
and \U$2927 ( \3232 , \3187 , \3192 );
and \U$2928 ( \3233 , \3183 , \3192 );
or \U$2929 ( \3234 , \3231 , \3232 , \3233 );
or \U$2930 ( \3235 , \3164 , \3177 );
xor \U$2931 ( \3236 , \3234 , \3235 );
and \U$2932 ( \3237 , \3131 , \3145 );
and \U$2933 ( \3238 , \3145 , \3159 );
and \U$2934 ( \3239 , \3131 , \3159 );
or \U$2935 ( \3240 , \3237 , \3238 , \3239 );
xor \U$2936 ( \3241 , \3236 , \3240 );
xor \U$2937 ( \3242 , \3230 , \3241 );
and \U$2938 ( \3243 , \3206 , \3210 );
and \U$2939 ( \3244 , \3210 , \3215 );
and \U$2940 ( \3245 , \3206 , \3215 );
or \U$2941 ( \3246 , \3243 , \3244 , \3245 );
and \U$2942 ( \3247 , \3160 , \3178 );
and \U$2943 ( \3248 , \3178 , \3193 );
and \U$2944 ( \3249 , \3160 , \3193 );
or \U$2945 ( \3250 , \3247 , \3248 , \3249 );
xor \U$2946 ( \3251 , \3246 , \3250 );
and \U$2947 ( \3252 , \676 , \887 );
and \U$2948 ( \3253 , \1053 , \885 );
nor \U$2949 ( \3254 , \3252 , \3253 );
xnor \U$2950 ( \3255 , \3254 , \894 );
and \U$2951 ( \3256 , \699 , \912 );
and \U$2952 ( \3257 , \629 , \910 );
nor \U$2953 ( \3258 , \3256 , \3257 );
xnor \U$2954 ( \3259 , \3258 , \919 );
xor \U$2955 ( \3260 , \3255 , \3259 );
and \U$2956 ( \3261 , \727 , \938 );
and \U$2957 ( \3262 , \681 , \936 );
nor \U$2958 ( \3263 , \3261 , \3262 );
xnor \U$2959 ( \3264 , \3263 , \945 );
xor \U$2960 ( \3265 , \3260 , \3264 );
not \U$2961 ( \3266 , \812 );
and \U$2962 ( \3267 , \568 , \830 );
and \U$2963 ( \3268 , \227 , \828 );
nor \U$2964 ( \3269 , \3267 , \3268 );
xnor \U$2965 ( \3270 , \3269 , \837 );
xor \U$2966 ( \3271 , \3266 , \3270 );
and \U$2967 ( \3272 , \1055 , \856 );
and \U$2968 ( \3273 , \601 , \854 );
nor \U$2969 ( \3274 , \3272 , \3273 );
xnor \U$2970 ( \3275 , \3274 , \863 );
xor \U$2971 ( \3276 , \3271 , \3275 );
xor \U$2972 ( \3277 , \3265 , \3276 );
and \U$2973 ( \3278 , \3168 , \3172 );
and \U$2974 ( \3279 , \3172 , \3176 );
and \U$2975 ( \3280 , \3168 , \3176 );
or \U$2976 ( \3281 , \3278 , \3279 , \3280 );
and \U$2977 ( \3282 , \832 , \1233 );
and \U$2978 ( \3283 , \789 , \1114 );
nor \U$2979 ( \3284 , \3282 , \3283 );
xnor \U$2980 ( \3285 , \3284 , \594 );
and \U$2981 ( \3286 , \858 , \561 );
and \U$2982 ( \3287 , \814 , \559 );
nor \U$2983 ( \3288 , \3286 , \3287 );
xnor \U$2984 ( \3289 , \3288 , \566 );
xor \U$2985 ( \3290 , \3285 , \3289 );
and \U$2987 ( \3291 , \840 , \569 );
nor \U$2988 ( \3292 , 1'b0 , \3291 );
not \U$2989 ( \3293 , \3292 );
xor \U$2990 ( \3294 , \3290 , \3293 );
xor \U$2991 ( \3295 , \3281 , \3294 );
and \U$2992 ( \3296 , \752 , \966 );
and \U$2993 ( \3297 , \709 , \964 );
nor \U$2994 ( \3298 , \3296 , \3297 );
xnor \U$2995 ( \3299 , \3298 , \973 );
and \U$2996 ( \3300 , \778 , \985 );
and \U$2997 ( \3301 , \734 , \983 );
nor \U$2998 ( \3302 , \3300 , \3301 );
xnor \U$2999 ( \3303 , \3302 , \992 );
xor \U$3000 ( \3304 , \3299 , \3303 );
and \U$3001 ( \3305 , \807 , \1013 );
and \U$3002 ( \3306 , \760 , \996 );
nor \U$3003 ( \3307 , \3305 , \3306 );
xnor \U$3004 ( \3308 , \3307 , \628 );
xor \U$3005 ( \3309 , \3304 , \3308 );
xor \U$3006 ( \3310 , \3295 , \3309 );
xor \U$3007 ( \3311 , \3277 , \3310 );
and \U$3008 ( \3312 , \3149 , \3153 );
and \U$3009 ( \3313 , \3153 , \3158 );
and \U$3010 ( \3314 , \3149 , \3158 );
or \U$3011 ( \3315 , \3312 , \3313 , \3314 );
and \U$3012 ( \3316 , \3135 , \3139 );
and \U$3013 ( \3317 , \3139 , \3144 );
and \U$3014 ( \3318 , \3135 , \3144 );
or \U$3015 ( \3319 , \3316 , \3317 , \3318 );
xor \U$3016 ( \3320 , \3315 , \3319 );
and \U$3017 ( \3321 , \3121 , \3125 );
and \U$3018 ( \3322 , \3125 , \3130 );
and \U$3019 ( \3323 , \3121 , \3130 );
or \U$3020 ( \3324 , \3321 , \3322 , \3323 );
xor \U$3021 ( \3325 , \3320 , \3324 );
xor \U$3022 ( \3326 , \3311 , \3325 );
xor \U$3023 ( \3327 , \3251 , \3326 );
xor \U$3024 ( \3328 , \3242 , \3327 );
xor \U$3025 ( \3329 , \3226 , \3328 );
and \U$3026 ( \3330 , \3108 , \3195 );
and \U$3027 ( \3331 , \3195 , \3217 );
and \U$3028 ( \3332 , \3108 , \3217 );
or \U$3029 ( \3333 , \3330 , \3331 , \3332 );
nor \U$3030 ( \3334 , \3329 , \3333 );
and \U$3031 ( \3335 , \3230 , \3241 );
and \U$3032 ( \3336 , \3241 , \3327 );
and \U$3033 ( \3337 , \3230 , \3327 );
or \U$3034 ( \3338 , \3335 , \3336 , \3337 );
and \U$3035 ( \3339 , \3246 , \3250 );
and \U$3036 ( \3340 , \3250 , \3326 );
and \U$3037 ( \3341 , \3246 , \3326 );
or \U$3038 ( \3342 , \3339 , \3340 , \3341 );
and \U$3039 ( \3343 , \3315 , \3319 );
and \U$3040 ( \3344 , \3319 , \3324 );
and \U$3041 ( \3345 , \3315 , \3324 );
or \U$3042 ( \3346 , \3343 , \3344 , \3345 );
and \U$3043 ( \3347 , \3281 , \3294 );
and \U$3044 ( \3348 , \3294 , \3309 );
and \U$3045 ( \3349 , \3281 , \3309 );
or \U$3046 ( \3350 , \3347 , \3348 , \3349 );
xor \U$3047 ( \3351 , \3346 , \3350 );
and \U$3048 ( \3352 , \3265 , \3276 );
xor \U$3049 ( \3353 , \3351 , \3352 );
xor \U$3050 ( \3354 , \3342 , \3353 );
and \U$3051 ( \3355 , \3234 , \3235 );
and \U$3052 ( \3356 , \3235 , \3240 );
and \U$3053 ( \3357 , \3234 , \3240 );
or \U$3054 ( \3358 , \3355 , \3356 , \3357 );
and \U$3055 ( \3359 , \3277 , \3310 );
and \U$3056 ( \3360 , \3310 , \3325 );
and \U$3057 ( \3361 , \3277 , \3325 );
or \U$3058 ( \3362 , \3359 , \3360 , \3361 );
xor \U$3059 ( \3363 , \3358 , \3362 );
and \U$3060 ( \3364 , \629 , \912 );
and \U$3061 ( \3365 , \676 , \910 );
nor \U$3062 ( \3366 , \3364 , \3365 );
xnor \U$3063 ( \3367 , \3366 , \919 );
and \U$3064 ( \3368 , \681 , \938 );
and \U$3065 ( \3369 , \699 , \936 );
nor \U$3066 ( \3370 , \3368 , \3369 );
xnor \U$3067 ( \3371 , \3370 , \945 );
xor \U$3068 ( \3372 , \3367 , \3371 );
and \U$3069 ( \3373 , \709 , \966 );
and \U$3070 ( \3374 , \727 , \964 );
nor \U$3071 ( \3375 , \3373 , \3374 );
xnor \U$3072 ( \3376 , \3375 , \973 );
xor \U$3073 ( \3377 , \3372 , \3376 );
and \U$3074 ( \3378 , \227 , \830 );
not \U$3075 ( \3379 , \3378 );
xnor \U$3076 ( \3380 , \3379 , \837 );
and \U$3077 ( \3381 , \601 , \856 );
and \U$3078 ( \3382 , \568 , \854 );
nor \U$3079 ( \3383 , \3381 , \3382 );
xnor \U$3080 ( \3384 , \3383 , \863 );
xor \U$3081 ( \3385 , \3380 , \3384 );
and \U$3082 ( \3386 , \1053 , \887 );
and \U$3083 ( \3387 , \1055 , \885 );
nor \U$3084 ( \3388 , \3386 , \3387 );
xnor \U$3085 ( \3389 , \3388 , \894 );
xor \U$3086 ( \3390 , \3385 , \3389 );
xor \U$3087 ( \3391 , \3377 , \3390 );
and \U$3088 ( \3392 , \3285 , \3289 );
and \U$3089 ( \3393 , \3289 , \3293 );
and \U$3090 ( \3394 , \3285 , \3293 );
or \U$3091 ( \3395 , \3392 , \3393 , \3394 );
and \U$3092 ( \3396 , \814 , \561 );
and \U$3093 ( \3397 , \832 , \559 );
nor \U$3094 ( \3398 , \3396 , \3397 );
xnor \U$3095 ( \3399 , \3398 , \566 );
and \U$3097 ( \3400 , \858 , \569 );
nor \U$3098 ( \3401 , 1'b0 , \3400 );
not \U$3099 ( \3402 , \3401 );
xnor \U$3100 ( \3403 , \3399 , \3402 );
xor \U$3101 ( \3404 , \3395 , \3403 );
and \U$3102 ( \3405 , \734 , \985 );
and \U$3103 ( \3406 , \752 , \983 );
nor \U$3104 ( \3407 , \3405 , \3406 );
xnor \U$3105 ( \3408 , \3407 , \992 );
and \U$3106 ( \3409 , \760 , \1013 );
and \U$3107 ( \3410 , \778 , \996 );
nor \U$3108 ( \3411 , \3409 , \3410 );
xnor \U$3109 ( \3412 , \3411 , \628 );
xor \U$3110 ( \3413 , \3408 , \3412 );
and \U$3111 ( \3414 , \789 , \1233 );
and \U$3112 ( \3415 , \807 , \1114 );
nor \U$3113 ( \3416 , \3414 , \3415 );
xnor \U$3114 ( \3417 , \3416 , \594 );
xor \U$3115 ( \3418 , \3413 , \3417 );
xor \U$3116 ( \3419 , \3404 , \3418 );
xor \U$3117 ( \3420 , \3391 , \3419 );
and \U$3118 ( \3421 , \3266 , \3270 );
and \U$3119 ( \3422 , \3270 , \3275 );
and \U$3120 ( \3423 , \3266 , \3275 );
or \U$3121 ( \3424 , \3421 , \3422 , \3423 );
and \U$3122 ( \3425 , \3255 , \3259 );
and \U$3123 ( \3426 , \3259 , \3264 );
and \U$3124 ( \3427 , \3255 , \3264 );
or \U$3125 ( \3428 , \3425 , \3426 , \3427 );
xor \U$3126 ( \3429 , \3424 , \3428 );
and \U$3127 ( \3430 , \3299 , \3303 );
and \U$3128 ( \3431 , \3303 , \3308 );
and \U$3129 ( \3432 , \3299 , \3308 );
or \U$3130 ( \3433 , \3430 , \3431 , \3432 );
xor \U$3131 ( \3434 , \3429 , \3433 );
xor \U$3132 ( \3435 , \3420 , \3434 );
xor \U$3133 ( \3436 , \3363 , \3435 );
xor \U$3134 ( \3437 , \3354 , \3436 );
xor \U$3135 ( \3438 , \3338 , \3437 );
and \U$3136 ( \3439 , \3226 , \3328 );
nor \U$3137 ( \3440 , \3438 , \3439 );
nor \U$3138 ( \3441 , \3334 , \3440 );
and \U$3139 ( \3442 , \3342 , \3353 );
and \U$3140 ( \3443 , \3353 , \3436 );
and \U$3141 ( \3444 , \3342 , \3436 );
or \U$3142 ( \3445 , \3442 , \3443 , \3444 );
and \U$3143 ( \3446 , \3358 , \3362 );
and \U$3144 ( \3447 , \3362 , \3435 );
and \U$3145 ( \3448 , \3358 , \3435 );
or \U$3146 ( \3449 , \3446 , \3447 , \3448 );
and \U$3147 ( \3450 , \3424 , \3428 );
and \U$3148 ( \3451 , \3428 , \3433 );
and \U$3149 ( \3452 , \3424 , \3433 );
or \U$3150 ( \3453 , \3450 , \3451 , \3452 );
and \U$3151 ( \3454 , \3395 , \3403 );
and \U$3152 ( \3455 , \3403 , \3418 );
and \U$3153 ( \3456 , \3395 , \3418 );
or \U$3154 ( \3457 , \3454 , \3455 , \3456 );
xor \U$3155 ( \3458 , \3453 , \3457 );
and \U$3156 ( \3459 , \3377 , \3390 );
xor \U$3157 ( \3460 , \3458 , \3459 );
xor \U$3158 ( \3461 , \3449 , \3460 );
and \U$3159 ( \3462 , \3346 , \3350 );
and \U$3160 ( \3463 , \3350 , \3352 );
and \U$3161 ( \3464 , \3346 , \3352 );
or \U$3162 ( \3465 , \3462 , \3463 , \3464 );
and \U$3163 ( \3466 , \3391 , \3419 );
and \U$3164 ( \3467 , \3419 , \3434 );
and \U$3165 ( \3468 , \3391 , \3434 );
or \U$3166 ( \3469 , \3466 , \3467 , \3468 );
xor \U$3167 ( \3470 , \3465 , \3469 );
and \U$3168 ( \3471 , \752 , \985 );
and \U$3169 ( \3472 , \709 , \983 );
nor \U$3170 ( \3473 , \3471 , \3472 );
xnor \U$3171 ( \3474 , \3473 , \992 );
and \U$3172 ( \3475 , \778 , \1013 );
and \U$3173 ( \3476 , \734 , \996 );
nor \U$3174 ( \3477 , \3475 , \3476 );
xnor \U$3175 ( \3478 , \3477 , \628 );
xor \U$3176 ( \3479 , \3474 , \3478 );
and \U$3177 ( \3480 , \807 , \1233 );
and \U$3178 ( \3481 , \760 , \1114 );
nor \U$3179 ( \3482 , \3480 , \3481 );
xnor \U$3180 ( \3483 , \3482 , \594 );
xor \U$3181 ( \3484 , \3479 , \3483 );
and \U$3182 ( \3485 , \676 , \912 );
and \U$3183 ( \3486 , \1053 , \910 );
nor \U$3184 ( \3487 , \3485 , \3486 );
xnor \U$3185 ( \3488 , \3487 , \919 );
and \U$3186 ( \3489 , \699 , \938 );
and \U$3187 ( \3490 , \629 , \936 );
nor \U$3188 ( \3491 , \3489 , \3490 );
xnor \U$3189 ( \3492 , \3491 , \945 );
xor \U$3190 ( \3493 , \3488 , \3492 );
and \U$3191 ( \3494 , \727 , \966 );
and \U$3192 ( \3495 , \681 , \964 );
nor \U$3193 ( \3496 , \3494 , \3495 );
xnor \U$3194 ( \3497 , \3496 , \973 );
xor \U$3195 ( \3498 , \3493 , \3497 );
xor \U$3196 ( \3499 , \3484 , \3498 );
not \U$3197 ( \3500 , \837 );
and \U$3198 ( \3501 , \568 , \856 );
and \U$3199 ( \3502 , \227 , \854 );
nor \U$3200 ( \3503 , \3501 , \3502 );
xnor \U$3201 ( \3504 , \3503 , \863 );
xor \U$3202 ( \3505 , \3500 , \3504 );
and \U$3203 ( \3506 , \1055 , \887 );
and \U$3204 ( \3507 , \601 , \885 );
nor \U$3205 ( \3508 , \3506 , \3507 );
xnor \U$3206 ( \3509 , \3508 , \894 );
xor \U$3207 ( \3510 , \3505 , \3509 );
xor \U$3208 ( \3511 , \3499 , \3510 );
or \U$3209 ( \3512 , \3399 , \3402 );
and \U$3210 ( \3513 , \832 , \561 );
and \U$3211 ( \3514 , \789 , \559 );
nor \U$3212 ( \3515 , \3513 , \3514 );
xnor \U$3213 ( \3516 , \3515 , \566 );
xor \U$3214 ( \3517 , \3512 , \3516 );
and \U$3216 ( \3518 , \814 , \569 );
nor \U$3217 ( \3519 , 1'b0 , \3518 );
not \U$3218 ( \3520 , \3519 );
xor \U$3219 ( \3521 , \3517 , \3520 );
xor \U$3220 ( \3522 , \3511 , \3521 );
and \U$3221 ( \3523 , \3380 , \3384 );
and \U$3222 ( \3524 , \3384 , \3389 );
and \U$3223 ( \3525 , \3380 , \3389 );
or \U$3224 ( \3526 , \3523 , \3524 , \3525 );
and \U$3225 ( \3527 , \3367 , \3371 );
and \U$3226 ( \3528 , \3371 , \3376 );
and \U$3227 ( \3529 , \3367 , \3376 );
or \U$3228 ( \3530 , \3527 , \3528 , \3529 );
xor \U$3229 ( \3531 , \3526 , \3530 );
and \U$3230 ( \3532 , \3408 , \3412 );
and \U$3231 ( \3533 , \3412 , \3417 );
and \U$3232 ( \3534 , \3408 , \3417 );
or \U$3233 ( \3535 , \3532 , \3533 , \3534 );
xor \U$3234 ( \3536 , \3531 , \3535 );
xor \U$3235 ( \3537 , \3522 , \3536 );
xor \U$3236 ( \3538 , \3470 , \3537 );
xor \U$3237 ( \3539 , \3461 , \3538 );
xor \U$3238 ( \3540 , \3445 , \3539 );
and \U$3239 ( \3541 , \3338 , \3437 );
nor \U$3240 ( \3542 , \3540 , \3541 );
and \U$3241 ( \3543 , \3449 , \3460 );
and \U$3242 ( \3544 , \3460 , \3538 );
and \U$3243 ( \3545 , \3449 , \3538 );
or \U$3244 ( \3546 , \3543 , \3544 , \3545 );
and \U$3245 ( \3547 , \3465 , \3469 );
and \U$3246 ( \3548 , \3469 , \3537 );
and \U$3247 ( \3549 , \3465 , \3537 );
or \U$3248 ( \3550 , \3547 , \3548 , \3549 );
and \U$3249 ( \3551 , \3526 , \3530 );
and \U$3250 ( \3552 , \3530 , \3535 );
and \U$3251 ( \3553 , \3526 , \3535 );
or \U$3252 ( \3554 , \3551 , \3552 , \3553 );
and \U$3253 ( \3555 , \3512 , \3516 );
and \U$3254 ( \3556 , \3516 , \3520 );
and \U$3255 ( \3557 , \3512 , \3520 );
or \U$3256 ( \3558 , \3555 , \3556 , \3557 );
xor \U$3257 ( \3559 , \3554 , \3558 );
and \U$3258 ( \3560 , \3484 , \3498 );
and \U$3259 ( \3561 , \3498 , \3510 );
and \U$3260 ( \3562 , \3484 , \3510 );
or \U$3261 ( \3563 , \3560 , \3561 , \3562 );
xor \U$3262 ( \3564 , \3559 , \3563 );
xor \U$3263 ( \3565 , \3550 , \3564 );
and \U$3264 ( \3566 , \3453 , \3457 );
and \U$3265 ( \3567 , \3457 , \3459 );
and \U$3266 ( \3568 , \3453 , \3459 );
or \U$3267 ( \3569 , \3566 , \3567 , \3568 );
and \U$3268 ( \3570 , \3511 , \3521 );
and \U$3269 ( \3571 , \3521 , \3536 );
and \U$3270 ( \3572 , \3511 , \3536 );
or \U$3271 ( \3573 , \3570 , \3571 , \3572 );
xor \U$3272 ( \3574 , \3569 , \3573 );
and \U$3273 ( \3575 , \629 , \938 );
and \U$3274 ( \3576 , \676 , \936 );
nor \U$3275 ( \3577 , \3575 , \3576 );
xnor \U$3276 ( \3578 , \3577 , \945 );
and \U$3277 ( \3579 , \681 , \966 );
and \U$3278 ( \3580 , \699 , \964 );
nor \U$3279 ( \3581 , \3579 , \3580 );
xnor \U$3280 ( \3582 , \3581 , \973 );
xor \U$3281 ( \3583 , \3578 , \3582 );
and \U$3282 ( \3584 , \709 , \985 );
and \U$3283 ( \3585 , \727 , \983 );
nor \U$3284 ( \3586 , \3584 , \3585 );
xnor \U$3285 ( \3587 , \3586 , \992 );
xor \U$3286 ( \3588 , \3583 , \3587 );
and \U$3287 ( \3589 , \227 , \856 );
not \U$3288 ( \3590 , \3589 );
xnor \U$3289 ( \3591 , \3590 , \863 );
and \U$3290 ( \3592 , \601 , \887 );
and \U$3291 ( \3593 , \568 , \885 );
nor \U$3292 ( \3594 , \3592 , \3593 );
xnor \U$3293 ( \3595 , \3594 , \894 );
xor \U$3294 ( \3596 , \3591 , \3595 );
and \U$3295 ( \3597 , \1053 , \912 );
and \U$3296 ( \3598 , \1055 , \910 );
nor \U$3297 ( \3599 , \3597 , \3598 );
xnor \U$3298 ( \3600 , \3599 , \919 );
xor \U$3299 ( \3601 , \3596 , \3600 );
xor \U$3300 ( \3602 , \3588 , \3601 );
and \U$3302 ( \3603 , \832 , \569 );
nor \U$3303 ( \3604 , 1'b0 , \3603 );
not \U$3304 ( \3605 , \3604 );
and \U$3305 ( \3606 , \734 , \1013 );
and \U$3306 ( \3607 , \752 , \996 );
nor \U$3307 ( \3608 , \3606 , \3607 );
xnor \U$3308 ( \3609 , \3608 , \628 );
and \U$3309 ( \3610 , \760 , \1233 );
and \U$3310 ( \3611 , \778 , \1114 );
nor \U$3311 ( \3612 , \3610 , \3611 );
xnor \U$3312 ( \3613 , \3612 , \594 );
xor \U$3313 ( \3614 , \3609 , \3613 );
and \U$3314 ( \3615 , \789 , \561 );
and \U$3315 ( \3616 , \807 , \559 );
nor \U$3316 ( \3617 , \3615 , \3616 );
xnor \U$3317 ( \3618 , \3617 , \566 );
xor \U$3318 ( \3619 , \3614 , \3618 );
xnor \U$3319 ( \3620 , \3605 , \3619 );
xor \U$3320 ( \3621 , \3602 , \3620 );
and \U$3321 ( \3622 , \3500 , \3504 );
and \U$3322 ( \3623 , \3504 , \3509 );
and \U$3323 ( \3624 , \3500 , \3509 );
or \U$3324 ( \3625 , \3622 , \3623 , \3624 );
and \U$3325 ( \3626 , \3488 , \3492 );
and \U$3326 ( \3627 , \3492 , \3497 );
and \U$3327 ( \3628 , \3488 , \3497 );
or \U$3328 ( \3629 , \3626 , \3627 , \3628 );
xor \U$3329 ( \3630 , \3625 , \3629 );
and \U$3330 ( \3631 , \3474 , \3478 );
and \U$3331 ( \3632 , \3478 , \3483 );
and \U$3332 ( \3633 , \3474 , \3483 );
or \U$3333 ( \3634 , \3631 , \3632 , \3633 );
xor \U$3334 ( \3635 , \3630 , \3634 );
xor \U$3335 ( \3636 , \3621 , \3635 );
xor \U$3336 ( \3637 , \3574 , \3636 );
xor \U$3337 ( \3638 , \3565 , \3637 );
xor \U$3338 ( \3639 , \3546 , \3638 );
and \U$3339 ( \3640 , \3445 , \3539 );
nor \U$3340 ( \3641 , \3639 , \3640 );
nor \U$3341 ( \3642 , \3542 , \3641 );
nand \U$3342 ( \3643 , \3441 , \3642 );
nor \U$3343 ( \3644 , \3222 , \3643 );
nand \U$3344 ( \3645 , \2726 , \3644 );
and \U$3345 ( \3646 , \3550 , \3564 );
and \U$3346 ( \3647 , \3564 , \3637 );
and \U$3347 ( \3648 , \3550 , \3637 );
or \U$3348 ( \3649 , \3646 , \3647 , \3648 );
and \U$3349 ( \3650 , \3569 , \3573 );
and \U$3350 ( \3651 , \3573 , \3636 );
and \U$3351 ( \3652 , \3569 , \3636 );
or \U$3352 ( \3653 , \3650 , \3651 , \3652 );
and \U$3353 ( \3654 , \3625 , \3629 );
and \U$3354 ( \3655 , \3629 , \3634 );
and \U$3355 ( \3656 , \3625 , \3634 );
or \U$3356 ( \3657 , \3654 , \3655 , \3656 );
or \U$3357 ( \3658 , \3605 , \3619 );
xor \U$3358 ( \3659 , \3657 , \3658 );
and \U$3359 ( \3660 , \3588 , \3601 );
xor \U$3360 ( \3661 , \3659 , \3660 );
xor \U$3361 ( \3662 , \3653 , \3661 );
and \U$3362 ( \3663 , \3554 , \3558 );
and \U$3363 ( \3664 , \3558 , \3563 );
and \U$3364 ( \3665 , \3554 , \3563 );
or \U$3365 ( \3666 , \3663 , \3664 , \3665 );
and \U$3366 ( \3667 , \3602 , \3620 );
and \U$3367 ( \3668 , \3620 , \3635 );
and \U$3368 ( \3669 , \3602 , \3635 );
or \U$3369 ( \3670 , \3667 , \3668 , \3669 );
xor \U$3370 ( \3671 , \3666 , \3670 );
not \U$3371 ( \3672 , \863 );
and \U$3372 ( \3673 , \568 , \887 );
and \U$3373 ( \3674 , \227 , \885 );
nor \U$3374 ( \3675 , \3673 , \3674 );
xnor \U$3375 ( \3676 , \3675 , \894 );
xor \U$3376 ( \3677 , \3672 , \3676 );
and \U$3377 ( \3678 , \1055 , \912 );
and \U$3378 ( \3679 , \601 , \910 );
nor \U$3379 ( \3680 , \3678 , \3679 );
xnor \U$3380 ( \3681 , \3680 , \919 );
xor \U$3381 ( \3682 , \3677 , \3681 );
and \U$3383 ( \3683 , \789 , \569 );
nor \U$3384 ( \3684 , 1'b0 , \3683 );
not \U$3385 ( \3685 , \3684 );
and \U$3386 ( \3686 , \752 , \1013 );
and \U$3387 ( \3687 , \709 , \996 );
nor \U$3388 ( \3688 , \3686 , \3687 );
xnor \U$3389 ( \3689 , \3688 , \628 );
and \U$3390 ( \3690 , \778 , \1233 );
and \U$3391 ( \3691 , \734 , \1114 );
nor \U$3392 ( \3692 , \3690 , \3691 );
xnor \U$3393 ( \3693 , \3692 , \594 );
xor \U$3394 ( \3694 , \3689 , \3693 );
and \U$3395 ( \3695 , \807 , \561 );
and \U$3396 ( \3696 , \760 , \559 );
nor \U$3397 ( \3697 , \3695 , \3696 );
xnor \U$3398 ( \3698 , \3697 , \566 );
xor \U$3399 ( \3699 , \3694 , \3698 );
xor \U$3400 ( \3700 , \3685 , \3699 );
and \U$3401 ( \3701 , \676 , \938 );
and \U$3402 ( \3702 , \1053 , \936 );
nor \U$3403 ( \3703 , \3701 , \3702 );
xnor \U$3404 ( \3704 , \3703 , \945 );
and \U$3405 ( \3705 , \699 , \966 );
and \U$3406 ( \3706 , \629 , \964 );
nor \U$3407 ( \3707 , \3705 , \3706 );
xnor \U$3408 ( \3708 , \3707 , \973 );
xor \U$3409 ( \3709 , \3704 , \3708 );
and \U$3410 ( \3710 , \727 , \985 );
and \U$3411 ( \3711 , \681 , \983 );
nor \U$3412 ( \3712 , \3710 , \3711 );
xnor \U$3413 ( \3713 , \3712 , \992 );
xor \U$3414 ( \3714 , \3709 , \3713 );
xor \U$3415 ( \3715 , \3700 , \3714 );
xor \U$3416 ( \3716 , \3682 , \3715 );
and \U$3417 ( \3717 , \3591 , \3595 );
and \U$3418 ( \3718 , \3595 , \3600 );
and \U$3419 ( \3719 , \3591 , \3600 );
or \U$3420 ( \3720 , \3717 , \3718 , \3719 );
and \U$3421 ( \3721 , \3578 , \3582 );
and \U$3422 ( \3722 , \3582 , \3587 );
and \U$3423 ( \3723 , \3578 , \3587 );
or \U$3424 ( \3724 , \3721 , \3722 , \3723 );
xor \U$3425 ( \3725 , \3720 , \3724 );
and \U$3426 ( \3726 , \3609 , \3613 );
and \U$3427 ( \3727 , \3613 , \3618 );
and \U$3428 ( \3728 , \3609 , \3618 );
or \U$3429 ( \3729 , \3726 , \3727 , \3728 );
xor \U$3430 ( \3730 , \3725 , \3729 );
xor \U$3431 ( \3731 , \3716 , \3730 );
xor \U$3432 ( \3732 , \3671 , \3731 );
xor \U$3433 ( \3733 , \3662 , \3732 );
xor \U$3434 ( \3734 , \3649 , \3733 );
and \U$3435 ( \3735 , \3546 , \3638 );
nor \U$3436 ( \3736 , \3734 , \3735 );
and \U$3437 ( \3737 , \3653 , \3661 );
and \U$3438 ( \3738 , \3661 , \3732 );
and \U$3439 ( \3739 , \3653 , \3732 );
or \U$3440 ( \3740 , \3737 , \3738 , \3739 );
and \U$3441 ( \3741 , \3666 , \3670 );
and \U$3442 ( \3742 , \3670 , \3731 );
and \U$3443 ( \3743 , \3666 , \3731 );
or \U$3444 ( \3744 , \3741 , \3742 , \3743 );
and \U$3445 ( \3745 , \3672 , \3676 );
and \U$3446 ( \3746 , \3676 , \3681 );
and \U$3447 ( \3747 , \3672 , \3681 );
or \U$3448 ( \3748 , \3745 , \3746 , \3747 );
and \U$3449 ( \3749 , \3704 , \3708 );
and \U$3450 ( \3750 , \3708 , \3713 );
and \U$3451 ( \3751 , \3704 , \3713 );
or \U$3452 ( \3752 , \3749 , \3750 , \3751 );
xor \U$3453 ( \3753 , \3748 , \3752 );
and \U$3454 ( \3754 , \3689 , \3693 );
and \U$3455 ( \3755 , \3693 , \3698 );
and \U$3456 ( \3756 , \3689 , \3698 );
or \U$3457 ( \3757 , \3754 , \3755 , \3756 );
xor \U$3458 ( \3758 , \3753 , \3757 );
and \U$3459 ( \3759 , \3720 , \3724 );
and \U$3460 ( \3760 , \3724 , \3729 );
and \U$3461 ( \3761 , \3720 , \3729 );
or \U$3462 ( \3762 , \3759 , \3760 , \3761 );
and \U$3463 ( \3763 , \3685 , \3699 );
and \U$3464 ( \3764 , \3699 , \3714 );
and \U$3465 ( \3765 , \3685 , \3714 );
or \U$3466 ( \3766 , \3763 , \3764 , \3765 );
xor \U$3467 ( \3767 , \3762 , \3766 );
and \U$3468 ( \3768 , \227 , \887 );
not \U$3469 ( \3769 , \3768 );
xnor \U$3470 ( \3770 , \3769 , \894 );
and \U$3471 ( \3771 , \601 , \912 );
and \U$3472 ( \3772 , \568 , \910 );
nor \U$3473 ( \3773 , \3771 , \3772 );
xnor \U$3474 ( \3774 , \3773 , \919 );
xor \U$3475 ( \3775 , \3770 , \3774 );
and \U$3476 ( \3776 , \1053 , \938 );
and \U$3477 ( \3777 , \1055 , \936 );
nor \U$3478 ( \3778 , \3776 , \3777 );
xnor \U$3479 ( \3779 , \3778 , \945 );
xor \U$3480 ( \3780 , \3775 , \3779 );
xor \U$3481 ( \3781 , \3767 , \3780 );
xor \U$3482 ( \3782 , \3758 , \3781 );
xor \U$3483 ( \3783 , \3744 , \3782 );
and \U$3484 ( \3784 , \3657 , \3658 );
and \U$3485 ( \3785 , \3658 , \3660 );
and \U$3486 ( \3786 , \3657 , \3660 );
or \U$3487 ( \3787 , \3784 , \3785 , \3786 );
and \U$3488 ( \3788 , \3682 , \3715 );
and \U$3489 ( \3789 , \3715 , \3730 );
and \U$3490 ( \3790 , \3682 , \3730 );
or \U$3491 ( \3791 , \3788 , \3789 , \3790 );
xor \U$3492 ( \3792 , \3787 , \3791 );
and \U$3493 ( \3793 , \734 , \1233 );
and \U$3494 ( \3794 , \752 , \1114 );
nor \U$3495 ( \3795 , \3793 , \3794 );
xnor \U$3496 ( \3796 , \3795 , \594 );
and \U$3497 ( \3797 , \760 , \561 );
and \U$3498 ( \3798 , \778 , \559 );
nor \U$3499 ( \3799 , \3797 , \3798 );
xnor \U$3500 ( \3800 , \3799 , \566 );
xor \U$3501 ( \3801 , \3796 , \3800 );
and \U$3503 ( \3802 , \807 , \569 );
nor \U$3504 ( \3803 , 1'b0 , \3802 );
not \U$3505 ( \3804 , \3803 );
xor \U$3506 ( \3805 , \3801 , \3804 );
and \U$3507 ( \3806 , \629 , \966 );
and \U$3508 ( \3807 , \676 , \964 );
nor \U$3509 ( \3808 , \3806 , \3807 );
xnor \U$3510 ( \3809 , \3808 , \973 );
and \U$3511 ( \3810 , \681 , \985 );
and \U$3512 ( \3811 , \699 , \983 );
nor \U$3513 ( \3812 , \3810 , \3811 );
xnor \U$3514 ( \3813 , \3812 , \992 );
xor \U$3515 ( \3814 , \3809 , \3813 );
and \U$3516 ( \3815 , \709 , \1013 );
and \U$3517 ( \3816 , \727 , \996 );
nor \U$3518 ( \3817 , \3815 , \3816 );
xnor \U$3519 ( \3818 , \3817 , \628 );
xor \U$3520 ( \3819 , \3814 , \3818 );
xnor \U$3521 ( \3820 , \3805 , \3819 );
xor \U$3522 ( \3821 , \3792 , \3820 );
xor \U$3523 ( \3822 , \3783 , \3821 );
xor \U$3524 ( \3823 , \3740 , \3822 );
and \U$3525 ( \3824 , \3649 , \3733 );
nor \U$3526 ( \3825 , \3823 , \3824 );
nor \U$3527 ( \3826 , \3736 , \3825 );
and \U$3528 ( \3827 , \3744 , \3782 );
and \U$3529 ( \3828 , \3782 , \3821 );
and \U$3530 ( \3829 , \3744 , \3821 );
or \U$3531 ( \3830 , \3827 , \3828 , \3829 );
and \U$3532 ( \3831 , \3787 , \3791 );
and \U$3533 ( \3832 , \3791 , \3820 );
and \U$3534 ( \3833 , \3787 , \3820 );
or \U$3535 ( \3834 , \3831 , \3832 , \3833 );
and \U$3536 ( \3835 , \3758 , \3781 );
xor \U$3537 ( \3836 , \3834 , \3835 );
and \U$3538 ( \3837 , \3762 , \3766 );
and \U$3539 ( \3838 , \3766 , \3780 );
and \U$3540 ( \3839 , \3762 , \3780 );
or \U$3541 ( \3840 , \3837 , \3838 , \3839 );
and \U$3542 ( \3841 , \3770 , \3774 );
and \U$3543 ( \3842 , \3774 , \3779 );
and \U$3544 ( \3843 , \3770 , \3779 );
or \U$3545 ( \3844 , \3841 , \3842 , \3843 );
and \U$3546 ( \3845 , \3809 , \3813 );
and \U$3547 ( \3846 , \3813 , \3818 );
and \U$3548 ( \3847 , \3809 , \3818 );
or \U$3549 ( \3848 , \3845 , \3846 , \3847 );
xor \U$3550 ( \3849 , \3844 , \3848 );
and \U$3551 ( \3850 , \3796 , \3800 );
and \U$3552 ( \3851 , \3800 , \3804 );
and \U$3553 ( \3852 , \3796 , \3804 );
or \U$3554 ( \3853 , \3850 , \3851 , \3852 );
xor \U$3555 ( \3854 , \3849 , \3853 );
xor \U$3556 ( \3855 , \3840 , \3854 );
and \U$3557 ( \3856 , \3748 , \3752 );
and \U$3558 ( \3857 , \3752 , \3757 );
and \U$3559 ( \3858 , \3748 , \3757 );
or \U$3560 ( \3859 , \3856 , \3857 , \3858 );
or \U$3561 ( \3860 , \3805 , \3819 );
xor \U$3562 ( \3861 , \3859 , \3860 );
and \U$3563 ( \3862 , \752 , \1233 );
and \U$3564 ( \3863 , \709 , \1114 );
nor \U$3565 ( \3864 , \3862 , \3863 );
xnor \U$3566 ( \3865 , \3864 , \594 );
and \U$3567 ( \3866 , \778 , \561 );
and \U$3568 ( \3867 , \734 , \559 );
nor \U$3569 ( \3868 , \3866 , \3867 );
xnor \U$3570 ( \3869 , \3868 , \566 );
xor \U$3571 ( \3870 , \3865 , \3869 );
and \U$3573 ( \3871 , \760 , \569 );
nor \U$3574 ( \3872 , 1'b0 , \3871 );
not \U$3575 ( \3873 , \3872 );
xor \U$3576 ( \3874 , \3870 , \3873 );
and \U$3577 ( \3875 , \676 , \966 );
and \U$3578 ( \3876 , \1053 , \964 );
nor \U$3579 ( \3877 , \3875 , \3876 );
xnor \U$3580 ( \3878 , \3877 , \973 );
and \U$3581 ( \3879 , \699 , \985 );
and \U$3582 ( \3880 , \629 , \983 );
nor \U$3583 ( \3881 , \3879 , \3880 );
xnor \U$3584 ( \3882 , \3881 , \992 );
xor \U$3585 ( \3883 , \3878 , \3882 );
and \U$3586 ( \3884 , \727 , \1013 );
and \U$3587 ( \3885 , \681 , \996 );
nor \U$3588 ( \3886 , \3884 , \3885 );
xnor \U$3589 ( \3887 , \3886 , \628 );
xor \U$3590 ( \3888 , \3883 , \3887 );
xor \U$3591 ( \3889 , \3874 , \3888 );
not \U$3592 ( \3890 , \894 );
and \U$3593 ( \3891 , \568 , \912 );
and \U$3594 ( \3892 , \227 , \910 );
nor \U$3595 ( \3893 , \3891 , \3892 );
xnor \U$3596 ( \3894 , \3893 , \919 );
xor \U$3597 ( \3895 , \3890 , \3894 );
and \U$3598 ( \3896 , \1055 , \938 );
and \U$3599 ( \3897 , \601 , \936 );
nor \U$3600 ( \3898 , \3896 , \3897 );
xnor \U$3601 ( \3899 , \3898 , \945 );
xor \U$3602 ( \3900 , \3895 , \3899 );
xor \U$3603 ( \3901 , \3889 , \3900 );
xor \U$3604 ( \3902 , \3861 , \3901 );
xor \U$3605 ( \3903 , \3855 , \3902 );
xor \U$3606 ( \3904 , \3836 , \3903 );
xor \U$3607 ( \3905 , \3830 , \3904 );
and \U$3608 ( \3906 , \3740 , \3822 );
nor \U$3609 ( \3907 , \3905 , \3906 );
and \U$3610 ( \3908 , \3834 , \3835 );
and \U$3611 ( \3909 , \3835 , \3903 );
and \U$3612 ( \3910 , \3834 , \3903 );
or \U$3613 ( \3911 , \3908 , \3909 , \3910 );
and \U$3614 ( \3912 , \3840 , \3854 );
and \U$3615 ( \3913 , \3854 , \3902 );
and \U$3616 ( \3914 , \3840 , \3902 );
or \U$3617 ( \3915 , \3912 , \3913 , \3914 );
xor \U$3618 ( \3916 , \3911 , \3915 );
and \U$3619 ( \3917 , \3859 , \3860 );
and \U$3620 ( \3918 , \3860 , \3901 );
and \U$3621 ( \3919 , \3859 , \3901 );
or \U$3622 ( \3920 , \3917 , \3918 , \3919 );
and \U$3623 ( \3921 , \3890 , \3894 );
and \U$3624 ( \3922 , \3894 , \3899 );
and \U$3625 ( \3923 , \3890 , \3899 );
or \U$3626 ( \3924 , \3921 , \3922 , \3923 );
and \U$3627 ( \3925 , \3878 , \3882 );
and \U$3628 ( \3926 , \3882 , \3887 );
and \U$3629 ( \3927 , \3878 , \3887 );
or \U$3630 ( \3928 , \3925 , \3926 , \3927 );
xor \U$3631 ( \3929 , \3924 , \3928 );
and \U$3632 ( \3930 , \3865 , \3869 );
and \U$3633 ( \3931 , \3869 , \3873 );
and \U$3634 ( \3932 , \3865 , \3873 );
or \U$3635 ( \3933 , \3930 , \3931 , \3932 );
xor \U$3636 ( \3934 , \3929 , \3933 );
xor \U$3637 ( \3935 , \3920 , \3934 );
and \U$3638 ( \3936 , \3844 , \3848 );
and \U$3639 ( \3937 , \3848 , \3853 );
and \U$3640 ( \3938 , \3844 , \3853 );
or \U$3641 ( \3939 , \3936 , \3937 , \3938 );
and \U$3642 ( \3940 , \3874 , \3888 );
and \U$3643 ( \3941 , \3888 , \3900 );
and \U$3644 ( \3942 , \3874 , \3900 );
or \U$3645 ( \3943 , \3940 , \3941 , \3942 );
xor \U$3646 ( \3944 , \3939 , \3943 );
and \U$3647 ( \3945 , \734 , \561 );
and \U$3648 ( \3946 , \752 , \559 );
nor \U$3649 ( \3947 , \3945 , \3946 );
xnor \U$3650 ( \3948 , \3947 , \566 );
and \U$3652 ( \3949 , \778 , \569 );
nor \U$3653 ( \3950 , 1'b0 , \3949 );
not \U$3654 ( \3951 , \3950 );
xnor \U$3655 ( \3952 , \3948 , \3951 );
and \U$3656 ( \3953 , \629 , \985 );
and \U$3657 ( \3954 , \676 , \983 );
nor \U$3658 ( \3955 , \3953 , \3954 );
xnor \U$3659 ( \3956 , \3955 , \992 );
and \U$3660 ( \3957 , \681 , \1013 );
and \U$3661 ( \3958 , \699 , \996 );
nor \U$3662 ( \3959 , \3957 , \3958 );
xnor \U$3663 ( \3960 , \3959 , \628 );
xor \U$3664 ( \3961 , \3956 , \3960 );
and \U$3665 ( \3962 , \709 , \1233 );
and \U$3666 ( \3963 , \727 , \1114 );
nor \U$3667 ( \3964 , \3962 , \3963 );
xnor \U$3668 ( \3965 , \3964 , \594 );
xor \U$3669 ( \3966 , \3961 , \3965 );
xor \U$3670 ( \3967 , \3952 , \3966 );
and \U$3671 ( \3968 , \227 , \912 );
not \U$3672 ( \3969 , \3968 );
xnor \U$3673 ( \3970 , \3969 , \919 );
and \U$3674 ( \3971 , \601 , \938 );
and \U$3675 ( \3972 , \568 , \936 );
nor \U$3676 ( \3973 , \3971 , \3972 );
xnor \U$3677 ( \3974 , \3973 , \945 );
xor \U$3678 ( \3975 , \3970 , \3974 );
and \U$3679 ( \3976 , \1053 , \966 );
and \U$3680 ( \3977 , \1055 , \964 );
nor \U$3681 ( \3978 , \3976 , \3977 );
xnor \U$3682 ( \3979 , \3978 , \973 );
xor \U$3683 ( \3980 , \3975 , \3979 );
xor \U$3684 ( \3981 , \3967 , \3980 );
xor \U$3685 ( \3982 , \3944 , \3981 );
xor \U$3686 ( \3983 , \3935 , \3982 );
xor \U$3687 ( \3984 , \3916 , \3983 );
and \U$3688 ( \3985 , \3830 , \3904 );
nor \U$3689 ( \3986 , \3984 , \3985 );
nor \U$3690 ( \3987 , \3907 , \3986 );
nand \U$3691 ( \3988 , \3826 , \3987 );
and \U$3692 ( \3989 , \3920 , \3934 );
and \U$3693 ( \3990 , \3934 , \3982 );
and \U$3694 ( \3991 , \3920 , \3982 );
or \U$3695 ( \3992 , \3989 , \3990 , \3991 );
and \U$3696 ( \3993 , \3939 , \3943 );
and \U$3697 ( \3994 , \3943 , \3981 );
and \U$3698 ( \3995 , \3939 , \3981 );
or \U$3699 ( \3996 , \3993 , \3994 , \3995 );
and \U$3700 ( \3997 , \3970 , \3974 );
and \U$3701 ( \3998 , \3974 , \3979 );
and \U$3702 ( \3999 , \3970 , \3979 );
or \U$3703 ( \4000 , \3997 , \3998 , \3999 );
and \U$3704 ( \4001 , \3956 , \3960 );
and \U$3705 ( \4002 , \3960 , \3965 );
and \U$3706 ( \4003 , \3956 , \3965 );
or \U$3707 ( \4004 , \4001 , \4002 , \4003 );
xor \U$3708 ( \4005 , \4000 , \4004 );
or \U$3709 ( \4006 , \3948 , \3951 );
xor \U$3710 ( \4007 , \4005 , \4006 );
xor \U$3711 ( \4008 , \3996 , \4007 );
and \U$3712 ( \4009 , \3924 , \3928 );
and \U$3713 ( \4010 , \3928 , \3933 );
and \U$3714 ( \4011 , \3924 , \3933 );
or \U$3715 ( \4012 , \4009 , \4010 , \4011 );
and \U$3716 ( \4013 , \3952 , \3966 );
and \U$3717 ( \4014 , \3966 , \3980 );
and \U$3718 ( \4015 , \3952 , \3980 );
or \U$3719 ( \4016 , \4013 , \4014 , \4015 );
xor \U$3720 ( \4017 , \4012 , \4016 );
and \U$3721 ( \4018 , \752 , \561 );
and \U$3722 ( \4019 , \709 , \559 );
nor \U$3723 ( \4020 , \4018 , \4019 );
xnor \U$3724 ( \4021 , \4020 , \566 );
and \U$3726 ( \4022 , \734 , \569 );
nor \U$3727 ( \4023 , 1'b0 , \4022 );
not \U$3728 ( \4024 , \4023 );
xor \U$3729 ( \4025 , \4021 , \4024 );
and \U$3730 ( \4026 , \676 , \985 );
and \U$3731 ( \4027 , \1053 , \983 );
nor \U$3732 ( \4028 , \4026 , \4027 );
xnor \U$3733 ( \4029 , \4028 , \992 );
and \U$3734 ( \4030 , \699 , \1013 );
and \U$3735 ( \4031 , \629 , \996 );
nor \U$3736 ( \4032 , \4030 , \4031 );
xnor \U$3737 ( \4033 , \4032 , \628 );
xor \U$3738 ( \4034 , \4029 , \4033 );
and \U$3739 ( \4035 , \727 , \1233 );
and \U$3740 ( \4036 , \681 , \1114 );
nor \U$3741 ( \4037 , \4035 , \4036 );
xnor \U$3742 ( \4038 , \4037 , \594 );
xor \U$3743 ( \4039 , \4034 , \4038 );
xor \U$3744 ( \4040 , \4025 , \4039 );
not \U$3745 ( \4041 , \919 );
and \U$3746 ( \4042 , \568 , \938 );
and \U$3747 ( \4043 , \227 , \936 );
nor \U$3748 ( \4044 , \4042 , \4043 );
xnor \U$3749 ( \4045 , \4044 , \945 );
xor \U$3750 ( \4046 , \4041 , \4045 );
and \U$3751 ( \4047 , \1055 , \966 );
and \U$3752 ( \4048 , \601 , \964 );
nor \U$3753 ( \4049 , \4047 , \4048 );
xnor \U$3754 ( \4050 , \4049 , \973 );
xor \U$3755 ( \4051 , \4046 , \4050 );
xor \U$3756 ( \4052 , \4040 , \4051 );
xor \U$3757 ( \4053 , \4017 , \4052 );
xor \U$3758 ( \4054 , \4008 , \4053 );
xor \U$3759 ( \4055 , \3992 , \4054 );
and \U$3760 ( \4056 , \3911 , \3915 );
and \U$3761 ( \4057 , \3915 , \3983 );
and \U$3762 ( \4058 , \3911 , \3983 );
or \U$3763 ( \4059 , \4056 , \4057 , \4058 );
nor \U$3764 ( \4060 , \4055 , \4059 );
and \U$3765 ( \4061 , \3996 , \4007 );
and \U$3766 ( \4062 , \4007 , \4053 );
and \U$3767 ( \4063 , \3996 , \4053 );
or \U$3768 ( \4064 , \4061 , \4062 , \4063 );
and \U$3769 ( \4065 , \4012 , \4016 );
and \U$3770 ( \4066 , \4016 , \4052 );
and \U$3771 ( \4067 , \4012 , \4052 );
or \U$3772 ( \4068 , \4065 , \4066 , \4067 );
and \U$3773 ( \4069 , \4041 , \4045 );
and \U$3774 ( \4070 , \4045 , \4050 );
and \U$3775 ( \4071 , \4041 , \4050 );
or \U$3776 ( \4072 , \4069 , \4070 , \4071 );
and \U$3777 ( \4073 , \4029 , \4033 );
and \U$3778 ( \4074 , \4033 , \4038 );
and \U$3779 ( \4075 , \4029 , \4038 );
or \U$3780 ( \4076 , \4073 , \4074 , \4075 );
xor \U$3781 ( \4077 , \4072 , \4076 );
and \U$3782 ( \4078 , \4021 , \4024 );
xor \U$3783 ( \4079 , \4077 , \4078 );
xor \U$3784 ( \4080 , \4068 , \4079 );
and \U$3785 ( \4081 , \4000 , \4004 );
and \U$3786 ( \4082 , \4004 , \4006 );
and \U$3787 ( \4083 , \4000 , \4006 );
or \U$3788 ( \4084 , \4081 , \4082 , \4083 );
and \U$3789 ( \4085 , \4025 , \4039 );
and \U$3790 ( \4086 , \4039 , \4051 );
and \U$3791 ( \4087 , \4025 , \4051 );
or \U$3792 ( \4088 , \4085 , \4086 , \4087 );
xor \U$3793 ( \4089 , \4084 , \4088 );
and \U$3795 ( \4090 , \752 , \569 );
nor \U$3796 ( \4091 , 1'b0 , \4090 );
and \U$3797 ( \4092 , \629 , \1013 );
and \U$3798 ( \4093 , \676 , \996 );
nor \U$3799 ( \4094 , \4092 , \4093 );
xnor \U$3800 ( \4095 , \4094 , \628 );
and \U$3801 ( \4096 , \681 , \1233 );
and \U$3802 ( \4097 , \699 , \1114 );
nor \U$3803 ( \4098 , \4096 , \4097 );
xnor \U$3804 ( \4099 , \4098 , \594 );
xor \U$3805 ( \4100 , \4095 , \4099 );
and \U$3806 ( \4101 , \709 , \561 );
and \U$3807 ( \4102 , \727 , \559 );
nor \U$3808 ( \4103 , \4101 , \4102 );
xnor \U$3809 ( \4104 , \4103 , \566 );
xor \U$3810 ( \4105 , \4100 , \4104 );
xor \U$3811 ( \4106 , \4091 , \4105 );
and \U$3812 ( \4107 , \227 , \938 );
not \U$3813 ( \4108 , \4107 );
xnor \U$3814 ( \4109 , \4108 , \945 );
and \U$3815 ( \4110 , \601 , \966 );
and \U$3816 ( \4111 , \568 , \964 );
nor \U$3817 ( \4112 , \4110 , \4111 );
xnor \U$3818 ( \4113 , \4112 , \973 );
xor \U$3819 ( \4114 , \4109 , \4113 );
and \U$3820 ( \4115 , \1053 , \985 );
and \U$3821 ( \4116 , \1055 , \983 );
nor \U$3822 ( \4117 , \4115 , \4116 );
xnor \U$3823 ( \4118 , \4117 , \992 );
xor \U$3824 ( \4119 , \4114 , \4118 );
xor \U$3825 ( \4120 , \4106 , \4119 );
xor \U$3826 ( \4121 , \4089 , \4120 );
xor \U$3827 ( \4122 , \4080 , \4121 );
xor \U$3828 ( \4123 , \4064 , \4122 );
and \U$3829 ( \4124 , \3992 , \4054 );
nor \U$3830 ( \4125 , \4123 , \4124 );
nor \U$3831 ( \4126 , \4060 , \4125 );
and \U$3832 ( \4127 , \4068 , \4079 );
and \U$3833 ( \4128 , \4079 , \4121 );
and \U$3834 ( \4129 , \4068 , \4121 );
or \U$3835 ( \4130 , \4127 , \4128 , \4129 );
and \U$3836 ( \4131 , \4084 , \4088 );
and \U$3837 ( \4132 , \4088 , \4120 );
and \U$3838 ( \4133 , \4084 , \4120 );
or \U$3839 ( \4134 , \4131 , \4132 , \4133 );
and \U$3840 ( \4135 , \4109 , \4113 );
and \U$3841 ( \4136 , \4113 , \4118 );
and \U$3842 ( \4137 , \4109 , \4118 );
or \U$3843 ( \4138 , \4135 , \4136 , \4137 );
and \U$3844 ( \4139 , \4095 , \4099 );
and \U$3845 ( \4140 , \4099 , \4104 );
and \U$3846 ( \4141 , \4095 , \4104 );
or \U$3847 ( \4142 , \4139 , \4140 , \4141 );
xor \U$3848 ( \4143 , \4138 , \4142 );
not \U$3849 ( \4144 , \4091 );
xor \U$3850 ( \4145 , \4143 , \4144 );
xor \U$3851 ( \4146 , \4134 , \4145 );
and \U$3852 ( \4147 , \4072 , \4076 );
and \U$3853 ( \4148 , \4076 , \4078 );
and \U$3854 ( \4149 , \4072 , \4078 );
or \U$3855 ( \4150 , \4147 , \4148 , \4149 );
and \U$3856 ( \4151 , \4091 , \4105 );
and \U$3857 ( \4152 , \4105 , \4119 );
and \U$3858 ( \4153 , \4091 , \4119 );
or \U$3859 ( \4154 , \4151 , \4152 , \4153 );
xor \U$3860 ( \4155 , \4150 , \4154 );
and \U$3862 ( \4156 , \709 , \569 );
nor \U$3863 ( \4157 , 1'b0 , \4156 );
not \U$3864 ( \4158 , \4157 );
and \U$3865 ( \4159 , \676 , \1013 );
and \U$3866 ( \4160 , \1053 , \996 );
nor \U$3867 ( \4161 , \4159 , \4160 );
xnor \U$3868 ( \4162 , \4161 , \628 );
and \U$3869 ( \4163 , \699 , \1233 );
and \U$3870 ( \4164 , \629 , \1114 );
nor \U$3871 ( \4165 , \4163 , \4164 );
xnor \U$3872 ( \4166 , \4165 , \594 );
xor \U$3873 ( \4167 , \4162 , \4166 );
and \U$3874 ( \4168 , \727 , \561 );
and \U$3875 ( \4169 , \681 , \559 );
nor \U$3876 ( \4170 , \4168 , \4169 );
xnor \U$3877 ( \4171 , \4170 , \566 );
xor \U$3878 ( \4172 , \4167 , \4171 );
xor \U$3879 ( \4173 , \4158 , \4172 );
not \U$3880 ( \4174 , \945 );
and \U$3881 ( \4175 , \568 , \966 );
and \U$3882 ( \4176 , \227 , \964 );
nor \U$3883 ( \4177 , \4175 , \4176 );
xnor \U$3884 ( \4178 , \4177 , \973 );
xor \U$3885 ( \4179 , \4174 , \4178 );
and \U$3886 ( \4180 , \1055 , \985 );
and \U$3887 ( \4181 , \601 , \983 );
nor \U$3888 ( \4182 , \4180 , \4181 );
xnor \U$3889 ( \4183 , \4182 , \992 );
xor \U$3890 ( \4184 , \4179 , \4183 );
xor \U$3891 ( \4185 , \4173 , \4184 );
xor \U$3892 ( \4186 , \4155 , \4185 );
xor \U$3893 ( \4187 , \4146 , \4186 );
xor \U$3894 ( \4188 , \4130 , \4187 );
and \U$3895 ( \4189 , \4064 , \4122 );
nor \U$3896 ( \4190 , \4188 , \4189 );
and \U$3897 ( \4191 , \4134 , \4145 );
and \U$3898 ( \4192 , \4145 , \4186 );
and \U$3899 ( \4193 , \4134 , \4186 );
or \U$3900 ( \4194 , \4191 , \4192 , \4193 );
and \U$3901 ( \4195 , \4150 , \4154 );
and \U$3902 ( \4196 , \4154 , \4185 );
and \U$3903 ( \4197 , \4150 , \4185 );
or \U$3904 ( \4198 , \4195 , \4196 , \4197 );
and \U$3905 ( \4199 , \227 , \966 );
not \U$3906 ( \4200 , \4199 );
xnor \U$3907 ( \4201 , \4200 , \973 );
and \U$3908 ( \4202 , \601 , \985 );
and \U$3909 ( \4203 , \568 , \983 );
nor \U$3910 ( \4204 , \4202 , \4203 );
xnor \U$3911 ( \4205 , \4204 , \992 );
xor \U$3912 ( \4206 , \4201 , \4205 );
and \U$3913 ( \4207 , \1053 , \1013 );
and \U$3914 ( \4208 , \1055 , \996 );
nor \U$3915 ( \4209 , \4207 , \4208 );
xnor \U$3916 ( \4210 , \4209 , \628 );
xor \U$3917 ( \4211 , \4206 , \4210 );
and \U$3918 ( \4212 , \4174 , \4178 );
and \U$3919 ( \4213 , \4178 , \4183 );
and \U$3920 ( \4214 , \4174 , \4183 );
or \U$3921 ( \4215 , \4212 , \4213 , \4214 );
and \U$3922 ( \4216 , \4162 , \4166 );
and \U$3923 ( \4217 , \4166 , \4171 );
and \U$3924 ( \4218 , \4162 , \4171 );
or \U$3925 ( \4219 , \4216 , \4217 , \4218 );
xnor \U$3926 ( \4220 , \4215 , \4219 );
xor \U$3927 ( \4221 , \4211 , \4220 );
xor \U$3928 ( \4222 , \4198 , \4221 );
and \U$3929 ( \4223 , \4138 , \4142 );
and \U$3930 ( \4224 , \4142 , \4144 );
and \U$3931 ( \4225 , \4138 , \4144 );
or \U$3932 ( \4226 , \4223 , \4224 , \4225 );
and \U$3933 ( \4227 , \4158 , \4172 );
and \U$3934 ( \4228 , \4172 , \4184 );
and \U$3935 ( \4229 , \4158 , \4184 );
or \U$3936 ( \4230 , \4227 , \4228 , \4229 );
xor \U$3937 ( \4231 , \4226 , \4230 );
and \U$3938 ( \4232 , \629 , \1233 );
and \U$3939 ( \4233 , \676 , \1114 );
nor \U$3940 ( \4234 , \4232 , \4233 );
xnor \U$3941 ( \4235 , \4234 , \594 );
and \U$3942 ( \4236 , \681 , \561 );
and \U$3943 ( \4237 , \699 , \559 );
nor \U$3944 ( \4238 , \4236 , \4237 );
xnor \U$3945 ( \4239 , \4238 , \566 );
xor \U$3946 ( \4240 , \4235 , \4239 );
and \U$3948 ( \4241 , \727 , \569 );
nor \U$3949 ( \4242 , 1'b0 , \4241 );
not \U$3950 ( \4243 , \4242 );
xor \U$3951 ( \4244 , \4240 , \4243 );
xor \U$3952 ( \4245 , \4231 , \4244 );
xor \U$3953 ( \4246 , \4222 , \4245 );
xor \U$3954 ( \4247 , \4194 , \4246 );
and \U$3955 ( \4248 , \4130 , \4187 );
nor \U$3956 ( \4249 , \4247 , \4248 );
nor \U$3957 ( \4250 , \4190 , \4249 );
nand \U$3958 ( \4251 , \4126 , \4250 );
nor \U$3959 ( \4252 , \3988 , \4251 );
and \U$3960 ( \4253 , \4198 , \4221 );
and \U$3961 ( \4254 , \4221 , \4245 );
and \U$3962 ( \4255 , \4198 , \4245 );
or \U$3963 ( \4256 , \4253 , \4254 , \4255 );
and \U$3964 ( \4257 , \4226 , \4230 );
and \U$3965 ( \4258 , \4230 , \4244 );
and \U$3966 ( \4259 , \4226 , \4244 );
or \U$3967 ( \4260 , \4257 , \4258 , \4259 );
and \U$3968 ( \4261 , \4211 , \4220 );
xor \U$3969 ( \4262 , \4260 , \4261 );
or \U$3970 ( \4263 , \4215 , \4219 );
not \U$3971 ( \4264 , \973 );
and \U$3972 ( \4265 , \568 , \985 );
and \U$3973 ( \4266 , \227 , \983 );
nor \U$3974 ( \4267 , \4265 , \4266 );
xnor \U$3975 ( \4268 , \4267 , \992 );
xor \U$3976 ( \4269 , \4264 , \4268 );
and \U$3977 ( \4270 , \1055 , \1013 );
and \U$3978 ( \4271 , \601 , \996 );
nor \U$3979 ( \4272 , \4270 , \4271 );
xnor \U$3980 ( \4273 , \4272 , \628 );
xor \U$3981 ( \4274 , \4269 , \4273 );
xor \U$3982 ( \4275 , \4263 , \4274 );
and \U$3983 ( \4276 , \4201 , \4205 );
and \U$3984 ( \4277 , \4205 , \4210 );
and \U$3985 ( \4278 , \4201 , \4210 );
or \U$3986 ( \4279 , \4276 , \4277 , \4278 );
and \U$3987 ( \4280 , \4235 , \4239 );
and \U$3988 ( \4281 , \4239 , \4243 );
and \U$3989 ( \4282 , \4235 , \4243 );
or \U$3990 ( \4283 , \4280 , \4281 , \4282 );
xor \U$3991 ( \4284 , \4279 , \4283 );
and \U$3992 ( \4285 , \676 , \1233 );
and \U$3993 ( \4286 , \1053 , \1114 );
nor \U$3994 ( \4287 , \4285 , \4286 );
xnor \U$3995 ( \4288 , \4287 , \594 );
and \U$3996 ( \4289 , \699 , \561 );
and \U$3997 ( \4290 , \629 , \559 );
nor \U$3998 ( \4291 , \4289 , \4290 );
xnor \U$3999 ( \4292 , \4291 , \566 );
xor \U$4000 ( \4293 , \4288 , \4292 );
and \U$4002 ( \4294 , \681 , \569 );
nor \U$4003 ( \4295 , 1'b0 , \4294 );
not \U$4004 ( \4296 , \4295 );
xor \U$4005 ( \4297 , \4293 , \4296 );
xor \U$4006 ( \4298 , \4284 , \4297 );
xor \U$4007 ( \4299 , \4275 , \4298 );
xor \U$4008 ( \4300 , \4262 , \4299 );
xor \U$4009 ( \4301 , \4256 , \4300 );
and \U$4010 ( \4302 , \4194 , \4246 );
nor \U$4011 ( \4303 , \4301 , \4302 );
and \U$4012 ( \4304 , \4260 , \4261 );
and \U$4013 ( \4305 , \4261 , \4299 );
and \U$4014 ( \4306 , \4260 , \4299 );
or \U$4015 ( \4307 , \4304 , \4305 , \4306 );
and \U$4016 ( \4308 , \4263 , \4274 );
and \U$4017 ( \4309 , \4274 , \4298 );
and \U$4018 ( \4310 , \4263 , \4298 );
or \U$4019 ( \4311 , \4308 , \4309 , \4310 );
xor \U$4020 ( \4312 , \4307 , \4311 );
and \U$4021 ( \4313 , \4279 , \4283 );
and \U$4022 ( \4314 , \4283 , \4297 );
and \U$4023 ( \4315 , \4279 , \4297 );
or \U$4024 ( \4316 , \4313 , \4314 , \4315 );
and \U$4025 ( \4317 , \227 , \985 );
not \U$4026 ( \4318 , \4317 );
xnor \U$4027 ( \4319 , \4318 , \992 );
and \U$4028 ( \4320 , \601 , \1013 );
and \U$4029 ( \4321 , \568 , \996 );
nor \U$4030 ( \4322 , \4320 , \4321 );
xnor \U$4031 ( \4323 , \4322 , \628 );
xor \U$4032 ( \4324 , \4319 , \4323 );
and \U$4033 ( \4325 , \1053 , \1233 );
and \U$4034 ( \4326 , \1055 , \1114 );
nor \U$4035 ( \4327 , \4325 , \4326 );
xnor \U$4036 ( \4328 , \4327 , \594 );
xor \U$4037 ( \4329 , \4324 , \4328 );
xor \U$4038 ( \4330 , \4316 , \4329 );
and \U$4039 ( \4331 , \4264 , \4268 );
and \U$4040 ( \4332 , \4268 , \4273 );
and \U$4041 ( \4333 , \4264 , \4273 );
or \U$4042 ( \4334 , \4331 , \4332 , \4333 );
and \U$4043 ( \4335 , \4288 , \4292 );
and \U$4044 ( \4336 , \4292 , \4296 );
and \U$4045 ( \4337 , \4288 , \4296 );
or \U$4046 ( \4338 , \4335 , \4336 , \4337 );
xor \U$4047 ( \4339 , \4334 , \4338 );
and \U$4048 ( \4340 , \629 , \561 );
and \U$4049 ( \4341 , \676 , \559 );
nor \U$4050 ( \4342 , \4340 , \4341 );
xnor \U$4051 ( \4343 , \4342 , \566 );
and \U$4053 ( \4344 , \699 , \569 );
nor \U$4054 ( \4345 , 1'b0 , \4344 );
not \U$4055 ( \4346 , \4345 );
xnor \U$4056 ( \4347 , \4343 , \4346 );
xor \U$4057 ( \4348 , \4339 , \4347 );
xor \U$4058 ( \4349 , \4330 , \4348 );
xor \U$4059 ( \4350 , \4312 , \4349 );
and \U$4060 ( \4351 , \4256 , \4300 );
nor \U$4061 ( \4352 , \4350 , \4351 );
nor \U$4062 ( \4353 , \4303 , \4352 );
and \U$4063 ( \4354 , \4316 , \4329 );
and \U$4064 ( \4355 , \4329 , \4348 );
and \U$4065 ( \4356 , \4316 , \4348 );
or \U$4066 ( \4357 , \4354 , \4355 , \4356 );
and \U$4067 ( \4358 , \4334 , \4338 );
and \U$4068 ( \4359 , \4338 , \4347 );
and \U$4069 ( \4360 , \4334 , \4347 );
or \U$4070 ( \4361 , \4358 , \4359 , \4360 );
and \U$4072 ( \4362 , \629 , \569 );
nor \U$4073 ( \4363 , 1'b0 , \4362 );
not \U$4074 ( \4364 , \4363 );
not \U$4075 ( \4365 , \992 );
and \U$4076 ( \4366 , \568 , \1013 );
and \U$4077 ( \4367 , \227 , \996 );
nor \U$4078 ( \4368 , \4366 , \4367 );
xnor \U$4079 ( \4369 , \4368 , \628 );
xor \U$4080 ( \4370 , \4365 , \4369 );
and \U$4081 ( \4371 , \1055 , \1233 );
and \U$4082 ( \4372 , \601 , \1114 );
nor \U$4083 ( \4373 , \4371 , \4372 );
xnor \U$4084 ( \4374 , \4373 , \594 );
xor \U$4085 ( \4375 , \4370 , \4374 );
xor \U$4086 ( \4376 , \4364 , \4375 );
xor \U$4087 ( \4377 , \4361 , \4376 );
and \U$4088 ( \4378 , \4319 , \4323 );
and \U$4089 ( \4379 , \4323 , \4328 );
and \U$4090 ( \4380 , \4319 , \4328 );
or \U$4091 ( \4381 , \4378 , \4379 , \4380 );
or \U$4092 ( \4382 , \4343 , \4346 );
xor \U$4093 ( \4383 , \4381 , \4382 );
and \U$4094 ( \4384 , \676 , \561 );
and \U$4095 ( \4385 , \1053 , \559 );
nor \U$4096 ( \4386 , \4384 , \4385 );
xnor \U$4097 ( \4387 , \4386 , \566 );
xor \U$4098 ( \4388 , \4383 , \4387 );
xor \U$4099 ( \4389 , \4377 , \4388 );
xor \U$4100 ( \4390 , \4357 , \4389 );
and \U$4101 ( \4391 , \4307 , \4311 );
and \U$4102 ( \4392 , \4311 , \4349 );
and \U$4103 ( \4393 , \4307 , \4349 );
or \U$4104 ( \4394 , \4391 , \4392 , \4393 );
nor \U$4105 ( \4395 , \4390 , \4394 );
and \U$4106 ( \4396 , \4361 , \4376 );
and \U$4107 ( \4397 , \4376 , \4388 );
and \U$4108 ( \4398 , \4361 , \4388 );
or \U$4109 ( \4399 , \4396 , \4397 , \4398 );
and \U$4110 ( \4400 , \4381 , \4382 );
and \U$4111 ( \4401 , \4382 , \4387 );
and \U$4112 ( \4402 , \4381 , \4387 );
or \U$4113 ( \4403 , \4400 , \4401 , \4402 );
and \U$4114 ( \4404 , \4364 , \4375 );
xor \U$4115 ( \4405 , \4403 , \4404 );
and \U$4116 ( \4406 , \4365 , \4369 );
and \U$4117 ( \4407 , \4369 , \4374 );
and \U$4118 ( \4408 , \4365 , \4374 );
or \U$4119 ( \4409 , \4406 , \4407 , \4408 );
and \U$4121 ( \4410 , \676 , \569 );
nor \U$4122 ( \4411 , 1'b0 , \4410 );
xor \U$4123 ( \4412 , \4409 , \4411 );
and \U$4124 ( \4413 , \227 , \1013 );
not \U$4125 ( \4414 , \4413 );
xnor \U$4126 ( \4415 , \4414 , \628 );
and \U$4127 ( \4416 , \601 , \1233 );
and \U$4128 ( \4417 , \568 , \1114 );
nor \U$4129 ( \4418 , \4416 , \4417 );
xnor \U$4130 ( \4419 , \4418 , \594 );
xor \U$4131 ( \4420 , \4415 , \4419 );
and \U$4132 ( \4421 , \1053 , \561 );
and \U$4133 ( \4422 , \1055 , \559 );
nor \U$4134 ( \4423 , \4421 , \4422 );
xnor \U$4135 ( \4424 , \4423 , \566 );
xor \U$4136 ( \4425 , \4420 , \4424 );
xor \U$4137 ( \4426 , \4412 , \4425 );
xor \U$4138 ( \4427 , \4405 , \4426 );
xor \U$4139 ( \4428 , \4399 , \4427 );
and \U$4140 ( \4429 , \4357 , \4389 );
nor \U$4141 ( \4430 , \4428 , \4429 );
nor \U$4142 ( \4431 , \4395 , \4430 );
nand \U$4143 ( \4432 , \4353 , \4431 );
and \U$4144 ( \4433 , \4403 , \4404 );
and \U$4145 ( \4434 , \4404 , \4426 );
and \U$4146 ( \4435 , \4403 , \4426 );
or \U$4147 ( \4436 , \4433 , \4434 , \4435 );
and \U$4148 ( \4437 , \4409 , \4411 );
and \U$4149 ( \4438 , \4411 , \4425 );
and \U$4150 ( \4439 , \4409 , \4425 );
or \U$4151 ( \4440 , \4437 , \4438 , \4439 );
not \U$4152 ( \4441 , \628 );
and \U$4153 ( \4442 , \568 , \1233 );
and \U$4154 ( \4443 , \227 , \1114 );
nor \U$4155 ( \4444 , \4442 , \4443 );
xnor \U$4156 ( \4445 , \4444 , \594 );
xor \U$4157 ( \4446 , \4441 , \4445 );
and \U$4158 ( \4447 , \1055 , \561 );
and \U$4159 ( \4448 , \601 , \559 );
nor \U$4160 ( \4449 , \4447 , \4448 );
xnor \U$4161 ( \4450 , \4449 , \566 );
xor \U$4162 ( \4451 , \4446 , \4450 );
xor \U$4163 ( \4452 , \4440 , \4451 );
and \U$4164 ( \4453 , \4415 , \4419 );
and \U$4165 ( \4454 , \4419 , \4424 );
and \U$4166 ( \4455 , \4415 , \4424 );
or \U$4167 ( \4456 , \4453 , \4454 , \4455 );
not \U$4168 ( \4457 , \4411 );
xor \U$4169 ( \4458 , \4456 , \4457 );
and \U$4171 ( \4459 , \1053 , \569 );
nor \U$4172 ( \4460 , 1'b0 , \4459 );
not \U$4173 ( \4461 , \4460 );
xor \U$4174 ( \4462 , \4458 , \4461 );
xor \U$4175 ( \4463 , \4452 , \4462 );
xor \U$4176 ( \4464 , \4436 , \4463 );
and \U$4177 ( \4465 , \4399 , \4427 );
nor \U$4178 ( \4466 , \4464 , \4465 );
and \U$4179 ( \4467 , \4440 , \4451 );
and \U$4180 ( \4468 , \4451 , \4462 );
and \U$4181 ( \4469 , \4440 , \4462 );
or \U$4182 ( \4470 , \4467 , \4468 , \4469 );
and \U$4183 ( \4471 , \4456 , \4457 );
and \U$4184 ( \4472 , \4457 , \4461 );
and \U$4185 ( \4473 , \4456 , \4461 );
or \U$4186 ( \4474 , \4471 , \4472 , \4473 );
xor \U$4187 ( \4475 , \4470 , \4474 );
and \U$4188 ( \4476 , \4441 , \4445 );
and \U$4189 ( \4477 , \4445 , \4450 );
and \U$4190 ( \4478 , \4441 , \4450 );
or \U$4191 ( \4479 , \4476 , \4477 , \4478 );
and \U$4192 ( \4480 , \227 , \1233 );
not \U$4193 ( \4481 , \4480 );
xnor \U$4194 ( \4482 , \4481 , \594 );
and \U$4195 ( \4483 , \601 , \561 );
and \U$4196 ( \4484 , \568 , \559 );
nor \U$4197 ( \4485 , \4483 , \4484 );
xnor \U$4198 ( \4486 , \4485 , \566 );
xor \U$4199 ( \4487 , \4482 , \4486 );
and \U$4201 ( \4488 , \1055 , \569 );
nor \U$4202 ( \4489 , 1'b0 , \4488 );
not \U$4203 ( \4490 , \4489 );
xor \U$4204 ( \4491 , \4487 , \4490 );
xnor \U$4205 ( \4492 , \4479 , \4491 );
xor \U$4206 ( \4493 , \4475 , \4492 );
and \U$4207 ( \4494 , \4436 , \4463 );
nor \U$4208 ( \4495 , \4493 , \4494 );
nor \U$4209 ( \4496 , \4466 , \4495 );
or \U$4210 ( \4497 , \4479 , \4491 );
and \U$4211 ( \4498 , \4482 , \4486 );
and \U$4212 ( \4499 , \4486 , \4490 );
and \U$4213 ( \4500 , \4482 , \4490 );
or \U$4214 ( \4501 , \4498 , \4499 , \4500 );
xor \U$4215 ( \4502 , \4497 , \4501 );
xor \U$4216 ( \4503 , \595 , \599 );
xor \U$4217 ( \4504 , \4503 , \604 );
xor \U$4218 ( \4505 , \4502 , \4504 );
and \U$4219 ( \4506 , \4470 , \4474 );
and \U$4220 ( \4507 , \4474 , \4492 );
and \U$4221 ( \4508 , \4470 , \4492 );
or \U$4222 ( \4509 , \4506 , \4507 , \4508 );
nor \U$4223 ( \4510 , \4505 , \4509 );
xor \U$4224 ( \4511 , \607 , \608 );
and \U$4225 ( \4512 , \4497 , \4501 );
and \U$4226 ( \4513 , \4501 , \4504 );
and \U$4227 ( \4514 , \4497 , \4504 );
or \U$4228 ( \4515 , \4512 , \4513 , \4514 );
nor \U$4229 ( \4516 , \4511 , \4515 );
nor \U$4230 ( \4517 , \4510 , \4516 );
nand \U$4231 ( \4518 , \4496 , \4517 );
nor \U$4232 ( \4519 , \4432 , \4518 );
nand \U$4233 ( \4520 , \4252 , \4519 );
nor \U$4234 ( \4521 , \3645 , \4520 );
and \U$4235 ( \4522 , \840 , \674 );
and \U$4236 ( \4523 , \858 , \671 );
nor \U$4237 ( \4524 , \4522 , \4523 );
xnor \U$4238 ( \4525 , \4524 , \635 );
and \U$4239 ( \4526 , \837 , \4525 );
and \U$4240 ( \4527 , \871 , \697 );
and \U$4241 ( \4528 , \889 , \695 );
nor \U$4242 ( \4529 , \4527 , \4528 );
xnor \U$4243 ( \4530 , \4529 , \704 );
and \U$4244 ( \4531 , \4525 , \4530 );
and \U$4245 ( \4532 , \837 , \4530 );
or \U$4246 ( \4533 , \4526 , \4531 , \4532 );
and \U$4247 ( \4534 , \896 , \725 );
and \U$4248 ( \4535 , \914 , \723 );
nor \U$4249 ( \4536 , \4534 , \4535 );
xnor \U$4250 ( \4537 , \4536 , \732 );
and \U$4251 ( \4538 , \922 , \750 );
and \U$4252 ( \4539 , \940 , \748 );
nor \U$4253 ( \4540 , \4538 , \4539 );
xnor \U$4254 ( \4541 , \4540 , \757 );
and \U$4255 ( \4542 , \4537 , \4541 );
and \U$4256 ( \4543 , \950 , \776 );
and \U$4257 ( \4544 , \968 , \774 );
nor \U$4258 ( \4545 , \4543 , \4544 );
xnor \U$4259 ( \4546 , \4545 , \783 );
and \U$4260 ( \4547 , \4541 , \4546 );
and \U$4261 ( \4548 , \4537 , \4546 );
or \U$4262 ( \4549 , \4542 , \4547 , \4548 );
and \U$4263 ( \4550 , \4533 , \4549 );
and \U$4264 ( \4551 , \995 , \830 );
and \U$4265 ( \4552 , \975 , \828 );
nor \U$4266 ( \4553 , \4551 , \4552 );
xnor \U$4267 ( \4554 , \4553 , \837 );
and \U$4268 ( \4555 , \4549 , \4554 );
and \U$4269 ( \4556 , \4533 , \4554 );
or \U$4270 ( \4557 , \4550 , \4555 , \4556 );
and \U$4271 ( \4558 , \871 , \725 );
and \U$4272 ( \4559 , \889 , \723 );
nor \U$4273 ( \4560 , \4558 , \4559 );
xnor \U$4274 ( \4561 , \4560 , \732 );
and \U$4275 ( \4562 , \896 , \750 );
and \U$4276 ( \4563 , \914 , \748 );
nor \U$4277 ( \4564 , \4562 , \4563 );
xnor \U$4278 ( \4565 , \4564 , \757 );
xor \U$4279 ( \4566 , \4561 , \4565 );
and \U$4280 ( \4567 , \922 , \776 );
and \U$4281 ( \4568 , \940 , \774 );
nor \U$4282 ( \4569 , \4567 , \4568 );
xnor \U$4283 ( \4570 , \4569 , \783 );
xor \U$4284 ( \4571 , \4566 , \4570 );
and \U$4285 ( \4572 , \814 , \674 );
and \U$4286 ( \4573 , \832 , \671 );
nor \U$4287 ( \4574 , \4572 , \4573 );
xnor \U$4288 ( \4575 , \4574 , \635 );
xor \U$4289 ( \4576 , \863 , \4575 );
and \U$4290 ( \4577 , \840 , \697 );
and \U$4291 ( \4578 , \858 , \695 );
nor \U$4292 ( \4579 , \4577 , \4578 );
xnor \U$4293 ( \4580 , \4579 , \704 );
xor \U$4294 ( \4581 , \4576 , \4580 );
xor \U$4295 ( \4582 , \4571 , \4581 );
and \U$4296 ( \4583 , \4557 , \4582 );
and \U$4297 ( \4584 , \858 , \674 );
and \U$4298 ( \4585 , \814 , \671 );
nor \U$4299 ( \4586 , \4584 , \4585 );
xnor \U$4300 ( \4587 , \4586 , \635 );
and \U$4301 ( \4588 , \889 , \697 );
and \U$4302 ( \4589 , \840 , \695 );
nor \U$4303 ( \4590 , \4588 , \4589 );
xnor \U$4304 ( \4591 , \4590 , \704 );
and \U$4305 ( \4592 , \4587 , \4591 );
and \U$4306 ( \4593 , \914 , \725 );
and \U$4307 ( \4594 , \871 , \723 );
nor \U$4308 ( \4595 , \4593 , \4594 );
xnor \U$4309 ( \4596 , \4595 , \732 );
and \U$4310 ( \4597 , \4591 , \4596 );
and \U$4311 ( \4598 , \4587 , \4596 );
or \U$4312 ( \4599 , \4592 , \4597 , \4598 );
and \U$4313 ( \4600 , \940 , \750 );
and \U$4314 ( \4601 , \896 , \748 );
nor \U$4315 ( \4602 , \4600 , \4601 );
xnor \U$4316 ( \4603 , \4602 , \757 );
and \U$4317 ( \4604 , \968 , \776 );
and \U$4318 ( \4605 , \922 , \774 );
nor \U$4319 ( \4606 , \4604 , \4605 );
xnor \U$4320 ( \4607 , \4606 , \783 );
and \U$4321 ( \4608 , \4603 , \4607 );
and \U$4322 ( \4609 , \987 , \805 );
and \U$4323 ( \4610 , \950 , \803 );
nor \U$4324 ( \4611 , \4609 , \4610 );
xnor \U$4325 ( \4612 , \4611 , \812 );
and \U$4326 ( \4613 , \4607 , \4612 );
and \U$4327 ( \4614 , \4603 , \4612 );
or \U$4328 ( \4615 , \4608 , \4613 , \4614 );
xor \U$4329 ( \4616 , \4599 , \4615 );
and \U$4330 ( \4617 , \950 , \805 );
and \U$4331 ( \4618 , \968 , \803 );
nor \U$4332 ( \4619 , \4617 , \4618 );
xnor \U$4333 ( \4620 , \4619 , \812 );
and \U$4334 ( \4621 , \975 , \830 );
and \U$4335 ( \4622 , \987 , \828 );
nor \U$4336 ( \4623 , \4621 , \4622 );
xnor \U$4337 ( \4624 , \4623 , \837 );
xor \U$4338 ( \4625 , \4620 , \4624 );
nand \U$4339 ( \4626 , \995 , \854 );
xnor \U$4340 ( \4627 , \4626 , \863 );
xor \U$4341 ( \4628 , \4625 , \4627 );
xor \U$4342 ( \4629 , \4616 , \4628 );
and \U$4343 ( \4630 , \4582 , \4629 );
and \U$4344 ( \4631 , \4557 , \4629 );
or \U$4345 ( \4632 , \4583 , \4630 , \4631 );
and \U$4346 ( \4633 , \863 , \4575 );
and \U$4347 ( \4634 , \4575 , \4580 );
and \U$4348 ( \4635 , \863 , \4580 );
or \U$4349 ( \4636 , \4633 , \4634 , \4635 );
and \U$4350 ( \4637 , \4561 , \4565 );
and \U$4351 ( \4638 , \4565 , \4570 );
and \U$4352 ( \4639 , \4561 , \4570 );
or \U$4353 ( \4640 , \4637 , \4638 , \4639 );
xor \U$4354 ( \4641 , \4636 , \4640 );
and \U$4355 ( \4642 , \4620 , \4624 );
and \U$4356 ( \4643 , \4624 , \4627 );
and \U$4357 ( \4644 , \4620 , \4627 );
or \U$4358 ( \4645 , \4642 , \4643 , \4644 );
xor \U$4359 ( \4646 , \4641 , \4645 );
xor \U$4360 ( \4647 , \4632 , \4646 );
and \U$4361 ( \4648 , \4599 , \4615 );
and \U$4362 ( \4649 , \4615 , \4628 );
and \U$4363 ( \4650 , \4599 , \4628 );
or \U$4364 ( \4651 , \4648 , \4649 , \4650 );
and \U$4365 ( \4652 , \4571 , \4581 );
xor \U$4366 ( \4653 , \4651 , \4652 );
and \U$4367 ( \4654 , \987 , \830 );
and \U$4368 ( \4655 , \950 , \828 );
nor \U$4369 ( \4656 , \4654 , \4655 );
xnor \U$4370 ( \4657 , \4656 , \837 );
and \U$4371 ( \4658 , \995 , \856 );
and \U$4372 ( \4659 , \975 , \854 );
nor \U$4373 ( \4660 , \4658 , \4659 );
xnor \U$4374 ( \4661 , \4660 , \863 );
xor \U$4375 ( \4662 , \4657 , \4661 );
and \U$4376 ( \4663 , \914 , \750 );
and \U$4377 ( \4664 , \871 , \748 );
nor \U$4378 ( \4665 , \4663 , \4664 );
xnor \U$4379 ( \4666 , \4665 , \757 );
and \U$4380 ( \4667 , \940 , \776 );
and \U$4381 ( \4668 , \896 , \774 );
nor \U$4382 ( \4669 , \4667 , \4668 );
xnor \U$4383 ( \4670 , \4669 , \783 );
xor \U$4384 ( \4671 , \4666 , \4670 );
and \U$4385 ( \4672 , \968 , \805 );
and \U$4386 ( \4673 , \922 , \803 );
nor \U$4387 ( \4674 , \4672 , \4673 );
xnor \U$4388 ( \4675 , \4674 , \812 );
xor \U$4389 ( \4676 , \4671 , \4675 );
xor \U$4390 ( \4677 , \4662 , \4676 );
and \U$4391 ( \4678 , \832 , \674 );
and \U$4392 ( \4679 , \789 , \671 );
nor \U$4393 ( \4680 , \4678 , \4679 );
xnor \U$4394 ( \4681 , \4680 , \635 );
and \U$4395 ( \4682 , \858 , \697 );
and \U$4396 ( \4683 , \814 , \695 );
nor \U$4397 ( \4684 , \4682 , \4683 );
xnor \U$4398 ( \4685 , \4684 , \704 );
xor \U$4399 ( \4686 , \4681 , \4685 );
and \U$4400 ( \4687 , \889 , \725 );
and \U$4401 ( \4688 , \840 , \723 );
nor \U$4402 ( \4689 , \4687 , \4688 );
xnor \U$4403 ( \4690 , \4689 , \732 );
xor \U$4404 ( \4691 , \4686 , \4690 );
xor \U$4405 ( \4692 , \4677 , \4691 );
xor \U$4406 ( \4693 , \4653 , \4692 );
xor \U$4407 ( \4694 , \4647 , \4693 );
and \U$4408 ( \4695 , \889 , \674 );
and \U$4409 ( \4696 , \840 , \671 );
nor \U$4410 ( \4697 , \4695 , \4696 );
xnor \U$4411 ( \4698 , \4697 , \635 );
and \U$4412 ( \4699 , \914 , \697 );
and \U$4413 ( \4700 , \871 , \695 );
nor \U$4414 ( \4701 , \4699 , \4700 );
xnor \U$4415 ( \4702 , \4701 , \704 );
and \U$4416 ( \4703 , \4698 , \4702 );
and \U$4417 ( \4704 , \940 , \725 );
and \U$4418 ( \4705 , \896 , \723 );
nor \U$4419 ( \4706 , \4704 , \4705 );
xnor \U$4420 ( \4707 , \4706 , \732 );
and \U$4421 ( \4708 , \4702 , \4707 );
and \U$4422 ( \4709 , \4698 , \4707 );
or \U$4423 ( \4710 , \4703 , \4708 , \4709 );
and \U$4424 ( \4711 , \968 , \750 );
and \U$4425 ( \4712 , \922 , \748 );
nor \U$4426 ( \4713 , \4711 , \4712 );
xnor \U$4427 ( \4714 , \4713 , \757 );
and \U$4428 ( \4715 , \987 , \776 );
and \U$4429 ( \4716 , \950 , \774 );
nor \U$4430 ( \4717 , \4715 , \4716 );
xnor \U$4431 ( \4718 , \4717 , \783 );
and \U$4432 ( \4719 , \4714 , \4718 );
and \U$4433 ( \4720 , \995 , \805 );
and \U$4434 ( \4721 , \975 , \803 );
nor \U$4435 ( \4722 , \4720 , \4721 );
xnor \U$4436 ( \4723 , \4722 , \812 );
and \U$4437 ( \4724 , \4718 , \4723 );
and \U$4438 ( \4725 , \4714 , \4723 );
or \U$4439 ( \4726 , \4719 , \4724 , \4725 );
and \U$4440 ( \4727 , \4710 , \4726 );
and \U$4441 ( \4728 , \975 , \805 );
and \U$4442 ( \4729 , \987 , \803 );
nor \U$4443 ( \4730 , \4728 , \4729 );
xnor \U$4444 ( \4731 , \4730 , \812 );
and \U$4445 ( \4732 , \4726 , \4731 );
and \U$4446 ( \4733 , \4710 , \4731 );
or \U$4447 ( \4734 , \4727 , \4732 , \4733 );
nand \U$4448 ( \4735 , \995 , \828 );
xnor \U$4449 ( \4736 , \4735 , \837 );
xor \U$4450 ( \4737 , \4537 , \4541 );
xor \U$4451 ( \4738 , \4737 , \4546 );
and \U$4452 ( \4739 , \4736 , \4738 );
xor \U$4453 ( \4740 , \837 , \4525 );
xor \U$4454 ( \4741 , \4740 , \4530 );
and \U$4455 ( \4742 , \4738 , \4741 );
and \U$4456 ( \4743 , \4736 , \4741 );
or \U$4457 ( \4744 , \4739 , \4742 , \4743 );
and \U$4458 ( \4745 , \4734 , \4744 );
xor \U$4459 ( \4746 , \4603 , \4607 );
xor \U$4460 ( \4747 , \4746 , \4612 );
and \U$4461 ( \4748 , \4744 , \4747 );
and \U$4462 ( \4749 , \4734 , \4747 );
or \U$4463 ( \4750 , \4745 , \4748 , \4749 );
xor \U$4464 ( \4751 , \4587 , \4591 );
xor \U$4465 ( \4752 , \4751 , \4596 );
xor \U$4466 ( \4753 , \4533 , \4549 );
xor \U$4467 ( \4754 , \4753 , \4554 );
and \U$4468 ( \4755 , \4752 , \4754 );
and \U$4469 ( \4756 , \4750 , \4755 );
xor \U$4470 ( \4757 , \4557 , \4582 );
xor \U$4471 ( \4758 , \4757 , \4629 );
and \U$4472 ( \4759 , \4755 , \4758 );
and \U$4473 ( \4760 , \4750 , \4758 );
or \U$4474 ( \4761 , \4756 , \4759 , \4760 );
nor \U$4475 ( \4762 , \4694 , \4761 );
and \U$4476 ( \4763 , \4651 , \4652 );
and \U$4477 ( \4764 , \4652 , \4692 );
and \U$4478 ( \4765 , \4651 , \4692 );
or \U$4479 ( \4766 , \4763 , \4764 , \4765 );
nand \U$4480 ( \4767 , \995 , \885 );
xnor \U$4481 ( \4768 , \4767 , \894 );
and \U$4482 ( \4769 , \922 , \805 );
and \U$4483 ( \4770 , \940 , \803 );
nor \U$4484 ( \4771 , \4769 , \4770 );
xnor \U$4485 ( \4772 , \4771 , \812 );
and \U$4486 ( \4773 , \950 , \830 );
and \U$4487 ( \4774 , \968 , \828 );
nor \U$4488 ( \4775 , \4773 , \4774 );
xnor \U$4489 ( \4776 , \4775 , \837 );
xor \U$4490 ( \4777 , \4772 , \4776 );
and \U$4491 ( \4778 , \975 , \856 );
and \U$4492 ( \4779 , \987 , \854 );
nor \U$4493 ( \4780 , \4778 , \4779 );
xnor \U$4494 ( \4781 , \4780 , \863 );
xor \U$4495 ( \4782 , \4777 , \4781 );
xor \U$4496 ( \4783 , \4768 , \4782 );
and \U$4497 ( \4784 , \840 , \725 );
and \U$4498 ( \4785 , \858 , \723 );
nor \U$4499 ( \4786 , \4784 , \4785 );
xnor \U$4500 ( \4787 , \4786 , \732 );
and \U$4501 ( \4788 , \871 , \750 );
and \U$4502 ( \4789 , \889 , \748 );
nor \U$4503 ( \4790 , \4788 , \4789 );
xnor \U$4504 ( \4791 , \4790 , \757 );
xor \U$4505 ( \4792 , \4787 , \4791 );
and \U$4506 ( \4793 , \896 , \776 );
and \U$4507 ( \4794 , \914 , \774 );
nor \U$4508 ( \4795 , \4793 , \4794 );
xnor \U$4509 ( \4796 , \4795 , \783 );
xor \U$4510 ( \4797 , \4792 , \4796 );
xor \U$4511 ( \4798 , \4783 , \4797 );
and \U$4512 ( \4799 , \4681 , \4685 );
and \U$4513 ( \4800 , \4685 , \4690 );
and \U$4514 ( \4801 , \4681 , \4690 );
or \U$4515 ( \4802 , \4799 , \4800 , \4801 );
and \U$4516 ( \4803 , \4666 , \4670 );
and \U$4517 ( \4804 , \4670 , \4675 );
and \U$4518 ( \4805 , \4666 , \4675 );
or \U$4519 ( \4806 , \4803 , \4804 , \4805 );
xor \U$4520 ( \4807 , \4802 , \4806 );
and \U$4521 ( \4808 , \4657 , \4661 );
xor \U$4522 ( \4809 , \4807 , \4808 );
xor \U$4523 ( \4810 , \4798 , \4809 );
xor \U$4524 ( \4811 , \4766 , \4810 );
and \U$4525 ( \4812 , \4636 , \4640 );
and \U$4526 ( \4813 , \4640 , \4645 );
and \U$4527 ( \4814 , \4636 , \4645 );
or \U$4528 ( \4815 , \4812 , \4813 , \4814 );
and \U$4529 ( \4816 , \4662 , \4676 );
and \U$4530 ( \4817 , \4676 , \4691 );
and \U$4531 ( \4818 , \4662 , \4691 );
or \U$4532 ( \4819 , \4816 , \4817 , \4818 );
xor \U$4533 ( \4820 , \4815 , \4819 );
and \U$4534 ( \4821 , \789 , \674 );
and \U$4535 ( \4822 , \807 , \671 );
nor \U$4536 ( \4823 , \4821 , \4822 );
xnor \U$4537 ( \4824 , \4823 , \635 );
xor \U$4538 ( \4825 , \894 , \4824 );
and \U$4539 ( \4826 , \814 , \697 );
and \U$4540 ( \4827 , \832 , \695 );
nor \U$4541 ( \4828 , \4826 , \4827 );
xnor \U$4542 ( \4829 , \4828 , \704 );
xor \U$4543 ( \4830 , \4825 , \4829 );
xor \U$4544 ( \4831 , \4820 , \4830 );
xor \U$4545 ( \4832 , \4811 , \4831 );
and \U$4546 ( \4833 , \4632 , \4646 );
and \U$4547 ( \4834 , \4646 , \4693 );
and \U$4548 ( \4835 , \4632 , \4693 );
or \U$4549 ( \4836 , \4833 , \4834 , \4835 );
nor \U$4550 ( \4837 , \4832 , \4836 );
nor \U$4551 ( \4838 , \4762 , \4837 );
and \U$4552 ( \4839 , \4802 , \4806 );
and \U$4553 ( \4840 , \4806 , \4808 );
and \U$4554 ( \4841 , \4802 , \4808 );
or \U$4555 ( \4842 , \4839 , \4840 , \4841 );
and \U$4556 ( \4843 , \4768 , \4782 );
and \U$4557 ( \4844 , \4782 , \4797 );
and \U$4558 ( \4845 , \4768 , \4797 );
or \U$4559 ( \4846 , \4843 , \4844 , \4845 );
xor \U$4560 ( \4847 , \4842 , \4846 );
and \U$4561 ( \4848 , \968 , \830 );
and \U$4562 ( \4849 , \922 , \828 );
nor \U$4563 ( \4850 , \4848 , \4849 );
xnor \U$4564 ( \4851 , \4850 , \837 );
and \U$4565 ( \4852 , \987 , \856 );
and \U$4566 ( \4853 , \950 , \854 );
nor \U$4567 ( \4854 , \4852 , \4853 );
xnor \U$4568 ( \4855 , \4854 , \863 );
xor \U$4569 ( \4856 , \4851 , \4855 );
and \U$4570 ( \4857 , \995 , \887 );
and \U$4571 ( \4858 , \975 , \885 );
nor \U$4572 ( \4859 , \4857 , \4858 );
xnor \U$4573 ( \4860 , \4859 , \894 );
xor \U$4574 ( \4861 , \4856 , \4860 );
and \U$4575 ( \4862 , \889 , \750 );
and \U$4576 ( \4863 , \840 , \748 );
nor \U$4577 ( \4864 , \4862 , \4863 );
xnor \U$4578 ( \4865 , \4864 , \757 );
and \U$4579 ( \4866 , \914 , \776 );
and \U$4580 ( \4867 , \871 , \774 );
nor \U$4581 ( \4868 , \4866 , \4867 );
xnor \U$4582 ( \4869 , \4868 , \783 );
xor \U$4583 ( \4870 , \4865 , \4869 );
and \U$4584 ( \4871 , \940 , \805 );
and \U$4585 ( \4872 , \896 , \803 );
nor \U$4586 ( \4873 , \4871 , \4872 );
xnor \U$4587 ( \4874 , \4873 , \812 );
xor \U$4588 ( \4875 , \4870 , \4874 );
xor \U$4589 ( \4876 , \4861 , \4875 );
and \U$4590 ( \4877 , \807 , \674 );
and \U$4591 ( \4878 , \760 , \671 );
nor \U$4592 ( \4879 , \4877 , \4878 );
xnor \U$4593 ( \4880 , \4879 , \635 );
and \U$4594 ( \4881 , \832 , \697 );
and \U$4595 ( \4882 , \789 , \695 );
nor \U$4596 ( \4883 , \4881 , \4882 );
xnor \U$4597 ( \4884 , \4883 , \704 );
xor \U$4598 ( \4885 , \4880 , \4884 );
and \U$4599 ( \4886 , \858 , \725 );
and \U$4600 ( \4887 , \814 , \723 );
nor \U$4601 ( \4888 , \4886 , \4887 );
xnor \U$4602 ( \4889 , \4888 , \732 );
xor \U$4603 ( \4890 , \4885 , \4889 );
xor \U$4604 ( \4891 , \4876 , \4890 );
xor \U$4605 ( \4892 , \4847 , \4891 );
and \U$4606 ( \4893 , \4815 , \4819 );
and \U$4607 ( \4894 , \4819 , \4830 );
and \U$4608 ( \4895 , \4815 , \4830 );
or \U$4609 ( \4896 , \4893 , \4894 , \4895 );
and \U$4610 ( \4897 , \4798 , \4809 );
xor \U$4611 ( \4898 , \4896 , \4897 );
and \U$4612 ( \4899 , \894 , \4824 );
and \U$4613 ( \4900 , \4824 , \4829 );
and \U$4614 ( \4901 , \894 , \4829 );
or \U$4615 ( \4902 , \4899 , \4900 , \4901 );
and \U$4616 ( \4903 , \4787 , \4791 );
and \U$4617 ( \4904 , \4791 , \4796 );
and \U$4618 ( \4905 , \4787 , \4796 );
or \U$4619 ( \4906 , \4903 , \4904 , \4905 );
xor \U$4620 ( \4907 , \4902 , \4906 );
and \U$4621 ( \4908 , \4772 , \4776 );
and \U$4622 ( \4909 , \4776 , \4781 );
and \U$4623 ( \4910 , \4772 , \4781 );
or \U$4624 ( \4911 , \4908 , \4909 , \4910 );
xor \U$4625 ( \4912 , \4907 , \4911 );
xor \U$4626 ( \4913 , \4898 , \4912 );
xor \U$4627 ( \4914 , \4892 , \4913 );
and \U$4628 ( \4915 , \4766 , \4810 );
and \U$4629 ( \4916 , \4810 , \4831 );
and \U$4630 ( \4917 , \4766 , \4831 );
or \U$4631 ( \4918 , \4915 , \4916 , \4917 );
nor \U$4632 ( \4919 , \4914 , \4918 );
and \U$4633 ( \4920 , \4896 , \4897 );
and \U$4634 ( \4921 , \4897 , \4912 );
and \U$4635 ( \4922 , \4896 , \4912 );
or \U$4636 ( \4923 , \4920 , \4921 , \4922 );
and \U$4637 ( \4924 , \4842 , \4846 );
and \U$4638 ( \4925 , \4846 , \4891 );
and \U$4639 ( \4926 , \4842 , \4891 );
or \U$4640 ( \4927 , \4924 , \4925 , \4926 );
and \U$4641 ( \4928 , \760 , \674 );
and \U$4642 ( \4929 , \778 , \671 );
nor \U$4643 ( \4930 , \4928 , \4929 );
xnor \U$4644 ( \4931 , \4930 , \635 );
xor \U$4645 ( \4932 , \919 , \4931 );
and \U$4646 ( \4933 , \789 , \697 );
and \U$4647 ( \4934 , \807 , \695 );
nor \U$4648 ( \4935 , \4933 , \4934 );
xnor \U$4649 ( \4936 , \4935 , \704 );
xor \U$4650 ( \4937 , \4932 , \4936 );
and \U$4651 ( \4938 , \975 , \887 );
and \U$4652 ( \4939 , \987 , \885 );
nor \U$4653 ( \4940 , \4938 , \4939 );
xnor \U$4654 ( \4941 , \4940 , \894 );
nand \U$4655 ( \4942 , \995 , \910 );
xnor \U$4656 ( \4943 , \4942 , \919 );
xor \U$4657 ( \4944 , \4941 , \4943 );
and \U$4658 ( \4945 , \896 , \805 );
and \U$4659 ( \4946 , \914 , \803 );
nor \U$4660 ( \4947 , \4945 , \4946 );
xnor \U$4661 ( \4948 , \4947 , \812 );
and \U$4662 ( \4949 , \922 , \830 );
and \U$4663 ( \4950 , \940 , \828 );
nor \U$4664 ( \4951 , \4949 , \4950 );
xnor \U$4665 ( \4952 , \4951 , \837 );
xor \U$4666 ( \4953 , \4948 , \4952 );
and \U$4667 ( \4954 , \950 , \856 );
and \U$4668 ( \4955 , \968 , \854 );
nor \U$4669 ( \4956 , \4954 , \4955 );
xnor \U$4670 ( \4957 , \4956 , \863 );
xor \U$4671 ( \4958 , \4953 , \4957 );
xor \U$4672 ( \4959 , \4944 , \4958 );
xor \U$4673 ( \4960 , \4937 , \4959 );
and \U$4674 ( \4961 , \4880 , \4884 );
and \U$4675 ( \4962 , \4884 , \4889 );
and \U$4676 ( \4963 , \4880 , \4889 );
or \U$4677 ( \4964 , \4961 , \4962 , \4963 );
and \U$4678 ( \4965 , \4865 , \4869 );
and \U$4679 ( \4966 , \4869 , \4874 );
and \U$4680 ( \4967 , \4865 , \4874 );
or \U$4681 ( \4968 , \4965 , \4966 , \4967 );
xor \U$4682 ( \4969 , \4964 , \4968 );
and \U$4683 ( \4970 , \4851 , \4855 );
and \U$4684 ( \4971 , \4855 , \4860 );
and \U$4685 ( \4972 , \4851 , \4860 );
or \U$4686 ( \4973 , \4970 , \4971 , \4972 );
xor \U$4687 ( \4974 , \4969 , \4973 );
xor \U$4688 ( \4975 , \4960 , \4974 );
xor \U$4689 ( \4976 , \4927 , \4975 );
and \U$4690 ( \4977 , \4902 , \4906 );
and \U$4691 ( \4978 , \4906 , \4911 );
and \U$4692 ( \4979 , \4902 , \4911 );
or \U$4693 ( \4980 , \4977 , \4978 , \4979 );
and \U$4694 ( \4981 , \4861 , \4875 );
and \U$4695 ( \4982 , \4875 , \4890 );
and \U$4696 ( \4983 , \4861 , \4890 );
or \U$4697 ( \4984 , \4981 , \4982 , \4983 );
xor \U$4698 ( \4985 , \4980 , \4984 );
and \U$4699 ( \4986 , \814 , \725 );
and \U$4700 ( \4987 , \832 , \723 );
nor \U$4701 ( \4988 , \4986 , \4987 );
xnor \U$4702 ( \4989 , \4988 , \732 );
and \U$4703 ( \4990 , \840 , \750 );
and \U$4704 ( \4991 , \858 , \748 );
nor \U$4705 ( \4992 , \4990 , \4991 );
xnor \U$4706 ( \4993 , \4992 , \757 );
xor \U$4707 ( \4994 , \4989 , \4993 );
and \U$4708 ( \4995 , \871 , \776 );
and \U$4709 ( \4996 , \889 , \774 );
nor \U$4710 ( \4997 , \4995 , \4996 );
xnor \U$4711 ( \4998 , \4997 , \783 );
xor \U$4712 ( \4999 , \4994 , \4998 );
xor \U$4713 ( \5000 , \4985 , \4999 );
xor \U$4714 ( \5001 , \4976 , \5000 );
xor \U$4715 ( \5002 , \4923 , \5001 );
and \U$4716 ( \5003 , \4892 , \4913 );
nor \U$4717 ( \5004 , \5002 , \5003 );
nor \U$4718 ( \5005 , \4919 , \5004 );
nand \U$4719 ( \5006 , \4838 , \5005 );
and \U$4720 ( \5007 , \4927 , \4975 );
and \U$4721 ( \5008 , \4975 , \5000 );
and \U$4722 ( \5009 , \4927 , \5000 );
or \U$4723 ( \5010 , \5007 , \5008 , \5009 );
and \U$4724 ( \5011 , \919 , \4931 );
and \U$4725 ( \5012 , \4931 , \4936 );
and \U$4726 ( \5013 , \919 , \4936 );
or \U$4727 ( \5014 , \5011 , \5012 , \5013 );
and \U$4728 ( \5015 , \4989 , \4993 );
and \U$4729 ( \5016 , \4993 , \4998 );
and \U$4730 ( \5017 , \4989 , \4998 );
or \U$4731 ( \5018 , \5015 , \5016 , \5017 );
xor \U$4732 ( \5019 , \5014 , \5018 );
and \U$4733 ( \5020 , \4948 , \4952 );
and \U$4734 ( \5021 , \4952 , \4957 );
and \U$4735 ( \5022 , \4948 , \4957 );
or \U$4736 ( \5023 , \5020 , \5021 , \5022 );
xor \U$4737 ( \5024 , \5019 , \5023 );
and \U$4738 ( \5025 , \4964 , \4968 );
and \U$4739 ( \5026 , \4968 , \4973 );
and \U$4740 ( \5027 , \4964 , \4973 );
or \U$4741 ( \5028 , \5025 , \5026 , \5027 );
and \U$4742 ( \5029 , \4941 , \4943 );
and \U$4743 ( \5030 , \4943 , \4958 );
and \U$4744 ( \5031 , \4941 , \4958 );
or \U$4745 ( \5032 , \5029 , \5030 , \5031 );
xor \U$4746 ( \5033 , \5028 , \5032 );
and \U$4747 ( \5034 , \778 , \674 );
and \U$4748 ( \5035 , \734 , \671 );
nor \U$4749 ( \5036 , \5034 , \5035 );
xnor \U$4750 ( \5037 , \5036 , \635 );
and \U$4751 ( \5038 , \807 , \697 );
and \U$4752 ( \5039 , \760 , \695 );
nor \U$4753 ( \5040 , \5038 , \5039 );
xnor \U$4754 ( \5041 , \5040 , \704 );
xor \U$4755 ( \5042 , \5037 , \5041 );
and \U$4756 ( \5043 , \832 , \725 );
and \U$4757 ( \5044 , \789 , \723 );
nor \U$4758 ( \5045 , \5043 , \5044 );
xnor \U$4759 ( \5046 , \5045 , \732 );
xor \U$4760 ( \5047 , \5042 , \5046 );
xor \U$4761 ( \5048 , \5033 , \5047 );
xor \U$4762 ( \5049 , \5024 , \5048 );
xor \U$4763 ( \5050 , \5010 , \5049 );
and \U$4764 ( \5051 , \4980 , \4984 );
and \U$4765 ( \5052 , \4984 , \4999 );
and \U$4766 ( \5053 , \4980 , \4999 );
or \U$4767 ( \5054 , \5051 , \5052 , \5053 );
and \U$4768 ( \5055 , \4937 , \4959 );
and \U$4769 ( \5056 , \4959 , \4974 );
and \U$4770 ( \5057 , \4937 , \4974 );
or \U$4771 ( \5058 , \5055 , \5056 , \5057 );
xor \U$4772 ( \5059 , \5054 , \5058 );
and \U$4773 ( \5060 , \995 , \912 );
and \U$4774 ( \5061 , \975 , \910 );
nor \U$4775 ( \5062 , \5060 , \5061 );
xnor \U$4776 ( \5063 , \5062 , \919 );
and \U$4777 ( \5064 , \940 , \830 );
and \U$4778 ( \5065 , \896 , \828 );
nor \U$4779 ( \5066 , \5064 , \5065 );
xnor \U$4780 ( \5067 , \5066 , \837 );
and \U$4781 ( \5068 , \968 , \856 );
and \U$4782 ( \5069 , \922 , \854 );
nor \U$4783 ( \5070 , \5068 , \5069 );
xnor \U$4784 ( \5071 , \5070 , \863 );
xor \U$4785 ( \5072 , \5067 , \5071 );
and \U$4786 ( \5073 , \987 , \887 );
and \U$4787 ( \5074 , \950 , \885 );
nor \U$4788 ( \5075 , \5073 , \5074 );
xnor \U$4789 ( \5076 , \5075 , \894 );
xor \U$4790 ( \5077 , \5072 , \5076 );
xor \U$4791 ( \5078 , \5063 , \5077 );
and \U$4792 ( \5079 , \858 , \750 );
and \U$4793 ( \5080 , \814 , \748 );
nor \U$4794 ( \5081 , \5079 , \5080 );
xnor \U$4795 ( \5082 , \5081 , \757 );
and \U$4796 ( \5083 , \889 , \776 );
and \U$4797 ( \5084 , \840 , \774 );
nor \U$4798 ( \5085 , \5083 , \5084 );
xnor \U$4799 ( \5086 , \5085 , \783 );
xor \U$4800 ( \5087 , \5082 , \5086 );
and \U$4801 ( \5088 , \914 , \805 );
and \U$4802 ( \5089 , \871 , \803 );
nor \U$4803 ( \5090 , \5088 , \5089 );
xnor \U$4804 ( \5091 , \5090 , \812 );
xor \U$4805 ( \5092 , \5087 , \5091 );
xor \U$4806 ( \5093 , \5078 , \5092 );
xor \U$4807 ( \5094 , \5059 , \5093 );
xor \U$4808 ( \5095 , \5050 , \5094 );
and \U$4809 ( \5096 , \4923 , \5001 );
nor \U$4810 ( \5097 , \5095 , \5096 );
and \U$4811 ( \5098 , \5054 , \5058 );
and \U$4812 ( \5099 , \5058 , \5093 );
and \U$4813 ( \5100 , \5054 , \5093 );
or \U$4814 ( \5101 , \5098 , \5099 , \5100 );
and \U$4815 ( \5102 , \5024 , \5048 );
xor \U$4816 ( \5103 , \5101 , \5102 );
and \U$4817 ( \5104 , \5028 , \5032 );
and \U$4818 ( \5105 , \5032 , \5047 );
and \U$4819 ( \5106 , \5028 , \5047 );
or \U$4820 ( \5107 , \5104 , \5105 , \5106 );
and \U$4821 ( \5108 , \950 , \887 );
and \U$4822 ( \5109 , \968 , \885 );
nor \U$4823 ( \5110 , \5108 , \5109 );
xnor \U$4824 ( \5111 , \5110 , \894 );
and \U$4825 ( \5112 , \975 , \912 );
and \U$4826 ( \5113 , \987 , \910 );
nor \U$4827 ( \5114 , \5112 , \5113 );
xnor \U$4828 ( \5115 , \5114 , \919 );
xor \U$4829 ( \5116 , \5111 , \5115 );
nand \U$4830 ( \5117 , \995 , \936 );
xnor \U$4831 ( \5118 , \5117 , \945 );
xor \U$4832 ( \5119 , \5116 , \5118 );
and \U$4833 ( \5120 , \871 , \805 );
and \U$4834 ( \5121 , \889 , \803 );
nor \U$4835 ( \5122 , \5120 , \5121 );
xnor \U$4836 ( \5123 , \5122 , \812 );
and \U$4837 ( \5124 , \896 , \830 );
and \U$4838 ( \5125 , \914 , \828 );
nor \U$4839 ( \5126 , \5124 , \5125 );
xnor \U$4840 ( \5127 , \5126 , \837 );
xor \U$4841 ( \5128 , \5123 , \5127 );
and \U$4842 ( \5129 , \922 , \856 );
and \U$4843 ( \5130 , \940 , \854 );
nor \U$4844 ( \5131 , \5129 , \5130 );
xnor \U$4845 ( \5132 , \5131 , \863 );
xor \U$4846 ( \5133 , \5128 , \5132 );
xor \U$4847 ( \5134 , \5119 , \5133 );
and \U$4848 ( \5135 , \789 , \725 );
and \U$4849 ( \5136 , \807 , \723 );
nor \U$4850 ( \5137 , \5135 , \5136 );
xnor \U$4851 ( \5138 , \5137 , \732 );
and \U$4852 ( \5139 , \814 , \750 );
and \U$4853 ( \5140 , \832 , \748 );
nor \U$4854 ( \5141 , \5139 , \5140 );
xnor \U$4855 ( \5142 , \5141 , \757 );
xor \U$4856 ( \5143 , \5138 , \5142 );
and \U$4857 ( \5144 , \840 , \776 );
and \U$4858 ( \5145 , \858 , \774 );
nor \U$4859 ( \5146 , \5144 , \5145 );
xnor \U$4860 ( \5147 , \5146 , \783 );
xor \U$4861 ( \5148 , \5143 , \5147 );
xor \U$4862 ( \5149 , \5134 , \5148 );
and \U$4863 ( \5150 , \5037 , \5041 );
and \U$4864 ( \5151 , \5041 , \5046 );
and \U$4865 ( \5152 , \5037 , \5046 );
or \U$4866 ( \5153 , \5150 , \5151 , \5152 );
and \U$4867 ( \5154 , \5082 , \5086 );
and \U$4868 ( \5155 , \5086 , \5091 );
and \U$4869 ( \5156 , \5082 , \5091 );
or \U$4870 ( \5157 , \5154 , \5155 , \5156 );
xor \U$4871 ( \5158 , \5153 , \5157 );
and \U$4872 ( \5159 , \5067 , \5071 );
and \U$4873 ( \5160 , \5071 , \5076 );
and \U$4874 ( \5161 , \5067 , \5076 );
or \U$4875 ( \5162 , \5159 , \5160 , \5161 );
xor \U$4876 ( \5163 , \5158 , \5162 );
xor \U$4877 ( \5164 , \5149 , \5163 );
xor \U$4878 ( \5165 , \5107 , \5164 );
and \U$4879 ( \5166 , \5014 , \5018 );
and \U$4880 ( \5167 , \5018 , \5023 );
and \U$4881 ( \5168 , \5014 , \5023 );
or \U$4882 ( \5169 , \5166 , \5167 , \5168 );
and \U$4883 ( \5170 , \5063 , \5077 );
and \U$4884 ( \5171 , \5077 , \5092 );
and \U$4885 ( \5172 , \5063 , \5092 );
or \U$4886 ( \5173 , \5170 , \5171 , \5172 );
xor \U$4887 ( \5174 , \5169 , \5173 );
and \U$4888 ( \5175 , \734 , \674 );
and \U$4889 ( \5176 , \752 , \671 );
nor \U$4890 ( \5177 , \5175 , \5176 );
xnor \U$4891 ( \5178 , \5177 , \635 );
xor \U$4892 ( \5179 , \945 , \5178 );
and \U$4893 ( \5180 , \760 , \697 );
and \U$4894 ( \5181 , \778 , \695 );
nor \U$4895 ( \5182 , \5180 , \5181 );
xnor \U$4896 ( \5183 , \5182 , \704 );
xor \U$4897 ( \5184 , \5179 , \5183 );
xor \U$4898 ( \5185 , \5174 , \5184 );
xor \U$4899 ( \5186 , \5165 , \5185 );
xor \U$4900 ( \5187 , \5103 , \5186 );
and \U$4901 ( \5188 , \5010 , \5049 );
and \U$4902 ( \5189 , \5049 , \5094 );
and \U$4903 ( \5190 , \5010 , \5094 );
or \U$4904 ( \5191 , \5188 , \5189 , \5190 );
nor \U$4905 ( \5192 , \5187 , \5191 );
nor \U$4906 ( \5193 , \5097 , \5192 );
and \U$4907 ( \5194 , \5107 , \5164 );
and \U$4908 ( \5195 , \5164 , \5185 );
and \U$4909 ( \5196 , \5107 , \5185 );
or \U$4910 ( \5197 , \5194 , \5195 , \5196 );
and \U$4911 ( \5198 , \945 , \5178 );
and \U$4912 ( \5199 , \5178 , \5183 );
and \U$4913 ( \5200 , \945 , \5183 );
or \U$4914 ( \5201 , \5198 , \5199 , \5200 );
and \U$4915 ( \5202 , \5138 , \5142 );
and \U$4916 ( \5203 , \5142 , \5147 );
and \U$4917 ( \5204 , \5138 , \5147 );
or \U$4918 ( \5205 , \5202 , \5203 , \5204 );
xor \U$4919 ( \5206 , \5201 , \5205 );
and \U$4920 ( \5207 , \5123 , \5127 );
and \U$4921 ( \5208 , \5127 , \5132 );
and \U$4922 ( \5209 , \5123 , \5132 );
or \U$4923 ( \5210 , \5207 , \5208 , \5209 );
xor \U$4924 ( \5211 , \5206 , \5210 );
and \U$4925 ( \5212 , \5153 , \5157 );
and \U$4926 ( \5213 , \5157 , \5162 );
and \U$4927 ( \5214 , \5153 , \5162 );
or \U$4928 ( \5215 , \5212 , \5213 , \5214 );
and \U$4929 ( \5216 , \5119 , \5133 );
and \U$4930 ( \5217 , \5133 , \5148 );
and \U$4931 ( \5218 , \5119 , \5148 );
or \U$4932 ( \5219 , \5216 , \5217 , \5218 );
xor \U$4933 ( \5220 , \5215 , \5219 );
and \U$4934 ( \5221 , \914 , \830 );
and \U$4935 ( \5222 , \871 , \828 );
nor \U$4936 ( \5223 , \5221 , \5222 );
xnor \U$4937 ( \5224 , \5223 , \837 );
and \U$4938 ( \5225 , \940 , \856 );
and \U$4939 ( \5226 , \896 , \854 );
nor \U$4940 ( \5227 , \5225 , \5226 );
xnor \U$4941 ( \5228 , \5227 , \863 );
xor \U$4942 ( \5229 , \5224 , \5228 );
and \U$4943 ( \5230 , \968 , \887 );
and \U$4944 ( \5231 , \922 , \885 );
nor \U$4945 ( \5232 , \5230 , \5231 );
xnor \U$4946 ( \5233 , \5232 , \894 );
xor \U$4947 ( \5234 , \5229 , \5233 );
and \U$4948 ( \5235 , \832 , \750 );
and \U$4949 ( \5236 , \789 , \748 );
nor \U$4950 ( \5237 , \5235 , \5236 );
xnor \U$4951 ( \5238 , \5237 , \757 );
and \U$4952 ( \5239 , \858 , \776 );
and \U$4953 ( \5240 , \814 , \774 );
nor \U$4954 ( \5241 , \5239 , \5240 );
xnor \U$4955 ( \5242 , \5241 , \783 );
xor \U$4956 ( \5243 , \5238 , \5242 );
and \U$4957 ( \5244 , \889 , \805 );
and \U$4958 ( \5245 , \840 , \803 );
nor \U$4959 ( \5246 , \5244 , \5245 );
xnor \U$4960 ( \5247 , \5246 , \812 );
xor \U$4961 ( \5248 , \5243 , \5247 );
xor \U$4962 ( \5249 , \5234 , \5248 );
and \U$4963 ( \5250 , \752 , \674 );
and \U$4964 ( \5251 , \709 , \671 );
nor \U$4965 ( \5252 , \5250 , \5251 );
xnor \U$4966 ( \5253 , \5252 , \635 );
and \U$4967 ( \5254 , \778 , \697 );
and \U$4968 ( \5255 , \734 , \695 );
nor \U$4969 ( \5256 , \5254 , \5255 );
xnor \U$4970 ( \5257 , \5256 , \704 );
xor \U$4971 ( \5258 , \5253 , \5257 );
and \U$4972 ( \5259 , \807 , \725 );
and \U$4973 ( \5260 , \760 , \723 );
nor \U$4974 ( \5261 , \5259 , \5260 );
xnor \U$4975 ( \5262 , \5261 , \732 );
xor \U$4976 ( \5263 , \5258 , \5262 );
xor \U$4977 ( \5264 , \5249 , \5263 );
xor \U$4978 ( \5265 , \5220 , \5264 );
xor \U$4979 ( \5266 , \5211 , \5265 );
xor \U$4980 ( \5267 , \5197 , \5266 );
and \U$4981 ( \5268 , \5169 , \5173 );
and \U$4982 ( \5269 , \5173 , \5184 );
and \U$4983 ( \5270 , \5169 , \5184 );
or \U$4984 ( \5271 , \5268 , \5269 , \5270 );
and \U$4985 ( \5272 , \5149 , \5163 );
xor \U$4986 ( \5273 , \5271 , \5272 );
and \U$4987 ( \5274 , \5111 , \5115 );
and \U$4988 ( \5275 , \5115 , \5118 );
and \U$4989 ( \5276 , \5111 , \5118 );
or \U$4990 ( \5277 , \5274 , \5275 , \5276 );
and \U$4991 ( \5278 , \987 , \912 );
and \U$4992 ( \5279 , \950 , \910 );
nor \U$4993 ( \5280 , \5278 , \5279 );
xnor \U$4994 ( \5281 , \5280 , \919 );
xor \U$4995 ( \5282 , \5277 , \5281 );
and \U$4996 ( \5283 , \995 , \938 );
and \U$4997 ( \5284 , \975 , \936 );
nor \U$4998 ( \5285 , \5283 , \5284 );
xnor \U$4999 ( \5286 , \5285 , \945 );
xor \U$5000 ( \5287 , \5282 , \5286 );
xor \U$5001 ( \5288 , \5273 , \5287 );
xor \U$5002 ( \5289 , \5267 , \5288 );
and \U$5003 ( \5290 , \5101 , \5102 );
and \U$5004 ( \5291 , \5102 , \5186 );
and \U$5005 ( \5292 , \5101 , \5186 );
or \U$5006 ( \5293 , \5290 , \5291 , \5292 );
nor \U$5007 ( \5294 , \5289 , \5293 );
and \U$5008 ( \5295 , \5271 , \5272 );
and \U$5009 ( \5296 , \5272 , \5287 );
and \U$5010 ( \5297 , \5271 , \5287 );
or \U$5011 ( \5298 , \5295 , \5296 , \5297 );
and \U$5012 ( \5299 , \5211 , \5265 );
xor \U$5013 ( \5300 , \5298 , \5299 );
and \U$5014 ( \5301 , \5215 , \5219 );
and \U$5015 ( \5302 , \5219 , \5264 );
and \U$5016 ( \5303 , \5215 , \5264 );
or \U$5017 ( \5304 , \5301 , \5302 , \5303 );
and \U$5018 ( \5305 , \760 , \725 );
and \U$5019 ( \5306 , \778 , \723 );
nor \U$5020 ( \5307 , \5305 , \5306 );
xnor \U$5021 ( \5308 , \5307 , \732 );
and \U$5022 ( \5309 , \789 , \750 );
and \U$5023 ( \5310 , \807 , \748 );
nor \U$5024 ( \5311 , \5309 , \5310 );
xnor \U$5025 ( \5312 , \5311 , \757 );
xor \U$5026 ( \5313 , \5308 , \5312 );
and \U$5027 ( \5314 , \814 , \776 );
and \U$5028 ( \5315 , \832 , \774 );
nor \U$5029 ( \5316 , \5314 , \5315 );
xnor \U$5030 ( \5317 , \5316 , \783 );
xor \U$5031 ( \5318 , \5313 , \5317 );
and \U$5032 ( \5319 , \709 , \674 );
and \U$5033 ( \5320 , \727 , \671 );
nor \U$5034 ( \5321 , \5319 , \5320 );
xnor \U$5035 ( \5322 , \5321 , \635 );
xor \U$5036 ( \5323 , \973 , \5322 );
and \U$5037 ( \5324 , \734 , \697 );
and \U$5038 ( \5325 , \752 , \695 );
nor \U$5039 ( \5326 , \5324 , \5325 );
xnor \U$5040 ( \5327 , \5326 , \704 );
xor \U$5041 ( \5328 , \5323 , \5327 );
xor \U$5042 ( \5329 , \5318 , \5328 );
nand \U$5043 ( \5330 , \995 , \964 );
xnor \U$5044 ( \5331 , \5330 , \973 );
and \U$5045 ( \5332 , \922 , \887 );
and \U$5046 ( \5333 , \940 , \885 );
nor \U$5047 ( \5334 , \5332 , \5333 );
xnor \U$5048 ( \5335 , \5334 , \894 );
and \U$5049 ( \5336 , \950 , \912 );
and \U$5050 ( \5337 , \968 , \910 );
nor \U$5051 ( \5338 , \5336 , \5337 );
xnor \U$5052 ( \5339 , \5338 , \919 );
xor \U$5053 ( \5340 , \5335 , \5339 );
and \U$5054 ( \5341 , \975 , \938 );
and \U$5055 ( \5342 , \987 , \936 );
nor \U$5056 ( \5343 , \5341 , \5342 );
xnor \U$5057 ( \5344 , \5343 , \945 );
xor \U$5058 ( \5345 , \5340 , \5344 );
xor \U$5059 ( \5346 , \5331 , \5345 );
and \U$5060 ( \5347 , \840 , \805 );
and \U$5061 ( \5348 , \858 , \803 );
nor \U$5062 ( \5349 , \5347 , \5348 );
xnor \U$5063 ( \5350 , \5349 , \812 );
and \U$5064 ( \5351 , \871 , \830 );
and \U$5065 ( \5352 , \889 , \828 );
nor \U$5066 ( \5353 , \5351 , \5352 );
xnor \U$5067 ( \5354 , \5353 , \837 );
xor \U$5068 ( \5355 , \5350 , \5354 );
and \U$5069 ( \5356 , \896 , \856 );
and \U$5070 ( \5357 , \914 , \854 );
nor \U$5071 ( \5358 , \5356 , \5357 );
xnor \U$5072 ( \5359 , \5358 , \863 );
xor \U$5073 ( \5360 , \5355 , \5359 );
xor \U$5074 ( \5361 , \5346 , \5360 );
xor \U$5075 ( \5362 , \5329 , \5361 );
and \U$5076 ( \5363 , \5253 , \5257 );
and \U$5077 ( \5364 , \5257 , \5262 );
and \U$5078 ( \5365 , \5253 , \5262 );
or \U$5079 ( \5366 , \5363 , \5364 , \5365 );
and \U$5080 ( \5367 , \5238 , \5242 );
and \U$5081 ( \5368 , \5242 , \5247 );
and \U$5082 ( \5369 , \5238 , \5247 );
or \U$5083 ( \5370 , \5367 , \5368 , \5369 );
xor \U$5084 ( \5371 , \5366 , \5370 );
and \U$5085 ( \5372 , \5224 , \5228 );
and \U$5086 ( \5373 , \5228 , \5233 );
and \U$5087 ( \5374 , \5224 , \5233 );
or \U$5088 ( \5375 , \5372 , \5373 , \5374 );
xor \U$5089 ( \5376 , \5371 , \5375 );
xor \U$5090 ( \5377 , \5362 , \5376 );
xor \U$5091 ( \5378 , \5304 , \5377 );
and \U$5092 ( \5379 , \5201 , \5205 );
and \U$5093 ( \5380 , \5205 , \5210 );
and \U$5094 ( \5381 , \5201 , \5210 );
or \U$5095 ( \5382 , \5379 , \5380 , \5381 );
and \U$5096 ( \5383 , \5277 , \5281 );
and \U$5097 ( \5384 , \5281 , \5286 );
and \U$5098 ( \5385 , \5277 , \5286 );
or \U$5099 ( \5386 , \5383 , \5384 , \5385 );
xor \U$5100 ( \5387 , \5382 , \5386 );
and \U$5101 ( \5388 , \5234 , \5248 );
and \U$5102 ( \5389 , \5248 , \5263 );
and \U$5103 ( \5390 , \5234 , \5263 );
or \U$5104 ( \5391 , \5388 , \5389 , \5390 );
xor \U$5105 ( \5392 , \5387 , \5391 );
xor \U$5106 ( \5393 , \5378 , \5392 );
xor \U$5107 ( \5394 , \5300 , \5393 );
and \U$5108 ( \5395 , \5197 , \5266 );
and \U$5109 ( \5396 , \5266 , \5288 );
and \U$5110 ( \5397 , \5197 , \5288 );
or \U$5111 ( \5398 , \5395 , \5396 , \5397 );
nor \U$5112 ( \5399 , \5394 , \5398 );
nor \U$5113 ( \5400 , \5294 , \5399 );
nand \U$5114 ( \5401 , \5193 , \5400 );
nor \U$5115 ( \5402 , \5006 , \5401 );
and \U$5116 ( \5403 , \5304 , \5377 );
and \U$5117 ( \5404 , \5377 , \5392 );
and \U$5118 ( \5405 , \5304 , \5392 );
or \U$5119 ( \5406 , \5403 , \5404 , \5405 );
and \U$5120 ( \5407 , \5366 , \5370 );
and \U$5121 ( \5408 , \5370 , \5375 );
and \U$5122 ( \5409 , \5366 , \5375 );
or \U$5123 ( \5410 , \5407 , \5408 , \5409 );
and \U$5124 ( \5411 , \5331 , \5345 );
and \U$5125 ( \5412 , \5345 , \5360 );
and \U$5126 ( \5413 , \5331 , \5360 );
or \U$5127 ( \5414 , \5411 , \5412 , \5413 );
xor \U$5128 ( \5415 , \5410 , \5414 );
and \U$5129 ( \5416 , \5318 , \5328 );
xor \U$5130 ( \5417 , \5415 , \5416 );
xor \U$5131 ( \5418 , \5406 , \5417 );
and \U$5132 ( \5419 , \5382 , \5386 );
and \U$5133 ( \5420 , \5386 , \5391 );
and \U$5134 ( \5421 , \5382 , \5391 );
or \U$5135 ( \5422 , \5419 , \5420 , \5421 );
and \U$5136 ( \5423 , \5329 , \5361 );
and \U$5137 ( \5424 , \5361 , \5376 );
and \U$5138 ( \5425 , \5329 , \5376 );
or \U$5139 ( \5426 , \5423 , \5424 , \5425 );
xor \U$5140 ( \5427 , \5422 , \5426 );
and \U$5141 ( \5428 , \807 , \750 );
and \U$5142 ( \5429 , \760 , \748 );
nor \U$5143 ( \5430 , \5428 , \5429 );
xnor \U$5144 ( \5431 , \5430 , \757 );
and \U$5145 ( \5432 , \832 , \776 );
and \U$5146 ( \5433 , \789 , \774 );
nor \U$5147 ( \5434 , \5432 , \5433 );
xnor \U$5148 ( \5435 , \5434 , \783 );
xor \U$5149 ( \5436 , \5431 , \5435 );
and \U$5150 ( \5437 , \858 , \805 );
and \U$5151 ( \5438 , \814 , \803 );
nor \U$5152 ( \5439 , \5437 , \5438 );
xnor \U$5153 ( \5440 , \5439 , \812 );
xor \U$5154 ( \5441 , \5436 , \5440 );
and \U$5155 ( \5442 , \727 , \674 );
and \U$5156 ( \5443 , \681 , \671 );
nor \U$5157 ( \5444 , \5442 , \5443 );
xnor \U$5158 ( \5445 , \5444 , \635 );
and \U$5159 ( \5446 , \752 , \697 );
and \U$5160 ( \5447 , \709 , \695 );
nor \U$5161 ( \5448 , \5446 , \5447 );
xnor \U$5162 ( \5449 , \5448 , \704 );
xor \U$5163 ( \5450 , \5445 , \5449 );
and \U$5164 ( \5451 , \778 , \725 );
and \U$5165 ( \5452 , \734 , \723 );
nor \U$5166 ( \5453 , \5451 , \5452 );
xnor \U$5167 ( \5454 , \5453 , \732 );
xor \U$5168 ( \5455 , \5450 , \5454 );
xor \U$5169 ( \5456 , \5441 , \5455 );
and \U$5170 ( \5457 , \5335 , \5339 );
and \U$5171 ( \5458 , \5339 , \5344 );
and \U$5172 ( \5459 , \5335 , \5344 );
or \U$5173 ( \5460 , \5457 , \5458 , \5459 );
and \U$5174 ( \5461 , \968 , \912 );
and \U$5175 ( \5462 , \922 , \910 );
nor \U$5176 ( \5463 , \5461 , \5462 );
xnor \U$5177 ( \5464 , \5463 , \919 );
and \U$5178 ( \5465 , \987 , \938 );
and \U$5179 ( \5466 , \950 , \936 );
nor \U$5180 ( \5467 , \5465 , \5466 );
xnor \U$5181 ( \5468 , \5467 , \945 );
xor \U$5182 ( \5469 , \5464 , \5468 );
and \U$5183 ( \5470 , \995 , \966 );
and \U$5184 ( \5471 , \975 , \964 );
nor \U$5185 ( \5472 , \5470 , \5471 );
xnor \U$5186 ( \5473 , \5472 , \973 );
xor \U$5187 ( \5474 , \5469 , \5473 );
xor \U$5188 ( \5475 , \5460 , \5474 );
and \U$5189 ( \5476 , \889 , \830 );
and \U$5190 ( \5477 , \840 , \828 );
nor \U$5191 ( \5478 , \5476 , \5477 );
xnor \U$5192 ( \5479 , \5478 , \837 );
and \U$5193 ( \5480 , \914 , \856 );
and \U$5194 ( \5481 , \871 , \854 );
nor \U$5195 ( \5482 , \5480 , \5481 );
xnor \U$5196 ( \5483 , \5482 , \863 );
xor \U$5197 ( \5484 , \5479 , \5483 );
and \U$5198 ( \5485 , \940 , \887 );
and \U$5199 ( \5486 , \896 , \885 );
nor \U$5200 ( \5487 , \5485 , \5486 );
xnor \U$5201 ( \5488 , \5487 , \894 );
xor \U$5202 ( \5489 , \5484 , \5488 );
xor \U$5203 ( \5490 , \5475 , \5489 );
xor \U$5204 ( \5491 , \5456 , \5490 );
and \U$5205 ( \5492 , \973 , \5322 );
and \U$5206 ( \5493 , \5322 , \5327 );
and \U$5207 ( \5494 , \973 , \5327 );
or \U$5208 ( \5495 , \5492 , \5493 , \5494 );
and \U$5209 ( \5496 , \5308 , \5312 );
and \U$5210 ( \5497 , \5312 , \5317 );
and \U$5211 ( \5498 , \5308 , \5317 );
or \U$5212 ( \5499 , \5496 , \5497 , \5498 );
xor \U$5213 ( \5500 , \5495 , \5499 );
and \U$5214 ( \5501 , \5350 , \5354 );
and \U$5215 ( \5502 , \5354 , \5359 );
and \U$5216 ( \5503 , \5350 , \5359 );
or \U$5217 ( \5504 , \5501 , \5502 , \5503 );
xor \U$5218 ( \5505 , \5500 , \5504 );
xor \U$5219 ( \5506 , \5491 , \5505 );
xor \U$5220 ( \5507 , \5427 , \5506 );
xor \U$5221 ( \5508 , \5418 , \5507 );
and \U$5222 ( \5509 , \5298 , \5299 );
and \U$5223 ( \5510 , \5299 , \5393 );
and \U$5224 ( \5511 , \5298 , \5393 );
or \U$5225 ( \5512 , \5509 , \5510 , \5511 );
nor \U$5226 ( \5513 , \5508 , \5512 );
and \U$5227 ( \5514 , \5422 , \5426 );
and \U$5228 ( \5515 , \5426 , \5506 );
and \U$5229 ( \5516 , \5422 , \5506 );
or \U$5230 ( \5517 , \5514 , \5515 , \5516 );
and \U$5231 ( \5518 , \5495 , \5499 );
and \U$5232 ( \5519 , \5499 , \5504 );
and \U$5233 ( \5520 , \5495 , \5504 );
or \U$5234 ( \5521 , \5518 , \5519 , \5520 );
and \U$5235 ( \5522 , \5460 , \5474 );
and \U$5236 ( \5523 , \5474 , \5489 );
and \U$5237 ( \5524 , \5460 , \5489 );
or \U$5238 ( \5525 , \5522 , \5523 , \5524 );
xor \U$5239 ( \5526 , \5521 , \5525 );
and \U$5240 ( \5527 , \5441 , \5455 );
xor \U$5241 ( \5528 , \5526 , \5527 );
xor \U$5242 ( \5529 , \5517 , \5528 );
and \U$5243 ( \5530 , \5410 , \5414 );
and \U$5244 ( \5531 , \5414 , \5416 );
and \U$5245 ( \5532 , \5410 , \5416 );
or \U$5246 ( \5533 , \5530 , \5531 , \5532 );
and \U$5247 ( \5534 , \5456 , \5490 );
and \U$5248 ( \5535 , \5490 , \5505 );
and \U$5249 ( \5536 , \5456 , \5505 );
or \U$5250 ( \5537 , \5534 , \5535 , \5536 );
xor \U$5251 ( \5538 , \5533 , \5537 );
and \U$5252 ( \5539 , \814 , \805 );
and \U$5253 ( \5540 , \832 , \803 );
nor \U$5254 ( \5541 , \5539 , \5540 );
xnor \U$5255 ( \5542 , \5541 , \812 );
and \U$5256 ( \5543 , \840 , \830 );
and \U$5257 ( \5544 , \858 , \828 );
nor \U$5258 ( \5545 , \5543 , \5544 );
xnor \U$5259 ( \5546 , \5545 , \837 );
xor \U$5260 ( \5547 , \5542 , \5546 );
and \U$5261 ( \5548 , \871 , \856 );
and \U$5262 ( \5549 , \889 , \854 );
nor \U$5263 ( \5550 , \5548 , \5549 );
xnor \U$5264 ( \5551 , \5550 , \863 );
xor \U$5265 ( \5552 , \5547 , \5551 );
and \U$5266 ( \5553 , \734 , \725 );
and \U$5267 ( \5554 , \752 , \723 );
nor \U$5268 ( \5555 , \5553 , \5554 );
xnor \U$5269 ( \5556 , \5555 , \732 );
and \U$5270 ( \5557 , \760 , \750 );
and \U$5271 ( \5558 , \778 , \748 );
nor \U$5272 ( \5559 , \5557 , \5558 );
xnor \U$5273 ( \5560 , \5559 , \757 );
xor \U$5274 ( \5561 , \5556 , \5560 );
and \U$5275 ( \5562 , \789 , \776 );
and \U$5276 ( \5563 , \807 , \774 );
nor \U$5277 ( \5564 , \5562 , \5563 );
xnor \U$5278 ( \5565 , \5564 , \783 );
xor \U$5279 ( \5566 , \5561 , \5565 );
xor \U$5280 ( \5567 , \5552 , \5566 );
and \U$5281 ( \5568 , \681 , \674 );
and \U$5282 ( \5569 , \699 , \671 );
nor \U$5283 ( \5570 , \5568 , \5569 );
xnor \U$5284 ( \5571 , \5570 , \635 );
xor \U$5285 ( \5572 , \992 , \5571 );
and \U$5286 ( \5573 , \709 , \697 );
and \U$5287 ( \5574 , \727 , \695 );
nor \U$5288 ( \5575 , \5573 , \5574 );
xnor \U$5289 ( \5576 , \5575 , \704 );
xor \U$5290 ( \5577 , \5572 , \5576 );
xor \U$5291 ( \5578 , \5567 , \5577 );
and \U$5292 ( \5579 , \5464 , \5468 );
and \U$5293 ( \5580 , \5468 , \5473 );
and \U$5294 ( \5581 , \5464 , \5473 );
or \U$5295 ( \5582 , \5579 , \5580 , \5581 );
and \U$5296 ( \5583 , \975 , \966 );
and \U$5297 ( \5584 , \987 , \964 );
nor \U$5298 ( \5585 , \5583 , \5584 );
xnor \U$5299 ( \5586 , \5585 , \973 );
nand \U$5300 ( \5587 , \995 , \983 );
xnor \U$5301 ( \5588 , \5587 , \992 );
xor \U$5302 ( \5589 , \5586 , \5588 );
xor \U$5303 ( \5590 , \5582 , \5589 );
and \U$5304 ( \5591 , \896 , \887 );
and \U$5305 ( \5592 , \914 , \885 );
nor \U$5306 ( \5593 , \5591 , \5592 );
xnor \U$5307 ( \5594 , \5593 , \894 );
and \U$5308 ( \5595 , \922 , \912 );
and \U$5309 ( \5596 , \940 , \910 );
nor \U$5310 ( \5597 , \5595 , \5596 );
xnor \U$5311 ( \5598 , \5597 , \919 );
xor \U$5312 ( \5599 , \5594 , \5598 );
and \U$5313 ( \5600 , \950 , \938 );
and \U$5314 ( \5601 , \968 , \936 );
nor \U$5315 ( \5602 , \5600 , \5601 );
xnor \U$5316 ( \5603 , \5602 , \945 );
xor \U$5317 ( \5604 , \5599 , \5603 );
xor \U$5318 ( \5605 , \5590 , \5604 );
xor \U$5319 ( \5606 , \5578 , \5605 );
and \U$5320 ( \5607 , \5445 , \5449 );
and \U$5321 ( \5608 , \5449 , \5454 );
and \U$5322 ( \5609 , \5445 , \5454 );
or \U$5323 ( \5610 , \5607 , \5608 , \5609 );
and \U$5324 ( \5611 , \5431 , \5435 );
and \U$5325 ( \5612 , \5435 , \5440 );
and \U$5326 ( \5613 , \5431 , \5440 );
or \U$5327 ( \5614 , \5611 , \5612 , \5613 );
xor \U$5328 ( \5615 , \5610 , \5614 );
and \U$5329 ( \5616 , \5479 , \5483 );
and \U$5330 ( \5617 , \5483 , \5488 );
and \U$5331 ( \5618 , \5479 , \5488 );
or \U$5332 ( \5619 , \5616 , \5617 , \5618 );
xor \U$5333 ( \5620 , \5615 , \5619 );
xor \U$5334 ( \5621 , \5606 , \5620 );
xor \U$5335 ( \5622 , \5538 , \5621 );
xor \U$5336 ( \5623 , \5529 , \5622 );
and \U$5337 ( \5624 , \5406 , \5417 );
and \U$5338 ( \5625 , \5417 , \5507 );
and \U$5339 ( \5626 , \5406 , \5507 );
or \U$5340 ( \5627 , \5624 , \5625 , \5626 );
nor \U$5341 ( \5628 , \5623 , \5627 );
nor \U$5342 ( \5629 , \5513 , \5628 );
and \U$5343 ( \5630 , \5533 , \5537 );
and \U$5344 ( \5631 , \5537 , \5621 );
and \U$5345 ( \5632 , \5533 , \5621 );
or \U$5346 ( \5633 , \5630 , \5631 , \5632 );
xor \U$5347 ( \5634 , \1567 , \1571 );
xor \U$5348 ( \5635 , \5634 , \1576 );
xor \U$5349 ( \5636 , \1619 , \1623 );
xor \U$5350 ( \5637 , \5636 , \1628 );
xor \U$5351 ( \5638 , \1600 , \1604 );
xor \U$5352 ( \5639 , \5638 , \1609 );
xor \U$5353 ( \5640 , \5637 , \5639 );
xor \U$5354 ( \5641 , \1583 , \1587 );
xor \U$5355 ( \5642 , \5641 , \1592 );
xor \U$5356 ( \5643 , \5640 , \5642 );
xor \U$5357 ( \5644 , \5635 , \5643 );
and \U$5358 ( \5645 , \5594 , \5598 );
and \U$5359 ( \5646 , \5598 , \5603 );
and \U$5360 ( \5647 , \5594 , \5603 );
or \U$5361 ( \5648 , \5645 , \5646 , \5647 );
and \U$5362 ( \5649 , \5586 , \5588 );
xor \U$5363 ( \5650 , \5648 , \5649 );
and \U$5364 ( \5651 , \995 , \985 );
and \U$5365 ( \5652 , \975 , \983 );
nor \U$5366 ( \5653 , \5651 , \5652 );
xnor \U$5367 ( \5654 , \5653 , \992 );
xor \U$5368 ( \5655 , \5650 , \5654 );
xor \U$5369 ( \5656 , \5644 , \5655 );
and \U$5370 ( \5657 , \5610 , \5614 );
and \U$5371 ( \5658 , \5614 , \5619 );
and \U$5372 ( \5659 , \5610 , \5619 );
or \U$5373 ( \5660 , \5657 , \5658 , \5659 );
and \U$5374 ( \5661 , \5582 , \5589 );
and \U$5375 ( \5662 , \5589 , \5604 );
and \U$5376 ( \5663 , \5582 , \5604 );
or \U$5377 ( \5664 , \5661 , \5662 , \5663 );
xor \U$5378 ( \5665 , \5660 , \5664 );
and \U$5379 ( \5666 , \5552 , \5566 );
and \U$5380 ( \5667 , \5566 , \5577 );
and \U$5381 ( \5668 , \5552 , \5577 );
or \U$5382 ( \5669 , \5666 , \5667 , \5668 );
xor \U$5383 ( \5670 , \5665 , \5669 );
xor \U$5384 ( \5671 , \5656 , \5670 );
xor \U$5385 ( \5672 , \5633 , \5671 );
and \U$5386 ( \5673 , \5521 , \5525 );
and \U$5387 ( \5674 , \5525 , \5527 );
and \U$5388 ( \5675 , \5521 , \5527 );
or \U$5389 ( \5676 , \5673 , \5674 , \5675 );
and \U$5390 ( \5677 , \5578 , \5605 );
and \U$5391 ( \5678 , \5605 , \5620 );
and \U$5392 ( \5679 , \5578 , \5620 );
or \U$5393 ( \5680 , \5677 , \5678 , \5679 );
xor \U$5394 ( \5681 , \5676 , \5680 );
and \U$5395 ( \5682 , \992 , \5571 );
and \U$5396 ( \5683 , \5571 , \5576 );
and \U$5397 ( \5684 , \992 , \5576 );
or \U$5398 ( \5685 , \5682 , \5683 , \5684 );
and \U$5399 ( \5686 , \5556 , \5560 );
and \U$5400 ( \5687 , \5560 , \5565 );
and \U$5401 ( \5688 , \5556 , \5565 );
or \U$5402 ( \5689 , \5686 , \5687 , \5688 );
xor \U$5403 ( \5690 , \5685 , \5689 );
and \U$5404 ( \5691 , \5542 , \5546 );
and \U$5405 ( \5692 , \5546 , \5551 );
and \U$5406 ( \5693 , \5542 , \5551 );
or \U$5407 ( \5694 , \5691 , \5692 , \5693 );
xor \U$5408 ( \5695 , \5690 , \5694 );
xor \U$5409 ( \5696 , \5681 , \5695 );
xor \U$5410 ( \5697 , \5672 , \5696 );
and \U$5411 ( \5698 , \5517 , \5528 );
and \U$5412 ( \5699 , \5528 , \5622 );
and \U$5413 ( \5700 , \5517 , \5622 );
or \U$5414 ( \5701 , \5698 , \5699 , \5700 );
nor \U$5415 ( \5702 , \5697 , \5701 );
and \U$5416 ( \5703 , \5660 , \5664 );
and \U$5417 ( \5704 , \5664 , \5669 );
and \U$5418 ( \5705 , \5660 , \5669 );
or \U$5419 ( \5706 , \5703 , \5704 , \5705 );
and \U$5420 ( \5707 , \5635 , \5643 );
and \U$5421 ( \5708 , \5643 , \5655 );
and \U$5422 ( \5709 , \5635 , \5655 );
or \U$5423 ( \5710 , \5707 , \5708 , \5709 );
xor \U$5424 ( \5711 , \5706 , \5710 );
xor \U$5425 ( \5712 , \1642 , \1644 );
xor \U$5426 ( \5713 , \5712 , \1647 );
xor \U$5427 ( \5714 , \1631 , \1633 );
xor \U$5428 ( \5715 , \5714 , \1636 );
xor \U$5429 ( \5716 , \5713 , \5715 );
xor \U$5430 ( \5717 , \1579 , \1595 );
xor \U$5431 ( \5718 , \5717 , \1612 );
xor \U$5432 ( \5719 , \5716 , \5718 );
xor \U$5433 ( \5720 , \5711 , \5719 );
and \U$5434 ( \5721 , \5676 , \5680 );
and \U$5435 ( \5722 , \5680 , \5695 );
and \U$5436 ( \5723 , \5676 , \5695 );
or \U$5437 ( \5724 , \5721 , \5722 , \5723 );
and \U$5438 ( \5725 , \5656 , \5670 );
xor \U$5439 ( \5726 , \5724 , \5725 );
and \U$5440 ( \5727 , \5685 , \5689 );
and \U$5441 ( \5728 , \5689 , \5694 );
and \U$5442 ( \5729 , \5685 , \5694 );
or \U$5443 ( \5730 , \5727 , \5728 , \5729 );
and \U$5444 ( \5731 , \5648 , \5649 );
and \U$5445 ( \5732 , \5649 , \5654 );
and \U$5446 ( \5733 , \5648 , \5654 );
or \U$5447 ( \5734 , \5731 , \5732 , \5733 );
xor \U$5448 ( \5735 , \5730 , \5734 );
and \U$5449 ( \5736 , \5637 , \5639 );
and \U$5450 ( \5737 , \5639 , \5642 );
and \U$5451 ( \5738 , \5637 , \5642 );
or \U$5452 ( \5739 , \5736 , \5737 , \5738 );
xor \U$5453 ( \5740 , \5735 , \5739 );
xor \U$5454 ( \5741 , \5726 , \5740 );
xor \U$5455 ( \5742 , \5720 , \5741 );
and \U$5456 ( \5743 , \5633 , \5671 );
and \U$5457 ( \5744 , \5671 , \5696 );
and \U$5458 ( \5745 , \5633 , \5696 );
or \U$5459 ( \5746 , \5743 , \5744 , \5745 );
nor \U$5460 ( \5747 , \5742 , \5746 );
nor \U$5461 ( \5748 , \5702 , \5747 );
nand \U$5462 ( \5749 , \5629 , \5748 );
and \U$5463 ( \5750 , \5724 , \5725 );
and \U$5464 ( \5751 , \5725 , \5740 );
and \U$5465 ( \5752 , \5724 , \5740 );
or \U$5466 ( \5753 , \5750 , \5751 , \5752 );
and \U$5467 ( \5754 , \5706 , \5710 );
and \U$5468 ( \5755 , \5710 , \5719 );
and \U$5469 ( \5756 , \5706 , \5719 );
or \U$5470 ( \5757 , \5754 , \5755 , \5756 );
xor \U$5471 ( \5758 , \708 , \787 );
xor \U$5472 ( \5759 , \5758 , \867 );
xor \U$5473 ( \5760 , \1655 , \1657 );
xor \U$5474 ( \5761 , \5760 , \1660 );
xor \U$5475 ( \5762 , \5759 , \5761 );
xor \U$5476 ( \5763 , \1615 , \1639 );
xor \U$5477 ( \5764 , \5763 , \1650 );
xor \U$5478 ( \5765 , \5762 , \5764 );
xor \U$5479 ( \5766 , \5757 , \5765 );
and \U$5480 ( \5767 , \5730 , \5734 );
and \U$5481 ( \5768 , \5734 , \5739 );
and \U$5482 ( \5769 , \5730 , \5739 );
or \U$5483 ( \5770 , \5767 , \5768 , \5769 );
and \U$5484 ( \5771 , \5713 , \5715 );
and \U$5485 ( \5772 , \5715 , \5718 );
and \U$5486 ( \5773 , \5713 , \5718 );
or \U$5487 ( \5774 , \5771 , \5772 , \5773 );
xor \U$5488 ( \5775 , \5770 , \5774 );
xor \U$5489 ( \5776 , \949 , \1001 );
xor \U$5490 ( \5777 , \5776 , \1006 );
xor \U$5491 ( \5778 , \5775 , \5777 );
xor \U$5492 ( \5779 , \5766 , \5778 );
xor \U$5493 ( \5780 , \5753 , \5779 );
and \U$5494 ( \5781 , \5720 , \5741 );
nor \U$5495 ( \5782 , \5780 , \5781 );
and \U$5496 ( \5783 , \5757 , \5765 );
and \U$5497 ( \5784 , \5765 , \5778 );
and \U$5498 ( \5785 , \5757 , \5778 );
or \U$5499 ( \5786 , \5783 , \5784 , \5785 );
xor \U$5500 ( \5787 , \870 , \1009 );
xor \U$5501 ( \5788 , \5787 , \1049 );
xor \U$5502 ( \5789 , \1653 , \1663 );
xor \U$5503 ( \5790 , \5789 , \1666 );
xor \U$5504 ( \5791 , \5788 , \5790 );
xor \U$5505 ( \5792 , \5786 , \5791 );
and \U$5506 ( \5793 , \5770 , \5774 );
and \U$5507 ( \5794 , \5774 , \5777 );
and \U$5508 ( \5795 , \5770 , \5777 );
or \U$5509 ( \5796 , \5793 , \5794 , \5795 );
and \U$5510 ( \5797 , \5759 , \5761 );
and \U$5511 ( \5798 , \5761 , \5764 );
and \U$5512 ( \5799 , \5759 , \5764 );
or \U$5513 ( \5800 , \5797 , \5798 , \5799 );
xor \U$5514 ( \5801 , \5796 , \5800 );
xor \U$5515 ( \5802 , \1064 , \1108 );
xor \U$5516 ( \5803 , \5802 , \1132 );
xor \U$5517 ( \5804 , \5801 , \5803 );
xor \U$5518 ( \5805 , \5792 , \5804 );
and \U$5519 ( \5806 , \5753 , \5779 );
nor \U$5520 ( \5807 , \5805 , \5806 );
nor \U$5521 ( \5808 , \5782 , \5807 );
and \U$5522 ( \5809 , \5796 , \5800 );
and \U$5523 ( \5810 , \5800 , \5803 );
and \U$5524 ( \5811 , \5796 , \5803 );
or \U$5525 ( \5812 , \5809 , \5810 , \5811 );
and \U$5526 ( \5813 , \5788 , \5790 );
xor \U$5527 ( \5814 , \5812 , \5813 );
xor \U$5528 ( \5815 , \1669 , \1670 );
xor \U$5529 ( \5816 , \5815 , \1673 );
xor \U$5530 ( \5817 , \5814 , \5816 );
and \U$5531 ( \5818 , \5786 , \5791 );
and \U$5532 ( \5819 , \5791 , \5804 );
and \U$5533 ( \5820 , \5786 , \5804 );
or \U$5534 ( \5821 , \5818 , \5819 , \5820 );
nor \U$5535 ( \5822 , \5817 , \5821 );
xor \U$5536 ( \5823 , \1676 , \1677 );
xor \U$5537 ( \5824 , \5823 , \1680 );
and \U$5538 ( \5825 , \5812 , \5813 );
and \U$5539 ( \5826 , \5813 , \5816 );
and \U$5540 ( \5827 , \5812 , \5816 );
or \U$5541 ( \5828 , \5825 , \5826 , \5827 );
nor \U$5542 ( \5829 , \5824 , \5828 );
nor \U$5543 ( \5830 , \5822 , \5829 );
nand \U$5544 ( \5831 , \5808 , \5830 );
nor \U$5545 ( \5832 , \5749 , \5831 );
nand \U$5546 ( \5833 , \5402 , \5832 );
and \U$5547 ( \5834 , \940 , \674 );
and \U$5548 ( \5835 , \896 , \671 );
nor \U$5549 ( \5836 , \5834 , \5835 );
xnor \U$5550 ( \5837 , \5836 , \635 );
and \U$5551 ( \5838 , \968 , \697 );
and \U$5552 ( \5839 , \922 , \695 );
nor \U$5553 ( \5840 , \5838 , \5839 );
xnor \U$5554 ( \5841 , \5840 , \704 );
xor \U$5555 ( \5842 , \5837 , \5841 );
and \U$5556 ( \5843 , \987 , \725 );
and \U$5557 ( \5844 , \950 , \723 );
nor \U$5558 ( \5845 , \5843 , \5844 );
xnor \U$5559 ( \5846 , \5845 , \732 );
xor \U$5560 ( \5847 , \5842 , \5846 );
and \U$5561 ( \5848 , \922 , \674 );
and \U$5562 ( \5849 , \940 , \671 );
nor \U$5563 ( \5850 , \5848 , \5849 );
xnor \U$5564 ( \5851 , \5850 , \635 );
and \U$5565 ( \5852 , \757 , \5851 );
and \U$5566 ( \5853 , \950 , \697 );
and \U$5567 ( \5854 , \968 , \695 );
nor \U$5568 ( \5855 , \5853 , \5854 );
xnor \U$5569 ( \5856 , \5855 , \704 );
and \U$5570 ( \5857 , \5851 , \5856 );
and \U$5571 ( \5858 , \757 , \5856 );
or \U$5572 ( \5859 , \5852 , \5857 , \5858 );
and \U$5573 ( \5860 , \975 , \725 );
and \U$5574 ( \5861 , \987 , \723 );
nor \U$5575 ( \5862 , \5860 , \5861 );
xnor \U$5576 ( \5863 , \5862 , \732 );
nand \U$5577 ( \5864 , \995 , \748 );
xnor \U$5578 ( \5865 , \5864 , \757 );
and \U$5579 ( \5866 , \5863 , \5865 );
xor \U$5580 ( \5867 , \5859 , \5866 );
and \U$5581 ( \5868 , \995 , \750 );
and \U$5582 ( \5869 , \975 , \748 );
nor \U$5583 ( \5870 , \5868 , \5869 );
xnor \U$5584 ( \5871 , \5870 , \757 );
xor \U$5585 ( \5872 , \5867 , \5871 );
xor \U$5586 ( \5873 , \5847 , \5872 );
and \U$5587 ( \5874 , \968 , \674 );
and \U$5588 ( \5875 , \922 , \671 );
nor \U$5589 ( \5876 , \5874 , \5875 );
xnor \U$5590 ( \5877 , \5876 , \635 );
and \U$5591 ( \5878 , \987 , \697 );
and \U$5592 ( \5879 , \950 , \695 );
nor \U$5593 ( \5880 , \5878 , \5879 );
xnor \U$5594 ( \5881 , \5880 , \704 );
and \U$5595 ( \5882 , \5877 , \5881 );
and \U$5596 ( \5883 , \995 , \725 );
and \U$5597 ( \5884 , \975 , \723 );
nor \U$5598 ( \5885 , \5883 , \5884 );
xnor \U$5599 ( \5886 , \5885 , \732 );
and \U$5600 ( \5887 , \5881 , \5886 );
and \U$5601 ( \5888 , \5877 , \5886 );
or \U$5602 ( \5889 , \5882 , \5887 , \5888 );
xor \U$5603 ( \5890 , \5863 , \5865 );
and \U$5604 ( \5891 , \5889 , \5890 );
xor \U$5605 ( \5892 , \757 , \5851 );
xor \U$5606 ( \5893 , \5892 , \5856 );
and \U$5607 ( \5894 , \5890 , \5893 );
and \U$5608 ( \5895 , \5889 , \5893 );
or \U$5609 ( \5896 , \5891 , \5894 , \5895 );
nor \U$5610 ( \5897 , \5873 , \5896 );
and \U$5611 ( \5898 , \5859 , \5866 );
and \U$5612 ( \5899 , \5866 , \5871 );
and \U$5613 ( \5900 , \5859 , \5871 );
or \U$5614 ( \5901 , \5898 , \5899 , \5900 );
and \U$5615 ( \5902 , \5837 , \5841 );
and \U$5616 ( \5903 , \5841 , \5846 );
and \U$5617 ( \5904 , \5837 , \5846 );
or \U$5618 ( \5905 , \5902 , \5903 , \5904 );
and \U$5619 ( \5906 , \950 , \725 );
and \U$5620 ( \5907 , \968 , \723 );
nor \U$5621 ( \5908 , \5906 , \5907 );
xnor \U$5622 ( \5909 , \5908 , \732 );
and \U$5623 ( \5910 , \975 , \750 );
and \U$5624 ( \5911 , \987 , \748 );
nor \U$5625 ( \5912 , \5910 , \5911 );
xnor \U$5626 ( \5913 , \5912 , \757 );
xor \U$5627 ( \5914 , \5909 , \5913 );
nand \U$5628 ( \5915 , \995 , \774 );
xnor \U$5629 ( \5916 , \5915 , \783 );
xor \U$5630 ( \5917 , \5914 , \5916 );
xor \U$5631 ( \5918 , \5905 , \5917 );
and \U$5632 ( \5919 , \896 , \674 );
and \U$5633 ( \5920 , \914 , \671 );
nor \U$5634 ( \5921 , \5919 , \5920 );
xnor \U$5635 ( \5922 , \5921 , \635 );
xor \U$5636 ( \5923 , \783 , \5922 );
and \U$5637 ( \5924 , \922 , \697 );
and \U$5638 ( \5925 , \940 , \695 );
nor \U$5639 ( \5926 , \5924 , \5925 );
xnor \U$5640 ( \5927 , \5926 , \704 );
xor \U$5641 ( \5928 , \5923 , \5927 );
xor \U$5642 ( \5929 , \5918 , \5928 );
xor \U$5643 ( \5930 , \5901 , \5929 );
and \U$5644 ( \5931 , \5847 , \5872 );
nor \U$5645 ( \5932 , \5930 , \5931 );
nor \U$5646 ( \5933 , \5897 , \5932 );
and \U$5647 ( \5934 , \5905 , \5917 );
and \U$5648 ( \5935 , \5917 , \5928 );
and \U$5649 ( \5936 , \5905 , \5928 );
or \U$5650 ( \5937 , \5934 , \5935 , \5936 );
and \U$5651 ( \5938 , \995 , \776 );
and \U$5652 ( \5939 , \975 , \774 );
nor \U$5653 ( \5940 , \5938 , \5939 );
xnor \U$5654 ( \5941 , \5940 , \783 );
and \U$5655 ( \5942 , \914 , \674 );
and \U$5656 ( \5943 , \871 , \671 );
nor \U$5657 ( \5944 , \5942 , \5943 );
xnor \U$5658 ( \5945 , \5944 , \635 );
and \U$5659 ( \5946 , \940 , \697 );
and \U$5660 ( \5947 , \896 , \695 );
nor \U$5661 ( \5948 , \5946 , \5947 );
xnor \U$5662 ( \5949 , \5948 , \704 );
xor \U$5663 ( \5950 , \5945 , \5949 );
and \U$5664 ( \5951 , \968 , \725 );
and \U$5665 ( \5952 , \922 , \723 );
nor \U$5666 ( \5953 , \5951 , \5952 );
xnor \U$5667 ( \5954 , \5953 , \732 );
xor \U$5668 ( \5955 , \5950 , \5954 );
xor \U$5669 ( \5956 , \5941 , \5955 );
xor \U$5670 ( \5957 , \5937 , \5956 );
and \U$5671 ( \5958 , \783 , \5922 );
and \U$5672 ( \5959 , \5922 , \5927 );
and \U$5673 ( \5960 , \783 , \5927 );
or \U$5674 ( \5961 , \5958 , \5959 , \5960 );
and \U$5675 ( \5962 , \5909 , \5913 );
and \U$5676 ( \5963 , \5913 , \5916 );
and \U$5677 ( \5964 , \5909 , \5916 );
or \U$5678 ( \5965 , \5962 , \5963 , \5964 );
xor \U$5679 ( \5966 , \5961 , \5965 );
and \U$5680 ( \5967 , \987 , \750 );
and \U$5681 ( \5968 , \950 , \748 );
nor \U$5682 ( \5969 , \5967 , \5968 );
xnor \U$5683 ( \5970 , \5969 , \757 );
xor \U$5684 ( \5971 , \5966 , \5970 );
xor \U$5685 ( \5972 , \5957 , \5971 );
and \U$5686 ( \5973 , \5901 , \5929 );
nor \U$5687 ( \5974 , \5972 , \5973 );
and \U$5688 ( \5975 , \5945 , \5949 );
and \U$5689 ( \5976 , \5949 , \5954 );
and \U$5690 ( \5977 , \5945 , \5954 );
or \U$5691 ( \5978 , \5975 , \5976 , \5977 );
nand \U$5692 ( \5979 , \995 , \803 );
xnor \U$5693 ( \5980 , \5979 , \812 );
xor \U$5694 ( \5981 , \5978 , \5980 );
and \U$5695 ( \5982 , \922 , \725 );
and \U$5696 ( \5983 , \940 , \723 );
nor \U$5697 ( \5984 , \5982 , \5983 );
xnor \U$5698 ( \5985 , \5984 , \732 );
and \U$5699 ( \5986 , \950 , \750 );
and \U$5700 ( \5987 , \968 , \748 );
nor \U$5701 ( \5988 , \5986 , \5987 );
xnor \U$5702 ( \5989 , \5988 , \757 );
xor \U$5703 ( \5990 , \5985 , \5989 );
and \U$5704 ( \5991 , \975 , \776 );
and \U$5705 ( \5992 , \987 , \774 );
nor \U$5706 ( \5993 , \5991 , \5992 );
xnor \U$5707 ( \5994 , \5993 , \783 );
xor \U$5708 ( \5995 , \5990 , \5994 );
xor \U$5709 ( \5996 , \5981 , \5995 );
and \U$5710 ( \5997 , \5961 , \5965 );
and \U$5711 ( \5998 , \5965 , \5970 );
and \U$5712 ( \5999 , \5961 , \5970 );
or \U$5713 ( \6000 , \5997 , \5998 , \5999 );
and \U$5714 ( \6001 , \5941 , \5955 );
xor \U$5715 ( \6002 , \6000 , \6001 );
and \U$5716 ( \6003 , \871 , \674 );
and \U$5717 ( \6004 , \889 , \671 );
nor \U$5718 ( \6005 , \6003 , \6004 );
xnor \U$5719 ( \6006 , \6005 , \635 );
xor \U$5720 ( \6007 , \812 , \6006 );
and \U$5721 ( \6008 , \896 , \697 );
and \U$5722 ( \6009 , \914 , \695 );
nor \U$5723 ( \6010 , \6008 , \6009 );
xnor \U$5724 ( \6011 , \6010 , \704 );
xor \U$5725 ( \6012 , \6007 , \6011 );
xor \U$5726 ( \6013 , \6002 , \6012 );
xor \U$5727 ( \6014 , \5996 , \6013 );
and \U$5728 ( \6015 , \5937 , \5956 );
and \U$5729 ( \6016 , \5956 , \5971 );
and \U$5730 ( \6017 , \5937 , \5971 );
or \U$5731 ( \6018 , \6015 , \6016 , \6017 );
nor \U$5732 ( \6019 , \6014 , \6018 );
nor \U$5733 ( \6020 , \5974 , \6019 );
nand \U$5734 ( \6021 , \5933 , \6020 );
and \U$5735 ( \6022 , \6000 , \6001 );
and \U$5736 ( \6023 , \6001 , \6012 );
and \U$5737 ( \6024 , \6000 , \6012 );
or \U$5738 ( \6025 , \6022 , \6023 , \6024 );
and \U$5739 ( \6026 , \5978 , \5980 );
and \U$5740 ( \6027 , \5980 , \5995 );
and \U$5741 ( \6028 , \5978 , \5995 );
or \U$5742 ( \6029 , \6026 , \6027 , \6028 );
xor \U$5743 ( \6030 , \4698 , \4702 );
xor \U$5744 ( \6031 , \6030 , \4707 );
xor \U$5745 ( \6032 , \6029 , \6031 );
and \U$5746 ( \6033 , \812 , \6006 );
and \U$5747 ( \6034 , \6006 , \6011 );
and \U$5748 ( \6035 , \812 , \6011 );
or \U$5749 ( \6036 , \6033 , \6034 , \6035 );
and \U$5750 ( \6037 , \5985 , \5989 );
and \U$5751 ( \6038 , \5989 , \5994 );
and \U$5752 ( \6039 , \5985 , \5994 );
or \U$5753 ( \6040 , \6037 , \6038 , \6039 );
xor \U$5754 ( \6041 , \6036 , \6040 );
xor \U$5755 ( \6042 , \4714 , \4718 );
xor \U$5756 ( \6043 , \6042 , \4723 );
xor \U$5757 ( \6044 , \6041 , \6043 );
xor \U$5758 ( \6045 , \6032 , \6044 );
xor \U$5759 ( \6046 , \6025 , \6045 );
and \U$5760 ( \6047 , \5996 , \6013 );
nor \U$5761 ( \6048 , \6046 , \6047 );
and \U$5762 ( \6049 , \6029 , \6031 );
and \U$5763 ( \6050 , \6031 , \6044 );
and \U$5764 ( \6051 , \6029 , \6044 );
or \U$5765 ( \6052 , \6049 , \6050 , \6051 );
and \U$5766 ( \6053 , \6036 , \6040 );
and \U$5767 ( \6054 , \6040 , \6043 );
and \U$5768 ( \6055 , \6036 , \6043 );
or \U$5769 ( \6056 , \6053 , \6054 , \6055 );
xor \U$5770 ( \6057 , \4736 , \4738 );
xor \U$5771 ( \6058 , \6057 , \4741 );
xor \U$5772 ( \6059 , \6056 , \6058 );
xor \U$5773 ( \6060 , \4710 , \4726 );
xor \U$5774 ( \6061 , \6060 , \4731 );
xor \U$5775 ( \6062 , \6059 , \6061 );
xor \U$5776 ( \6063 , \6052 , \6062 );
and \U$5777 ( \6064 , \6025 , \6045 );
nor \U$5778 ( \6065 , \6063 , \6064 );
nor \U$5779 ( \6066 , \6048 , \6065 );
and \U$5780 ( \6067 , \6056 , \6058 );
and \U$5781 ( \6068 , \6058 , \6061 );
and \U$5782 ( \6069 , \6056 , \6061 );
or \U$5783 ( \6070 , \6067 , \6068 , \6069 );
xor \U$5784 ( \6071 , \4752 , \4754 );
xor \U$5785 ( \6072 , \6070 , \6071 );
xor \U$5786 ( \6073 , \4734 , \4744 );
xor \U$5787 ( \6074 , \6073 , \4747 );
xor \U$5788 ( \6075 , \6072 , \6074 );
and \U$5789 ( \6076 , \6052 , \6062 );
nor \U$5790 ( \6077 , \6075 , \6076 );
xor \U$5791 ( \6078 , \4750 , \4755 );
xor \U$5792 ( \6079 , \6078 , \4758 );
and \U$5793 ( \6080 , \6070 , \6071 );
and \U$5794 ( \6081 , \6071 , \6074 );
and \U$5795 ( \6082 , \6070 , \6074 );
or \U$5796 ( \6083 , \6080 , \6081 , \6082 );
nor \U$5797 ( \6084 , \6079 , \6083 );
nor \U$5798 ( \6085 , \6077 , \6084 );
nand \U$5799 ( \6086 , \6066 , \6085 );
nor \U$5800 ( \6087 , \6021 , \6086 );
and \U$5801 ( \6088 , \987 , \674 );
and \U$5802 ( \6089 , \950 , \671 );
nor \U$5803 ( \6090 , \6088 , \6089 );
xnor \U$5804 ( \6091 , \6090 , \635 );
and \U$5805 ( \6092 , \995 , \697 );
and \U$5806 ( \6093 , \975 , \695 );
nor \U$5807 ( \6094 , \6092 , \6093 );
xnor \U$5808 ( \6095 , \6094 , \704 );
xor \U$5809 ( \6096 , \6091 , \6095 );
and \U$5810 ( \6097 , \975 , \674 );
and \U$5811 ( \6098 , \987 , \671 );
nor \U$5812 ( \6099 , \6097 , \6098 );
xnor \U$5813 ( \6100 , \6099 , \635 );
and \U$5814 ( \6101 , \6100 , \704 );
nor \U$5815 ( \6102 , \6096 , \6101 );
nand \U$5816 ( \6103 , \995 , \723 );
xnor \U$5817 ( \6104 , \6103 , \732 );
and \U$5818 ( \6105 , \950 , \674 );
and \U$5819 ( \6106 , \968 , \671 );
nor \U$5820 ( \6107 , \6105 , \6106 );
xnor \U$5821 ( \6108 , \6107 , \635 );
xor \U$5822 ( \6109 , \732 , \6108 );
and \U$5823 ( \6110 , \975 , \697 );
and \U$5824 ( \6111 , \987 , \695 );
nor \U$5825 ( \6112 , \6110 , \6111 );
xnor \U$5826 ( \6113 , \6112 , \704 );
xor \U$5827 ( \6114 , \6109 , \6113 );
xor \U$5828 ( \6115 , \6104 , \6114 );
and \U$5829 ( \6116 , \6091 , \6095 );
nor \U$5830 ( \6117 , \6115 , \6116 );
nor \U$5831 ( \6118 , \6102 , \6117 );
and \U$5832 ( \6119 , \732 , \6108 );
and \U$5833 ( \6120 , \6108 , \6113 );
and \U$5834 ( \6121 , \732 , \6113 );
or \U$5835 ( \6122 , \6119 , \6120 , \6121 );
xor \U$5836 ( \6123 , \5877 , \5881 );
xor \U$5837 ( \6124 , \6123 , \5886 );
xor \U$5838 ( \6125 , \6122 , \6124 );
and \U$5839 ( \6126 , \6104 , \6114 );
nor \U$5840 ( \6127 , \6125 , \6126 );
xor \U$5841 ( \6128 , \5889 , \5890 );
xor \U$5842 ( \6129 , \6128 , \5893 );
and \U$5843 ( \6130 , \6122 , \6124 );
nor \U$5844 ( \6131 , \6129 , \6130 );
nor \U$5845 ( \6132 , \6127 , \6131 );
nand \U$5846 ( \6133 , \6118 , \6132 );
xor \U$5847 ( \6134 , \6100 , \704 );
nand \U$5848 ( \6135 , \995 , \695 );
xnor \U$5849 ( \6136 , \6135 , \704 );
nor \U$5850 ( \6137 , \6134 , \6136 );
and \U$5851 ( \6138 , \995 , \674 );
and \U$5852 ( \6139 , \975 , \671 );
nor \U$5853 ( \6140 , \6138 , \6139 );
xnor \U$5854 ( \6141 , \6140 , \635 );
nand \U$5855 ( \6142 , \995 , \671 );
xnor \U$5856 ( \6143 , \6142 , \635 );
and \U$5857 ( \6144 , \6143 , \635 );
nand \U$5858 ( \6145 , \6141 , \6144 );
or \U$5859 ( \6146 , \6137 , \6145 );
nand \U$5860 ( \6147 , \6134 , \6136 );
nand \U$5861 ( \6148 , \6146 , \6147 );
not \U$5862 ( \6149 , \6148 );
or \U$5863 ( \6150 , \6133 , \6149 );
nand \U$5864 ( \6151 , \6096 , \6101 );
or \U$5865 ( \6152 , \6117 , \6151 );
nand \U$5866 ( \6153 , \6115 , \6116 );
nand \U$5867 ( \6154 , \6152 , \6153 );
and \U$5868 ( \6155 , \6132 , \6154 );
nand \U$5869 ( \6156 , \6125 , \6126 );
or \U$5870 ( \6157 , \6131 , \6156 );
nand \U$5871 ( \6158 , \6129 , \6130 );
nand \U$5872 ( \6159 , \6157 , \6158 );
nor \U$5873 ( \6160 , \6155 , \6159 );
nand \U$5874 ( \6161 , \6150 , \6160 );
and \U$5875 ( \6162 , \6087 , \6161 );
nand \U$5876 ( \6163 , \5873 , \5896 );
or \U$5877 ( \6164 , \5932 , \6163 );
nand \U$5878 ( \6165 , \5930 , \5931 );
nand \U$5879 ( \6166 , \6164 , \6165 );
and \U$5880 ( \6167 , \6020 , \6166 );
nand \U$5881 ( \6168 , \5972 , \5973 );
or \U$5882 ( \6169 , \6019 , \6168 );
nand \U$5883 ( \6170 , \6014 , \6018 );
nand \U$5884 ( \6171 , \6169 , \6170 );
nor \U$5885 ( \6172 , \6167 , \6171 );
or \U$5886 ( \6173 , \6086 , \6172 );
nand \U$5887 ( \6174 , \6046 , \6047 );
or \U$5888 ( \6175 , \6065 , \6174 );
nand \U$5889 ( \6176 , \6063 , \6064 );
nand \U$5890 ( \6177 , \6175 , \6176 );
and \U$5891 ( \6178 , \6085 , \6177 );
nand \U$5892 ( \6179 , \6075 , \6076 );
or \U$5893 ( \6180 , \6084 , \6179 );
nand \U$5894 ( \6181 , \6079 , \6083 );
nand \U$5895 ( \6182 , \6180 , \6181 );
nor \U$5896 ( \6183 , \6178 , \6182 );
nand \U$5897 ( \6184 , \6173 , \6183 );
nor \U$5898 ( \6185 , \6162 , \6184 );
or \U$5899 ( \6186 , \5833 , \6185 );
nand \U$5900 ( \6187 , \4694 , \4761 );
or \U$5901 ( \6188 , \4837 , \6187 );
nand \U$5902 ( \6189 , \4832 , \4836 );
nand \U$5903 ( \6190 , \6188 , \6189 );
and \U$5904 ( \6191 , \5005 , \6190 );
nand \U$5905 ( \6192 , \4914 , \4918 );
or \U$5906 ( \6193 , \5004 , \6192 );
nand \U$5907 ( \6194 , \5002 , \5003 );
nand \U$5908 ( \6195 , \6193 , \6194 );
nor \U$5909 ( \6196 , \6191 , \6195 );
or \U$5910 ( \6197 , \5401 , \6196 );
nand \U$5911 ( \6198 , \5095 , \5096 );
or \U$5912 ( \6199 , \5192 , \6198 );
nand \U$5913 ( \6200 , \5187 , \5191 );
nand \U$5914 ( \6201 , \6199 , \6200 );
and \U$5915 ( \6202 , \5400 , \6201 );
nand \U$5916 ( \6203 , \5289 , \5293 );
or \U$5917 ( \6204 , \5399 , \6203 );
nand \U$5918 ( \6205 , \5394 , \5398 );
nand \U$5919 ( \6206 , \6204 , \6205 );
nor \U$5920 ( \6207 , \6202 , \6206 );
nand \U$5921 ( \6208 , \6197 , \6207 );
and \U$5922 ( \6209 , \5832 , \6208 );
nand \U$5923 ( \6210 , \5508 , \5512 );
or \U$5924 ( \6211 , \5628 , \6210 );
nand \U$5925 ( \6212 , \5623 , \5627 );
nand \U$5926 ( \6213 , \6211 , \6212 );
and \U$5927 ( \6214 , \5748 , \6213 );
nand \U$5928 ( \6215 , \5697 , \5701 );
or \U$5929 ( \6216 , \5747 , \6215 );
nand \U$5930 ( \6217 , \5742 , \5746 );
nand \U$5931 ( \6218 , \6216 , \6217 );
nor \U$5932 ( \6219 , \6214 , \6218 );
or \U$5933 ( \6220 , \5831 , \6219 );
nand \U$5934 ( \6221 , \5780 , \5781 );
or \U$5935 ( \6222 , \5807 , \6221 );
nand \U$5936 ( \6223 , \5805 , \5806 );
nand \U$5937 ( \6224 , \6222 , \6223 );
and \U$5938 ( \6225 , \5830 , \6224 );
nand \U$5939 ( \6226 , \5817 , \5821 );
or \U$5940 ( \6227 , \5829 , \6226 );
nand \U$5941 ( \6228 , \5824 , \5828 );
nand \U$5942 ( \6229 , \6227 , \6228 );
nor \U$5943 ( \6230 , \6225 , \6229 );
nand \U$5944 ( \6231 , \6220 , \6230 );
nor \U$5945 ( \6232 , \6209 , \6231 );
nand \U$5946 ( \6233 , \6186 , \6232 );
and \U$5947 ( \6234 , \4521 , \6233 );
nand \U$5948 ( \6235 , \1563 , \1683 );
or \U$5949 ( \6236 , \1837 , \6235 );
nand \U$5950 ( \6237 , \1832 , \1836 );
nand \U$5951 ( \6238 , \6236 , \6237 );
and \U$5952 ( \6239 , \2146 , \6238 );
nand \U$5953 ( \6240 , \1987 , \1991 );
or \U$5954 ( \6241 , \2145 , \6240 );
nand \U$5955 ( \6242 , \2140 , \2144 );
nand \U$5956 ( \6243 , \6241 , \6242 );
nor \U$5957 ( \6244 , \6239 , \6243 );
or \U$5958 ( \6245 , \2725 , \6244 );
nand \U$5959 ( \6246 , \2294 , \2298 );
or \U$5960 ( \6247 , \2446 , \6246 );
nand \U$5961 ( \6248 , \2441 , \2445 );
nand \U$5962 ( \6249 , \6247 , \6248 );
and \U$5963 ( \6250 , \2724 , \6249 );
nand \U$5964 ( \6251 , \2581 , \2585 );
or \U$5965 ( \6252 , \2723 , \6251 );
nand \U$5966 ( \6253 , \2718 , \2722 );
nand \U$5967 ( \6254 , \6252 , \6253 );
nor \U$5968 ( \6255 , \6250 , \6254 );
nand \U$5969 ( \6256 , \6245 , \6255 );
and \U$5970 ( \6257 , \3644 , \6256 );
nand \U$5971 ( \6258 , \2850 , \2854 );
or \U$5972 ( \6259 , \2981 , \6258 );
nand \U$5973 ( \6260 , \2976 , \2980 );
nand \U$5974 ( \6261 , \6259 , \6260 );
and \U$5975 ( \6262 , \3221 , \6261 );
nand \U$5976 ( \6263 , \3099 , \3103 );
or \U$5977 ( \6264 , \3220 , \6263 );
nand \U$5978 ( \6265 , \3218 , \3219 );
nand \U$5979 ( \6266 , \6264 , \6265 );
nor \U$5980 ( \6267 , \6262 , \6266 );
or \U$5981 ( \6268 , \3643 , \6267 );
nand \U$5982 ( \6269 , \3329 , \3333 );
or \U$5983 ( \6270 , \3440 , \6269 );
nand \U$5984 ( \6271 , \3438 , \3439 );
nand \U$5985 ( \6272 , \6270 , \6271 );
and \U$5986 ( \6273 , \3642 , \6272 );
nand \U$5987 ( \6274 , \3540 , \3541 );
or \U$5988 ( \6275 , \3641 , \6274 );
nand \U$5989 ( \6276 , \3639 , \3640 );
nand \U$5990 ( \6277 , \6275 , \6276 );
nor \U$5991 ( \6278 , \6273 , \6277 );
nand \U$5992 ( \6279 , \6268 , \6278 );
nor \U$5993 ( \6280 , \6257 , \6279 );
or \U$5994 ( \6281 , \4520 , \6280 );
nand \U$5995 ( \6282 , \3734 , \3735 );
or \U$5996 ( \6283 , \3825 , \6282 );
nand \U$5997 ( \6284 , \3823 , \3824 );
nand \U$5998 ( \6285 , \6283 , \6284 );
and \U$5999 ( \6286 , \3987 , \6285 );
nand \U$6000 ( \6287 , \3905 , \3906 );
or \U$6001 ( \6288 , \3986 , \6287 );
nand \U$6002 ( \6289 , \3984 , \3985 );
nand \U$6003 ( \6290 , \6288 , \6289 );
nor \U$6004 ( \6291 , \6286 , \6290 );
or \U$6005 ( \6292 , \4251 , \6291 );
nand \U$6006 ( \6293 , \4055 , \4059 );
or \U$6007 ( \6294 , \4125 , \6293 );
nand \U$6008 ( \6295 , \4123 , \4124 );
nand \U$6009 ( \6296 , \6294 , \6295 );
and \U$6010 ( \6297 , \4250 , \6296 );
nand \U$6011 ( \6298 , \4188 , \4189 );
or \U$6012 ( \6299 , \4249 , \6298 );
nand \U$6013 ( \6300 , \4247 , \4248 );
nand \U$6014 ( \6301 , \6299 , \6300 );
nor \U$6015 ( \6302 , \6297 , \6301 );
nand \U$6016 ( \6303 , \6292 , \6302 );
and \U$6017 ( \6304 , \4519 , \6303 );
nand \U$6018 ( \6305 , \4301 , \4302 );
or \U$6019 ( \6306 , \4352 , \6305 );
nand \U$6020 ( \6307 , \4350 , \4351 );
nand \U$6021 ( \6308 , \6306 , \6307 );
and \U$6022 ( \6309 , \4431 , \6308 );
nand \U$6023 ( \6310 , \4390 , \4394 );
or \U$6024 ( \6311 , \4430 , \6310 );
nand \U$6025 ( \6312 , \4428 , \4429 );
nand \U$6026 ( \6313 , \6311 , \6312 );
nor \U$6027 ( \6314 , \6309 , \6313 );
or \U$6028 ( \6315 , \4518 , \6314 );
nand \U$6029 ( \6316 , \4464 , \4465 );
or \U$6030 ( \6317 , \4495 , \6316 );
nand \U$6031 ( \6318 , \4493 , \4494 );
nand \U$6032 ( \6319 , \6317 , \6318 );
and \U$6033 ( \6320 , \4517 , \6319 );
nand \U$6034 ( \6321 , \4505 , \4509 );
or \U$6035 ( \6322 , \4516 , \6321 );
nand \U$6036 ( \6323 , \4511 , \4515 );
nand \U$6037 ( \6324 , \6322 , \6323 );
nor \U$6038 ( \6325 , \6320 , \6324 );
nand \U$6039 ( \6326 , \6315 , \6325 );
nor \U$6040 ( \6327 , \6304 , \6326 );
nand \U$6041 ( \6328 , \6281 , \6327 );
nor \U$6042 ( \6329 , \6234 , \6328 );
not \U$6043 ( \6330 , \6329 );
xnor \U$6044 ( \6331 , \613 , \6330 );
buf g18bf ( \6332_nG18bf , \6331 );
buf \U$6045 ( \6333 , \6332_nG18bf );
not \U$6046 ( \6334 , \4516 );
nand \U$6047 ( \6335 , \6323 , \6334 );
nor \U$6048 ( \6336 , \5829 , \1684 );
nor \U$6049 ( \6337 , \1837 , \1992 );
nand \U$6050 ( \6338 , \6336 , \6337 );
nor \U$6051 ( \6339 , \2145 , \2299 );
nor \U$6052 ( \6340 , \2446 , \2586 );
nand \U$6053 ( \6341 , \6339 , \6340 );
nor \U$6054 ( \6342 , \6338 , \6341 );
nor \U$6055 ( \6343 , \2723 , \2855 );
nor \U$6056 ( \6344 , \2981 , \3104 );
nand \U$6057 ( \6345 , \6343 , \6344 );
nor \U$6058 ( \6346 , \3220 , \3334 );
nor \U$6059 ( \6347 , \3440 , \3542 );
nand \U$6060 ( \6348 , \6346 , \6347 );
nor \U$6061 ( \6349 , \6345 , \6348 );
nand \U$6062 ( \6350 , \6342 , \6349 );
nor \U$6063 ( \6351 , \3641 , \3736 );
nor \U$6064 ( \6352 , \3825 , \3907 );
nand \U$6065 ( \6353 , \6351 , \6352 );
nor \U$6066 ( \6354 , \3986 , \4060 );
nor \U$6067 ( \6355 , \4125 , \4190 );
nand \U$6068 ( \6356 , \6354 , \6355 );
nor \U$6069 ( \6357 , \6353 , \6356 );
nor \U$6070 ( \6358 , \4249 , \4303 );
nor \U$6071 ( \6359 , \4352 , \4395 );
nand \U$6072 ( \6360 , \6358 , \6359 );
nor \U$6073 ( \6361 , \4430 , \4466 );
nor \U$6074 ( \6362 , \4495 , \4510 );
nand \U$6075 ( \6363 , \6361 , \6362 );
nor \U$6076 ( \6364 , \6360 , \6363 );
nand \U$6077 ( \6365 , \6357 , \6364 );
nor \U$6078 ( \6366 , \6350 , \6365 );
nor \U$6079 ( \6367 , \6084 , \4762 );
nor \U$6080 ( \6368 , \4837 , \4919 );
nand \U$6081 ( \6369 , \6367 , \6368 );
nor \U$6082 ( \6370 , \5004 , \5097 );
nor \U$6083 ( \6371 , \5192 , \5294 );
nand \U$6084 ( \6372 , \6370 , \6371 );
nor \U$6085 ( \6373 , \6369 , \6372 );
nor \U$6086 ( \6374 , \5399 , \5513 );
nor \U$6087 ( \6375 , \5628 , \5702 );
nand \U$6088 ( \6376 , \6374 , \6375 );
nor \U$6089 ( \6377 , \5747 , \5782 );
nor \U$6090 ( \6378 , \5807 , \5822 );
nand \U$6091 ( \6379 , \6377 , \6378 );
nor \U$6092 ( \6380 , \6376 , \6379 );
nand \U$6093 ( \6381 , \6373 , \6380 );
nor \U$6094 ( \6382 , \6131 , \5897 );
nor \U$6095 ( \6383 , \5932 , \5974 );
nand \U$6096 ( \6384 , \6382 , \6383 );
nor \U$6097 ( \6385 , \6019 , \6048 );
nor \U$6098 ( \6386 , \6065 , \6077 );
nand \U$6099 ( \6387 , \6385 , \6386 );
nor \U$6100 ( \6388 , \6384 , \6387 );
nor \U$6101 ( \6389 , \6137 , \6102 );
nor \U$6102 ( \6390 , \6117 , \6127 );
nand \U$6103 ( \6391 , \6389 , \6390 );
or \U$6104 ( \6392 , \6391 , \6145 );
or \U$6105 ( \6393 , \6102 , \6147 );
nand \U$6106 ( \6394 , \6393 , \6151 );
and \U$6107 ( \6395 , \6390 , \6394 );
or \U$6108 ( \6396 , \6127 , \6153 );
nand \U$6109 ( \6397 , \6396 , \6156 );
nor \U$6110 ( \6398 , \6395 , \6397 );
nand \U$6111 ( \6399 , \6392 , \6398 );
and \U$6112 ( \6400 , \6388 , \6399 );
or \U$6113 ( \6401 , \5897 , \6158 );
nand \U$6114 ( \6402 , \6401 , \6163 );
and \U$6115 ( \6403 , \6383 , \6402 );
or \U$6116 ( \6404 , \5974 , \6165 );
nand \U$6117 ( \6405 , \6404 , \6168 );
nor \U$6118 ( \6406 , \6403 , \6405 );
or \U$6119 ( \6407 , \6387 , \6406 );
or \U$6120 ( \6408 , \6048 , \6170 );
nand \U$6121 ( \6409 , \6408 , \6174 );
and \U$6122 ( \6410 , \6386 , \6409 );
or \U$6123 ( \6411 , \6077 , \6176 );
nand \U$6124 ( \6412 , \6411 , \6179 );
nor \U$6125 ( \6413 , \6410 , \6412 );
nand \U$6126 ( \6414 , \6407 , \6413 );
nor \U$6127 ( \6415 , \6400 , \6414 );
or \U$6128 ( \6416 , \6381 , \6415 );
or \U$6129 ( \6417 , \4762 , \6181 );
nand \U$6130 ( \6418 , \6417 , \6187 );
and \U$6131 ( \6419 , \6368 , \6418 );
or \U$6132 ( \6420 , \4919 , \6189 );
nand \U$6133 ( \6421 , \6420 , \6192 );
nor \U$6134 ( \6422 , \6419 , \6421 );
or \U$6135 ( \6423 , \6372 , \6422 );
or \U$6136 ( \6424 , \5097 , \6194 );
nand \U$6137 ( \6425 , \6424 , \6198 );
and \U$6138 ( \6426 , \6371 , \6425 );
or \U$6139 ( \6427 , \5294 , \6200 );
nand \U$6140 ( \6428 , \6427 , \6203 );
nor \U$6141 ( \6429 , \6426 , \6428 );
nand \U$6142 ( \6430 , \6423 , \6429 );
and \U$6143 ( \6431 , \6380 , \6430 );
or \U$6144 ( \6432 , \5513 , \6205 );
nand \U$6145 ( \6433 , \6432 , \6210 );
and \U$6146 ( \6434 , \6375 , \6433 );
or \U$6147 ( \6435 , \5702 , \6212 );
nand \U$6148 ( \6436 , \6435 , \6215 );
nor \U$6149 ( \6437 , \6434 , \6436 );
or \U$6150 ( \6438 , \6379 , \6437 );
or \U$6151 ( \6439 , \5782 , \6217 );
nand \U$6152 ( \6440 , \6439 , \6221 );
and \U$6153 ( \6441 , \6378 , \6440 );
or \U$6154 ( \6442 , \5822 , \6223 );
nand \U$6155 ( \6443 , \6442 , \6226 );
nor \U$6156 ( \6444 , \6441 , \6443 );
nand \U$6157 ( \6445 , \6438 , \6444 );
nor \U$6158 ( \6446 , \6431 , \6445 );
nand \U$6159 ( \6447 , \6416 , \6446 );
and \U$6160 ( \6448 , \6366 , \6447 );
or \U$6161 ( \6449 , \1684 , \6228 );
nand \U$6162 ( \6450 , \6449 , \6235 );
and \U$6163 ( \6451 , \6337 , \6450 );
or \U$6164 ( \6452 , \1992 , \6237 );
nand \U$6165 ( \6453 , \6452 , \6240 );
nor \U$6166 ( \6454 , \6451 , \6453 );
or \U$6167 ( \6455 , \6341 , \6454 );
or \U$6168 ( \6456 , \2299 , \6242 );
nand \U$6169 ( \6457 , \6456 , \6246 );
and \U$6170 ( \6458 , \6340 , \6457 );
or \U$6171 ( \6459 , \2586 , \6248 );
nand \U$6172 ( \6460 , \6459 , \6251 );
nor \U$6173 ( \6461 , \6458 , \6460 );
nand \U$6174 ( \6462 , \6455 , \6461 );
and \U$6175 ( \6463 , \6349 , \6462 );
or \U$6176 ( \6464 , \2855 , \6253 );
nand \U$6177 ( \6465 , \6464 , \6258 );
and \U$6178 ( \6466 , \6344 , \6465 );
or \U$6179 ( \6467 , \3104 , \6260 );
nand \U$6180 ( \6468 , \6467 , \6263 );
nor \U$6181 ( \6469 , \6466 , \6468 );
or \U$6182 ( \6470 , \6348 , \6469 );
or \U$6183 ( \6471 , \3334 , \6265 );
nand \U$6184 ( \6472 , \6471 , \6269 );
and \U$6185 ( \6473 , \6347 , \6472 );
or \U$6186 ( \6474 , \3542 , \6271 );
nand \U$6187 ( \6475 , \6474 , \6274 );
nor \U$6188 ( \6476 , \6473 , \6475 );
nand \U$6189 ( \6477 , \6470 , \6476 );
nor \U$6190 ( \6478 , \6463 , \6477 );
or \U$6191 ( \6479 , \6365 , \6478 );
or \U$6192 ( \6480 , \3736 , \6276 );
nand \U$6193 ( \6481 , \6480 , \6282 );
and \U$6194 ( \6482 , \6352 , \6481 );
or \U$6195 ( \6483 , \3907 , \6284 );
nand \U$6196 ( \6484 , \6483 , \6287 );
nor \U$6197 ( \6485 , \6482 , \6484 );
or \U$6198 ( \6486 , \6356 , \6485 );
or \U$6199 ( \6487 , \4060 , \6289 );
nand \U$6200 ( \6488 , \6487 , \6293 );
and \U$6201 ( \6489 , \6355 , \6488 );
or \U$6202 ( \6490 , \4190 , \6295 );
nand \U$6203 ( \6491 , \6490 , \6298 );
nor \U$6204 ( \6492 , \6489 , \6491 );
nand \U$6205 ( \6493 , \6486 , \6492 );
and \U$6206 ( \6494 , \6364 , \6493 );
or \U$6207 ( \6495 , \4303 , \6300 );
nand \U$6208 ( \6496 , \6495 , \6305 );
and \U$6209 ( \6497 , \6359 , \6496 );
or \U$6210 ( \6498 , \4395 , \6307 );
nand \U$6211 ( \6499 , \6498 , \6310 );
nor \U$6212 ( \6500 , \6497 , \6499 );
or \U$6213 ( \6501 , \6363 , \6500 );
or \U$6214 ( \6502 , \4466 , \6312 );
nand \U$6215 ( \6503 , \6502 , \6316 );
and \U$6216 ( \6504 , \6362 , \6503 );
or \U$6217 ( \6505 , \4510 , \6318 );
nand \U$6218 ( \6506 , \6505 , \6321 );
nor \U$6219 ( \6507 , \6504 , \6506 );
nand \U$6220 ( \6508 , \6501 , \6507 );
nor \U$6221 ( \6509 , \6494 , \6508 );
nand \U$6222 ( \6510 , \6479 , \6509 );
nor \U$6223 ( \6511 , \6448 , \6510 );
not \U$6224 ( \6512 , \6511 );
xnor \U$6225 ( \6513 , \6335 , \6512 );
buf g1974 ( \6514_nG1974 , \6513 );
buf \U$6226 ( \6515 , \6514_nG1974 );
not \U$6227 ( \6516 , \4510 );
nand \U$6228 ( \6517 , \6321 , \6516 );
nand \U$6229 ( \6518 , \5830 , \1838 );
nand \U$6230 ( \6519 , \2146 , \2447 );
nor \U$6231 ( \6520 , \6518 , \6519 );
nand \U$6232 ( \6521 , \2724 , \2982 );
nand \U$6233 ( \6522 , \3221 , \3441 );
nor \U$6234 ( \6523 , \6521 , \6522 );
nand \U$6235 ( \6524 , \6520 , \6523 );
nand \U$6236 ( \6525 , \3642 , \3826 );
nand \U$6237 ( \6526 , \3987 , \4126 );
nor \U$6238 ( \6527 , \6525 , \6526 );
nand \U$6239 ( \6528 , \4250 , \4353 );
nand \U$6240 ( \6529 , \4431 , \4496 );
nor \U$6241 ( \6530 , \6528 , \6529 );
nand \U$6242 ( \6531 , \6527 , \6530 );
nor \U$6243 ( \6532 , \6524 , \6531 );
nand \U$6244 ( \6533 , \6085 , \4838 );
nand \U$6245 ( \6534 , \5005 , \5193 );
nor \U$6246 ( \6535 , \6533 , \6534 );
nand \U$6247 ( \6536 , \5400 , \5629 );
nand \U$6248 ( \6537 , \5748 , \5808 );
nor \U$6249 ( \6538 , \6536 , \6537 );
nand \U$6250 ( \6539 , \6535 , \6538 );
nand \U$6251 ( \6540 , \6132 , \5933 );
nand \U$6252 ( \6541 , \6020 , \6066 );
nor \U$6253 ( \6542 , \6540 , \6541 );
and \U$6254 ( \6543 , \6118 , \6148 );
nor \U$6255 ( \6544 , \6543 , \6154 );
not \U$6256 ( \6545 , \6544 );
and \U$6257 ( \6546 , \6542 , \6545 );
and \U$6258 ( \6547 , \5933 , \6159 );
nor \U$6259 ( \6548 , \6547 , \6166 );
or \U$6260 ( \6549 , \6541 , \6548 );
and \U$6261 ( \6550 , \6066 , \6171 );
nor \U$6262 ( \6551 , \6550 , \6177 );
nand \U$6263 ( \6552 , \6549 , \6551 );
nor \U$6264 ( \6553 , \6546 , \6552 );
or \U$6265 ( \6554 , \6539 , \6553 );
and \U$6266 ( \6555 , \4838 , \6182 );
nor \U$6267 ( \6556 , \6555 , \6190 );
or \U$6268 ( \6557 , \6534 , \6556 );
and \U$6269 ( \6558 , \5193 , \6195 );
nor \U$6270 ( \6559 , \6558 , \6201 );
nand \U$6271 ( \6560 , \6557 , \6559 );
and \U$6272 ( \6561 , \6538 , \6560 );
and \U$6273 ( \6562 , \5629 , \6206 );
nor \U$6274 ( \6563 , \6562 , \6213 );
or \U$6275 ( \6564 , \6537 , \6563 );
and \U$6276 ( \6565 , \5808 , \6218 );
nor \U$6277 ( \6566 , \6565 , \6224 );
nand \U$6278 ( \6567 , \6564 , \6566 );
nor \U$6279 ( \6568 , \6561 , \6567 );
nand \U$6280 ( \6569 , \6554 , \6568 );
and \U$6281 ( \6570 , \6532 , \6569 );
and \U$6282 ( \6571 , \1838 , \6229 );
nor \U$6283 ( \6572 , \6571 , \6238 );
or \U$6284 ( \6573 , \6519 , \6572 );
and \U$6285 ( \6574 , \2447 , \6243 );
nor \U$6286 ( \6575 , \6574 , \6249 );
nand \U$6287 ( \6576 , \6573 , \6575 );
and \U$6288 ( \6577 , \6523 , \6576 );
and \U$6289 ( \6578 , \2982 , \6254 );
nor \U$6290 ( \6579 , \6578 , \6261 );
or \U$6291 ( \6580 , \6522 , \6579 );
and \U$6292 ( \6581 , \3441 , \6266 );
nor \U$6293 ( \6582 , \6581 , \6272 );
nand \U$6294 ( \6583 , \6580 , \6582 );
nor \U$6295 ( \6584 , \6577 , \6583 );
or \U$6296 ( \6585 , \6531 , \6584 );
and \U$6297 ( \6586 , \3826 , \6277 );
nor \U$6298 ( \6587 , \6586 , \6285 );
or \U$6299 ( \6588 , \6526 , \6587 );
and \U$6300 ( \6589 , \4126 , \6290 );
nor \U$6301 ( \6590 , \6589 , \6296 );
nand \U$6302 ( \6591 , \6588 , \6590 );
and \U$6303 ( \6592 , \6530 , \6591 );
and \U$6304 ( \6593 , \4353 , \6301 );
nor \U$6305 ( \6594 , \6593 , \6308 );
or \U$6306 ( \6595 , \6529 , \6594 );
and \U$6307 ( \6596 , \4496 , \6313 );
nor \U$6308 ( \6597 , \6596 , \6319 );
nand \U$6309 ( \6598 , \6595 , \6597 );
nor \U$6310 ( \6599 , \6592 , \6598 );
nand \U$6311 ( \6600 , \6585 , \6599 );
nor \U$6312 ( \6601 , \6570 , \6600 );
not \U$6313 ( \6602 , \6601 );
xnor \U$6314 ( \6603 , \6517 , \6602 );
buf g19cd ( \6604_nG19cd , \6603 );
buf \U$6315 ( \6605 , \6604_nG19cd );
not \U$6316 ( \6606 , \4495 );
nand \U$6317 ( \6607 , \6318 , \6606 );
nand \U$6318 ( \6608 , \6378 , \6336 );
nand \U$6319 ( \6609 , \6337 , \6339 );
nor \U$6320 ( \6610 , \6608 , \6609 );
nand \U$6321 ( \6611 , \6340 , \6343 );
nand \U$6322 ( \6612 , \6344 , \6346 );
nor \U$6323 ( \6613 , \6611 , \6612 );
nand \U$6324 ( \6614 , \6610 , \6613 );
nand \U$6325 ( \6615 , \6347 , \6351 );
nand \U$6326 ( \6616 , \6352 , \6354 );
nor \U$6327 ( \6617 , \6615 , \6616 );
nand \U$6328 ( \6618 , \6355 , \6358 );
nand \U$6329 ( \6619 , \6359 , \6361 );
nor \U$6330 ( \6620 , \6618 , \6619 );
nand \U$6331 ( \6621 , \6617 , \6620 );
nor \U$6332 ( \6622 , \6614 , \6621 );
nand \U$6333 ( \6623 , \6386 , \6367 );
nand \U$6334 ( \6624 , \6368 , \6370 );
nor \U$6335 ( \6625 , \6623 , \6624 );
nand \U$6336 ( \6626 , \6371 , \6374 );
nand \U$6337 ( \6627 , \6375 , \6377 );
nor \U$6338 ( \6628 , \6626 , \6627 );
nand \U$6339 ( \6629 , \6625 , \6628 );
nand \U$6340 ( \6630 , \6390 , \6382 );
nand \U$6341 ( \6631 , \6383 , \6385 );
nor \U$6342 ( \6632 , \6630 , \6631 );
not \U$6343 ( \6633 , \6145 );
and \U$6344 ( \6634 , \6389 , \6633 );
nor \U$6345 ( \6635 , \6634 , \6394 );
not \U$6346 ( \6636 , \6635 );
and \U$6347 ( \6637 , \6632 , \6636 );
and \U$6348 ( \6638 , \6382 , \6397 );
nor \U$6349 ( \6639 , \6638 , \6402 );
or \U$6350 ( \6640 , \6631 , \6639 );
and \U$6351 ( \6641 , \6385 , \6405 );
nor \U$6352 ( \6642 , \6641 , \6409 );
nand \U$6353 ( \6643 , \6640 , \6642 );
nor \U$6354 ( \6644 , \6637 , \6643 );
or \U$6355 ( \6645 , \6629 , \6644 );
and \U$6356 ( \6646 , \6367 , \6412 );
nor \U$6357 ( \6647 , \6646 , \6418 );
or \U$6358 ( \6648 , \6624 , \6647 );
and \U$6359 ( \6649 , \6370 , \6421 );
nor \U$6360 ( \6650 , \6649 , \6425 );
nand \U$6361 ( \6651 , \6648 , \6650 );
and \U$6362 ( \6652 , \6628 , \6651 );
and \U$6363 ( \6653 , \6374 , \6428 );
nor \U$6364 ( \6654 , \6653 , \6433 );
or \U$6365 ( \6655 , \6627 , \6654 );
and \U$6366 ( \6656 , \6377 , \6436 );
nor \U$6367 ( \6657 , \6656 , \6440 );
nand \U$6368 ( \6658 , \6655 , \6657 );
nor \U$6369 ( \6659 , \6652 , \6658 );
nand \U$6370 ( \6660 , \6645 , \6659 );
and \U$6371 ( \6661 , \6622 , \6660 );
and \U$6372 ( \6662 , \6336 , \6443 );
nor \U$6373 ( \6663 , \6662 , \6450 );
or \U$6374 ( \6664 , \6609 , \6663 );
and \U$6375 ( \6665 , \6339 , \6453 );
nor \U$6376 ( \6666 , \6665 , \6457 );
nand \U$6377 ( \6667 , \6664 , \6666 );
and \U$6378 ( \6668 , \6613 , \6667 );
and \U$6379 ( \6669 , \6343 , \6460 );
nor \U$6380 ( \6670 , \6669 , \6465 );
or \U$6381 ( \6671 , \6612 , \6670 );
and \U$6382 ( \6672 , \6346 , \6468 );
nor \U$6383 ( \6673 , \6672 , \6472 );
nand \U$6384 ( \6674 , \6671 , \6673 );
nor \U$6385 ( \6675 , \6668 , \6674 );
or \U$6386 ( \6676 , \6621 , \6675 );
and \U$6387 ( \6677 , \6351 , \6475 );
nor \U$6388 ( \6678 , \6677 , \6481 );
or \U$6389 ( \6679 , \6616 , \6678 );
and \U$6390 ( \6680 , \6354 , \6484 );
nor \U$6391 ( \6681 , \6680 , \6488 );
nand \U$6392 ( \6682 , \6679 , \6681 );
and \U$6393 ( \6683 , \6620 , \6682 );
and \U$6394 ( \6684 , \6358 , \6491 );
nor \U$6395 ( \6685 , \6684 , \6496 );
or \U$6396 ( \6686 , \6619 , \6685 );
and \U$6397 ( \6687 , \6361 , \6499 );
nor \U$6398 ( \6688 , \6687 , \6503 );
nand \U$6399 ( \6689 , \6686 , \6688 );
nor \U$6400 ( \6690 , \6683 , \6689 );
nand \U$6401 ( \6691 , \6676 , \6690 );
nor \U$6402 ( \6692 , \6661 , \6691 );
not \U$6403 ( \6693 , \6692 );
xnor \U$6404 ( \6694 , \6607 , \6693 );
buf g1a27 ( \6695_nG1a27 , \6694 );
buf \U$6405 ( \6696 , \6695_nG1a27 );
not \U$6406 ( \6697 , \4466 );
nand \U$6407 ( \6698 , \6316 , \6697 );
nor \U$6408 ( \6699 , \5831 , \2147 );
nor \U$6409 ( \6700 , \2725 , \3222 );
nand \U$6410 ( \6701 , \6699 , \6700 );
nor \U$6411 ( \6702 , \3643 , \3988 );
nor \U$6412 ( \6703 , \4251 , \4432 );
nand \U$6413 ( \6704 , \6702 , \6703 );
nor \U$6414 ( \6705 , \6701 , \6704 );
nor \U$6415 ( \6706 , \6086 , \5006 );
nor \U$6416 ( \6707 , \5401 , \5749 );
nand \U$6417 ( \6708 , \6706 , \6707 );
nor \U$6418 ( \6709 , \6133 , \6021 );
and \U$6419 ( \6710 , \6709 , \6148 );
or \U$6420 ( \6711 , \6021 , \6160 );
nand \U$6421 ( \6712 , \6711 , \6172 );
nor \U$6422 ( \6713 , \6710 , \6712 );
or \U$6423 ( \6714 , \6708 , \6713 );
or \U$6424 ( \6715 , \5006 , \6183 );
nand \U$6425 ( \6716 , \6715 , \6196 );
and \U$6426 ( \6717 , \6707 , \6716 );
or \U$6427 ( \6718 , \5749 , \6207 );
nand \U$6428 ( \6719 , \6718 , \6219 );
nor \U$6429 ( \6720 , \6717 , \6719 );
nand \U$6430 ( \6721 , \6714 , \6720 );
and \U$6431 ( \6722 , \6705 , \6721 );
or \U$6432 ( \6723 , \2147 , \6230 );
nand \U$6433 ( \6724 , \6723 , \6244 );
and \U$6434 ( \6725 , \6700 , \6724 );
or \U$6435 ( \6726 , \3222 , \6255 );
nand \U$6436 ( \6727 , \6726 , \6267 );
nor \U$6437 ( \6728 , \6725 , \6727 );
or \U$6438 ( \6729 , \6704 , \6728 );
or \U$6439 ( \6730 , \3988 , \6278 );
nand \U$6440 ( \6731 , \6730 , \6291 );
and \U$6441 ( \6732 , \6703 , \6731 );
or \U$6442 ( \6733 , \4432 , \6302 );
nand \U$6443 ( \6734 , \6733 , \6314 );
nor \U$6444 ( \6735 , \6732 , \6734 );
nand \U$6445 ( \6736 , \6729 , \6735 );
nor \U$6446 ( \6737 , \6722 , \6736 );
not \U$6447 ( \6738 , \6737 );
xnor \U$6448 ( \6739 , \6698 , \6738 );
buf g1a53 ( \6740_nG1a53 , \6739 );
buf \U$6449 ( \6741 , \6740_nG1a53 );
not \U$6450 ( \6742 , \4430 );
nand \U$6451 ( \6743 , \6312 , \6742 );
nor \U$6452 ( \6744 , \6379 , \6338 );
nor \U$6453 ( \6745 , \6341 , \6345 );
nand \U$6454 ( \6746 , \6744 , \6745 );
nor \U$6455 ( \6747 , \6348 , \6353 );
nor \U$6456 ( \6748 , \6356 , \6360 );
nand \U$6457 ( \6749 , \6747 , \6748 );
nor \U$6458 ( \6750 , \6746 , \6749 );
nor \U$6459 ( \6751 , \6387 , \6369 );
nor \U$6460 ( \6752 , \6372 , \6376 );
nand \U$6461 ( \6753 , \6751 , \6752 );
nor \U$6462 ( \6754 , \6391 , \6384 );
and \U$6463 ( \6755 , \6754 , \6633 );
or \U$6464 ( \6756 , \6384 , \6398 );
nand \U$6465 ( \6757 , \6756 , \6406 );
nor \U$6466 ( \6758 , \6755 , \6757 );
or \U$6467 ( \6759 , \6753 , \6758 );
or \U$6468 ( \6760 , \6369 , \6413 );
nand \U$6469 ( \6761 , \6760 , \6422 );
and \U$6470 ( \6762 , \6752 , \6761 );
or \U$6471 ( \6763 , \6376 , \6429 );
nand \U$6472 ( \6764 , \6763 , \6437 );
nor \U$6473 ( \6765 , \6762 , \6764 );
nand \U$6474 ( \6766 , \6759 , \6765 );
and \U$6475 ( \6767 , \6750 , \6766 );
or \U$6476 ( \6768 , \6338 , \6444 );
nand \U$6477 ( \6769 , \6768 , \6454 );
and \U$6478 ( \6770 , \6745 , \6769 );
or \U$6479 ( \6771 , \6345 , \6461 );
nand \U$6480 ( \6772 , \6771 , \6469 );
nor \U$6481 ( \6773 , \6770 , \6772 );
or \U$6482 ( \6774 , \6749 , \6773 );
or \U$6483 ( \6775 , \6353 , \6476 );
nand \U$6484 ( \6776 , \6775 , \6485 );
and \U$6485 ( \6777 , \6748 , \6776 );
or \U$6486 ( \6778 , \6360 , \6492 );
nand \U$6487 ( \6779 , \6778 , \6500 );
nor \U$6488 ( \6780 , \6777 , \6779 );
nand \U$6489 ( \6781 , \6774 , \6780 );
nor \U$6490 ( \6782 , \6767 , \6781 );
not \U$6491 ( \6783 , \6782 );
xnor \U$6492 ( \6784 , \6743 , \6783 );
buf g1a7f ( \6785_nG1a7f , \6784 );
buf \U$6493 ( \6786 , \6785_nG1a7f );
not \U$6494 ( \6787 , \4395 );
nand \U$6495 ( \6788 , \6310 , \6787 );
nor \U$6496 ( \6789 , \6537 , \6518 );
nor \U$6497 ( \6790 , \6519 , \6521 );
nand \U$6498 ( \6791 , \6789 , \6790 );
nor \U$6499 ( \6792 , \6522 , \6525 );
nor \U$6500 ( \6793 , \6526 , \6528 );
nand \U$6501 ( \6794 , \6792 , \6793 );
nor \U$6502 ( \6795 , \6791 , \6794 );
nor \U$6503 ( \6796 , \6541 , \6533 );
nor \U$6504 ( \6797 , \6534 , \6536 );
nand \U$6505 ( \6798 , \6796 , \6797 );
or \U$6506 ( \6799 , \6540 , \6544 );
nand \U$6507 ( \6800 , \6799 , \6548 );
not \U$6508 ( \6801 , \6800 );
or \U$6509 ( \6802 , \6798 , \6801 );
or \U$6510 ( \6803 , \6533 , \6551 );
nand \U$6511 ( \6804 , \6803 , \6556 );
and \U$6512 ( \6805 , \6797 , \6804 );
or \U$6513 ( \6806 , \6536 , \6559 );
nand \U$6514 ( \6807 , \6806 , \6563 );
nor \U$6515 ( \6808 , \6805 , \6807 );
nand \U$6516 ( \6809 , \6802 , \6808 );
and \U$6517 ( \6810 , \6795 , \6809 );
or \U$6518 ( \6811 , \6518 , \6566 );
nand \U$6519 ( \6812 , \6811 , \6572 );
and \U$6520 ( \6813 , \6790 , \6812 );
or \U$6521 ( \6814 , \6521 , \6575 );
nand \U$6522 ( \6815 , \6814 , \6579 );
nor \U$6523 ( \6816 , \6813 , \6815 );
or \U$6524 ( \6817 , \6794 , \6816 );
or \U$6525 ( \6818 , \6525 , \6582 );
nand \U$6526 ( \6819 , \6818 , \6587 );
and \U$6527 ( \6820 , \6793 , \6819 );
or \U$6528 ( \6821 , \6528 , \6590 );
nand \U$6529 ( \6822 , \6821 , \6594 );
nor \U$6530 ( \6823 , \6820 , \6822 );
nand \U$6531 ( \6824 , \6817 , \6823 );
nor \U$6532 ( \6825 , \6810 , \6824 );
not \U$6533 ( \6826 , \6825 );
xnor \U$6534 ( \6827 , \6788 , \6826 );
buf g1aa9 ( \6828_nG1aa9 , \6827 );
buf \U$6535 ( \6829 , \6828_nG1aa9 );
not \U$6536 ( \6830 , \4352 );
nand \U$6537 ( \6831 , \6307 , \6830 );
nor \U$6538 ( \6832 , \6627 , \6608 );
nor \U$6539 ( \6833 , \6609 , \6611 );
nand \U$6540 ( \6834 , \6832 , \6833 );
nor \U$6541 ( \6835 , \6612 , \6615 );
nor \U$6542 ( \6836 , \6616 , \6618 );
nand \U$6543 ( \6837 , \6835 , \6836 );
nor \U$6544 ( \6838 , \6834 , \6837 );
nor \U$6545 ( \6839 , \6631 , \6623 );
nor \U$6546 ( \6840 , \6624 , \6626 );
nand \U$6547 ( \6841 , \6839 , \6840 );
or \U$6548 ( \6842 , \6630 , \6635 );
nand \U$6549 ( \6843 , \6842 , \6639 );
not \U$6550 ( \6844 , \6843 );
or \U$6551 ( \6845 , \6841 , \6844 );
or \U$6552 ( \6846 , \6623 , \6642 );
nand \U$6553 ( \6847 , \6846 , \6647 );
and \U$6554 ( \6848 , \6840 , \6847 );
or \U$6555 ( \6849 , \6626 , \6650 );
nand \U$6556 ( \6850 , \6849 , \6654 );
nor \U$6557 ( \6851 , \6848 , \6850 );
nand \U$6558 ( \6852 , \6845 , \6851 );
and \U$6559 ( \6853 , \6838 , \6852 );
or \U$6560 ( \6854 , \6608 , \6657 );
nand \U$6561 ( \6855 , \6854 , \6663 );
and \U$6562 ( \6856 , \6833 , \6855 );
or \U$6563 ( \6857 , \6611 , \6666 );
nand \U$6564 ( \6858 , \6857 , \6670 );
nor \U$6565 ( \6859 , \6856 , \6858 );
or \U$6566 ( \6860 , \6837 , \6859 );
or \U$6567 ( \6861 , \6615 , \6673 );
nand \U$6568 ( \6862 , \6861 , \6678 );
and \U$6569 ( \6863 , \6836 , \6862 );
or \U$6570 ( \6864 , \6618 , \6681 );
nand \U$6571 ( \6865 , \6864 , \6685 );
nor \U$6572 ( \6866 , \6863 , \6865 );
nand \U$6573 ( \6867 , \6860 , \6866 );
nor \U$6574 ( \6868 , \6853 , \6867 );
not \U$6575 ( \6869 , \6868 );
xnor \U$6576 ( \6870 , \6831 , \6869 );
buf g1ad3 ( \6871_nG1ad3 , \6870 );
buf \U$6577 ( \6872 , \6871_nG1ad3 );
not \U$6578 ( \6873 , \4303 );
nand \U$6579 ( \6874 , \6305 , \6873 );
nand \U$6580 ( \6875 , \5832 , \2726 );
nand \U$6581 ( \6876 , \3644 , \4252 );
nor \U$6582 ( \6877 , \6875 , \6876 );
nand \U$6583 ( \6878 , \6087 , \5402 );
not \U$6584 ( \6879 , \6161 );
or \U$6585 ( \6880 , \6878 , \6879 );
and \U$6586 ( \6881 , \5402 , \6184 );
nor \U$6587 ( \6882 , \6881 , \6208 );
nand \U$6588 ( \6883 , \6880 , \6882 );
and \U$6589 ( \6884 , \6877 , \6883 );
and \U$6590 ( \6885 , \2726 , \6231 );
nor \U$6591 ( \6886 , \6885 , \6256 );
or \U$6592 ( \6887 , \6876 , \6886 );
and \U$6593 ( \6888 , \4252 , \6279 );
nor \U$6594 ( \6889 , \6888 , \6303 );
nand \U$6595 ( \6890 , \6887 , \6889 );
nor \U$6596 ( \6891 , \6884 , \6890 );
not \U$6597 ( \6892 , \6891 );
xnor \U$6598 ( \6893 , \6874 , \6892 );
buf g1ae9 ( \6894_nG1ae9 , \6893 );
buf \U$6599 ( \6895 , \6894_nG1ae9 );
not \U$6600 ( \6896 , \4249 );
nand \U$6601 ( \6897 , \6300 , \6896 );
nand \U$6602 ( \6898 , \6380 , \6342 );
nand \U$6603 ( \6899 , \6349 , \6357 );
nor \U$6604 ( \6900 , \6898 , \6899 );
nand \U$6605 ( \6901 , \6388 , \6373 );
not \U$6606 ( \6902 , \6399 );
or \U$6607 ( \6903 , \6901 , \6902 );
and \U$6608 ( \6904 , \6373 , \6414 );
nor \U$6609 ( \6905 , \6904 , \6430 );
nand \U$6610 ( \6906 , \6903 , \6905 );
and \U$6611 ( \6907 , \6900 , \6906 );
and \U$6612 ( \6908 , \6342 , \6445 );
nor \U$6613 ( \6909 , \6908 , \6462 );
or \U$6614 ( \6910 , \6899 , \6909 );
and \U$6615 ( \6911 , \6357 , \6477 );
nor \U$6616 ( \6912 , \6911 , \6493 );
nand \U$6617 ( \6913 , \6910 , \6912 );
nor \U$6618 ( \6914 , \6907 , \6913 );
not \U$6619 ( \6915 , \6914 );
xnor \U$6620 ( \6916 , \6897 , \6915 );
buf g1aff ( \6917_nG1aff , \6916 );
buf \U$6621 ( \6918 , \6917_nG1aff );
not \U$6622 ( \6919 , \4190 );
nand \U$6623 ( \6920 , \6298 , \6919 );
nand \U$6624 ( \6921 , \6538 , \6520 );
nand \U$6625 ( \6922 , \6523 , \6527 );
nor \U$6626 ( \6923 , \6921 , \6922 );
nand \U$6627 ( \6924 , \6542 , \6535 );
or \U$6628 ( \6925 , \6924 , \6544 );
and \U$6629 ( \6926 , \6535 , \6552 );
nor \U$6630 ( \6927 , \6926 , \6560 );
nand \U$6631 ( \6928 , \6925 , \6927 );
and \U$6632 ( \6929 , \6923 , \6928 );
and \U$6633 ( \6930 , \6520 , \6567 );
nor \U$6634 ( \6931 , \6930 , \6576 );
or \U$6635 ( \6932 , \6922 , \6931 );
and \U$6636 ( \6933 , \6527 , \6583 );
nor \U$6637 ( \6934 , \6933 , \6591 );
nand \U$6638 ( \6935 , \6932 , \6934 );
nor \U$6639 ( \6936 , \6929 , \6935 );
not \U$6640 ( \6937 , \6936 );
xnor \U$6641 ( \6938 , \6920 , \6937 );
buf g1b14 ( \6939_nG1b14 , \6938 );
buf \U$6642 ( \6940 , \6939_nG1b14 );
not \U$6643 ( \6941 , \4125 );
nand \U$6644 ( \6942 , \6295 , \6941 );
nand \U$6645 ( \6943 , \6628 , \6610 );
nand \U$6646 ( \6944 , \6613 , \6617 );
nor \U$6647 ( \6945 , \6943 , \6944 );
nand \U$6648 ( \6946 , \6632 , \6625 );
or \U$6649 ( \6947 , \6946 , \6635 );
and \U$6650 ( \6948 , \6625 , \6643 );
nor \U$6651 ( \6949 , \6948 , \6651 );
nand \U$6652 ( \6950 , \6947 , \6949 );
and \U$6653 ( \6951 , \6945 , \6950 );
and \U$6654 ( \6952 , \6610 , \6658 );
nor \U$6655 ( \6953 , \6952 , \6667 );
or \U$6656 ( \6954 , \6944 , \6953 );
and \U$6657 ( \6955 , \6617 , \6674 );
nor \U$6658 ( \6956 , \6955 , \6682 );
nand \U$6659 ( \6957 , \6954 , \6956 );
nor \U$6660 ( \6958 , \6951 , \6957 );
not \U$6661 ( \6959 , \6958 );
xnor \U$6662 ( \6960 , \6942 , \6959 );
buf g1b29 ( \6961_nG1b29 , \6960 );
buf \U$6663 ( \6962 , \6961_nG1b29 );
not \U$6664 ( \6963 , \4060 );
nand \U$6665 ( \6964 , \6293 , \6963 );
nand \U$6666 ( \6965 , \6707 , \6699 );
nand \U$6667 ( \6966 , \6700 , \6702 );
nor \U$6668 ( \6967 , \6965 , \6966 );
nand \U$6669 ( \6968 , \6709 , \6706 );
or \U$6670 ( \6969 , \6968 , \6149 );
and \U$6671 ( \6970 , \6706 , \6712 );
nor \U$6672 ( \6971 , \6970 , \6716 );
nand \U$6673 ( \6972 , \6969 , \6971 );
and \U$6674 ( \6973 , \6967 , \6972 );
and \U$6675 ( \6974 , \6699 , \6719 );
nor \U$6676 ( \6975 , \6974 , \6724 );
or \U$6677 ( \6976 , \6966 , \6975 );
and \U$6678 ( \6977 , \6702 , \6727 );
nor \U$6679 ( \6978 , \6977 , \6731 );
nand \U$6680 ( \6979 , \6976 , \6978 );
nor \U$6681 ( \6980 , \6973 , \6979 );
not \U$6682 ( \6981 , \6980 );
xnor \U$6683 ( \6982 , \6964 , \6981 );
buf g1b3e ( \6983_nG1b3e , \6982 );
buf \U$6684 ( \6984 , \6983_nG1b3e );
not \U$6685 ( \6985 , \3986 );
nand \U$6686 ( \6986 , \6289 , \6985 );
nand \U$6687 ( \6987 , \6752 , \6744 );
nand \U$6688 ( \6988 , \6745 , \6747 );
nor \U$6689 ( \6989 , \6987 , \6988 );
nand \U$6690 ( \6990 , \6754 , \6751 );
or \U$6691 ( \6991 , \6990 , \6145 );
and \U$6692 ( \6992 , \6751 , \6757 );
nor \U$6693 ( \6993 , \6992 , \6761 );
nand \U$6694 ( \6994 , \6991 , \6993 );
and \U$6695 ( \6995 , \6989 , \6994 );
and \U$6696 ( \6996 , \6744 , \6764 );
nor \U$6697 ( \6997 , \6996 , \6769 );
or \U$6698 ( \6998 , \6988 , \6997 );
and \U$6699 ( \6999 , \6747 , \6772 );
nor \U$6700 ( \7000 , \6999 , \6776 );
nand \U$6701 ( \7001 , \6998 , \7000 );
nor \U$6702 ( \7002 , \6995 , \7001 );
not \U$6703 ( \7003 , \7002 );
xnor \U$6704 ( \7004 , \6986 , \7003 );
buf g1b53 ( \7005_nG1b53 , \7004 );
buf \U$6705 ( \7006 , \7005_nG1b53 );
not \U$6706 ( \7007 , \3907 );
nand \U$6707 ( \7008 , \6287 , \7007 );
nand \U$6708 ( \7009 , \6797 , \6789 );
nand \U$6709 ( \7010 , \6790 , \6792 );
nor \U$6710 ( \7011 , \7009 , \7010 );
and \U$6711 ( \7012 , \6796 , \6800 );
nor \U$6712 ( \7013 , \7012 , \6804 );
not \U$6713 ( \7014 , \7013 );
and \U$6714 ( \7015 , \7011 , \7014 );
and \U$6715 ( \7016 , \6789 , \6807 );
nor \U$6716 ( \7017 , \7016 , \6812 );
or \U$6717 ( \7018 , \7010 , \7017 );
and \U$6718 ( \7019 , \6792 , \6815 );
nor \U$6719 ( \7020 , \7019 , \6819 );
nand \U$6720 ( \7021 , \7018 , \7020 );
nor \U$6721 ( \7022 , \7015 , \7021 );
not \U$6722 ( \7023 , \7022 );
xnor \U$6723 ( \7024 , \7008 , \7023 );
buf g1b66 ( \7025_nG1b66 , \7024 );
buf \U$6724 ( \7026 , \7025_nG1b66 );
not \U$6725 ( \7027 , \3825 );
nand \U$6726 ( \7028 , \6284 , \7027 );
nand \U$6727 ( \7029 , \6840 , \6832 );
nand \U$6728 ( \7030 , \6833 , \6835 );
nor \U$6729 ( \7031 , \7029 , \7030 );
and \U$6730 ( \7032 , \6839 , \6843 );
nor \U$6731 ( \7033 , \7032 , \6847 );
not \U$6732 ( \7034 , \7033 );
and \U$6733 ( \7035 , \7031 , \7034 );
and \U$6734 ( \7036 , \6832 , \6850 );
nor \U$6735 ( \7037 , \7036 , \6855 );
or \U$6736 ( \7038 , \7030 , \7037 );
and \U$6737 ( \7039 , \6835 , \6858 );
nor \U$6738 ( \7040 , \7039 , \6862 );
nand \U$6739 ( \7041 , \7038 , \7040 );
nor \U$6740 ( \7042 , \7035 , \7041 );
not \U$6741 ( \7043 , \7042 );
xnor \U$6742 ( \7044 , \7028 , \7043 );
buf g1b79 ( \7045_nG1b79 , \7044 );
buf \U$6743 ( \7046 , \7045_nG1b79 );
not \U$6744 ( \7047 , \3736 );
nand \U$6745 ( \7048 , \6282 , \7047 );
nor \U$6746 ( \7049 , \5833 , \3645 );
not \U$6747 ( \7050 , \6185 );
and \U$6748 ( \7051 , \7049 , \7050 );
or \U$6749 ( \7052 , \3645 , \6232 );
nand \U$6750 ( \7053 , \7052 , \6280 );
nor \U$6751 ( \7054 , \7051 , \7053 );
not \U$6752 ( \7055 , \7054 );
xnor \U$6753 ( \7056 , \7048 , \7055 );
buf g1b84 ( \7057_nG1b84 , \7056 );
buf \U$6754 ( \7058 , \7057_nG1b84 );
not \U$6755 ( \7059 , \3641 );
nand \U$6756 ( \7060 , \6276 , \7059 );
nor \U$6757 ( \7061 , \6381 , \6350 );
not \U$6758 ( \7062 , \6415 );
and \U$6759 ( \7063 , \7061 , \7062 );
or \U$6760 ( \7064 , \6350 , \6446 );
nand \U$6761 ( \7065 , \7064 , \6478 );
nor \U$6762 ( \7066 , \7063 , \7065 );
not \U$6763 ( \7067 , \7066 );
xnor \U$6764 ( \7068 , \7060 , \7067 );
buf g1b8f ( \7069_nG1b8f , \7068 );
buf \U$6765 ( \7070 , \7069_nG1b8f );
not \U$6766 ( \7071 , \3542 );
nand \U$6767 ( \7072 , \6274 , \7071 );
nor \U$6768 ( \7073 , \6539 , \6524 );
not \U$6769 ( \7074 , \6553 );
and \U$6770 ( \7075 , \7073 , \7074 );
or \U$6771 ( \7076 , \6524 , \6568 );
nand \U$6772 ( \7077 , \7076 , \6584 );
nor \U$6773 ( \7078 , \7075 , \7077 );
not \U$6774 ( \7079 , \7078 );
xnor \U$6775 ( \7080 , \7072 , \7079 );
buf g1b9a ( \7081_nG1b9a , \7080 );
buf \U$6776 ( \7082 , \7081_nG1b9a );
not \U$6777 ( \7083 , \3440 );
nand \U$6778 ( \7084 , \6271 , \7083 );
nor \U$6779 ( \7085 , \6629 , \6614 );
not \U$6780 ( \7086 , \6644 );
and \U$6781 ( \7087 , \7085 , \7086 );
or \U$6782 ( \7088 , \6614 , \6659 );
nand \U$6783 ( \7089 , \7088 , \6675 );
nor \U$6784 ( \7090 , \7087 , \7089 );
not \U$6785 ( \7091 , \7090 );
xnor \U$6786 ( \7092 , \7084 , \7091 );
buf g1ba5 ( \7093_nG1ba5 , \7092 );
buf \U$6787 ( \7094 , \7093_nG1ba5 );
not \U$6788 ( \7095 , \3334 );
nand \U$6789 ( \7096 , \6269 , \7095 );
nor \U$6790 ( \7097 , \6708 , \6701 );
not \U$6791 ( \7098 , \6713 );
and \U$6792 ( \7099 , \7097 , \7098 );
or \U$6793 ( \7100 , \6701 , \6720 );
nand \U$6794 ( \7101 , \7100 , \6728 );
nor \U$6795 ( \7102 , \7099 , \7101 );
not \U$6796 ( \7103 , \7102 );
xnor \U$6797 ( \7104 , \7096 , \7103 );
buf g1bb0 ( \7105_nG1bb0 , \7104 );
buf \U$6798 ( \7106 , \7105_nG1bb0 );
not \U$6799 ( \7107 , \3220 );
nand \U$6800 ( \7108 , \6265 , \7107 );
nor \U$6801 ( \7109 , \6753 , \6746 );
not \U$6802 ( \7110 , \6758 );
and \U$6803 ( \7111 , \7109 , \7110 );
or \U$6804 ( \7112 , \6746 , \6765 );
nand \U$6805 ( \7113 , \7112 , \6773 );
nor \U$6806 ( \7114 , \7111 , \7113 );
not \U$6807 ( \7115 , \7114 );
xnor \U$6808 ( \7116 , \7108 , \7115 );
buf g1bbb ( \7117_nG1bbb , \7116 );
buf \U$6809 ( \7118 , \7117_nG1bbb );
not \U$6810 ( \7119 , \3104 );
nand \U$6811 ( \7120 , \6263 , \7119 );
nor \U$6812 ( \7121 , \6798 , \6791 );
and \U$6813 ( \7122 , \7121 , \6800 );
or \U$6814 ( \7123 , \6791 , \6808 );
nand \U$6815 ( \7124 , \7123 , \6816 );
nor \U$6816 ( \7125 , \7122 , \7124 );
not \U$6817 ( \7126 , \7125 );
xnor \U$6818 ( \7127 , \7120 , \7126 );
buf g1bc5 ( \7128_nG1bc5 , \7127 );
buf \U$6819 ( \7129 , \7128_nG1bc5 );
not \U$6820 ( \7130 , \2981 );
nand \U$6821 ( \7131 , \6260 , \7130 );
nor \U$6822 ( \7132 , \6841 , \6834 );
and \U$6823 ( \7133 , \7132 , \6843 );
or \U$6824 ( \7134 , \6834 , \6851 );
nand \U$6825 ( \7135 , \7134 , \6859 );
nor \U$6826 ( \7136 , \7133 , \7135 );
not \U$6827 ( \7137 , \7136 );
xnor \U$6828 ( \7138 , \7131 , \7137 );
buf g1bcf ( \7139_nG1bcf , \7138 );
buf \U$6829 ( \7140 , \7139_nG1bcf );
not \U$6830 ( \7141 , \2855 );
nand \U$6831 ( \7142 , \6258 , \7141 );
nor \U$6832 ( \7143 , \6878 , \6875 );
and \U$6833 ( \7144 , \7143 , \6161 );
or \U$6834 ( \7145 , \6875 , \6882 );
nand \U$6835 ( \7146 , \7145 , \6886 );
nor \U$6836 ( \7147 , \7144 , \7146 );
not \U$6837 ( \7148 , \7147 );
xnor \U$6838 ( \7149 , \7142 , \7148 );
buf g1bd9 ( \7150_nG1bd9 , \7149 );
buf \U$6839 ( \7151 , \7150_nG1bd9 );
not \U$6840 ( \7152 , \2723 );
nand \U$6841 ( \7153 , \6253 , \7152 );
nor \U$6842 ( \7154 , \6901 , \6898 );
and \U$6843 ( \7155 , \7154 , \6399 );
or \U$6844 ( \7156 , \6898 , \6905 );
nand \U$6845 ( \7157 , \7156 , \6909 );
nor \U$6846 ( \7158 , \7155 , \7157 );
not \U$6847 ( \7159 , \7158 );
xnor \U$6848 ( \7160 , \7153 , \7159 );
buf g1be3 ( \7161_nG1be3 , \7160 );
buf \U$6849 ( \7162 , \7161_nG1be3 );
not \U$6850 ( \7163 , \2586 );
nand \U$6851 ( \7164 , \6251 , \7163 );
nor \U$6852 ( \7165 , \6924 , \6921 );
and \U$6853 ( \7166 , \7165 , \6545 );
or \U$6854 ( \7167 , \6921 , \6927 );
nand \U$6855 ( \7168 , \7167 , \6931 );
nor \U$6856 ( \7169 , \7166 , \7168 );
not \U$6857 ( \7170 , \7169 );
xnor \U$6858 ( \7171 , \7164 , \7170 );
buf g1bed ( \7172_nG1bed , \7171 );
buf \U$6859 ( \7173 , \7172_nG1bed );
not \U$6860 ( \7174 , \2446 );
nand \U$6861 ( \7175 , \6248 , \7174 );
nor \U$6862 ( \7176 , \6946 , \6943 );
and \U$6863 ( \7177 , \7176 , \6636 );
or \U$6864 ( \7178 , \6943 , \6949 );
nand \U$6865 ( \7179 , \7178 , \6953 );
nor \U$6866 ( \7180 , \7177 , \7179 );
not \U$6867 ( \7181 , \7180 );
xnor \U$6868 ( \7182 , \7175 , \7181 );
buf g1bf7 ( \7183_nG1bf7 , \7182 );
buf \U$6869 ( \7184 , \7183_nG1bf7 );
not \U$6870 ( \7185 , \2299 );
nand \U$6871 ( \7186 , \6246 , \7185 );
nor \U$6872 ( \7187 , \6968 , \6965 );
and \U$6873 ( \7188 , \7187 , \6148 );
or \U$6874 ( \7189 , \6965 , \6971 );
nand \U$6875 ( \7190 , \7189 , \6975 );
nor \U$6876 ( \7191 , \7188 , \7190 );
not \U$6877 ( \7192 , \7191 );
xnor \U$6878 ( \7193 , \7186 , \7192 );
buf g1c01 ( \7194_nG1c01 , \7193 );
buf \U$6879 ( \7195 , \7194_nG1c01 );
not \U$6880 ( \7196 , \2145 );
nand \U$6881 ( \7197 , \6242 , \7196 );
nor \U$6882 ( \7198 , \6990 , \6987 );
and \U$6883 ( \7199 , \7198 , \6633 );
or \U$6884 ( \7200 , \6987 , \6993 );
nand \U$6885 ( \7201 , \7200 , \6997 );
nor \U$6886 ( \7202 , \7199 , \7201 );
not \U$6887 ( \7203 , \7202 );
xnor \U$6888 ( \7204 , \7197 , \7203 );
buf g1c0b ( \7205_nG1c0b , \7204 );
buf \U$6889 ( \7206 , \7205_nG1c0b );
not \U$6890 ( \7207 , \1992 );
nand \U$6891 ( \7208 , \6240 , \7207 );
or \U$6892 ( \7209 , \7009 , \7013 );
nand \U$6893 ( \7210 , \7209 , \7017 );
xnor \U$6894 ( \7211 , \7208 , \7210 );
buf g1c11 ( \7212_nG1c11 , \7211 );
buf \U$6895 ( \7213 , \7212_nG1c11 );
not \U$6896 ( \7214 , \1837 );
nand \U$6897 ( \7215 , \6237 , \7214 );
or \U$6898 ( \7216 , \7029 , \7033 );
nand \U$6899 ( \7217 , \7216 , \7037 );
xnor \U$6900 ( \7218 , \7215 , \7217 );
buf g1c17 ( \7219_nG1c17 , \7218 );
buf \U$6901 ( \7220 , \7219_nG1c17 );
not \U$6902 ( \7221 , \1684 );
nand \U$6903 ( \7222 , \6235 , \7221 );
xnor \U$6904 ( \7223 , \7222 , \6233 );
buf g1c1b ( \7224_nG1c1b , \7223 );
buf \U$6905 ( \7225 , \7224_nG1c1b );
not \U$6906 ( \7226 , \5829 );
nand \U$6907 ( \7227 , \6228 , \7226 );
xnor \U$6908 ( \7228 , \7227 , \6447 );
buf g1c1f ( \7229_nG1c1f , \7228 );
buf \U$6909 ( \7230 , \7229_nG1c1f );
not \U$6910 ( \7231 , \5822 );
nand \U$6911 ( \7232 , \6226 , \7231 );
xnor \U$6912 ( \7233 , \7232 , \6569 );
buf g1c23 ( \7234_nG1c23 , \7233 );
buf \U$6913 ( \7235 , \7234_nG1c23 );
not \U$6914 ( \7236 , \5807 );
nand \U$6915 ( \7237 , \6223 , \7236 );
xnor \U$6916 ( \7238 , \7237 , \6660 );
buf g1c27 ( \7239_nG1c27 , \7238 );
buf \U$6917 ( \7240 , \7239_nG1c27 );
not \U$6918 ( \7241 , \5782 );
nand \U$6919 ( \7242 , \6221 , \7241 );
xnor \U$6920 ( \7243 , \7242 , \6721 );
buf g1c2b ( \7244_nG1c2b , \7243 );
buf \U$6921 ( \7245 , \7244_nG1c2b );
not \U$6922 ( \7246 , \5747 );
nand \U$6923 ( \7247 , \6217 , \7246 );
xnor \U$6924 ( \7248 , \7247 , \6766 );
buf g1c2f ( \7249_nG1c2f , \7248 );
buf \U$6925 ( \7250 , \7249_nG1c2f );
not \U$6926 ( \7251 , \5702 );
nand \U$6927 ( \7252 , \6215 , \7251 );
xnor \U$6928 ( \7253 , \7252 , \6809 );
buf g1c33 ( \7254_nG1c33 , \7253 );
buf \U$6929 ( \7255 , \7254_nG1c33 );
not \U$6930 ( \7256 , \5628 );
nand \U$6931 ( \7257 , \6212 , \7256 );
xnor \U$6932 ( \7258 , \7257 , \6852 );
buf g1c37 ( \7259_nG1c37 , \7258 );
buf \U$6933 ( \7260 , \7259_nG1c37 );
not \U$6934 ( \7261 , \5513 );
nand \U$6935 ( \7262 , \6210 , \7261 );
xnor \U$6936 ( \7263 , \7262 , \6883 );
buf g1c3b ( \7264_nG1c3b , \7263 );
buf \U$6937 ( \7265 , \7264_nG1c3b );
not \U$6938 ( \7266 , \5399 );
nand \U$6939 ( \7267 , \6205 , \7266 );
xnor \U$6940 ( \7268 , \7267 , \6906 );
buf g1c3f ( \7269_nG1c3f , \7268 );
buf \U$6941 ( \7270 , \7269_nG1c3f );
not \U$6942 ( \7271 , \5294 );
nand \U$6943 ( \7272 , \6203 , \7271 );
xnor \U$6944 ( \7273 , \7272 , \6928 );
buf g1c43 ( \7274_nG1c43 , \7273 );
buf \U$6945 ( \7275 , \7274_nG1c43 );
not \U$6946 ( \7276 , \5192 );
nand \U$6947 ( \7277 , \6200 , \7276 );
xnor \U$6948 ( \7278 , \7277 , \6950 );
buf g1c47 ( \7279_nG1c47 , \7278 );
buf \U$6949 ( \7280 , \7279_nG1c47 );
not \U$6950 ( \7281 , \5097 );
nand \U$6951 ( \7282 , \6198 , \7281 );
xnor \U$6952 ( \7283 , \7282 , \6972 );
buf g1c4b ( \7284_nG1c4b , \7283 );
buf \U$6953 ( \7285 , \7284_nG1c4b );
not \U$6954 ( \7286 , \5004 );
nand \U$6955 ( \7287 , \6194 , \7286 );
xnor \U$6956 ( \7288 , \7287 , \6994 );
buf g1c4f ( \7289_nG1c4f , \7288 );
buf \U$6957 ( \7290 , \7289_nG1c4f );
not \U$6958 ( \7291 , \4919 );
nand \U$6959 ( \7292 , \6192 , \7291 );
xnor \U$6960 ( \7293 , \7292 , \7014 );
buf g1c53 ( \7294_nG1c53 , \7293 );
buf \U$6961 ( \7295 , \7294_nG1c53 );
not \U$6962 ( \7296 , \4837 );
nand \U$6963 ( \7297 , \6189 , \7296 );
xnor \U$6964 ( \7298 , \7297 , \7034 );
buf g1c57 ( \7299_nG1c57 , \7298 );
buf \U$6965 ( \7300 , \7299_nG1c57 );
not \U$6966 ( \7301 , \4762 );
nand \U$6967 ( \7302 , \6187 , \7301 );
xnor \U$6968 ( \7303 , \7302 , \7050 );
buf g1c5b ( \7304_nG1c5b , \7303 );
buf \U$6969 ( \7305 , \7304_nG1c5b );
not \U$6970 ( \7306 , \6084 );
nand \U$6971 ( \7307 , \6181 , \7306 );
xnor \U$6972 ( \7308 , \7307 , \7062 );
buf g1c5f ( \7309_nG1c5f , \7308 );
buf \U$6973 ( \7310 , \7309_nG1c5f );
not \U$6974 ( \7311 , \6077 );
nand \U$6975 ( \7312 , \6179 , \7311 );
xnor \U$6976 ( \7313 , \7312 , \7074 );
buf g1c63 ( \7314_nG1c63 , \7313 );
buf \U$6977 ( \7315 , \7314_nG1c63 );
not \U$6978 ( \7316 , \6065 );
nand \U$6979 ( \7317 , \6176 , \7316 );
xnor \U$6980 ( \7318 , \7317 , \7086 );
buf g1c67 ( \7319_nG1c67 , \7318 );
buf \U$6981 ( \7320 , \7319_nG1c67 );
not \U$6982 ( \7321 , \6048 );
nand \U$6983 ( \7322 , \6174 , \7321 );
xnor \U$6984 ( \7323 , \7322 , \7098 );
buf g1c6b ( \7324_nG1c6b , \7323 );
buf \U$6985 ( \7325 , \7324_nG1c6b );
not \U$6986 ( \7326 , \6019 );
nand \U$6987 ( \7327 , \6170 , \7326 );
xnor \U$6988 ( \7328 , \7327 , \7110 );
buf g1c6f ( \7329_nG1c6f , \7328 );
buf \U$6989 ( \7330 , \7329_nG1c6f );
not \U$6990 ( \7331 , \5974 );
nand \U$6991 ( \7332 , \6168 , \7331 );
xnor \U$6992 ( \7333 , \7332 , \6800 );
buf g1c73 ( \7334_nG1c73 , \7333 );
buf \U$6993 ( \7335 , \7334_nG1c73 );
not \U$6994 ( \7336 , \5932 );
nand \U$6995 ( \7337 , \6165 , \7336 );
xnor \U$6996 ( \7338 , \7337 , \6843 );
buf g1c77 ( \7339_nG1c77 , \7338 );
buf \U$6997 ( \7340 , \7339_nG1c77 );
not \U$6998 ( \7341 , \5897 );
nand \U$6999 ( \7342 , \6163 , \7341 );
xnor \U$7000 ( \7343 , \7342 , \6161 );
buf g1c7b ( \7344_nG1c7b , \7343 );
buf \U$7001 ( \7345 , \7344_nG1c7b );
not \U$7002 ( \7346 , \6131 );
nand \U$7003 ( \7347 , \6158 , \7346 );
xnor \U$7004 ( \7348 , \7347 , \6399 );
buf g1c7f ( \7349_nG1c7f , \7348 );
buf \U$7005 ( \7350 , \7349_nG1c7f );
not \U$7006 ( \7351 , \6127 );
nand \U$7007 ( \7352 , \6156 , \7351 );
xnor \U$7008 ( \7353 , \7352 , \6545 );
buf g1c83 ( \7354_nG1c83 , \7353 );
buf \U$7009 ( \7355 , \7354_nG1c83 );
endmodule

