//
// Conformal-LEC Version 20.10-d005 (29-Apr-2020)
//
module top(RIb4bfa38_65,RIb4c69c8_39,RIa167a08_1,RIb4ca3e8_33,RIa167990_2,RIb4c6c20_34,RIa167918_3,RIb4c6ba8_35,RIa1678a0_4,
        RIb4c6b30_36,RIa167828_5,RIb4c6ab8_37,RIa1677b0_6,RIb4c6a40_38,RIa167738_7,RIa1676c0_8,RIb4c6950_40,RIa167648_9,RIb4c68d8_41,
        RIa1675d0_10,RIb4c6860_42,RIa167558_11,RIb4c67e8_43,RIa1674e0_12,RIb4c6770_44,RIa167468_13,RIb4c3368_45,RIa1673f0_14,RIb4c32f0_46,
        RIa167378_15,RIb4c3278_47,RIa167300_16,RIb4c3200_48,RIa167288_17,RIb4c3188_49,RIa167210_18,RIb4c3110_50,RIa167198_19,RIb4c3098_51,
        RIa167120_20,RIb4c3020_52,RIa1670a8_21,RIb4c2fa8_53,RIa167030_22,RIb4c2f30_54,RIa166fb8_23,RIb4c2eb8_55,RIa166f40_24,RIb4c2e40_56,
        RIa166ec8_25,RIb4c2dc8_57,RIa166e50_26,RIb4c2d50_58,RIa166dd8_27,RIb4c2cd8_59,RIa166d60_28,RIb4c2c60_60,RIa166ce8_29,RIb4c2be8_61,
        RIa166c70_30,RIb4c2b70_62,RIb4ca4d8_31,RIb4c2af8_63,RIb4ca460_32,RIb4bfab0_64,RIb4bf948_67,RIb4bf9c0_66,RIb4bf858_69,RIb4bf8d0_68,
        RIb4bf768_71,RIb4bf7e0_70,RIb4bf6f0_72,RIb4bf678_73,RIb4bf600_74,RIb4bf588_75,RIb4bf510_76,RIb4bf498_77,RIb4bf420_78,RIb4bf3a8_79,
        RIb4bf330_80,RIb4bf2b8_81,RIb4bf240_82,RIb4bf1c8_83,RIb4bf150_84,RIb4bf0d8_85,RIb4bf060_86,RIb4befe8_87,RIb4bef70_88,RIb4beef8_89,
        RIb4bee80_90,RIb4bc1f8_91,RIb4bc180_92,RIb4bc108_93,RIb4bc090_94,RIb4bc018_95,RIb4bbfa0_96,R_61_85b54e8,R_62_85b5590,R_63_85b5638,
        R_64_85b56e0,R_65_85b5788,R_66_85b5830,R_67_85b58d8,R_68_85b5980,R_69_85b5a28,R_6a_85b5ad0,R_6b_85b5b78,R_6c_85b5c20,R_6d_85b5cc8,
        R_6e_85b5d70,R_6f_85b5e18,R_70_85b5ec0,R_71_85b5f68,R_72_85b6010,R_73_85b60b8,R_74_85b6160,R_75_85b6208,R_76_85b62b0,R_77_85b6358,
        R_78_85b6400,R_79_85b64a8,R_7a_85b6550,R_7b_85b65f8,R_7c_85b66a0,R_7d_85b6748,R_7e_85b67f0,R_7f_85b6898,R_80_85b6940,R_81_85b69e8,
        R_82_85b6a90,R_83_85b6b38,R_84_85b6be0,R_85_85b6c88,R_86_85b6d30,R_87_85b6dd8,R_88_85b6e80,R_89_85b6f28,R_8a_85b6fd0,R_8b_85b7078,
        R_8c_85b7120,R_8d_85b71c8,R_8e_85b7270,R_8f_85b7318,R_90_85b73c0,R_91_85b7468,R_92_85b7510,R_93_85b75b8,R_94_85b7660,R_95_85b7708,
        R_96_85b77b0,R_97_85b7858,R_98_85b7900,R_99_85b79a8,R_9a_85b7a50);
input RIb4bfa38_65,RIb4c69c8_39,RIa167a08_1,RIb4ca3e8_33,RIa167990_2,RIb4c6c20_34,RIa167918_3,RIb4c6ba8_35,RIa1678a0_4,
        RIb4c6b30_36,RIa167828_5,RIb4c6ab8_37,RIa1677b0_6,RIb4c6a40_38,RIa167738_7,RIa1676c0_8,RIb4c6950_40,RIa167648_9,RIb4c68d8_41,
        RIa1675d0_10,RIb4c6860_42,RIa167558_11,RIb4c67e8_43,RIa1674e0_12,RIb4c6770_44,RIa167468_13,RIb4c3368_45,RIa1673f0_14,RIb4c32f0_46,
        RIa167378_15,RIb4c3278_47,RIa167300_16,RIb4c3200_48,RIa167288_17,RIb4c3188_49,RIa167210_18,RIb4c3110_50,RIa167198_19,RIb4c3098_51,
        RIa167120_20,RIb4c3020_52,RIa1670a8_21,RIb4c2fa8_53,RIa167030_22,RIb4c2f30_54,RIa166fb8_23,RIb4c2eb8_55,RIa166f40_24,RIb4c2e40_56,
        RIa166ec8_25,RIb4c2dc8_57,RIa166e50_26,RIb4c2d50_58,RIa166dd8_27,RIb4c2cd8_59,RIa166d60_28,RIb4c2c60_60,RIa166ce8_29,RIb4c2be8_61,
        RIa166c70_30,RIb4c2b70_62,RIb4ca4d8_31,RIb4c2af8_63,RIb4ca460_32,RIb4bfab0_64,RIb4bf948_67,RIb4bf9c0_66,RIb4bf858_69,RIb4bf8d0_68,
        RIb4bf768_71,RIb4bf7e0_70,RIb4bf6f0_72,RIb4bf678_73,RIb4bf600_74,RIb4bf588_75,RIb4bf510_76,RIb4bf498_77,RIb4bf420_78,RIb4bf3a8_79,
        RIb4bf330_80,RIb4bf2b8_81,RIb4bf240_82,RIb4bf1c8_83,RIb4bf150_84,RIb4bf0d8_85,RIb4bf060_86,RIb4befe8_87,RIb4bef70_88,RIb4beef8_89,
        RIb4bee80_90,RIb4bc1f8_91,RIb4bc180_92,RIb4bc108_93,RIb4bc090_94,RIb4bc018_95,RIb4bbfa0_96;
output R_61_85b54e8,R_62_85b5590,R_63_85b5638,R_64_85b56e0,R_65_85b5788,R_66_85b5830,R_67_85b58d8,R_68_85b5980,R_69_85b5a28,
        R_6a_85b5ad0,R_6b_85b5b78,R_6c_85b5c20,R_6d_85b5cc8,R_6e_85b5d70,R_6f_85b5e18,R_70_85b5ec0,R_71_85b5f68,R_72_85b6010,R_73_85b60b8,
        R_74_85b6160,R_75_85b6208,R_76_85b62b0,R_77_85b6358,R_78_85b6400,R_79_85b64a8,R_7a_85b6550,R_7b_85b65f8,R_7c_85b66a0,R_7d_85b6748,
        R_7e_85b67f0,R_7f_85b6898,R_80_85b6940,R_81_85b69e8,R_82_85b6a90,R_83_85b6b38,R_84_85b6be0,R_85_85b6c88,R_86_85b6d30,R_87_85b6dd8,
        R_88_85b6e80,R_89_85b6f28,R_8a_85b6fd0,R_8b_85b7078,R_8c_85b7120,R_8d_85b71c8,R_8e_85b7270,R_8f_85b7318,R_90_85b73c0,R_91_85b7468,
        R_92_85b7510,R_93_85b75b8,R_94_85b7660,R_95_85b7708,R_96_85b77b0,R_97_85b7858,R_98_85b7900,R_99_85b79a8,R_9a_85b7a50;

wire \155 , \156_N$1 , \157_ZERO , \158_ONE , \159 , \160 , \161 , \162 , \163 ,
         \164 , \165 , \166 , \167 , \168 , \169 , \170 , \171 , \172 , \173 ,
         \174 , \175 , \176 , \177 , \178 , \179 , \180 , \181 , \182 , \183 ,
         \184 , \185 , \186 , \187 , \188 , \189 , \190 , \191 , \192 , \193 ,
         \194 , \195 , \196 , \197 , \198 , \199 , \200 , \201 , \202 , \203 ,
         \204 , \205 , \206 , \207 , \208 , \209 , \210 , \211 , \212 , \213 ,
         \214 , \215 , \216 , \217 , \218 , \219 , \220 , \221 , \222 , \223 ,
         \224 , \225 , \226 , \227 , \228 , \229 , \230 , \231 , \232 , \233 ,
         \234 , \235 , \236 , \237 , \238 , \239 , \240 , \241 , \242 , \243 ,
         \244 , \245 , \246 , \247 , \248 , \249 , \250 , \251 , \252 , \253 ,
         \254 , \255 , \256 , \257 , \258 , \259 , \260 , \261 , \262 , \263 ,
         \264 , \265 , \266 , \267 , \268 , \269 , \270 , \271 , \272 , \273 ,
         \274 , \275 , \276 , \277 , \278 , \279 , \280 , \281 , \282 , \283 ,
         \284 , \285 , \286 , \287 , \288 , \289_nR13d , \290 , \291_nR13c , \292 , \293 ,
         \294_nR13b , \295 , \296 , \297 , \298 , \299 , \300 , \301 , \302 , \303 ,
         \304 , \305 , \306_nR13f , \307 , \308_nR13e , \309 , \310 , \311 , \312 , \313 ,
         \314 , \315 , \316 , \317 , \318 , \319 , \320 , \321 , \322 , \323 ,
         \324_nR141 , \325 , \326_nR140 , \327 , \328 , \329 , \330 , \331 , \332 , \333 ,
         \334 , \335 , \336 , \337 , \338 , \339 , \340 , \341 , \342 , \343 ,
         \344_nR143 , \345 , \346_nR142 , \347 , \348 , \349 , \350 , \351 , \352 , \353 ,
         \354 , \355 , \356 , \357 , \358 , \359 , \360 , \361 , \362 , \363 ,
         \364 , \365 , \366 , \367 , \368 , \369 , \370 , \371 , \372 , \373 ,
         \374 , \375 , \376 , \377 , \378 , \379 , \380 , \381 , \382 , \383 ,
         \384 , \385 , \386 , \387 , \388 , \389 , \390 , \391 , \392 , \393 ,
         \394 , \395 , \396 , \397 , \398 , \399 , \400 , \401 , \402 , \403 ,
         \404 , \405 , \406 , \407 , \408 , \409 , \410 , \411 , \412 , \413 ,
         \414 , \415 , \416 , \417 , \418 , \419 , \420 , \421 , \422 , \423 ,
         \424 , \425 , \426 , \427 , \428 , \429 , \430 , \431 , \432 , \433 ,
         \434 , \435 , \436 , \437 , \438 , \439 , \440 , \441 , \442 , \443 ,
         \444 , \445 , \446 , \447 , \448 , \449_nR13a , \450 , \451_nR139 , \452 , \453 ,
         \454 , \455 , \456 , \457 , \458 , \459 , \460 , \461 , \462 , \463 ,
         \464 , \465 , \466 , \467 , \468 , \469 , \470 , \471 , \472 , \473 ,
         \474 , \475 , \476 , \477 , \478 , \479 , \480 , \481 , \482 , \483 ,
         \484 , \485 , \486 , \487 , \488 , \489 , \490 , \491 , \492 , \493 ,
         \494 , \495 , \496 , \497 , \498 , \499 , \500 , \501 , \502 , \503 ,
         \504 , \505 , \506 , \507 , \508 , \509 , \510 , \511 , \512 , \513 ,
         \514 , \515 , \516 , \517 , \518 , \519 , \520 , \521 , \522 , \523 ,
         \524 , \525 , \526 , \527 , \528 , \529 , \530 , \531 , \532 , \533 ,
         \534 , \535 , \536 , \537 , \538 , \539 , \540 , \541 , \542 , \543 ,
         \544 , \545 , \546 , \547 , \548 , \549 , \550 , \551 , \552 , \553 ,
         \554 , \555_nR138 , \556 , \557_nR137 , \558 , \559 , \560 , \561 , \562 , \563 ,
         \564 , \565 , \566 , \567 , \568 , \569 , \570 , \571 , \572 , \573 ,
         \574 , \575 , \576 , \577 , \578 , \579 , \580 , \581 , \582 , \583 ,
         \584 , \585 , \586 , \587 , \588 , \589 , \590 , \591 , \592 , \593 ,
         \594 , \595 , \596 , \597 , \598 , \599 , \600 , \601 , \602 , \603 ,
         \604 , \605 , \606 , \607 , \608 , \609 , \610 , \611 , \612 , \613 ,
         \614 , \615 , \616 , \617 , \618 , \619 , \620 , \621 , \622 , \623 ,
         \624 , \625 , \626 , \627 , \628 , \629 , \630 , \631 , \632 , \633 ,
         \634 , \635 , \636 , \637 , \638 , \639 , \640 , \641 , \642 , \643 ,
         \644 , \645 , \646 , \647 , \648 , \649 , \650 , \651 , \652 , \653 ,
         \654 , \655 , \656 , \657 , \658 , \659 , \660 , \661 , \662_nR136 , \663 ,
         \664_nR135 , \665 , \666 , \667 , \668 , \669 , \670 , \671 , \672 , \673 ,
         \674 , \675 , \676 , \677 , \678 , \679 , \680 , \681 , \682 , \683 ,
         \684 , \685 , \686 , \687 , \688 , \689 , \690 , \691 , \692 , \693 ,
         \694 , \695 , \696 , \697 , \698 , \699 , \700 , \701 , \702 , \703 ,
         \704 , \705 , \706 , \707 , \708 , \709 , \710 , \711 , \712 , \713 ,
         \714 , \715 , \716 , \717 , \718 , \719 , \720 , \721 , \722 , \723 ,
         \724 , \725 , \726 , \727 , \728 , \729 , \730 , \731 , \732 , \733 ,
         \734 , \735 , \736 , \737 , \738 , \739 , \740 , \741 , \742 , \743 ,
         \744 , \745 , \746 , \747 , \748 , \749 , \750 , \751 , \752 , \753 ,
         \754 , \755 , \756 , \757 , \758 , \759 , \760 , \761 , \762 , \763 ,
         \764 , \765 , \766 , \767 , \768 , \769 , \770 , \771 , \772 , \773 ,
         \774 , \775 , \776 , \777 , \778 , \779 , \780 , \781 , \782 , \783 ,
         \784 , \785 , \786 , \787 , \788 , \789 , \790 , \791 , \792 , \793 ,
         \794 , \795 , \796 , \797 , \798 , \799 , \800 , \801 , \802 , \803 ,
         \804 , \805 , \806 , \807 , \808 , \809 , \810 , \811 , \812_nR134 , \813 ,
         \814_nR133 , \815 , \816 , \817 , \818 , \819 , \820 , \821 , \822 , \823 ,
         \824 , \825 , \826 , \827 , \828 , \829 , \830 , \831 , \832 , \833 ,
         \834 , \835 , \836 , \837 , \838 , \839 , \840 , \841 , \842 , \843 ,
         \844 , \845 , \846 , \847 , \848 , \849 , \850 , \851 , \852 , \853 ,
         \854 , \855 , \856 , \857 , \858 , \859 , \860 , \861 , \862 , \863 ,
         \864 , \865 , \866 , \867 , \868 , \869 , \870 , \871 , \872 , \873 ,
         \874 , \875 , \876 , \877 , \878 , \879 , \880 , \881 , \882 , \883 ,
         \884 , \885 , \886 , \887 , \888 , \889 , \890 , \891 , \892 , \893 ,
         \894 , \895 , \896 , \897 , \898 , \899 , \900 , \901 , \902 , \903 ,
         \904 , \905 , \906 , \907 , \908 , \909 , \910 , \911 , \912 , \913 ,
         \914 , \915 , \916 , \917 , \918 , \919 , \920 , \921 , \922 , \923 ,
         \924 , \925 , \926 , \927 , \928 , \929 , \930 , \931 , \932 , \933 ,
         \934 , \935 , \936 , \937 , \938 , \939 , \940 , \941 , \942 , \943 ,
         \944 , \945 , \946 , \947 , \948 , \949 , \950 , \951 , \952 , \953 ,
         \954 , \955 , \956 , \957 , \958 , \959 , \960 , \961 , \962 , \963 ,
         \964 , \965 , \966 , \967 , \968 , \969 , \970 , \971 , \972 , \973 ,
         \974 , \975 , \976 , \977 , \978_nR132 , \979 , \980_nR131 , \981 , \982 , \983 ,
         \984 , \985 , \986 , \987 , \988 , \989 , \990 , \991 , \992 , \993 ,
         \994 , \995 , \996 , \997 , \998 , \999 , \1000 , \1001 , \1002 , \1003 ,
         \1004 , \1005 , \1006 , \1007 , \1008 , \1009 , \1010 , \1011 , \1012 , \1013 ,
         \1014 , \1015 , \1016 , \1017 , \1018 , \1019 , \1020 , \1021 , \1022 , \1023 ,
         \1024 , \1025 , \1026 , \1027 , \1028 , \1029 , \1030 , \1031 , \1032 , \1033 ,
         \1034 , \1035 , \1036 , \1037 , \1038 , \1039 , \1040 , \1041 , \1042 , \1043 ,
         \1044 , \1045 , \1046 , \1047 , \1048 , \1049 , \1050 , \1051 , \1052 , \1053 ,
         \1054 , \1055 , \1056 , \1057 , \1058 , \1059 , \1060 , \1061 , \1062 , \1063 ,
         \1064 , \1065 , \1066 , \1067 , \1068 , \1069 , \1070 , \1071 , \1072 , \1073 ,
         \1074 , \1075 , \1076 , \1077 , \1078 , \1079 , \1080 , \1081 , \1082 , \1083 ,
         \1084 , \1085 , \1086 , \1087 , \1088 , \1089 , \1090 , \1091 , \1092 , \1093 ,
         \1094 , \1095 , \1096 , \1097 , \1098 , \1099 , \1100 , \1101 , \1102 , \1103 ,
         \1104 , \1105 , \1106 , \1107 , \1108 , \1109 , \1110 , \1111 , \1112 , \1113 ,
         \1114 , \1115 , \1116 , \1117 , \1118 , \1119 , \1120 , \1121 , \1122 , \1123 ,
         \1124 , \1125 , \1126 , \1127 , \1128 , \1129 , \1130 , \1131 , \1132 , \1133 ,
         \1134 , \1135 , \1136 , \1137 , \1138 , \1139 , \1140 , \1141 , \1142 , \1143 ,
         \1144 , \1145 , \1146 , \1147 , \1148 , \1149 , \1150 , \1151 , \1152 , \1153 ,
         \1154 , \1155 , \1156 , \1157 , \1158 , \1159 , \1160 , \1161 , \1162 , \1163 ,
         \1164 , \1165 , \1166 , \1167 , \1168 , \1169 , \1170 , \1171_nR130 , \1172 , \1173_nR12f ,
         \1174 , \1175 , \1176 , \1177 , \1178 , \1179 , \1180 , \1181 , \1182 , \1183 ,
         \1184 , \1185 , \1186 , \1187 , \1188 , \1189 , \1190 , \1191 , \1192 , \1193 ,
         \1194 , \1195 , \1196 , \1197 , \1198 , \1199 , \1200 , \1201 , \1202 , \1203 ,
         \1204 , \1205 , \1206 , \1207 , \1208 , \1209 , \1210 , \1211 , \1212 , \1213 ,
         \1214 , \1215 , \1216 , \1217 , \1218 , \1219 , \1220 , \1221 , \1222 , \1223 ,
         \1224 , \1225 , \1226 , \1227 , \1228 , \1229 , \1230 , \1231 , \1232 , \1233 ,
         \1234 , \1235 , \1236 , \1237 , \1238 , \1239 , \1240 , \1241 , \1242 , \1243 ,
         \1244 , \1245 , \1246 , \1247 , \1248 , \1249 , \1250 , \1251 , \1252 , \1253 ,
         \1254 , \1255 , \1256 , \1257 , \1258 , \1259 , \1260 , \1261 , \1262 , \1263 ,
         \1264 , \1265 , \1266 , \1267 , \1268 , \1269 , \1270 , \1271 , \1272 , \1273 ,
         \1274 , \1275 , \1276 , \1277 , \1278 , \1279 , \1280 , \1281 , \1282 , \1283 ,
         \1284 , \1285 , \1286 , \1287 , \1288 , \1289 , \1290 , \1291 , \1292 , \1293 ,
         \1294 , \1295 , \1296 , \1297 , \1298 , \1299 , \1300 , \1301 , \1302 , \1303 ,
         \1304 , \1305 , \1306 , \1307 , \1308 , \1309 , \1310 , \1311 , \1312 , \1313 ,
         \1314 , \1315 , \1316 , \1317 , \1318 , \1319 , \1320 , \1321 , \1322 , \1323 ,
         \1324 , \1325 , \1326 , \1327 , \1328 , \1329 , \1330 , \1331 , \1332 , \1333 ,
         \1334 , \1335 , \1336 , \1337 , \1338 , \1339 , \1340 , \1341 , \1342 , \1343 ,
         \1344 , \1345 , \1346 , \1347 , \1348 , \1349 , \1350 , \1351 , \1352 , \1353 ,
         \1354 , \1355 , \1356 , \1357_nR12e , \1358 , \1359_nR12d , \1360 , \1361 , \1362 , \1363 ,
         \1364 , \1365 , \1366 , \1367 , \1368 , \1369 , \1370 , \1371 , \1372 , \1373 ,
         \1374 , \1375 , \1376 , \1377 , \1378 , \1379 , \1380 , \1381 , \1382 , \1383 ,
         \1384 , \1385 , \1386 , \1387 , \1388 , \1389 , \1390 , \1391 , \1392 , \1393 ,
         \1394 , \1395 , \1396 , \1397 , \1398 , \1399 , \1400 , \1401 , \1402 , \1403 ,
         \1404 , \1405 , \1406 , \1407 , \1408 , \1409 , \1410 , \1411 , \1412 , \1413 ,
         \1414 , \1415 , \1416 , \1417 , \1418 , \1419 , \1420 , \1421 , \1422 , \1423 ,
         \1424 , \1425 , \1426 , \1427 , \1428 , \1429 , \1430 , \1431 , \1432 , \1433 ,
         \1434 , \1435 , \1436 , \1437 , \1438 , \1439 , \1440 , \1441 , \1442 , \1443 ,
         \1444 , \1445 , \1446 , \1447 , \1448 , \1449 , \1450 , \1451 , \1452 , \1453 ,
         \1454 , \1455 , \1456 , \1457 , \1458 , \1459 , \1460 , \1461 , \1462 , \1463 ,
         \1464 , \1465 , \1466 , \1467 , \1468 , \1469 , \1470 , \1471 , \1472 , \1473 ,
         \1474 , \1475 , \1476 , \1477 , \1478 , \1479 , \1480 , \1481 , \1482 , \1483 ,
         \1484 , \1485 , \1486 , \1487 , \1488 , \1489 , \1490 , \1491 , \1492 , \1493 ,
         \1494 , \1495 , \1496 , \1497 , \1498 , \1499 , \1500 , \1501 , \1502 , \1503 ,
         \1504 , \1505 , \1506 , \1507 , \1508 , \1509 , \1510 , \1511 , \1512 , \1513 ,
         \1514 , \1515 , \1516 , \1517 , \1518 , \1519 , \1520 , \1521 , \1522 , \1523 ,
         \1524 , \1525 , \1526 , \1527 , \1528 , \1529 , \1530 , \1531 , \1532 , \1533 ,
         \1534 , \1535 , \1536 , \1537 , \1538 , \1539 , \1540 , \1541 , \1542 , \1543 ,
         \1544 , \1545 , \1546 , \1547 , \1548 , \1549 , \1550 , \1551 , \1552 , \1553 ,
         \1554 , \1555 , \1556 , \1557 , \1558 , \1559 , \1560 , \1561 , \1562 , \1563 ,
         \1564 , \1565 , \1566 , \1567 , \1568 , \1569 , \1570 , \1571 , \1572 , \1573 ,
         \1574 , \1575 , \1576 , \1577 , \1578 , \1579 , \1580 , \1581 , \1582 , \1583 ,
         \1584 , \1585 , \1586 , \1587 , \1588 , \1589 , \1590 , \1591 , \1592 , \1593 ,
         \1594 , \1595 , \1596 , \1597 , \1598 , \1599 , \1600 , \1601 , \1602 , \1603 ,
         \1604_nR12c , \1605 , \1606_nR12b , \1607 , \1608 , \1609 , \1610 , \1611 , \1612 , \1613 ,
         \1614 , \1615 , \1616 , \1617 , \1618 , \1619 , \1620 , \1621 , \1622 , \1623 ,
         \1624 , \1625 , \1626 , \1627 , \1628 , \1629 , \1630 , \1631 , \1632 , \1633 ,
         \1634 , \1635 , \1636 , \1637 , \1638 , \1639 , \1640 , \1641 , \1642 , \1643 ,
         \1644 , \1645 , \1646 , \1647 , \1648 , \1649 , \1650 , \1651 , \1652 , \1653 ,
         \1654 , \1655 , \1656 , \1657 , \1658 , \1659 , \1660 , \1661 , \1662 , \1663 ,
         \1664 , \1665 , \1666 , \1667 , \1668 , \1669 , \1670 , \1671 , \1672 , \1673 ,
         \1674 , \1675 , \1676 , \1677 , \1678 , \1679 , \1680 , \1681 , \1682 , \1683 ,
         \1684 , \1685 , \1686 , \1687 , \1688 , \1689 , \1690 , \1691 , \1692 , \1693 ,
         \1694 , \1695 , \1696 , \1697 , \1698 , \1699 , \1700 , \1701 , \1702 , \1703 ,
         \1704 , \1705 , \1706 , \1707 , \1708 , \1709 , \1710 , \1711 , \1712 , \1713 ,
         \1714 , \1715 , \1716 , \1717 , \1718 , \1719 , \1720 , \1721 , \1722 , \1723 ,
         \1724 , \1725 , \1726 , \1727 , \1728 , \1729 , \1730 , \1731 , \1732 , \1733 ,
         \1734 , \1735 , \1736 , \1737 , \1738 , \1739 , \1740 , \1741 , \1742 , \1743 ,
         \1744 , \1745 , \1746 , \1747 , \1748 , \1749 , \1750 , \1751 , \1752 , \1753 ,
         \1754 , \1755 , \1756 , \1757 , \1758 , \1759 , \1760 , \1761 , \1762 , \1763 ,
         \1764 , \1765 , \1766 , \1767 , \1768 , \1769 , \1770 , \1771 , \1772 , \1773 ,
         \1774 , \1775 , \1776 , \1777 , \1778 , \1779 , \1780 , \1781 , \1782 , \1783 ,
         \1784 , \1785 , \1786 , \1787 , \1788 , \1789 , \1790 , \1791 , \1792 , \1793 ,
         \1794 , \1795 , \1796 , \1797 , \1798 , \1799 , \1800 , \1801 , \1802 , \1803 ,
         \1804 , \1805 , \1806 , \1807 , \1808 , \1809 , \1810 , \1811 , \1812 , \1813 ,
         \1814 , \1815 , \1816 , \1817 , \1818 , \1819 , \1820 , \1821 , \1822 , \1823 ,
         \1824 , \1825 , \1826 , \1827 , \1828 , \1829_nR12a , \1830 , \1831_nR129 , \1832 , \1833 ,
         \1834 , \1835 , \1836 , \1837 , \1838 , \1839 , \1840 , \1841 , \1842 , \1843 ,
         \1844 , \1845 , \1846 , \1847 , \1848 , \1849 , \1850 , \1851 , \1852 , \1853 ,
         \1854 , \1855 , \1856 , \1857 , \1858 , \1859 , \1860 , \1861 , \1862 , \1863 ,
         \1864 , \1865 , \1866 , \1867 , \1868 , \1869 , \1870 , \1871 , \1872 , \1873 ,
         \1874 , \1875 , \1876 , \1877 , \1878 , \1879 , \1880 , \1881 , \1882 , \1883 ,
         \1884 , \1885 , \1886 , \1887 , \1888 , \1889 , \1890 , \1891 , \1892 , \1893 ,
         \1894 , \1895 , \1896 , \1897 , \1898 , \1899 , \1900 , \1901 , \1902 , \1903 ,
         \1904 , \1905 , \1906 , \1907 , \1908 , \1909 , \1910 , \1911 , \1912 , \1913 ,
         \1914 , \1915 , \1916 , \1917 , \1918 , \1919 , \1920 , \1921 , \1922 , \1923 ,
         \1924 , \1925 , \1926 , \1927 , \1928 , \1929 , \1930 , \1931 , \1932 , \1933 ,
         \1934 , \1935 , \1936 , \1937 , \1938 , \1939 , \1940 , \1941 , \1942 , \1943 ,
         \1944 , \1945 , \1946 , \1947 , \1948 , \1949 , \1950 , \1951 , \1952 , \1953 ,
         \1954 , \1955 , \1956 , \1957 , \1958 , \1959 , \1960 , \1961 , \1962 , \1963 ,
         \1964 , \1965 , \1966 , \1967 , \1968 , \1969 , \1970 , \1971 , \1972 , \1973 ,
         \1974 , \1975 , \1976 , \1977 , \1978 , \1979 , \1980 , \1981 , \1982 , \1983 ,
         \1984 , \1985 , \1986 , \1987 , \1988 , \1989 , \1990 , \1991 , \1992 , \1993 ,
         \1994 , \1995 , \1996 , \1997 , \1998 , \1999 , \2000 , \2001 , \2002 , \2003 ,
         \2004 , \2005 , \2006 , \2007 , \2008 , \2009 , \2010 , \2011 , \2012 , \2013 ,
         \2014 , \2015 , \2016 , \2017 , \2018 , \2019 , \2020 , \2021 , \2022 , \2023 ,
         \2024 , \2025 , \2026 , \2027 , \2028 , \2029 , \2030 , \2031 , \2032 , \2033 ,
         \2034 , \2035 , \2036 , \2037 , \2038 , \2039 , \2040 , \2041 , \2042 , \2043 ,
         \2044 , \2045 , \2046 , \2047 , \2048 , \2049 , \2050 , \2051 , \2052 , \2053 ,
         \2054 , \2055 , \2056 , \2057 , \2058 , \2059 , \2060 , \2061 , \2062 , \2063 ,
         \2064 , \2065 , \2066 , \2067 , \2068 , \2069 , \2070 , \2071 , \2072 , \2073 ,
         \2074 , \2075 , \2076 , \2077 , \2078 , \2079 , \2080 , \2081 , \2082 , \2083 ,
         \2084 , \2085 , \2086 , \2087 , \2088 , \2089 , \2090 , \2091 , \2092 , \2093 ,
         \2094 , \2095 , \2096 , \2097 , \2098 , \2099 , \2100 , \2101 , \2102 , \2103 ,
         \2104 , \2105 , \2106 , \2107 , \2108 , \2109 , \2110 , \2111 , \2112 , \2113 ,
         \2114 , \2115 , \2116 , \2117 , \2118_nR128 , \2119 , \2120_nR127 , \2121 , \2122 , \2123 ,
         \2124 , \2125 , \2126 , \2127 , \2128 , \2129 , \2130 , \2131 , \2132 , \2133 ,
         \2134 , \2135 , \2136 , \2137 , \2138 , \2139 , \2140 , \2141 , \2142 , \2143 ,
         \2144 , \2145 , \2146 , \2147 , \2148 , \2149 , \2150 , \2151 , \2152 , \2153 ,
         \2154 , \2155 , \2156 , \2157 , \2158 , \2159 , \2160 , \2161 , \2162 , \2163 ,
         \2164 , \2165 , \2166 , \2167 , \2168 , \2169 , \2170 , \2171 , \2172 , \2173 ,
         \2174 , \2175 , \2176 , \2177 , \2178 , \2179 , \2180 , \2181 , \2182 , \2183 ,
         \2184 , \2185 , \2186 , \2187 , \2188 , \2189 , \2190 , \2191 , \2192 , \2193 ,
         \2194 , \2195 , \2196 , \2197 , \2198 , \2199 , \2200 , \2201 , \2202 , \2203 ,
         \2204 , \2205 , \2206 , \2207 , \2208 , \2209 , \2210 , \2211 , \2212 , \2213 ,
         \2214 , \2215 , \2216 , \2217 , \2218 , \2219 , \2220 , \2221 , \2222 , \2223 ,
         \2224 , \2225 , \2226 , \2227 , \2228 , \2229 , \2230 , \2231 , \2232 , \2233 ,
         \2234 , \2235 , \2236 , \2237 , \2238 , \2239 , \2240 , \2241 , \2242 , \2243 ,
         \2244 , \2245 , \2246 , \2247 , \2248 , \2249 , \2250 , \2251 , \2252 , \2253 ,
         \2254 , \2255 , \2256 , \2257 , \2258 , \2259 , \2260 , \2261 , \2262 , \2263 ,
         \2264 , \2265 , \2266 , \2267 , \2268 , \2269 , \2270 , \2271 , \2272 , \2273 ,
         \2274 , \2275 , \2276 , \2277 , \2278 , \2279 , \2280 , \2281 , \2282 , \2283 ,
         \2284 , \2285 , \2286 , \2287 , \2288 , \2289 , \2290 , \2291 , \2292 , \2293 ,
         \2294 , \2295 , \2296 , \2297 , \2298 , \2299 , \2300 , \2301 , \2302 , \2303 ,
         \2304 , \2305 , \2306 , \2307 , \2308 , \2309 , \2310 , \2311 , \2312 , \2313 ,
         \2314 , \2315 , \2316 , \2317 , \2318 , \2319 , \2320 , \2321 , \2322 , \2323 ,
         \2324 , \2325 , \2326 , \2327 , \2328 , \2329 , \2330 , \2331 , \2332 , \2333 ,
         \2334 , \2335 , \2336 , \2337 , \2338 , \2339 , \2340 , \2341 , \2342 , \2343 ,
         \2344 , \2345 , \2346 , \2347 , \2348 , \2349 , \2350 , \2351 , \2352 , \2353 ,
         \2354 , \2355 , \2356 , \2357 , \2358 , \2359 , \2360 , \2361 , \2362 , \2363 ,
         \2364 , \2365 , \2366 , \2367 , \2368_nR126 , \2369 , \2370_nR125 , \2371 , \2372 , \2373 ,
         \2374 , \2375 , \2376 , \2377 , \2378 , \2379 , \2380 , \2381 , \2382 , \2383 ,
         \2384 , \2385 , \2386 , \2387 , \2388 , \2389 , \2390 , \2391 , \2392 , \2393 ,
         \2394 , \2395 , \2396 , \2397 , \2398 , \2399 , \2400 , \2401 , \2402 , \2403 ,
         \2404 , \2405 , \2406 , \2407 , \2408 , \2409 , \2410 , \2411 , \2412 , \2413 ,
         \2414 , \2415 , \2416 , \2417 , \2418 , \2419 , \2420 , \2421 , \2422 , \2423 ,
         \2424 , \2425 , \2426 , \2427 , \2428 , \2429 , \2430 , \2431 , \2432 , \2433 ,
         \2434 , \2435 , \2436 , \2437 , \2438 , \2439 , \2440 , \2441 , \2442 , \2443 ,
         \2444 , \2445 , \2446 , \2447 , \2448 , \2449 , \2450 , \2451 , \2452 , \2453 ,
         \2454 , \2455 , \2456 , \2457 , \2458 , \2459 , \2460 , \2461 , \2462 , \2463 ,
         \2464 , \2465 , \2466 , \2467 , \2468 , \2469 , \2470 , \2471 , \2472 , \2473 ,
         \2474 , \2475 , \2476 , \2477 , \2478 , \2479 , \2480 , \2481 , \2482 , \2483 ,
         \2484 , \2485 , \2486 , \2487 , \2488 , \2489 , \2490 , \2491 , \2492 , \2493 ,
         \2494 , \2495 , \2496 , \2497 , \2498 , \2499 , \2500 , \2501 , \2502 , \2503 ,
         \2504 , \2505 , \2506 , \2507 , \2508 , \2509 , \2510 , \2511 , \2512 , \2513 ,
         \2514 , \2515 , \2516 , \2517 , \2518 , \2519 , \2520 , \2521 , \2522 , \2523 ,
         \2524 , \2525 , \2526 , \2527 , \2528 , \2529 , \2530 , \2531 , \2532 , \2533 ,
         \2534 , \2535 , \2536 , \2537 , \2538 , \2539 , \2540 , \2541 , \2542 , \2543 ,
         \2544 , \2545 , \2546 , \2547 , \2548 , \2549 , \2550 , \2551 , \2552 , \2553 ,
         \2554 , \2555 , \2556 , \2557 , \2558 , \2559 , \2560 , \2561 , \2562 , \2563 ,
         \2564 , \2565 , \2566 , \2567 , \2568 , \2569 , \2570 , \2571 , \2572 , \2573 ,
         \2574 , \2575 , \2576 , \2577 , \2578 , \2579 , \2580 , \2581 , \2582 , \2583 ,
         \2584 , \2585 , \2586 , \2587 , \2588 , \2589 , \2590 , \2591 , \2592 , \2593 ,
         \2594 , \2595 , \2596 , \2597 , \2598 , \2599 , \2600 , \2601 , \2602 , \2603 ,
         \2604 , \2605 , \2606 , \2607 , \2608 , \2609 , \2610 , \2611 , \2612 , \2613 ,
         \2614 , \2615 , \2616 , \2617 , \2618 , \2619 , \2620 , \2621 , \2622 , \2623 ,
         \2624 , \2625 , \2626 , \2627 , \2628 , \2629 , \2630 , \2631 , \2632 , \2633 ,
         \2634 , \2635 , \2636 , \2637 , \2638 , \2639 , \2640 , \2641 , \2642 , \2643 ,
         \2644 , \2645 , \2646 , \2647 , \2648 , \2649 , \2650 , \2651 , \2652 , \2653 ,
         \2654 , \2655 , \2656 , \2657 , \2658 , \2659 , \2660 , \2661 , \2662 , \2663 ,
         \2664 , \2665 , \2666 , \2667 , \2668 , \2669 , \2670 , \2671 , \2672 , \2673 ,
         \2674 , \2675 , \2676 , \2677 , \2678 , \2679 , \2680 , \2681 , \2682 , \2683 ,
         \2684 , \2685 , \2686 , \2687 , \2688 , \2689 , \2690 , \2691 , \2692 , \2693 ,
         \2694 , \2695 , \2696 , \2697 , \2698 , \2699 , \2700 , \2701 , \2702 , \2703 ,
         \2704 , \2705 , \2706 , \2707 , \2708 , \2709 , \2710 , \2711 , \2712 , \2713 ,
         \2714 , \2715 , \2716 , \2717 , \2718 , \2719 , \2720 , \2721 , \2722 , \2723 ,
         \2724 , \2725 , \2726 , \2727 , \2728 , \2729 , \2730 , \2731 , \2732 , \2733 ,
         \2734 , \2735 , \2736 , \2737 , \2738 , \2739 , \2740 , \2741 , \2742 , \2743 ,
         \2744 , \2745 , \2746 , \2747 , \2748 , \2749 , \2750 , \2751 , \2752 , \2753 ,
         \2754 , \2755 , \2756 , \2757 , \2758 , \2759 , \2760 , \2761 , \2762 , \2763 ,
         \2764 , \2765 , \2766 , \2767 , \2768 , \2769 , \2770 , \2771 , \2772 , \2773 ,
         \2774 , \2775 , \2776 , \2777 , \2778 , \2779 , \2780 , \2781 , \2782 , \2783 ,
         \2784 , \2785 , \2786 , \2787 , \2788 , \2789 , \2790 , \2791 , \2792 , \2793 ,
         \2794 , \2795 , \2796 , \2797 , \2798 , \2799 , \2800 , \2801 , \2802 , \2803 ,
         \2804 , \2805 , \2806 , \2807 , \2808 , \2809 , \2810 , \2811 , \2812 , \2813 ,
         \2814 , \2815 , \2816 , \2817 , \2818 , \2819 , \2820 , \2821 , \2822 , \2823 ,
         \2824 , \2825 , \2826 , \2827 , \2828 , \2829 , \2830 , \2831 , \2832 , \2833 ,
         \2834 , \2835 , \2836 , \2837 , \2838 , \2839 , \2840 , \2841 , \2842 , \2843 ,
         \2844 , \2845 , \2846 , \2847 , \2848 , \2849 , \2850 , \2851 , \2852 , \2853 ,
         \2854 , \2855 , \2856 , \2857 , \2858 , \2859 , \2860 , \2861 , \2862 , \2863 ,
         \2864 , \2865 , \2866 , \2867 , \2868 , \2869 , \2870 , \2871 , \2872 , \2873 ,
         \2874 , \2875 , \2876 , \2877 , \2878 , \2879 , \2880 , \2881 , \2882 , \2883 ,
         \2884 , \2885 , \2886 , \2887 , \2888 , \2889 , \2890 , \2891 , \2892 , \2893 ,
         \2894 , \2895 , \2896 , \2897 , \2898 , \2899 , \2900 , \2901 , \2902 , \2903 ,
         \2904 , \2905 , \2906 , \2907 , \2908 , \2909_nR123 , \2910 , \2911 , \2912 , \2913 ,
         \2914 , \2915 , \2916 , \2917 , \2918 , \2919 , \2920 , \2921 , \2922 , \2923 ,
         \2924 , \2925 , \2926 , \2927 , \2928 , \2929 , \2930 , \2931 , \2932 , \2933 ,
         \2934 , \2935 , \2936 , \2937 , \2938 , \2939 , \2940 , \2941 , \2942 , \2943 ,
         \2944 , \2945 , \2946 , \2947 , \2948 , \2949 , \2950 , \2951 , \2952 , \2953 ,
         \2954 , \2955 , \2956 , \2957 , \2958 , \2959 , \2960 , \2961 , \2962 , \2963 ,
         \2964 , \2965 , \2966 , \2967 , \2968 , \2969 , \2970 , \2971 , \2972 , \2973 ,
         \2974 , \2975 , \2976 , \2977 , \2978 , \2979 , \2980 , \2981 , \2982 , \2983 ,
         \2984 , \2985 , \2986 , \2987 , \2988 , \2989 , \2990 , \2991 , \2992 , \2993 ,
         \2994 , \2995 , \2996 , \2997 , \2998 , \2999 , \3000 , \3001 , \3002 , \3003 ,
         \3004 , \3005 , \3006 , \3007 , \3008 , \3009 , \3010 , \3011 , \3012 , \3013 ,
         \3014 , \3015 , \3016 , \3017 , \3018 , \3019 , \3020 , \3021 , \3022 , \3023 ,
         \3024 , \3025 , \3026 , \3027 , \3028 , \3029 , \3030 , \3031 , \3032 , \3033 ,
         \3034 , \3035 , \3036 , \3037 , \3038 , \3039 , \3040 , \3041 , \3042 , \3043 ,
         \3044 , \3045 , \3046 , \3047 , \3048 , \3049 , \3050 , \3051 , \3052 , \3053 ,
         \3054 , \3055 , \3056 , \3057 , \3058 , \3059 , \3060 , \3061 , \3062 , \3063 ,
         \3064 , \3065 , \3066 , \3067 , \3068 , \3069 , \3070 , \3071 , \3072 , \3073 ,
         \3074 , \3075 , \3076 , \3077 , \3078 , \3079 , \3080 , \3081 , \3082 , \3083 ,
         \3084 , \3085 , \3086 , \3087 , \3088 , \3089 , \3090 , \3091 , \3092 , \3093 ,
         \3094 , \3095 , \3096 , \3097 , \3098 , \3099 , \3100 , \3101 , \3102 , \3103 ,
         \3104 , \3105 , \3106 , \3107 , \3108 , \3109 , \3110 , \3111 , \3112 , \3113 ,
         \3114 , \3115 , \3116 , \3117 , \3118 , \3119 , \3120 , \3121 , \3122 , \3123 ,
         \3124 , \3125 , \3126 , \3127 , \3128 , \3129 , \3130 , \3131 , \3132 , \3133 ,
         \3134 , \3135 , \3136 , \3137 , \3138 , \3139 , \3140 , \3141 , \3142 , \3143 ,
         \3144 , \3145 , \3146 , \3147 , \3148 , \3149 , \3150 , \3151 , \3152 , \3153 ,
         \3154 , \3155 , \3156 , \3157 , \3158 , \3159 , \3160 , \3161 , \3162 , \3163 ,
         \3164 , \3165 , \3166 , \3167 , \3168 , \3169 , \3170 , \3171 , \3172 , \3173 ,
         \3174 , \3175 , \3176 , \3177 , \3178 , \3179 , \3180 , \3181 , \3182 , \3183 ,
         \3184 , \3185 , \3186 , \3187 , \3188 , \3189 , \3190 , \3191 , \3192 , \3193 ,
         \3194 , \3195 , \3196 , \3197 , \3198 , \3199 , \3200 , \3201 , \3202 , \3203 ,
         \3204 , \3205 , \3206 , \3207 , \3208 , \3209 , \3210 , \3211 , \3212 , \3213 ,
         \3214 , \3215 , \3216 , \3217 , \3218 , \3219 , \3220 , \3221 , \3222 , \3223 ,
         \3224 , \3225 , \3226 , \3227 , \3228 , \3229 , \3230 , \3231 , \3232 , \3233 ,
         \3234 , \3235 , \3236 , \3237 , \3238 , \3239 , \3240 , \3241 , \3242 , \3243 ,
         \3244 , \3245 , \3246 , \3247 , \3248 , \3249 , \3250 , \3251 , \3252 , \3253 ,
         \3254 , \3255 , \3256 , \3257 , \3258 , \3259 , \3260 , \3261 , \3262 , \3263 ,
         \3264 , \3265 , \3266 , \3267 , \3268 , \3269 , \3270 , \3271 , \3272 , \3273 ,
         \3274 , \3275 , \3276 , \3277 , \3278 , \3279 , \3280 , \3281 , \3282 , \3283 ,
         \3284 , \3285 , \3286 , \3287 , \3288 , \3289 , \3290 , \3291 , \3292 , \3293 ,
         \3294 , \3295 , \3296 , \3297 , \3298 , \3299 , \3300 , \3301 , \3302 , \3303 ,
         \3304 , \3305 , \3306 , \3307 , \3308 , \3309 , \3310 , \3311 , \3312 , \3313 ,
         \3314 , \3315 , \3316 , \3317 , \3318 , \3319 , \3320 , \3321 , \3322 , \3323 ,
         \3324 , \3325 , \3326 , \3327 , \3328 , \3329 , \3330 , \3331 , \3332 , \3333 ,
         \3334 , \3335 , \3336 , \3337 , \3338 , \3339 , \3340 , \3341 , \3342 , \3343 ,
         \3344 , \3345 , \3346 , \3347 , \3348 , \3349 , \3350 , \3351 , \3352 , \3353 ,
         \3354 , \3355 , \3356 , \3357 , \3358 , \3359 , \3360 , \3361 , \3362 , \3363 ,
         \3364 , \3365 , \3366 , \3367 , \3368 , \3369 , \3370 , \3371 , \3372 , \3373 ,
         \3374 , \3375 , \3376 , \3377 , \3378 , \3379 , \3380 , \3381 , \3382 , \3383 ,
         \3384 , \3385 , \3386 , \3387 , \3388 , \3389 , \3390 , \3391 , \3392 , \3393 ,
         \3394 , \3395 , \3396 , \3397 , \3398 , \3399 , \3400 , \3401 , \3402 , \3403 ,
         \3404 , \3405 , \3406 , \3407 , \3408 , \3409 , \3410 , \3411 , \3412 , \3413 ,
         \3414 , \3415 , \3416 , \3417 , \3418 , \3419 , \3420 , \3421 , \3422 , \3423 ,
         \3424 , \3425 , \3426 , \3427 , \3428 , \3429 , \3430 , \3431 , \3432 , \3433 ,
         \3434 , \3435 , \3436 , \3437 , \3438 , \3439 , \3440 , \3441 , \3442 , \3443 ,
         \3444 , \3445 , \3446 , \3447 , \3448 , \3449 , \3450 , \3451 , \3452 , \3453 ,
         \3454 , \3455 , \3456 , \3457 , \3458 , \3459 , \3460 , \3461 , \3462 , \3463 ,
         \3464 , \3465 , \3466 , \3467 , \3468 , \3469 , \3470 , \3471 , \3472 , \3473 ,
         \3474 , \3475 , \3476 , \3477 , \3478 , \3479 , \3480 , \3481 , \3482 , \3483 ,
         \3484 , \3485 , \3486 , \3487 , \3488 , \3489 , \3490 , \3491 , \3492 , \3493 ,
         \3494 , \3495 , \3496 , \3497 , \3498 , \3499 , \3500 , \3501 , \3502 , \3503 ,
         \3504 , \3505 , \3506 , \3507 , \3508 , \3509 , \3510 , \3511 , \3512 , \3513 ,
         \3514 , \3515 , \3516 , \3517 , \3518 , \3519 , \3520 , \3521 , \3522 , \3523 ,
         \3524 , \3525 , \3526 , \3527 , \3528 , \3529 , \3530 , \3531 , \3532 , \3533 ,
         \3534 , \3535 , \3536 , \3537 , \3538 , \3539 , \3540 , \3541 , \3542 , \3543 ,
         \3544 , \3545 , \3546 , \3547 , \3548 , \3549 , \3550 , \3551 , \3552 , \3553 ,
         \3554 , \3555 , \3556 , \3557 , \3558 , \3559 , \3560 , \3561 , \3562 , \3563 ,
         \3564 , \3565 , \3566 , \3567 , \3568 , \3569 , \3570 , \3571 , \3572 , \3573 ,
         \3574 , \3575 , \3576 , \3577 , \3578 , \3579 , \3580 , \3581 , \3582 , \3583 ,
         \3584 , \3585 , \3586 , \3587 , \3588 , \3589 , \3590 , \3591 , \3592 , \3593 ,
         \3594 , \3595 , \3596 , \3597 , \3598 , \3599 , \3600 , \3601 , \3602 , \3603 ,
         \3604 , \3605 , \3606 , \3607 , \3608 , \3609 , \3610 , \3611 , \3612 , \3613 ,
         \3614 , \3615 , \3616 , \3617 , \3618 , \3619 , \3620 , \3621 , \3622 , \3623 ,
         \3624 , \3625 , \3626 , \3627 , \3628 , \3629 , \3630 , \3631 , \3632 , \3633 ,
         \3634 , \3635 , \3636 , \3637 , \3638 , \3639 , \3640 , \3641 , \3642 , \3643 ,
         \3644 , \3645 , \3646 , \3647 , \3648 , \3649 , \3650 , \3651 , \3652 , \3653 ,
         \3654 , \3655 , \3656 , \3657 , \3658 , \3659 , \3660 , \3661 , \3662 , \3663 ,
         \3664 , \3665 , \3666 , \3667 , \3668 , \3669 , \3670 , \3671 , \3672 , \3673 ,
         \3674 , \3675 , \3676 , \3677 , \3678 , \3679 , \3680 , \3681 , \3682 , \3683 ,
         \3684 , \3685 , \3686 , \3687 , \3688 , \3689 , \3690 , \3691 , \3692 , \3693 ,
         \3694 , \3695 , \3696 , \3697 , \3698 , \3699 , \3700 , \3701 , \3702 , \3703 ,
         \3704 , \3705 , \3706 , \3707 , \3708 , \3709 , \3710 , \3711 , \3712 , \3713 ,
         \3714 , \3715 , \3716 , \3717 , \3718 , \3719 , \3720 , \3721 , \3722 , \3723 ,
         \3724 , \3725 , \3726 , \3727 , \3728 , \3729 , \3730 , \3731 , \3732 , \3733 ,
         \3734 , \3735 , \3736 , \3737 , \3738 , \3739 , \3740 , \3741 , \3742 , \3743 ,
         \3744 , \3745 , \3746 , \3747 , \3748 , \3749 , \3750 , \3751 , \3752 , \3753 ,
         \3754 , \3755 , \3756 , \3757 , \3758 , \3759 , \3760 , \3761 , \3762 , \3763 ,
         \3764 , \3765 , \3766 , \3767 , \3768 , \3769 , \3770 , \3771 , \3772 , \3773 ,
         \3774 , \3775 , \3776 , \3777 , \3778 , \3779 , \3780 , \3781 , \3782 , \3783 ,
         \3784 , \3785 , \3786 , \3787 , \3788 , \3789 , \3790 , \3791 , \3792 , \3793 ,
         \3794 , \3795 , \3796 , \3797 , \3798 , \3799 , \3800 , \3801 , \3802 , \3803 ,
         \3804 , \3805 , \3806 , \3807 , \3808 , \3809 , \3810 , \3811 , \3812 , \3813 ,
         \3814 , \3815 , \3816 , \3817 , \3818 , \3819 , \3820 , \3821 , \3822 , \3823 ,
         \3824 , \3825 , \3826 , \3827 , \3828 , \3829 , \3830 , \3831 , \3832 , \3833 ,
         \3834 , \3835 , \3836 , \3837 , \3838 , \3839 , \3840 , \3841 , \3842 , \3843 ,
         \3844 , \3845 , \3846 , \3847 , \3848 , \3849 , \3850 , \3851 , \3852 , \3853 ,
         \3854 , \3855 , \3856 , \3857 , \3858 , \3859 , \3860 , \3861 , \3862 , \3863 ,
         \3864 , \3865 , \3866 , \3867 , \3868 , \3869 , \3870 , \3871 , \3872 , \3873 ,
         \3874 , \3875 , \3876 , \3877 , \3878 , \3879 , \3880 , \3881 , \3882 , \3883 ,
         \3884 , \3885 , \3886 , \3887 , \3888 , \3889 , \3890 , \3891 , \3892 , \3893 ,
         \3894 , \3895 , \3896 , \3897 , \3898 , \3899 , \3900 , \3901 , \3902 , \3903 ,
         \3904 , \3905 , \3906 , \3907 , \3908 , \3909 , \3910 , \3911 , \3912 , \3913 ,
         \3914 , \3915 , \3916 , \3917 , \3918 , \3919 , \3920 , \3921 , \3922 , \3923 ,
         \3924 , \3925 , \3926 , \3927 , \3928 , \3929 , \3930 , \3931 , \3932 , \3933 ,
         \3934 , \3935 , \3936 , \3937 , \3938 , \3939 , \3940 , \3941 , \3942 , \3943 ,
         \3944 , \3945 , \3946 , \3947 , \3948 , \3949 , \3950 , \3951 , \3952 , \3953 ,
         \3954 , \3955 , \3956 , \3957 , \3958 , \3959 , \3960 , \3961 , \3962 , \3963 ,
         \3964 , \3965 , \3966 , \3967 , \3968 , \3969 , \3970 , \3971 , \3972 , \3973 ,
         \3974 , \3975 , \3976 , \3977 , \3978 , \3979 , \3980 , \3981 , \3982 , \3983 ,
         \3984 , \3985 , \3986 , \3987 , \3988 , \3989 , \3990 , \3991 , \3992 , \3993 ,
         \3994 , \3995 , \3996 , \3997 , \3998 , \3999 , \4000 , \4001 , \4002 , \4003 ,
         \4004 , \4005 , \4006 , \4007 , \4008 , \4009 , \4010 , \4011 , \4012 , \4013 ,
         \4014 , \4015 , \4016 , \4017 , \4018 , \4019 , \4020 , \4021 , \4022 , \4023 ,
         \4024 , \4025 , \4026 , \4027 , \4028 , \4029 , \4030 , \4031 , \4032 , \4033 ,
         \4034 , \4035 , \4036 , \4037 , \4038 , \4039 , \4040 , \4041 , \4042 , \4043 ,
         \4044 , \4045 , \4046 , \4047 , \4048 , \4049 , \4050 , \4051 , \4052 , \4053 ,
         \4054 , \4055 , \4056 , \4057 , \4058 , \4059 , \4060 , \4061 , \4062 , \4063 ,
         \4064 , \4065 , \4066 , \4067 , \4068 , \4069 , \4070 , \4071 , \4072 , \4073 ,
         \4074 , \4075 , \4076 , \4077 , \4078 , \4079 , \4080 , \4081 , \4082 , \4083 ,
         \4084 , \4085 , \4086 , \4087 , \4088 , \4089 , \4090 , \4091 , \4092 , \4093 ,
         \4094 , \4095 , \4096 , \4097 , \4098 , \4099 , \4100 , \4101 , \4102 , \4103 ,
         \4104 , \4105 , \4106 , \4107 , \4108 , \4109 , \4110 , \4111 , \4112 , \4113 ,
         \4114 , \4115 , \4116 , \4117 , \4118 , \4119 , \4120 , \4121 , \4122 , \4123 ,
         \4124 , \4125 , \4126 , \4127 , \4128 , \4129 , \4130 , \4131 , \4132 , \4133 ,
         \4134 , \4135 , \4136 , \4137 , \4138 , \4139 , \4140 , \4141 , \4142 , \4143 ,
         \4144 , \4145 , \4146 , \4147 , \4148 , \4149 , \4150 , \4151 , \4152 , \4153 ,
         \4154 , \4155 , \4156 , \4157 , \4158 , \4159 , \4160 , \4161 , \4162 , \4163 ,
         \4164 , \4165 , \4166 , \4167 , \4168 , \4169 , \4170 , \4171 , \4172 , \4173 ,
         \4174 , \4175 , \4176 , \4177 , \4178 , \4179 , \4180 , \4181 , \4182 , \4183 ,
         \4184 , \4185 , \4186 , \4187 , \4188 , \4189 , \4190 , \4191 , \4192 , \4193 ,
         \4194 , \4195 , \4196 , \4197 , \4198 , \4199 , \4200 , \4201 , \4202 , \4203 ,
         \4204 , \4205 , \4206 , \4207 , \4208 , \4209 , \4210 , \4211 , \4212 , \4213 ,
         \4214 , \4215 , \4216 , \4217 , \4218 , \4219 , \4220 , \4221 , \4222 , \4223 ,
         \4224 , \4225 , \4226 , \4227 , \4228 , \4229 , \4230 , \4231 , \4232 , \4233 ,
         \4234 , \4235 , \4236 , \4237 , \4238 , \4239 , \4240 , \4241 , \4242 , \4243 ,
         \4244 , \4245 , \4246 , \4247 , \4248 , \4249 , \4250 , \4251 , \4252 , \4253 ,
         \4254 , \4255 , \4256 , \4257 , \4258 , \4259 , \4260 , \4261 , \4262 , \4263 ,
         \4264 , \4265 , \4266 , \4267 , \4268 , \4269 , \4270 , \4271 , \4272 , \4273 ,
         \4274 , \4275 , \4276 , \4277 , \4278 , \4279 , \4280 , \4281 , \4282 , \4283 ,
         \4284 , \4285 , \4286 , \4287 , \4288 , \4289 , \4290 , \4291 , \4292 , \4293 ,
         \4294 , \4295 , \4296 , \4297 , \4298 , \4299 , \4300 , \4301 , \4302 , \4303 ,
         \4304 , \4305 , \4306 , \4307 , \4308 , \4309 , \4310 , \4311 , \4312 , \4313 ,
         \4314 , \4315 , \4316 , \4317 , \4318 , \4319 , \4320 , \4321 , \4322 , \4323 ,
         \4324 , \4325 , \4326 , \4327 , \4328 , \4329 , \4330 , \4331 , \4332 , \4333 ,
         \4334 , \4335 , \4336 , \4337 , \4338 , \4339 , \4340 , \4341 , \4342 , \4343 ,
         \4344 , \4345 , \4346 , \4347 , \4348 , \4349 , \4350 , \4351 , \4352 , \4353 ,
         \4354 , \4355 , \4356 , \4357 , \4358 , \4359 , \4360 , \4361 , \4362 , \4363 ,
         \4364 , \4365 , \4366 , \4367 , \4368 , \4369 , \4370 , \4371 , \4372 , \4373 ,
         \4374 , \4375 , \4376 , \4377 , \4378 , \4379 , \4380 , \4381 , \4382 , \4383 ,
         \4384 , \4385 , \4386 , \4387 , \4388 , \4389 , \4390 , \4391 , \4392 , \4393 ,
         \4394 , \4395 , \4396 , \4397 , \4398 , \4399 , \4400 , \4401 , \4402 , \4403 ,
         \4404 , \4405 , \4406 , \4407 , \4408 , \4409 , \4410 , \4411 , \4412 , \4413 ,
         \4414 , \4415 , \4416 , \4417 , \4418 , \4419 , \4420 , \4421 , \4422 , \4423 ,
         \4424 , \4425 , \4426 , \4427 , \4428 , \4429 , \4430 , \4431 , \4432 , \4433 ,
         \4434 , \4435 , \4436 , \4437 , \4438 , \4439 , \4440 , \4441 , \4442 , \4443 ,
         \4444 , \4445 , \4446 , \4447 , \4448 , \4449 , \4450 , \4451 , \4452 , \4453 ,
         \4454 , \4455 , \4456 , \4457 , \4458 , \4459 , \4460 , \4461 , \4462 , \4463 ,
         \4464 , \4465 , \4466 , \4467 , \4468 , \4469 , \4470 , \4471 , \4472 , \4473 ,
         \4474 , \4475 , \4476 , \4477 , \4478 , \4479 , \4480 , \4481 , \4482 , \4483 ,
         \4484 , \4485 , \4486 , \4487 , \4488 , \4489 , \4490 , \4491 , \4492 , \4493 ,
         \4494 , \4495 , \4496 , \4497 , \4498 , \4499 , \4500 , \4501 , \4502 , \4503 ,
         \4504 , \4505 , \4506 , \4507 , \4508 , \4509 , \4510 , \4511 , \4512 , \4513 ,
         \4514 , \4515 , \4516 , \4517 , \4518 , \4519 , \4520 , \4521 , \4522 , \4523 ,
         \4524 , \4525 , \4526 , \4527 , \4528 , \4529 , \4530 , \4531 , \4532 , \4533 ,
         \4534 , \4535 , \4536 , \4537 , \4538 , \4539 , \4540 , \4541 , \4542 , \4543 ,
         \4544 , \4545 , \4546 , \4547 , \4548 , \4549 , \4550 , \4551 , \4552 , \4553 ,
         \4554 , \4555 , \4556 , \4557 , \4558 , \4559 , \4560 , \4561 , \4562 , \4563 ,
         \4564 , \4565 , \4566 , \4567 , \4568 , \4569 , \4570 , \4571 , \4572 , \4573 ,
         \4574 , \4575 , \4576 , \4577 , \4578 , \4579 , \4580 , \4581 , \4582 , \4583 ,
         \4584 , \4585 , \4586 , \4587 , \4588 , \4589 , \4590 , \4591 , \4592 , \4593 ,
         \4594 , \4595 , \4596 , \4597 , \4598 , \4599 , \4600 , \4601 , \4602 , \4603 ,
         \4604 , \4605 , \4606 , \4607 , \4608 , \4609 , \4610 , \4611 , \4612 , \4613 ,
         \4614 , \4615 , \4616 , \4617 , \4618 , \4619 , \4620 , \4621 , \4622 , \4623 ,
         \4624 , \4625 , \4626 , \4627 , \4628 , \4629 , \4630 , \4631 , \4632 , \4633 ,
         \4634 , \4635 , \4636 , \4637 , \4638 , \4639 , \4640 , \4641 , \4642 , \4643 ,
         \4644 , \4645 , \4646 , \4647 , \4648 , \4649 , \4650 , \4651 , \4652 , \4653 ,
         \4654 , \4655 , \4656 , \4657 , \4658 , \4659 , \4660 , \4661 , \4662 , \4663 ,
         \4664 , \4665 , \4666 , \4667 , \4668 , \4669 , \4670 , \4671 , \4672 , \4673 ,
         \4674 , \4675 , \4676 , \4677 , \4678 , \4679 , \4680 , \4681 , \4682 , \4683 ,
         \4684 , \4685 , \4686 , \4687 , \4688 , \4689 , \4690 , \4691 , \4692 , \4693 ,
         \4694 , \4695 , \4696 , \4697 , \4698 , \4699 , \4700 , \4701 , \4702 , \4703 ,
         \4704 , \4705 , \4706 , \4707 , \4708 , \4709 , \4710 , \4711 , \4712 , \4713 ,
         \4714 , \4715 , \4716 , \4717 , \4718 , \4719 , \4720 , \4721 , \4722 , \4723 ,
         \4724 , \4725 , \4726 , \4727 , \4728 , \4729 , \4730 , \4731 , \4732 , \4733 ,
         \4734 , \4735 , \4736 , \4737 , \4738 , \4739 , \4740 , \4741 , \4742 , \4743 ,
         \4744 , \4745 , \4746 , \4747 , \4748 , \4749 , \4750 , \4751 , \4752 , \4753 ,
         \4754 , \4755 , \4756 , \4757 , \4758 , \4759 , \4760 , \4761 , \4762 , \4763 ,
         \4764 , \4765 , \4766 , \4767 , \4768 , \4769 , \4770 , \4771 , \4772 , \4773 ,
         \4774 , \4775 , \4776 , \4777 , \4778 , \4779 , \4780 , \4781 , \4782 , \4783 ,
         \4784 , \4785 , \4786 , \4787 , \4788 , \4789 , \4790 , \4791 , \4792 , \4793 ,
         \4794 , \4795 , \4796 , \4797 , \4798 , \4799 , \4800 , \4801 , \4802 , \4803 ,
         \4804 , \4805 , \4806 , \4807 , \4808 , \4809 , \4810 , \4811 , \4812 , \4813 ,
         \4814 , \4815 , \4816 , \4817 , \4818 , \4819 , \4820 , \4821 , \4822 , \4823 ,
         \4824 , \4825 , \4826 , \4827 , \4828 , \4829 , \4830 , \4831 , \4832 , \4833 ,
         \4834 , \4835 , \4836 , \4837 , \4838 , \4839 , \4840 , \4841 , \4842 , \4843 ,
         \4844 , \4845 , \4846 , \4847 , \4848 , \4849 , \4850 , \4851 , \4852 , \4853 ,
         \4854 , \4855 , \4856 , \4857 , \4858 , \4859 , \4860 , \4861 , \4862 , \4863 ,
         \4864 , \4865 , \4866 , \4867 , \4868 , \4869 , \4870 , \4871 , \4872 , \4873 ,
         \4874 , \4875 , \4876 , \4877 , \4878 , \4879 , \4880 , \4881 , \4882 , \4883 ,
         \4884 , \4885 , \4886 , \4887 , \4888 , \4889 , \4890 , \4891 , \4892 , \4893 ,
         \4894 , \4895 , \4896 , \4897 , \4898 , \4899 , \4900 , \4901 , \4902 , \4903 ,
         \4904 , \4905 , \4906 , \4907 , \4908 , \4909 , \4910 , \4911 , \4912 , \4913 ,
         \4914 , \4915 , \4916 , \4917 , \4918 , \4919 , \4920 , \4921 , \4922 , \4923 ,
         \4924 , \4925 , \4926 , \4927 , \4928 , \4929 , \4930 , \4931 , \4932 , \4933 ,
         \4934 , \4935 , \4936 , \4937 , \4938 , \4939 , \4940 , \4941 , \4942 , \4943 ,
         \4944 , \4945 , \4946 , \4947 , \4948 , \4949 , \4950 , \4951 , \4952 , \4953 ,
         \4954 , \4955 , \4956 , \4957 , \4958 , \4959 , \4960 , \4961 , \4962 , \4963 ,
         \4964 , \4965 , \4966 , \4967 , \4968 , \4969 , \4970 , \4971 , \4972 , \4973 ,
         \4974 , \4975 , \4976 , \4977 , \4978 , \4979 , \4980 , \4981 , \4982 , \4983 ,
         \4984 , \4985 , \4986 , \4987 , \4988 , \4989 , \4990 , \4991 , \4992 , \4993 ,
         \4994 , \4995 , \4996 , \4997 , \4998 , \4999 , \5000 , \5001 , \5002 , \5003 ,
         \5004 , \5005 , \5006 , \5007 , \5008 , \5009 , \5010 , \5011 , \5012 , \5013 ,
         \5014 , \5015 , \5016 , \5017 , \5018 , \5019 , \5020 , \5021 , \5022 , \5023 ,
         \5024 , \5025 , \5026 , \5027 , \5028 , \5029 , \5030 , \5031 , \5032 , \5033 ,
         \5034 , \5035 , \5036 , \5037 , \5038 , \5039 , \5040 , \5041 , \5042 , \5043 ,
         \5044 , \5045 , \5046 , \5047 , \5048 , \5049 , \5050 , \5051 , \5052 , \5053 ,
         \5054 , \5055 , \5056 , \5057 , \5058 , \5059 , \5060 , \5061 , \5062 , \5063 ,
         \5064 , \5065 , \5066 , \5067 , \5068 , \5069 , \5070 , \5071 , \5072 , \5073 ,
         \5074 , \5075 , \5076 , \5077 , \5078 , \5079 , \5080 , \5081 , \5082 , \5083 ,
         \5084 , \5085 , \5086 , \5087 , \5088 , \5089 , \5090 , \5091 , \5092 , \5093 ,
         \5094 , \5095 , \5096 , \5097 , \5098 , \5099 , \5100 , \5101 , \5102 , \5103 ,
         \5104 , \5105 , \5106 , \5107 , \5108 , \5109 , \5110 , \5111 , \5112 , \5113 ,
         \5114 , \5115 , \5116 , \5117 , \5118 , \5119 , \5120 , \5121 , \5122 , \5123 ,
         \5124 , \5125 , \5126 , \5127 , \5128 , \5129 , \5130 , \5131 , \5132 , \5133 ,
         \5134 , \5135 , \5136 , \5137 , \5138 , \5139 , \5140 , \5141 , \5142 , \5143 ,
         \5144 , \5145 , \5146 , \5147 , \5148 , \5149 , \5150 , \5151 , \5152 , \5153 ,
         \5154 , \5155 , \5156 , \5157 , \5158 , \5159 , \5160 , \5161 , \5162 , \5163 ,
         \5164 , \5165 , \5166 , \5167 , \5168 , \5169 , \5170 , \5171 , \5172 , \5173 ,
         \5174 , \5175 , \5176 , \5177 , \5178 , \5179 , \5180 , \5181 , \5182 , \5183 ,
         \5184 , \5185 , \5186 , \5187 , \5188 , \5189 , \5190 , \5191 , \5192 , \5193 ,
         \5194 , \5195 , \5196 , \5197 , \5198 , \5199 , \5200 , \5201 , \5202 , \5203 ,
         \5204 , \5205 , \5206 , \5207 , \5208 , \5209 , \5210 , \5211 , \5212 , \5213 ,
         \5214 , \5215 , \5216 , \5217 , \5218 , \5219 , \5220 , \5221 , \5222 , \5223 ,
         \5224 , \5225 , \5226 , \5227 , \5228 , \5229 , \5230 , \5231 , \5232 , \5233 ,
         \5234 , \5235 , \5236 , \5237 , \5238 , \5239 , \5240 , \5241 , \5242 , \5243 ,
         \5244 , \5245 , \5246 , \5247 , \5248 , \5249 , \5250 , \5251 , \5252 , \5253 ,
         \5254 , \5255 , \5256 , \5257 , \5258 , \5259 , \5260 , \5261 , \5262 , \5263 ,
         \5264 , \5265 , \5266 , \5267 , \5268 , \5269 , \5270 , \5271 , \5272 , \5273 ,
         \5274 , \5275 , \5276 , \5277 , \5278 , \5279 , \5280 , \5281 , \5282 , \5283 ,
         \5284 , \5285 , \5286 , \5287 , \5288 , \5289 , \5290 , \5291 , \5292 , \5293 ,
         \5294 , \5295 , \5296 , \5297 , \5298 , \5299 , \5300 , \5301 , \5302 , \5303 ,
         \5304 , \5305 , \5306 , \5307 , \5308 , \5309 , \5310 , \5311 , \5312 , \5313 ,
         \5314 , \5315 , \5316 , \5317 , \5318 , \5319 , \5320 , \5321 , \5322 , \5323 ,
         \5324 , \5325 , \5326 , \5327 , \5328 , \5329 , \5330 , \5331 , \5332 , \5333 ,
         \5334 , \5335 , \5336 , \5337 , \5338 , \5339 , \5340 , \5341 , \5342 , \5343 ,
         \5344 , \5345 , \5346 , \5347 , \5348 , \5349 , \5350 , \5351 , \5352 , \5353 ,
         \5354 , \5355 , \5356 , \5357 , \5358 , \5359 , \5360 , \5361 , \5362 , \5363 ,
         \5364 , \5365 , \5366 , \5367 , \5368 , \5369 , \5370 , \5371 , \5372 , \5373 ,
         \5374 , \5375 , \5376 , \5377 , \5378 , \5379 , \5380 , \5381 , \5382 , \5383 ,
         \5384 , \5385 , \5386 , \5387 , \5388 , \5389 , \5390 , \5391 , \5392 , \5393 ,
         \5394 , \5395 , \5396 , \5397 , \5398 , \5399 , \5400 , \5401 , \5402 , \5403 ,
         \5404 , \5405 , \5406 , \5407 , \5408 , \5409 , \5410 , \5411 , \5412 , \5413 ,
         \5414 , \5415 , \5416 , \5417 , \5418 , \5419 , \5420 , \5421 , \5422 , \5423 ,
         \5424 , \5425 , \5426 , \5427 , \5428 , \5429 , \5430 , \5431 , \5432 , \5433 ,
         \5434 , \5435 , \5436 , \5437 , \5438 , \5439 , \5440 , \5441 , \5442 , \5443 ,
         \5444 , \5445 , \5446 , \5447 , \5448 , \5449 , \5450 , \5451 , \5452 , \5453 ,
         \5454 , \5455 , \5456 , \5457 , \5458 , \5459 , \5460 , \5461 , \5462 , \5463 ,
         \5464 , \5465 , \5466 , \5467 , \5468 , \5469 , \5470 , \5471 , \5472 , \5473 ,
         \5474 , \5475 , \5476 , \5477 , \5478 , \5479 , \5480 , \5481 , \5482 , \5483 ,
         \5484 , \5485 , \5486 , \5487 , \5488 , \5489 , \5490 , \5491 , \5492 , \5493 ,
         \5494 , \5495 , \5496 , \5497 , \5498 , \5499 , \5500 , \5501 , \5502 , \5503 ,
         \5504 , \5505 , \5506 , \5507 , \5508 , \5509 , \5510 , \5511 , \5512 , \5513 ,
         \5514 , \5515 , \5516 , \5517 , \5518 , \5519 , \5520 , \5521 , \5522 , \5523 ,
         \5524 , \5525 , \5526 , \5527 , \5528 , \5529 , \5530 , \5531 , \5532 , \5533 ,
         \5534 , \5535 , \5536 , \5537 , \5538 , \5539 , \5540 , \5541 , \5542 , \5543 ,
         \5544 , \5545 , \5546 , \5547 , \5548 , \5549 , \5550 , \5551 , \5552 , \5553 ,
         \5554 , \5555 , \5556 , \5557 , \5558 , \5559 , \5560 , \5561 , \5562 , \5563 ,
         \5564 , \5565 , \5566 , \5567 , \5568 , \5569 , \5570 , \5571 , \5572 , \5573 ,
         \5574 , \5575 , \5576 , \5577 , \5578 , \5579 , \5580 , \5581 , \5582 , \5583 ,
         \5584 , \5585 , \5586 , \5587 , \5588 , \5589 , \5590 , \5591 , \5592 , \5593 ,
         \5594 , \5595 , \5596 , \5597 , \5598 , \5599 , \5600 , \5601 , \5602 , \5603 ,
         \5604 , \5605 , \5606 , \5607 , \5608 , \5609 , \5610 , \5611 , \5612 , \5613 ,
         \5614 , \5615 , \5616 , \5617 , \5618 , \5619 , \5620 , \5621 , \5622 , \5623 ,
         \5624 , \5625 , \5626 , \5627 , \5628 , \5629 , \5630 , \5631 , \5632 , \5633 ,
         \5634 , \5635 , \5636 , \5637 , \5638 , \5639 , \5640 , \5641 , \5642 , \5643 ,
         \5644 , \5645 , \5646 , \5647 , \5648 , \5649 , \5650 , \5651 , \5652 , \5653 ,
         \5654 , \5655 , \5656 , \5657 , \5658 , \5659 , \5660 , \5661 , \5662 , \5663 ,
         \5664 , \5665 , \5666 , \5667 , \5668 , \5669 , \5670 , \5671 , \5672 , \5673 ,
         \5674 , \5675 , \5676 , \5677 , \5678 , \5679 , \5680 , \5681 , \5682 , \5683 ,
         \5684 , \5685 , \5686 , \5687 , \5688 , \5689 , \5690 , \5691 , \5692 , \5693 ,
         \5694 , \5695 , \5696 , \5697 , \5698 , \5699 , \5700 , \5701 , \5702 , \5703 ,
         \5704 , \5705 , \5706 , \5707 , \5708 , \5709 , \5710 , \5711 , \5712 , \5713 ,
         \5714 , \5715 , \5716 , \5717 , \5718 , \5719 , \5720 , \5721 , \5722 , \5723 ,
         \5724 , \5725 , \5726 , \5727 , \5728 , \5729 , \5730 , \5731 , \5732 , \5733 ,
         \5734 , \5735 , \5736 , \5737 , \5738 , \5739 , \5740 , \5741 , \5742 , \5743 ,
         \5744 , \5745 , \5746 , \5747 , \5748 , \5749 , \5750 , \5751 , \5752 , \5753 ,
         \5754 , \5755 , \5756 , \5757 , \5758 , \5759 , \5760 , \5761 , \5762 , \5763 ,
         \5764 , \5765 , \5766 , \5767 , \5768 , \5769 , \5770 , \5771 , \5772 , \5773 ,
         \5774 , \5775 , \5776 , \5777 , \5778 , \5779 , \5780 , \5781 , \5782 , \5783 ,
         \5784 , \5785 , \5786 , \5787 , \5788 , \5789 , \5790 , \5791 , \5792 , \5793 ,
         \5794 , \5795 , \5796 , \5797 , \5798 , \5799 , \5800 , \5801 , \5802 , \5803 ,
         \5804 , \5805 , \5806 , \5807 , \5808 , \5809 , \5810 , \5811 , \5812 , \5813 ,
         \5814 , \5815 , \5816 , \5817 , \5818 , \5819 , \5820 , \5821 , \5822 , \5823 ,
         \5824 , \5825 , \5826 , \5827 , \5828 , \5829 , \5830 , \5831 , \5832 , \5833 ,
         \5834 , \5835 , \5836 , \5837 , \5838 , \5839 , \5840 , \5841 , \5842 , \5843 ,
         \5844 , \5845 , \5846 , \5847 , \5848 , \5849 , \5850 , \5851 , \5852 , \5853 ,
         \5854 , \5855 , \5856 , \5857 , \5858 , \5859 , \5860 , \5861 , \5862 , \5863 ,
         \5864 , \5865 , \5866 , \5867 , \5868 , \5869 , \5870 , \5871 , \5872 , \5873 ,
         \5874 , \5875 , \5876 , \5877 , \5878 , \5879 , \5880 , \5881 , \5882 , \5883 ,
         \5884 , \5885 , \5886 , \5887 , \5888 , \5889 , \5890 , \5891 , \5892 , \5893 ,
         \5894 , \5895 , \5896 , \5897 , \5898 , \5899 , \5900 , \5901 , \5902 , \5903 ,
         \5904 , \5905 , \5906 , \5907 , \5908 , \5909 , \5910 , \5911 , \5912 , \5913 ,
         \5914 , \5915 , \5916 , \5917 , \5918 , \5919 , \5920 , \5921 , \5922 , \5923 ,
         \5924 , \5925 , \5926 , \5927 , \5928 , \5929 , \5930 , \5931 , \5932 , \5933 ,
         \5934 , \5935 , \5936 , \5937 , \5938 , \5939 , \5940 , \5941 , \5942 , \5943 ,
         \5944 , \5945 , \5946 , \5947 , \5948 , \5949 , \5950 , \5951 , \5952 , \5953 ,
         \5954 , \5955 , \5956 , \5957 , \5958 , \5959 , \5960 , \5961 , \5962 , \5963 ,
         \5964 , \5965 , \5966 , \5967 , \5968 , \5969 , \5970 , \5971 , \5972 , \5973 ,
         \5974 , \5975 , \5976 , \5977 , \5978 , \5979 , \5980 , \5981 , \5982 , \5983 ,
         \5984 , \5985 , \5986 , \5987 , \5988 , \5989 , \5990 , \5991 , \5992 , \5993 ,
         \5994 , \5995 , \5996 , \5997 , \5998 , \5999 , \6000 , \6001 , \6002 , \6003 ,
         \6004 , \6005 , \6006 , \6007 , \6008 , \6009 , \6010 , \6011 , \6012 , \6013 ,
         \6014 , \6015 , \6016 , \6017 , \6018 , \6019 , \6020 , \6021 , \6022 , \6023 ,
         \6024 , \6025 , \6026 , \6027 , \6028 , \6029 , \6030 , \6031 , \6032 , \6033 ,
         \6034 , \6035 , \6036 , \6037 , \6038 , \6039 , \6040 , \6041 , \6042 , \6043 ,
         \6044 , \6045 , \6046 , \6047 , \6048 , \6049 , \6050 , \6051 , \6052 , \6053 ,
         \6054 , \6055 , \6056 , \6057 , \6058 , \6059 , \6060 , \6061 , \6062 , \6063 ,
         \6064 , \6065 , \6066 , \6067 , \6068 , \6069 , \6070 , \6071 , \6072 , \6073 ,
         \6074 , \6075 , \6076 , \6077 , \6078 , \6079 , \6080 , \6081 , \6082 , \6083 ,
         \6084 , \6085 , \6086 , \6087 , \6088 , \6089 , \6090 , \6091 , \6092 , \6093 ,
         \6094 , \6095 , \6096 , \6097 , \6098 , \6099 , \6100 , \6101 , \6102 , \6103 ,
         \6104 , \6105 , \6106 , \6107 , \6108 , \6109 , \6110 , \6111 , \6112 , \6113 ,
         \6114 , \6115 , \6116 , \6117 , \6118 , \6119 , \6120 , \6121 , \6122 , \6123 ,
         \6124 , \6125 , \6126 , \6127 , \6128 , \6129 , \6130 , \6131 , \6132 , \6133 ,
         \6134 , \6135 , \6136 , \6137 , \6138 , \6139 , \6140 , \6141 , \6142 , \6143 ,
         \6144 , \6145 , \6146 , \6147 , \6148 , \6149 , \6150 , \6151 , \6152 , \6153 ,
         \6154 , \6155 , \6156 , \6157 , \6158 , \6159 , \6160 , \6161 , \6162 , \6163 ,
         \6164 , \6165 , \6166 , \6167 , \6168 , \6169 , \6170 , \6171 , \6172 , \6173 ,
         \6174 , \6175 , \6176 , \6177 , \6178 , \6179 , \6180 , \6181 , \6182 , \6183 ,
         \6184 , \6185 , \6186 , \6187 , \6188 , \6189 , \6190 , \6191 , \6192 , \6193 ,
         \6194 , \6195 , \6196 , \6197 , \6198 , \6199 , \6200 , \6201 , \6202 , \6203 ,
         \6204 , \6205 , \6206 , \6207 , \6208 , \6209 , \6210 , \6211 , \6212 , \6213 ,
         \6214 , \6215 , \6216 , \6217 , \6218 , \6219 , \6220 , \6221 , \6222 , \6223 ,
         \6224 , \6225 , \6226 , \6227 , \6228 , \6229 , \6230 , \6231 , \6232 , \6233 ,
         \6234 , \6235 , \6236 , \6237 , \6238 , \6239 , \6240 , \6241 , \6242 , \6243 ,
         \6244 , \6245 , \6246 , \6247 , \6248 , \6249 , \6250 , \6251 , \6252 , \6253 ,
         \6254 , \6255 , \6256 , \6257 , \6258 , \6259 , \6260 , \6261 , \6262 , \6263 ,
         \6264 , \6265 , \6266 , \6267 , \6268 , \6269 , \6270 , \6271 , \6272 , \6273 ,
         \6274 , \6275 , \6276 , \6277 , \6278 , \6279 , \6280 , \6281 , \6282 , \6283 ,
         \6284 , \6285 , \6286 , \6287 , \6288 , \6289 , \6290 , \6291 , \6292 , \6293 ,
         \6294 , \6295 , \6296 , \6297 , \6298 , \6299 , \6300 , \6301 , \6302 , \6303 ,
         \6304 , \6305 , \6306 , \6307 , \6308 , \6309 , \6310 , \6311 , \6312 , \6313 ,
         \6314 , \6315 , \6316 , \6317 , \6318 , \6319 , \6320 , \6321 , \6322 , \6323 ,
         \6324 , \6325 , \6326 , \6327 , \6328 , \6329 , \6330 , \6331 , \6332 , \6333 ,
         \6334 , \6335 , \6336 , \6337 , \6338 , \6339 , \6340 , \6341 , \6342 , \6343 ,
         \6344 , \6345 , \6346 , \6347 , \6348 , \6349 , \6350 , \6351 , \6352 , \6353 ,
         \6354 , \6355 , \6356 , \6357 , \6358 , \6359 , \6360 , \6361 , \6362 , \6363 ,
         \6364 , \6365 , \6366 , \6367 , \6368 , \6369 , \6370 , \6371 , \6372 , \6373 ,
         \6374 , \6375 , \6376 , \6377 , \6378 , \6379 , \6380 , \6381 , \6382 , \6383 ,
         \6384 , \6385 , \6386 , \6387 , \6388 , \6389 , \6390 , \6391 , \6392 , \6393 ,
         \6394 , \6395 , \6396 , \6397 , \6398 , \6399 , \6400 , \6401 , \6402 , \6403 ,
         \6404 , \6405 , \6406 , \6407 , \6408 , \6409 , \6410 , \6411 , \6412 , \6413 ,
         \6414 , \6415 , \6416 , \6417 , \6418 , \6419 , \6420 , \6421 , \6422 , \6423 ,
         \6424 , \6425 , \6426 , \6427 , \6428 , \6429 , \6430 , \6431 , \6432 , \6433 ,
         \6434 , \6435 , \6436 , \6437 , \6438 , \6439 , \6440 , \6441 , \6442 , \6443 ,
         \6444 , \6445 , \6446 , \6447 , \6448 , \6449 , \6450 , \6451 , \6452 , \6453 ,
         \6454 , \6455 , \6456 , \6457 , \6458 , \6459 , \6460 , \6461 , \6462 , \6463 ,
         \6464 , \6465 , \6466 , \6467 , \6468 , \6469 , \6470 , \6471 , \6472 , \6473 ,
         \6474 , \6475 , \6476 , \6477 , \6478 , \6479 , \6480 , \6481 , \6482 , \6483 ,
         \6484 , \6485 , \6486 , \6487 , \6488 , \6489 , \6490 , \6491 , \6492 , \6493 ,
         \6494 , \6495 , \6496 , \6497 , \6498 , \6499 , \6500 , \6501 , \6502 , \6503 ,
         \6504 , \6505 , \6506 , \6507 , \6508 , \6509 , \6510 , \6511 , \6512 , \6513 ,
         \6514 , \6515 , \6516 , \6517 , \6518 , \6519 , \6520 , \6521 , \6522 , \6523 ,
         \6524 , \6525 , \6526 , \6527 , \6528 , \6529 , \6530 , \6531 , \6532 , \6533 ,
         \6534 , \6535 , \6536 , \6537 , \6538 , \6539 , \6540 , \6541 , \6542 , \6543 ,
         \6544 , \6545 , \6546 , \6547 , \6548 , \6549 , \6550 , \6551 , \6552 , \6553 ,
         \6554 , \6555 , \6556 , \6557 , \6558 , \6559 , \6560 , \6561 , \6562 , \6563 ,
         \6564 , \6565 , \6566 , \6567 , \6568 , \6569 , \6570 , \6571 , \6572 , \6573 ,
         \6574 , \6575 , \6576 , \6577 , \6578 , \6579 , \6580 , \6581 , \6582 , \6583 ,
         \6584 , \6585 , \6586 , \6587 , \6588 , \6589 , \6590 , \6591 , \6592 , \6593 ,
         \6594 , \6595 , \6596 , \6597 , \6598 , \6599 , \6600 , \6601 , \6602 , \6603 ,
         \6604 , \6605 , \6606 , \6607 , \6608 , \6609 , \6610 , \6611 , \6612 , \6613 ,
         \6614 , \6615 , \6616 , \6617 , \6618 , \6619 , \6620 , \6621 , \6622 , \6623 ,
         \6624 , \6625 , \6626 , \6627 , \6628 , \6629 , \6630 , \6631 , \6632 , \6633 ,
         \6634 , \6635 , \6636 , \6637 , \6638 , \6639 , \6640 , \6641 , \6642 , \6643 ,
         \6644 , \6645 , \6646 , \6647 , \6648 , \6649 , \6650 , \6651 , \6652 , \6653 ,
         \6654 , \6655 , \6656 , \6657 , \6658 , \6659 , \6660 , \6661 , \6662 , \6663 ,
         \6664 , \6665 , \6666 , \6667 , \6668 , \6669 , \6670 , \6671 , \6672 , \6673 ,
         \6674 , \6675 , \6676 , \6677 , \6678 , \6679 , \6680 , \6681 , \6682 , \6683 ,
         \6684 , \6685 , \6686 , \6687 , \6688 , \6689 , \6690 , \6691 , \6692 , \6693 ,
         \6694 , \6695 , \6696 , \6697 , \6698 , \6699 , \6700 , \6701 , \6702 , \6703 ,
         \6704 , \6705 , \6706 , \6707 , \6708 , \6709 , \6710 , \6711 , \6712 , \6713 ,
         \6714 , \6715 , \6716 , \6717 , \6718 , \6719 , \6720 , \6721 , \6722 , \6723 ,
         \6724 , \6725 , \6726 , \6727 , \6728 , \6729 , \6730 , \6731 , \6732 , \6733 ,
         \6734 , \6735 , \6736 , \6737 , \6738 , \6739 , \6740 , \6741 , \6742 , \6743 ,
         \6744 , \6745 , \6746 , \6747 , \6748 , \6749 , \6750 , \6751 , \6752 , \6753 ,
         \6754 , \6755 , \6756 , \6757 , \6758 , \6759 , \6760 , \6761 , \6762 , \6763 ,
         \6764 , \6765 , \6766 , \6767 , \6768 , \6769 , \6770 , \6771 , \6772 , \6773 ,
         \6774 , \6775 , \6776 , \6777 , \6778 , \6779 , \6780 , \6781 , \6782 , \6783 ,
         \6784 , \6785 , \6786 , \6787 , \6788 , \6789 , \6790 , \6791 , \6792 , \6793 ,
         \6794 , \6795 , \6796 , \6797 , \6798 , \6799 , \6800 , \6801 , \6802 , \6803 ,
         \6804 , \6805 , \6806 , \6807 , \6808 , \6809 , \6810 , \6811 , \6812 , \6813 ,
         \6814 , \6815 , \6816 , \6817 , \6818 , \6819 , \6820 , \6821 , \6822 , \6823 ,
         \6824 , \6825 , \6826 , \6827 , \6828 , \6829 , \6830 , \6831 , \6832 , \6833 ,
         \6834 , \6835 , \6836 , \6837 , \6838 , \6839 , \6840 , \6841 , \6842 , \6843 ,
         \6844 , \6845 , \6846 , \6847 , \6848 , \6849 , \6850 , \6851 , \6852 , \6853 ,
         \6854 , \6855 , \6856 , \6857 , \6858 , \6859 , \6860 , \6861 , \6862 , \6863 ,
         \6864 , \6865 , \6866 , \6867 , \6868 , \6869 , \6870 , \6871 , \6872 , \6873 ,
         \6874 , \6875 , \6876 , \6877 , \6878 , \6879 , \6880 , \6881 , \6882 , \6883 ,
         \6884 , \6885 , \6886 , \6887 , \6888 , \6889 , \6890 , \6891 , \6892 , \6893 ,
         \6894 , \6895 , \6896 , \6897 , \6898 , \6899 , \6900 , \6901 , \6902 , \6903 ,
         \6904 , \6905 , \6906 , \6907 , \6908 , \6909 , \6910 , \6911 , \6912 , \6913 ,
         \6914 , \6915 , \6916 , \6917 , \6918 , \6919 , \6920 , \6921 , \6922 , \6923 ,
         \6924 , \6925 , \6926 , \6927 , \6928 , \6929 , \6930 , \6931 , \6932 , \6933 ,
         \6934 , \6935 , \6936 , \6937 , \6938 , \6939 , \6940 , \6941 , \6942 , \6943 ,
         \6944 , \6945 , \6946 , \6947 , \6948 , \6949 , \6950 , \6951 , \6952 , \6953 ,
         \6954 , \6955 , \6956 , \6957 , \6958 , \6959 , \6960 , \6961 , \6962 , \6963 ,
         \6964 , \6965 , \6966 , \6967 , \6968 , \6969 , \6970 , \6971 , \6972 , \6973 ,
         \6974 , \6975 , \6976 , \6977 , \6978 , \6979 , \6980 , \6981 , \6982 , \6983 ,
         \6984 , \6985 , \6986 , \6987 , \6988 , \6989 , \6990 , \6991 , \6992 , \6993 ,
         \6994 , \6995 , \6996 , \6997 , \6998 , \6999 , \7000 , \7001 , \7002 , \7003 ,
         \7004 , \7005 , \7006 , \7007 , \7008 , \7009 , \7010 , \7011 , \7012 , \7013 ,
         \7014 , \7015 , \7016 , \7017 , \7018 , \7019 , \7020 , \7021 , \7022 , \7023 ,
         \7024 , \7025 , \7026 , \7027 , \7028 , \7029 , \7030 , \7031 , \7032 , \7033 ,
         \7034 , \7035 , \7036 , \7037 , \7038 , \7039 , \7040 , \7041 , \7042 , \7043 ,
         \7044 , \7045 , \7046 , \7047 , \7048 , \7049 , \7050 , \7051 , \7052 , \7053 ,
         \7054 , \7055 , \7056 , \7057 , \7058 , \7059 , \7060 , \7061 , \7062 , \7063 ,
         \7064 , \7065 , \7066 , \7067 , \7068 , \7069 , \7070 , \7071 , \7072 , \7073 ,
         \7074 , \7075 , \7076 , \7077 , \7078 , \7079 , \7080 , \7081 , \7082 , \7083 ,
         \7084 , \7085 , \7086 , \7087 , \7088 , \7089 , \7090 , \7091 , \7092 , \7093 ,
         \7094 , \7095 , \7096 , \7097 , \7098 , \7099 , \7100 , \7101 , \7102 , \7103 ,
         \7104 , \7105 , \7106 , \7107 , \7108 , \7109 , \7110 , \7111 , \7112 , \7113 ,
         \7114 , \7115 , \7116 , \7117 , \7118 , \7119 , \7120 , \7121 , \7122 , \7123 ,
         \7124 , \7125 , \7126 , \7127 , \7128 , \7129 , \7130 , \7131 , \7132 , \7133 ,
         \7134 , \7135 , \7136 , \7137 , \7138 , \7139 , \7140 , \7141 , \7142 , \7143 ,
         \7144 , \7145 , \7146 , \7147 , \7148 , \7149 , \7150 , \7151 , \7152 , \7153 ,
         \7154 , \7155 , \7156 , \7157 , \7158 , \7159 , \7160 , \7161 , \7162 , \7163 ,
         \7164 , \7165 , \7166 , \7167 , \7168 , \7169 , \7170 , \7171 , \7172 , \7173 ,
         \7174 , \7175 , \7176 , \7177 , \7178 , \7179 , \7180 , \7181 , \7182 , \7183 ,
         \7184 , \7185 , \7186 , \7187 , \7188 , \7189 , \7190 , \7191 , \7192 , \7193 ,
         \7194 , \7195 , \7196 , \7197 , \7198 , \7199 , \7200 , \7201 , \7202 , \7203 ,
         \7204 , \7205 , \7206 , \7207 , \7208 , \7209 , \7210 , \7211 , \7212 , \7213 ,
         \7214 , \7215 , \7216 , \7217 , \7218 , \7219 , \7220 , \7221 , \7222 , \7223 ,
         \7224 , \7225 , \7226 , \7227 , \7228 , \7229 , \7230 , \7231 , \7232 , \7233 ,
         \7234 , \7235 , \7236 , \7237 , \7238 , \7239 , \7240 , \7241 , \7242 , \7243 ,
         \7244 , \7245 , \7246 , \7247 , \7248 , \7249 , \7250 , \7251 , \7252 , \7253 ,
         \7254 , \7255 , \7256 , \7257 , \7258 , \7259 , \7260 , \7261 , \7262 , \7263 ,
         \7264 , \7265 , \7266 , \7267 , \7268 , \7269 , \7270 , \7271 , \7272 , \7273 ,
         \7274 , \7275 , \7276 , \7277 , \7278 , \7279 , \7280 , \7281 , \7282 , \7283 ,
         \7284 , \7285 , \7286 , \7287 , \7288 , \7289 , \7290 , \7291 , \7292 , \7293 ,
         \7294 , \7295 , \7296 , \7297 , \7298 , \7299 , \7300 , \7301 , \7302 , \7303 ,
         \7304 , \7305 , \7306 , \7307 , \7308 , \7309 , \7310 , \7311 , \7312 , \7313 ,
         \7314 , \7315 , \7316 , \7317 , \7318 , \7319 , \7320 , \7321 , \7322 , \7323 ,
         \7324 , \7325 , \7326 , \7327 , \7328 , \7329 , \7330 , \7331 , \7332 , \7333 ,
         \7334 , \7335 , \7336 , \7337 , \7338 , \7339 , \7340 , \7341 , \7342 , \7343 ,
         \7344 , \7345 , \7346 , \7347 , \7348 , \7349 , \7350 , \7351 , \7352 , \7353 ,
         \7354 , \7355 , \7356 , \7357 , \7358 , \7359 , \7360 , \7361 , \7362 , \7363 ,
         \7364 , \7365 , \7366 , \7367 , \7368 , \7369 , \7370 , \7371 , \7372 , \7373 ,
         \7374 , \7375 , \7376 , \7377 , \7378 , \7379 , \7380 , \7381 , \7382 , \7383 ,
         \7384 , \7385 , \7386 , \7387 , \7388 , \7389 , \7390 , \7391 , \7392 , \7393 ,
         \7394 , \7395 , \7396 , \7397 , \7398 , \7399 , \7400 , \7401 , \7402 , \7403 ,
         \7404 , \7405 , \7406 , \7407 , \7408 , \7409 , \7410 , \7411 , \7412 , \7413 ,
         \7414 , \7415 , \7416 , \7417 , \7418 , \7419 , \7420 , \7421 , \7422 , \7423 ,
         \7424 , \7425 , \7426 , \7427 , \7428 , \7429 , \7430 , \7431 , \7432 , \7433 ,
         \7434 , \7435 , \7436 , \7437 , \7438 , \7439 , \7440 , \7441 , \7442 , \7443 ,
         \7444 , \7445 , \7446 , \7447 , \7448 , \7449 , \7450 , \7451 , \7452 , \7453 ,
         \7454 , \7455 , \7456 , \7457 , \7458 , \7459 , \7460 , \7461 , \7462 , \7463 ,
         \7464 , \7465 , \7466 , \7467 , \7468 , \7469 , \7470 , \7471 , \7472 , \7473 ,
         \7474 , \7475 , \7476 , \7477 , \7478 , \7479 , \7480 , \7481 , \7482 , \7483 ,
         \7484 , \7485 , \7486 , \7487 , \7488 , \7489 , \7490 , \7491 , \7492 , \7493 ,
         \7494 , \7495 , \7496 , \7497 , \7498 , \7499 , \7500 , \7501 , \7502 , \7503 ,
         \7504 , \7505 , \7506 , \7507 , \7508 , \7509 , \7510 , \7511 , \7512 , \7513 ,
         \7514 , \7515 , \7516 , \7517 , \7518 , \7519 , \7520 , \7521 , \7522 , \7523 ,
         \7524 , \7525 , \7526 , \7527 , \7528 , \7529 , \7530 , \7531 , \7532 , \7533 ,
         \7534 , \7535 , \7536 , \7537 , \7538 , \7539 , \7540 , \7541 , \7542 , \7543 ,
         \7544 , \7545 , \7546 , \7547 , \7548 , \7549 , \7550 , \7551 , \7552 , \7553 ,
         \7554 , \7555 , \7556 , \7557 , \7558 , \7559 , \7560 , \7561 , \7562 , \7563 ,
         \7564 , \7565 , \7566 , \7567 , \7568 , \7569 , \7570 , \7571 , \7572 , \7573 ,
         \7574 , \7575 , \7576 , \7577 , \7578 , \7579 , \7580 , \7581 , \7582 , \7583 ,
         \7584 , \7585 , \7586 , \7587 , \7588 , \7589 , \7590 , \7591 , \7592 , \7593 ,
         \7594 , \7595 , \7596 , \7597 , \7598 , \7599 , \7600 , \7601 , \7602 , \7603 ,
         \7604 , \7605 , \7606 , \7607 , \7608 , \7609 , \7610 , \7611 , \7612 , \7613 ,
         \7614 , \7615 , \7616 , \7617 , \7618 , \7619 , \7620 , \7621 , \7622 , \7623 ,
         \7624 , \7625 , \7626 , \7627 , \7628 , \7629 , \7630 , \7631 , \7632 , \7633 ,
         \7634 , \7635 , \7636 , \7637 , \7638 , \7639 , \7640 , \7641 , \7642 , \7643 ,
         \7644 , \7645 , \7646 , \7647 , \7648 , \7649 , \7650 , \7651 , \7652 , \7653 ,
         \7654 , \7655 , \7656 , \7657 , \7658 , \7659 , \7660 , \7661 , \7662 , \7663 ,
         \7664 , \7665 , \7666 , \7667 , \7668 , \7669 , \7670 , \7671 , \7672 , \7673 ,
         \7674 , \7675 , \7676 , \7677 , \7678 , \7679 , \7680 , \7681 , \7682 , \7683 ,
         \7684 , \7685 , \7686 , \7687 , \7688 , \7689 , \7690 , \7691 , \7692 , \7693 ,
         \7694 , \7695 , \7696 , \7697 , \7698 , \7699 , \7700 , \7701 , \7702 , \7703 ,
         \7704 , \7705 , \7706 , \7707 , \7708 , \7709 , \7710 , \7711 , \7712 , \7713 ,
         \7714 , \7715 , \7716 , \7717 , \7718 , \7719 , \7720 , \7721 , \7722 , \7723 ,
         \7724 , \7725 , \7726 , \7727 , \7728 , \7729 , \7730 , \7731 , \7732 , \7733 ,
         \7734 , \7735 , \7736 , \7737 , \7738 , \7739 , \7740 , \7741 , \7742 , \7743 ,
         \7744 , \7745 , \7746 , \7747 , \7748 , \7749 , \7750 , \7751 , \7752 , \7753 ,
         \7754 , \7755 , \7756 , \7757 , \7758 , \7759 , \7760 , \7761 , \7762 , \7763 ,
         \7764 , \7765 , \7766 , \7767 , \7768 , \7769 , \7770 , \7771 , \7772 , \7773 ,
         \7774 , \7775 , \7776 , \7777 , \7778 , \7779 , \7780 , \7781 , \7782 , \7783 ,
         \7784 , \7785 , \7786 , \7787 , \7788 , \7789 , \7790 , \7791 , \7792 , \7793 ,
         \7794 , \7795 , \7796 , \7797 , \7798 , \7799 , \7800 , \7801 , \7802 , \7803 ,
         \7804 , \7805 , \7806 , \7807 , \7808 , \7809 , \7810 , \7811 , \7812 , \7813 ,
         \7814 , \7815 , \7816 , \7817 , \7818 , \7819 , \7820 , \7821 , \7822 , \7823 ,
         \7824 , \7825 , \7826 , \7827 , \7828 , \7829 , \7830 , \7831 , \7832 , \7833 ,
         \7834 , \7835 , \7836 , \7837 , \7838 , \7839 , \7840 , \7841 , \7842 , \7843 ,
         \7844 , \7845 , \7846 , \7847 , \7848 , \7849 , \7850 , \7851 , \7852 , \7853 ,
         \7854 , \7855 , \7856 , \7857 , \7858 , \7859 , \7860 , \7861 , \7862 , \7863 ,
         \7864 , \7865 , \7866 , \7867 , \7868 , \7869 , \7870 , \7871 , \7872 , \7873 ,
         \7874 , \7875 , \7876 , \7877 , \7878 , \7879 , \7880 , \7881 , \7882 , \7883 ,
         \7884 , \7885 , \7886 , \7887 , \7888 , \7889 , \7890 , \7891 , \7892 , \7893 ,
         \7894 , \7895 , \7896 , \7897 , \7898 , \7899 , \7900 , \7901 , \7902 , \7903 ,
         \7904 , \7905 , \7906 , \7907 , \7908 , \7909 , \7910 , \7911 , \7912 , \7913 ,
         \7914 , \7915 , \7916 , \7917 , \7918 , \7919 , \7920 , \7921 , \7922 , \7923 ,
         \7924 , \7925 , \7926 , \7927 , \7928 , \7929 , \7930 , \7931 , \7932 , \7933 ,
         \7934 , \7935 , \7936 , \7937 , \7938 , \7939 , \7940 , \7941 , \7942 , \7943 ,
         \7944 , \7945 , \7946 , \7947 , \7948 , \7949 , \7950 , \7951 , \7952 , \7953 ,
         \7954 , \7955 , \7956 , \7957 , \7958 , \7959 , \7960 , \7961 , \7962 , \7963 ,
         \7964 , \7965 , \7966 , \7967 , \7968 , \7969 , \7970 , \7971 , \7972 , \7973 ,
         \7974 , \7975 , \7976 , \7977 , \7978 , \7979 , \7980 , \7981 , \7982 , \7983 ,
         \7984 , \7985 , \7986 , \7987 , \7988 , \7989 , \7990 , \7991 , \7992 , \7993 ,
         \7994 , \7995 , \7996 , \7997 , \7998 , \7999 , \8000 , \8001 , \8002 , \8003 ,
         \8004 , \8005 , \8006 , \8007 , \8008 , \8009 , \8010 , \8011 , \8012 , \8013 ,
         \8014 , \8015 , \8016 , \8017 , \8018 , \8019 , \8020 , \8021 , \8022 , \8023 ,
         \8024 , \8025 , \8026 , \8027 , \8028 , \8029 , \8030 , \8031 , \8032 , \8033 ,
         \8034 , \8035 , \8036 , \8037 , \8038 , \8039 , \8040 , \8041 , \8042 , \8043 ,
         \8044 , \8045 , \8046 , \8047 , \8048 , \8049 , \8050 , \8051 , \8052 , \8053 ,
         \8054 , \8055 , \8056 , \8057 , \8058 , \8059 , \8060 , \8061 , \8062 , \8063 ,
         \8064 , \8065 , \8066 , \8067 , \8068 , \8069 , \8070 , \8071 , \8072 , \8073 ,
         \8074 , \8075 , \8076 , \8077 , \8078 , \8079 , \8080 , \8081 , \8082 , \8083 ,
         \8084 , \8085 , \8086 , \8087 , \8088 , \8089 , \8090 , \8091 , \8092 , \8093 ,
         \8094 , \8095 , \8096 , \8097 , \8098 , \8099 , \8100 , \8101 , \8102 , \8103 ,
         \8104 , \8105 , \8106 , \8107 , \8108 , \8109 , \8110 , \8111 , \8112 , \8113 ,
         \8114 , \8115 , \8116 , \8117 , \8118 , \8119 , \8120 , \8121 , \8122 , \8123 ,
         \8124 , \8125 , \8126 , \8127 , \8128 , \8129 , \8130 , \8131 , \8132 , \8133 ,
         \8134 , \8135 , \8136 , \8137 , \8138 , \8139 , \8140 , \8141 , \8142 , \8143 ,
         \8144 , \8145 , \8146 , \8147 , \8148 , \8149 , \8150 , \8151 , \8152 , \8153 ,
         \8154 , \8155 , \8156 , \8157 , \8158 , \8159 , \8160 , \8161 , \8162 , \8163 ,
         \8164 , \8165 , \8166 , \8167 , \8168 , \8169 , \8170 , \8171 , \8172 , \8173 ,
         \8174 , \8175 , \8176 , \8177 , \8178 , \8179 , \8180 , \8181 , \8182 , \8183 ,
         \8184 , \8185 , \8186 , \8187 , \8188 , \8189 , \8190 , \8191 , \8192 , \8193 ,
         \8194 , \8195 , \8196 , \8197 , \8198 , \8199 , \8200 , \8201 , \8202 , \8203 ,
         \8204 , \8205 , \8206 , \8207 , \8208 , \8209 , \8210 , \8211 , \8212 , \8213 ,
         \8214 , \8215 , \8216 , \8217 , \8218 , \8219 , \8220 , \8221 , \8222 , \8223 ,
         \8224 , \8225 , \8226 , \8227 , \8228 , \8229 , \8230 , \8231 , \8232 , \8233 ,
         \8234 , \8235 , \8236 , \8237 , \8238 , \8239 , \8240 , \8241 , \8242 , \8243 ,
         \8244 , \8245 , \8246 , \8247 , \8248 , \8249 , \8250 , \8251 , \8252 , \8253 ,
         \8254 , \8255 , \8256 , \8257 , \8258 , \8259 , \8260 , \8261 , \8262 , \8263 ,
         \8264 , \8265 , \8266 , \8267 , \8268 , \8269 , \8270 , \8271 , \8272 , \8273 ,
         \8274 , \8275 , \8276 , \8277 , \8278 , \8279 , \8280 , \8281 , \8282 , \8283 ,
         \8284 , \8285 , \8286 , \8287 , \8288 , \8289 , \8290 , \8291 , \8292 , \8293 ,
         \8294 , \8295 , \8296 , \8297 , \8298 , \8299 , \8300 , \8301 , \8302 , \8303 ,
         \8304 , \8305 , \8306 , \8307 , \8308 , \8309 , \8310 , \8311 , \8312 , \8313 ,
         \8314 , \8315 , \8316 , \8317 , \8318 , \8319 , \8320 , \8321 , \8322 , \8323 ,
         \8324 , \8325 , \8326 , \8327 , \8328 , \8329 , \8330 , \8331 , \8332 , \8333 ,
         \8334 , \8335 , \8336 , \8337 , \8338 , \8339 , \8340 , \8341 , \8342 , \8343 ,
         \8344 , \8345 , \8346 , \8347 , \8348 , \8349 , \8350 , \8351 , \8352 , \8353 ,
         \8354 , \8355 , \8356 , \8357 , \8358 , \8359 , \8360 , \8361 , \8362 , \8363 ,
         \8364 , \8365 , \8366 , \8367 , \8368 , \8369 , \8370 , \8371 , \8372 , \8373 ,
         \8374 , \8375 , \8376 , \8377 , \8378 , \8379 , \8380 , \8381 , \8382 , \8383 ,
         \8384 , \8385 , \8386 , \8387 , \8388 , \8389 , \8390 , \8391 , \8392 , \8393 ,
         \8394 , \8395 , \8396 , \8397 , \8398 , \8399 , \8400 , \8401 , \8402 , \8403 ,
         \8404 , \8405 , \8406 , \8407 , \8408 , \8409 , \8410 , \8411 , \8412 , \8413 ,
         \8414 , \8415 , \8416 , \8417 , \8418 , \8419 , \8420 , \8421 , \8422 , \8423 ,
         \8424 , \8425 , \8426 , \8427 , \8428 , \8429 , \8430 , \8431 , \8432 , \8433 ,
         \8434 , \8435 , \8436 , \8437 , \8438 , \8439 , \8440 , \8441 , \8442 , \8443 ,
         \8444 , \8445 , \8446 , \8447 , \8448 , \8449 , \8450 , \8451 , \8452 , \8453 ,
         \8454 , \8455 , \8456 , \8457 , \8458 , \8459 , \8460 , \8461 , \8462 , \8463 ,
         \8464 , \8465 , \8466 , \8467 , \8468 , \8469 , \8470 , \8471 , \8472 , \8473 ,
         \8474 , \8475 , \8476 , \8477 , \8478 , \8479 , \8480 , \8481 , \8482 , \8483 ,
         \8484 , \8485 , \8486 , \8487 , \8488 , \8489 , \8490 , \8491 , \8492 , \8493 ,
         \8494 , \8495 , \8496 , \8497 , \8498 , \8499 , \8500 , \8501 , \8502 , \8503 ,
         \8504 , \8505 , \8506 , \8507 , \8508 , \8509 , \8510 , \8511 , \8512 , \8513 ,
         \8514 , \8515 , \8516 , \8517 , \8518 , \8519 , \8520 , \8521 , \8522 , \8523 ,
         \8524 , \8525 , \8526 , \8527 , \8528 , \8529 , \8530 , \8531 , \8532 , \8533 ,
         \8534 , \8535 , \8536 , \8537 , \8538 , \8539 , \8540 , \8541 , \8542 , \8543 ,
         \8544 , \8545 , \8546 , \8547 , \8548 , \8549 , \8550 , \8551 , \8552 , \8553 ,
         \8554 , \8555 , \8556 , \8557 , \8558 , \8559 , \8560 , \8561 , \8562 , \8563 ,
         \8564 , \8565 , \8566 , \8567 , \8568 , \8569 , \8570 , \8571 , \8572 , \8573 ,
         \8574 , \8575 , \8576 , \8577 , \8578 , \8579 , \8580 , \8581 , \8582 , \8583 ,
         \8584 , \8585 , \8586 , \8587 , \8588 , \8589 , \8590 , \8591 , \8592 , \8593 ,
         \8594 , \8595 , \8596 , \8597 , \8598 , \8599 , \8600 , \8601 , \8602 , \8603 ,
         \8604 , \8605 , \8606 , \8607 , \8608 , \8609 , \8610 , \8611 , \8612 , \8613 ,
         \8614 , \8615 , \8616 , \8617 , \8618 , \8619 , \8620 , \8621 , \8622 , \8623 ,
         \8624 , \8625 , \8626 , \8627 , \8628 , \8629 , \8630 , \8631 , \8632 , \8633 ,
         \8634 , \8635 , \8636 , \8637 , \8638 , \8639 , \8640 , \8641 , \8642 , \8643 ,
         \8644 , \8645 , \8646 , \8647 , \8648 , \8649 , \8650 , \8651 , \8652 , \8653 ,
         \8654 , \8655 , \8656 , \8657 , \8658 , \8659 , \8660 , \8661 , \8662 , \8663 ,
         \8664 , \8665 , \8666 , \8667 , \8668 , \8669 , \8670 , \8671 , \8672 , \8673 ,
         \8674 , \8675 , \8676 , \8677 , \8678 , \8679 , \8680 , \8681 , \8682 , \8683 ,
         \8684 , \8685 , \8686 , \8687 , \8688 , \8689 , \8690 , \8691 , \8692 , \8693 ,
         \8694 , \8695 , \8696 , \8697 , \8698 , \8699 , \8700 , \8701 , \8702 , \8703 ,
         \8704 , \8705 , \8706 , \8707 , \8708 , \8709 , \8710 , \8711 , \8712 , \8713 ,
         \8714 , \8715 , \8716 , \8717 , \8718 , \8719 , \8720 , \8721 , \8722 , \8723 ,
         \8724 , \8725 , \8726 , \8727 , \8728 , \8729 , \8730 , \8731 , \8732 , \8733 ,
         \8734 , \8735 , \8736 , \8737 , \8738 , \8739 , \8740 , \8741 , \8742 , \8743 ,
         \8744 , \8745 , \8746 , \8747 , \8748 , \8749 , \8750 , \8751 , \8752 , \8753 ,
         \8754 , \8755 , \8756 , \8757 , \8758 , \8759 , \8760 , \8761 , \8762 , \8763 ,
         \8764 , \8765 , \8766 , \8767 , \8768 , \8769 , \8770 , \8771 , \8772 , \8773 ,
         \8774 , \8775 , \8776 , \8777 , \8778 , \8779 , \8780 , \8781 , \8782 , \8783 ,
         \8784 , \8785 , \8786 , \8787 , \8788 , \8789 , \8790 , \8791 , \8792 , \8793 ,
         \8794 , \8795 , \8796 , \8797 , \8798 , \8799 , \8800 , \8801 , \8802 , \8803 ,
         \8804 , \8805 , \8806 , \8807 , \8808 , \8809 , \8810 , \8811 , \8812 , \8813 ,
         \8814 , \8815 , \8816 , \8817 , \8818 , \8819 , \8820 , \8821 , \8822 , \8823 ,
         \8824 , \8825 , \8826 , \8827 , \8828 , \8829 , \8830 , \8831 , \8832 , \8833 ,
         \8834 , \8835 , \8836 , \8837 , \8838 , \8839 , \8840 , \8841 , \8842 , \8843 ,
         \8844 , \8845 , \8846 , \8847 , \8848 , \8849 , \8850 , \8851 , \8852 , \8853 ,
         \8854 , \8855 , \8856 , \8857 , \8858 , \8859 , \8860 , \8861 , \8862 , \8863 ,
         \8864 , \8865 , \8866 , \8867 , \8868 , \8869 , \8870 , \8871 , \8872 , \8873 ,
         \8874 , \8875 , \8876 , \8877 , \8878 , \8879 , \8880 , \8881 , \8882 , \8883 ,
         \8884 , \8885 , \8886 , \8887 , \8888 , \8889 , \8890 , \8891 , \8892 , \8893 ,
         \8894 , \8895 , \8896 , \8897 , \8898 , \8899 , \8900 , \8901 , \8902 , \8903 ,
         \8904 , \8905 , \8906 , \8907 , \8908 , \8909 , \8910 , \8911 , \8912 , \8913 ,
         \8914 , \8915 , \8916 , \8917 , \8918 , \8919 , \8920 , \8921 , \8922 , \8923 ,
         \8924 , \8925 , \8926 , \8927 , \8928 , \8929 , \8930 , \8931 , \8932 , \8933 ,
         \8934 , \8935 , \8936 , \8937 , \8938 , \8939 , \8940 , \8941 , \8942 , \8943 ,
         \8944 , \8945 , \8946 , \8947 , \8948 , \8949 , \8950 , \8951 , \8952 , \8953 ,
         \8954 , \8955 , \8956 , \8957 , \8958 , \8959 , \8960 , \8961 , \8962 , \8963 ,
         \8964 , \8965 , \8966 , \8967 , \8968 , \8969 , \8970 , \8971 , \8972 , \8973 ,
         \8974 , \8975 , \8976 , \8977 , \8978 , \8979 , \8980 , \8981 , \8982 , \8983 ,
         \8984 , \8985 , \8986 , \8987 , \8988 , \8989 , \8990 , \8991 , \8992 , \8993 ,
         \8994 , \8995 , \8996 , \8997 , \8998 , \8999 , \9000 , \9001 , \9002 , \9003 ,
         \9004 , \9005 , \9006 , \9007 , \9008 , \9009 , \9010 , \9011 , \9012 , \9013 ,
         \9014 , \9015 , \9016 , \9017 , \9018 , \9019 , \9020 , \9021 , \9022 , \9023 ,
         \9024 , \9025 , \9026 , \9027 , \9028 , \9029 , \9030 , \9031 , \9032 , \9033 ,
         \9034 , \9035 , \9036 , \9037 , \9038 , \9039 , \9040 , \9041 , \9042 , \9043 ,
         \9044 , \9045 , \9046 , \9047 , \9048 , \9049 , \9050 , \9051 , \9052 , \9053 ,
         \9054 , \9055 , \9056 , \9057 , \9058 , \9059 , \9060 , \9061 , \9062 , \9063 ,
         \9064 , \9065 , \9066 , \9067 , \9068 , \9069 , \9070 , \9071 , \9072 , \9073 ,
         \9074 , \9075 , \9076 , \9077 , \9078 , \9079 , \9080 , \9081 , \9082 , \9083 ,
         \9084 , \9085 , \9086 , \9087 , \9088 , \9089 , \9090 , \9091 , \9092 , \9093 ,
         \9094 , \9095 , \9096 , \9097 , \9098 , \9099 , \9100 , \9101 , \9102 , \9103 ,
         \9104 , \9105 , \9106 , \9107 , \9108 , \9109 , \9110 , \9111 , \9112 , \9113 ,
         \9114 , \9115 , \9116 , \9117 , \9118 , \9119 , \9120 , \9121 , \9122 , \9123 ,
         \9124 , \9125 , \9126 , \9127 , \9128 , \9129 , \9130 , \9131 , \9132 , \9133 ,
         \9134 , \9135 , \9136 , \9137 , \9138 , \9139 , \9140 , \9141 , \9142 , \9143 ,
         \9144 , \9145 , \9146 , \9147 , \9148 , \9149 , \9150 , \9151 , \9152 , \9153 ,
         \9154 , \9155 , \9156 , \9157 , \9158 , \9159 , \9160 , \9161 , \9162 , \9163 ,
         \9164 , \9165 , \9166 , \9167 , \9168 , \9169 , \9170 , \9171 , \9172 , \9173 ,
         \9174 , \9175 , \9176 , \9177 , \9178 , \9179 , \9180 , \9181 , \9182 , \9183 ,
         \9184 , \9185 , \9186 , \9187 , \9188 , \9189 , \9190 , \9191 , \9192 , \9193 ,
         \9194 , \9195 , \9196 , \9197 , \9198 , \9199 , \9200 , \9201 , \9202 , \9203 ,
         \9204 , \9205 , \9206 , \9207 , \9208 , \9209 , \9210 , \9211 , \9212 , \9213 ,
         \9214 , \9215 , \9216 , \9217 , \9218 , \9219 , \9220 , \9221 , \9222 , \9223 ,
         \9224 , \9225 , \9226 , \9227 , \9228 , \9229 , \9230 , \9231 , \9232 , \9233 ,
         \9234 , \9235 , \9236 , \9237 , \9238 , \9239 , \9240 , \9241 , \9242 , \9243 ,
         \9244 , \9245 , \9246 , \9247 , \9248 , \9249 , \9250 , \9251 , \9252 , \9253 ,
         \9254 , \9255 , \9256 , \9257 , \9258 , \9259 , \9260 , \9261 , \9262 , \9263 ,
         \9264 , \9265 , \9266 , \9267 , \9268 , \9269 , \9270 , \9271 , \9272 , \9273 ,
         \9274 , \9275 , \9276 , \9277 , \9278 , \9279 , \9280 , \9281 , \9282 , \9283 ,
         \9284 , \9285 , \9286 , \9287 , \9288 , \9289 , \9290 , \9291 , \9292 , \9293 ,
         \9294 , \9295 , \9296 , \9297 , \9298 , \9299 , \9300 , \9301 , \9302 , \9303 ,
         \9304 , \9305 , \9306 , \9307 , \9308 , \9309 , \9310 , \9311 , \9312 , \9313 ,
         \9314 , \9315 , \9316 , \9317 , \9318 , \9319 , \9320 , \9321 , \9322 , \9323 ,
         \9324 , \9325 , \9326 , \9327 , \9328 , \9329 , \9330 , \9331 , \9332 , \9333 ,
         \9334 , \9335 , \9336 , \9337 , \9338 , \9339 , \9340 , \9341 , \9342 , \9343 ,
         \9344 , \9345 , \9346 , \9347 , \9348 , \9349 , \9350 , \9351 , \9352 , \9353 ,
         \9354 , \9355 , \9356 , \9357 , \9358 , \9359 , \9360 , \9361 , \9362 , \9363 ,
         \9364 , \9365 , \9366 , \9367 , \9368 , \9369 , \9370 , \9371 , \9372 , \9373 ,
         \9374 , \9375 , \9376 , \9377 , \9378 , \9379 , \9380 , \9381 , \9382 , \9383 ,
         \9384 , \9385 , \9386 , \9387 , \9388 , \9389 , \9390 , \9391 , \9392 , \9393 ,
         \9394 , \9395 , \9396 , \9397 , \9398 , \9399 , \9400 , \9401 , \9402 , \9403 ,
         \9404 , \9405 , \9406 , \9407 , \9408 , \9409 , \9410 , \9411 , \9412 , \9413 ,
         \9414 , \9415 , \9416 , \9417 , \9418 , \9419 , \9420 , \9421 , \9422 , \9423 ,
         \9424 , \9425 , \9426 , \9427 , \9428 , \9429 , \9430 , \9431 , \9432 , \9433 ,
         \9434 , \9435 , \9436 , \9437 , \9438 , \9439 , \9440 , \9441 , \9442 , \9443 ,
         \9444 , \9445 , \9446 , \9447 , \9448 , \9449 , \9450 , \9451 , \9452 , \9453 ,
         \9454 , \9455 , \9456 , \9457 , \9458 , \9459 , \9460 , \9461 , \9462 , \9463 ,
         \9464 , \9465 , \9466 , \9467 , \9468 , \9469 , \9470 , \9471 , \9472 , \9473 ,
         \9474 , \9475 , \9476 , \9477 , \9478 , \9479 , \9480 , \9481 , \9482 , \9483 ,
         \9484 , \9485 , \9486 , \9487 , \9488 , \9489 , \9490 , \9491 , \9492 , \9493 ,
         \9494 , \9495 , \9496 , \9497 , \9498 , \9499 , \9500 , \9501 , \9502 , \9503 ,
         \9504 , \9505 , \9506 , \9507 , \9508 , \9509 , \9510 , \9511 , \9512 , \9513 ,
         \9514 , \9515 , \9516 , \9517 , \9518 , \9519 , \9520 , \9521 , \9522 , \9523 ,
         \9524 , \9525 , \9526 , \9527 , \9528 , \9529 , \9530 , \9531 , \9532 , \9533 ,
         \9534 , \9535 , \9536 , \9537 , \9538 , \9539 , \9540 , \9541 , \9542 , \9543 ,
         \9544 , \9545 , \9546 , \9547 , \9548 , \9549 , \9550 , \9551 , \9552 , \9553 ,
         \9554 , \9555 , \9556 , \9557 , \9558 , \9559 , \9560 , \9561 , \9562 , \9563 ,
         \9564 , \9565 , \9566 , \9567 , \9568 , \9569 , \9570 , \9571 , \9572 , \9573 ,
         \9574 , \9575 , \9576 , \9577 , \9578 , \9579 , \9580 , \9581 , \9582 , \9583 ,
         \9584 , \9585 , \9586 , \9587 , \9588 , \9589 , \9590 , \9591 , \9592 , \9593 ,
         \9594 , \9595 , \9596 , \9597 , \9598 , \9599 , \9600 , \9601 , \9602 , \9603 ,
         \9604 , \9605 , \9606 , \9607 , \9608 , \9609 , \9610 , \9611 , \9612 , \9613 ,
         \9614 , \9615 , \9616 , \9617 , \9618 , \9619 , \9620 , \9621 , \9622 , \9623 ,
         \9624 , \9625 , \9626 , \9627 , \9628 , \9629 , \9630 , \9631 , \9632 , \9633 ,
         \9634 , \9635 , \9636 , \9637 , \9638 , \9639 , \9640 , \9641 , \9642 , \9643 ,
         \9644 , \9645 , \9646 , \9647 , \9648 , \9649 , \9650 , \9651 , \9652 , \9653 ,
         \9654 , \9655 , \9656 , \9657 , \9658 , \9659 , \9660 , \9661 , \9662 , \9663 ,
         \9664 , \9665 , \9666 , \9667 , \9668 , \9669 , \9670 , \9671 , \9672 , \9673 ,
         \9674 , \9675 , \9676 , \9677 , \9678 , \9679 , \9680 , \9681 , \9682 , \9683 ,
         \9684 , \9685 , \9686 , \9687 , \9688 , \9689 , \9690 , \9691 , \9692 , \9693 ,
         \9694 , \9695 , \9696 , \9697 , \9698 , \9699 , \9700 , \9701 , \9702 , \9703 ,
         \9704 , \9705 , \9706 , \9707 , \9708 , \9709 , \9710 , \9711 , \9712 , \9713 ,
         \9714 , \9715 , \9716 , \9717 , \9718 , \9719 , \9720 , \9721 , \9722 , \9723 ,
         \9724 , \9725 , \9726 , \9727 , \9728 , \9729 , \9730 , \9731 , \9732 , \9733 ,
         \9734 , \9735 , \9736 , \9737 , \9738 , \9739 , \9740 , \9741 , \9742 , \9743 ,
         \9744 , \9745 , \9746 , \9747 , \9748 , \9749 , \9750 , \9751 , \9752 , \9753 ,
         \9754 , \9755 , \9756 , \9757 , \9758 , \9759 , \9760 , \9761 , \9762 , \9763 ,
         \9764 , \9765 , \9766 , \9767 , \9768 , \9769 , \9770 , \9771 , \9772 , \9773 ,
         \9774 , \9775 , \9776 , \9777 , \9778 , \9779 , \9780 , \9781 , \9782 , \9783 ,
         \9784 , \9785 , \9786 , \9787 , \9788 , \9789 , \9790 , \9791 , \9792 , \9793 ,
         \9794 , \9795 , \9796 , \9797 , \9798 , \9799 , \9800 , \9801 , \9802 , \9803 ,
         \9804 , \9805 , \9806 , \9807 , \9808 , \9809 , \9810 , \9811 , \9812 , \9813 ,
         \9814 , \9815 , \9816 , \9817 , \9818 , \9819 , \9820 , \9821 , \9822 , \9823 ,
         \9824 , \9825 , \9826 , \9827 , \9828 , \9829 , \9830 , \9831 , \9832 , \9833 ,
         \9834 , \9835 , \9836 , \9837 , \9838 , \9839 , \9840 , \9841 , \9842 , \9843 ,
         \9844 , \9845 , \9846 , \9847 , \9848 , \9849 , \9850 , \9851 , \9852 , \9853 ,
         \9854 , \9855 , \9856 , \9857 , \9858 , \9859 , \9860 , \9861 , \9862 , \9863 ,
         \9864 , \9865 , \9866 , \9867 , \9868 , \9869 , \9870 , \9871 , \9872 , \9873 ,
         \9874 , \9875 , \9876 , \9877 , \9878 , \9879 , \9880 , \9881 , \9882 , \9883 ,
         \9884 , \9885 , \9886 , \9887 , \9888 , \9889 , \9890 , \9891 , \9892 , \9893 ,
         \9894 , \9895 , \9896 , \9897 , \9898 , \9899 , \9900 , \9901 , \9902 , \9903 ,
         \9904 , \9905 , \9906 , \9907 , \9908 , \9909 , \9910 , \9911 , \9912 , \9913 ,
         \9914 , \9915 , \9916 , \9917 , \9918 , \9919 , \9920 , \9921 , \9922 , \9923 ,
         \9924 , \9925 , \9926 , \9927 , \9928 , \9929 , \9930 , \9931 , \9932 , \9933 ,
         \9934 , \9935 , \9936 , \9937 , \9938 , \9939 , \9940 , \9941 , \9942 , \9943 ,
         \9944 , \9945 , \9946 , \9947 , \9948 , \9949 , \9950 , \9951 , \9952 , \9953 ,
         \9954 , \9955 , \9956 , \9957 , \9958 , \9959 , \9960 , \9961 , \9962 , \9963 ,
         \9964 , \9965 , \9966 , \9967 , \9968 , \9969 , \9970 , \9971 , \9972 , \9973 ,
         \9974 , \9975 , \9976 , \9977 , \9978 , \9979 , \9980 , \9981 , \9982 , \9983 ,
         \9984 , \9985 , \9986 , \9987 , \9988 , \9989 , \9990 , \9991 , \9992 , \9993 ,
         \9994 , \9995 , \9996 , \9997 , \9998 , \9999 , \10000 , \10001 , \10002 , \10003 ,
         \10004 , \10005 , \10006 , \10007 , \10008 , \10009 , \10010 , \10011 , \10012 , \10013 ,
         \10014 , \10015 , \10016 , \10017 , \10018 , \10019 , \10020 , \10021 , \10022 , \10023 ,
         \10024 , \10025 , \10026 , \10027 , \10028 , \10029 , \10030 , \10031 , \10032 , \10033 ,
         \10034 , \10035 , \10036 , \10037 , \10038 , \10039 , \10040 , \10041 , \10042 , \10043 ,
         \10044 , \10045 , \10046 , \10047 , \10048 , \10049 , \10050 , \10051 , \10052 , \10053 ,
         \10054 , \10055 , \10056 , \10057 , \10058 , \10059 , \10060 , \10061 , \10062 , \10063 ,
         \10064 , \10065 , \10066 , \10067 , \10068 , \10069 , \10070 , \10071 , \10072 , \10073 ,
         \10074 , \10075 , \10076 , \10077 , \10078 , \10079 , \10080 , \10081 , \10082 , \10083 ,
         \10084 , \10085 , \10086 , \10087 , \10088 , \10089 , \10090 , \10091 , \10092 , \10093 ,
         \10094 , \10095 , \10096 , \10097 , \10098 , \10099 , \10100 , \10101 , \10102 , \10103 ,
         \10104 , \10105 , \10106 , \10107 , \10108 , \10109 , \10110 , \10111 , \10112 , \10113 ,
         \10114 , \10115 , \10116 , \10117 , \10118 , \10119 , \10120 , \10121 , \10122 , \10123 ,
         \10124 , \10125 , \10126 , \10127 , \10128 , \10129 , \10130 , \10131 , \10132 , \10133 ,
         \10134 , \10135 , \10136 , \10137 , \10138 , \10139 , \10140 , \10141 , \10142 , \10143 ,
         \10144 , \10145 , \10146 , \10147 , \10148 , \10149 , \10150 , \10151 , \10152 , \10153 ,
         \10154 , \10155 , \10156 , \10157 , \10158 , \10159 , \10160 , \10161 , \10162 , \10163 ,
         \10164 , \10165 , \10166 , \10167 , \10168 , \10169 , \10170 , \10171 , \10172 , \10173 ,
         \10174 , \10175 , \10176 , \10177 , \10178 , \10179 , \10180 , \10181 , \10182 , \10183 ,
         \10184 , \10185 , \10186 , \10187 , \10188 , \10189 , \10190 , \10191 , \10192 , \10193 ,
         \10194 , \10195 , \10196 , \10197 , \10198 , \10199 , \10200 , \10201 , \10202 , \10203 ,
         \10204 , \10205 , \10206 , \10207 , \10208 , \10209 , \10210 , \10211 , \10212 , \10213 ,
         \10214 , \10215 , \10216 , \10217 , \10218 , \10219 , \10220 , \10221 , \10222 , \10223 ,
         \10224 , \10225 , \10226 , \10227 , \10228 , \10229 , \10230 , \10231 , \10232 , \10233 ,
         \10234 , \10235 , \10236 , \10237 , \10238 , \10239 , \10240 , \10241 , \10242 , \10243 ,
         \10244 , \10245 , \10246 , \10247 , \10248 , \10249 , \10250 , \10251 , \10252 , \10253 ,
         \10254 , \10255 , \10256 , \10257 , \10258 , \10259 , \10260 , \10261 , \10262 , \10263 ,
         \10264 , \10265 , \10266 , \10267 , \10268 , \10269 , \10270 , \10271 , \10272 , \10273 ,
         \10274 , \10275 , \10276 , \10277 , \10278 , \10279 , \10280 , \10281 , \10282 , \10283 ,
         \10284 , \10285 , \10286 , \10287 , \10288 , \10289 , \10290 , \10291 , \10292 , \10293 ,
         \10294 , \10295 , \10296 , \10297 , \10298 , \10299 , \10300 , \10301 , \10302 , \10303 ,
         \10304 , \10305 , \10306 , \10307 , \10308 , \10309 , \10310 , \10311 , \10312 , \10313 ,
         \10314 , \10315 , \10316 , \10317 , \10318 , \10319 , \10320 , \10321 , \10322 , \10323 ,
         \10324 , \10325 , \10326 , \10327 , \10328 , \10329 , \10330 , \10331 , \10332 , \10333 ,
         \10334 , \10335 , \10336 , \10337 , \10338 , \10339 , \10340 , \10341 , \10342 , \10343 ,
         \10344 , \10345 , \10346 , \10347 , \10348 , \10349 , \10350 , \10351 , \10352 , \10353 ,
         \10354 , \10355 , \10356 , \10357 , \10358 , \10359 , \10360 , \10361 , \10362 , \10363 ,
         \10364 , \10365 , \10366 , \10367 , \10368 , \10369 , \10370 , \10371 , \10372 , \10373 ,
         \10374 , \10375 , \10376 , \10377 , \10378 , \10379 , \10380 , \10381 , \10382 , \10383 ,
         \10384 , \10385 , \10386 , \10387 , \10388 , \10389 , \10390 , \10391 , \10392 , \10393 ,
         \10394 , \10395 , \10396 , \10397 , \10398 , \10399 , \10400 , \10401 , \10402 , \10403 ,
         \10404 , \10405 , \10406 , \10407 , \10408 , \10409 , \10410 , \10411 , \10412 , \10413 ,
         \10414 , \10415 , \10416 , \10417 , \10418 , \10419 , \10420 , \10421 , \10422 , \10423 ,
         \10424 , \10425 , \10426 , \10427 , \10428 , \10429 , \10430 , \10431 , \10432 , \10433 ,
         \10434 , \10435 , \10436 , \10437 , \10438 , \10439 , \10440 , \10441 , \10442 , \10443 ,
         \10444 , \10445 , \10446 , \10447 , \10448 , \10449 , \10450 , \10451 , \10452 , \10453 ,
         \10454 , \10455 , \10456 , \10457 , \10458 , \10459 , \10460 , \10461 , \10462 , \10463 ,
         \10464 , \10465 , \10466 , \10467 , \10468 , \10469 , \10470 , \10471 , \10472 , \10473 ,
         \10474 , \10475 , \10476 , \10477 , \10478 , \10479 , \10480 , \10481 , \10482 , \10483 ,
         \10484 , \10485 , \10486 , \10487 , \10488 , \10489 , \10490 , \10491 , \10492 , \10493 ,
         \10494 , \10495 , \10496 , \10497 , \10498 , \10499 , \10500 , \10501 , \10502 , \10503 ,
         \10504 , \10505 , \10506 , \10507 , \10508 , \10509 , \10510 , \10511 , \10512 , \10513 ,
         \10514 , \10515 , \10516 , \10517 , \10518 , \10519 , \10520 , \10521 , \10522 , \10523 ,
         \10524 , \10525 , \10526 , \10527 , \10528 , \10529 , \10530 , \10531 , \10532 , \10533 ,
         \10534 , \10535 , \10536 , \10537 , \10538 , \10539 , \10540 , \10541 , \10542 , \10543 ,
         \10544 , \10545 , \10546 , \10547 , \10548 , \10549 , \10550 , \10551 , \10552 , \10553 ,
         \10554 , \10555 , \10556 , \10557 , \10558 , \10559 , \10560 , \10561 , \10562 , \10563 ,
         \10564 , \10565 , \10566 , \10567 , \10568 , \10569 , \10570 , \10571 , \10572 , \10573 ,
         \10574 , \10575 , \10576 , \10577 , \10578 , \10579 , \10580 , \10581 , \10582 , \10583 ,
         \10584 , \10585 , \10586 , \10587 , \10588 , \10589 , \10590 , \10591 , \10592 , \10593 ,
         \10594 , \10595 , \10596 , \10597 , \10598 , \10599 , \10600 , \10601 , \10602 , \10603 ,
         \10604 , \10605 , \10606 , \10607 , \10608 , \10609 , \10610 , \10611 , \10612 , \10613 ,
         \10614 , \10615 , \10616 , \10617 , \10618 , \10619 , \10620 , \10621 , \10622 , \10623 ,
         \10624 , \10625 , \10626 , \10627 , \10628 , \10629 , \10630 , \10631 , \10632 , \10633 ,
         \10634 , \10635 , \10636 , \10637 , \10638 , \10639 , \10640 , \10641 , \10642 , \10643 ,
         \10644 , \10645 , \10646 , \10647 , \10648 , \10649 , \10650 , \10651 , \10652 , \10653 ,
         \10654 , \10655 , \10656 , \10657 , \10658 , \10659 , \10660 , \10661 , \10662 , \10663 ,
         \10664 , \10665 , \10666 , \10667 , \10668 , \10669 , \10670 , \10671 , \10672 , \10673 ,
         \10674 , \10675 , \10676 , \10677 , \10678 , \10679 , \10680 , \10681 , \10682 , \10683 ,
         \10684 , \10685 , \10686 , \10687 , \10688 , \10689 , \10690 , \10691 , \10692 , \10693 ,
         \10694 , \10695 , \10696 , \10697 , \10698 , \10699 , \10700 , \10701 , \10702 , \10703 ,
         \10704 , \10705 , \10706 , \10707 , \10708 , \10709 , \10710 , \10711 , \10712 , \10713 ,
         \10714 , \10715 , \10716 , \10717 , \10718 , \10719 , \10720 , \10721 , \10722 , \10723 ,
         \10724 , \10725 , \10726 , \10727 , \10728 , \10729 , \10730 , \10731 , \10732 , \10733 ,
         \10734 , \10735 , \10736 , \10737 , \10738 , \10739 , \10740 , \10741 , \10742 , \10743 ,
         \10744 , \10745 , \10746 , \10747 , \10748 , \10749 , \10750 , \10751 , \10752 , \10753 ,
         \10754 , \10755 , \10756 , \10757 , \10758 , \10759 , \10760 , \10761 , \10762 , \10763 ,
         \10764 , \10765 , \10766 , \10767 , \10768 , \10769 , \10770 , \10771 , \10772 , \10773 ,
         \10774 , \10775 , \10776 , \10777 , \10778 , \10779 , \10780 , \10781 , \10782 , \10783 ,
         \10784 , \10785 , \10786 , \10787 , \10788 , \10789 , \10790 , \10791 , \10792 , \10793 ,
         \10794 , \10795 , \10796 , \10797 , \10798 , \10799 , \10800 , \10801 , \10802 , \10803 ,
         \10804 , \10805 , \10806 , \10807 , \10808 , \10809 , \10810 , \10811 , \10812 , \10813 ,
         \10814 , \10815 , \10816 , \10817 , \10818 , \10819 , \10820 , \10821 , \10822 , \10823 ,
         \10824 , \10825 , \10826 , \10827 , \10828 , \10829 , \10830 , \10831 , \10832 , \10833 ,
         \10834 , \10835 , \10836 , \10837 , \10838 , \10839 , \10840 , \10841 , \10842 , \10843 ,
         \10844 , \10845 , \10846 , \10847 , \10848 , \10849 , \10850 , \10851 , \10852 , \10853 ,
         \10854 , \10855 , \10856 , \10857 , \10858 , \10859 , \10860 , \10861 , \10862 , \10863 ,
         \10864 , \10865 , \10866 , \10867 , \10868 , \10869 , \10870 , \10871 , \10872 , \10873 ,
         \10874 , \10875 , \10876 , \10877 , \10878 , \10879 , \10880 , \10881 , \10882 , \10883 ,
         \10884 , \10885 , \10886 , \10887 , \10888 , \10889 , \10890 , \10891 , \10892 , \10893 ,
         \10894 , \10895 , \10896 , \10897 , \10898 , \10899 , \10900 , \10901 , \10902 , \10903 ,
         \10904 , \10905 , \10906 , \10907 , \10908 , \10909 , \10910 , \10911 , \10912 , \10913 ,
         \10914 , \10915 , \10916 , \10917 , \10918 , \10919 , \10920 , \10921 , \10922 , \10923 ,
         \10924 , \10925 , \10926 , \10927 , \10928 , \10929 , \10930 , \10931 , \10932 , \10933 ,
         \10934 , \10935 , \10936 , \10937 , \10938 , \10939 , \10940 , \10941 , \10942 , \10943 ,
         \10944 , \10945 , \10946 , \10947 , \10948 , \10949 , \10950 , \10951 , \10952 , \10953 ,
         \10954 , \10955 , \10956 , \10957 , \10958 , \10959 , \10960 , \10961 , \10962 , \10963 ,
         \10964 , \10965 , \10966 , \10967 , \10968 , \10969 , \10970 , \10971 , \10972 , \10973 ,
         \10974 , \10975 , \10976 , \10977 , \10978 , \10979 , \10980 , \10981 , \10982 , \10983 ,
         \10984 , \10985 , \10986 , \10987 , \10988 , \10989 , \10990 , \10991 , \10992 , \10993 ,
         \10994 , \10995 , \10996 , \10997 , \10998 , \10999 , \11000 , \11001 , \11002 , \11003 ,
         \11004 , \11005 , \11006 , \11007 , \11008 , \11009 , \11010 , \11011 , \11012 , \11013 ,
         \11014 , \11015 , \11016 , \11017 , \11018 , \11019 , \11020 , \11021 , \11022 , \11023 ,
         \11024 , \11025 , \11026 , \11027 , \11028 , \11029 , \11030 , \11031 , \11032 , \11033 ,
         \11034 , \11035 , \11036 , \11037 , \11038 , \11039 , \11040 , \11041 , \11042 , \11043 ,
         \11044 , \11045 , \11046 , \11047 , \11048 , \11049 , \11050 , \11051 , \11052 , \11053 ,
         \11054 , \11055 , \11056 , \11057 , \11058 , \11059 , \11060 , \11061 , \11062 , \11063 ,
         \11064 , \11065 , \11066 , \11067 , \11068 , \11069 , \11070 , \11071 , \11072 , \11073 ,
         \11074 , \11075 , \11076 , \11077 , \11078 , \11079 , \11080 , \11081 , \11082 , \11083 ,
         \11084 , \11085 , \11086 , \11087 , \11088 , \11089 , \11090 , \11091 , \11092 , \11093 ,
         \11094 , \11095 , \11096 , \11097 , \11098 , \11099 , \11100 , \11101 , \11102 , \11103 ,
         \11104 , \11105 , \11106 , \11107 , \11108 , \11109 , \11110 , \11111 , \11112 , \11113 ,
         \11114 , \11115 , \11116 , \11117 , \11118 , \11119 , \11120 , \11121 , \11122 , \11123 ,
         \11124 , \11125 , \11126 , \11127 , \11128 , \11129 , \11130 , \11131 , \11132 , \11133 ,
         \11134 , \11135 , \11136 , \11137 , \11138 , \11139 , \11140 , \11141 , \11142 , \11143 ,
         \11144 , \11145 , \11146 , \11147 , \11148 , \11149 , \11150 , \11151 , \11152 , \11153 ,
         \11154 , \11155 , \11156 , \11157 , \11158 , \11159 , \11160 , \11161 , \11162 , \11163 ,
         \11164 , \11165 , \11166 , \11167 , \11168 , \11169 , \11170 , \11171 , \11172 , \11173 ,
         \11174 , \11175 , \11176 , \11177 , \11178 , \11179 , \11180 , \11181 , \11182 , \11183 ,
         \11184 , \11185 , \11186 , \11187 , \11188 , \11189 , \11190 , \11191 , \11192 , \11193 ,
         \11194 , \11195 , \11196 , \11197 , \11198 , \11199 , \11200 , \11201 , \11202 , \11203 ,
         \11204 , \11205 , \11206 , \11207 , \11208 , \11209 , \11210 , \11211 , \11212 , \11213 ,
         \11214 , \11215 , \11216 , \11217 , \11218 , \11219 , \11220 , \11221 , \11222 , \11223 ,
         \11224 , \11225 , \11226 , \11227 , \11228 , \11229 , \11230 , \11231 , \11232 , \11233 ,
         \11234 , \11235 , \11236 , \11237 , \11238 , \11239 , \11240 , \11241 , \11242 , \11243 ,
         \11244 , \11245 , \11246 , \11247 , \11248 , \11249 , \11250 , \11251 , \11252 , \11253 ,
         \11254 , \11255 , \11256 , \11257 , \11258 , \11259 , \11260 , \11261 , \11262 , \11263 ,
         \11264 , \11265 , \11266 , \11267 , \11268 , \11269 , \11270 , \11271 , \11272 , \11273 ,
         \11274 , \11275 , \11276 , \11277 , \11278 , \11279 , \11280 , \11281 , \11282 , \11283 ,
         \11284 , \11285 , \11286 , \11287 , \11288 , \11289 , \11290 , \11291 , \11292 , \11293 ,
         \11294 , \11295 , \11296 , \11297 , \11298 , \11299 , \11300 , \11301 , \11302 , \11303 ,
         \11304 , \11305 , \11306 , \11307 , \11308 , \11309 , \11310 , \11311 , \11312 , \11313 ,
         \11314 , \11315 , \11316 , \11317 , \11318 , \11319 , \11320 , \11321 , \11322 , \11323 ,
         \11324 , \11325 , \11326 , \11327 , \11328 , \11329 , \11330 , \11331 , \11332 , \11333 ,
         \11334 , \11335 , \11336 , \11337 , \11338 , \11339 , \11340 , \11341 , \11342 , \11343 ,
         \11344 , \11345 , \11346 , \11347 , \11348 , \11349 , \11350 , \11351 , \11352 , \11353 ,
         \11354 , \11355 , \11356 , \11357 , \11358 , \11359 , \11360 , \11361 , \11362 , \11363 ,
         \11364 , \11365 , \11366 , \11367 , \11368 , \11369 , \11370 , \11371 , \11372 , \11373 ,
         \11374 , \11375 , \11376 , \11377 , \11378 , \11379 , \11380 , \11381 , \11382 , \11383 ,
         \11384 , \11385 , \11386 , \11387 , \11388 , \11389 , \11390 , \11391 , \11392 , \11393 ,
         \11394 , \11395 , \11396 , \11397 , \11398 , \11399 , \11400 , \11401 , \11402 , \11403 ,
         \11404 , \11405 , \11406 , \11407 , \11408 , \11409 , \11410 , \11411 , \11412 , \11413 ,
         \11414 , \11415 , \11416 , \11417 , \11418 , \11419 , \11420 , \11421 , \11422 , \11423 ,
         \11424 , \11425 , \11426 , \11427 , \11428 , \11429 , \11430 , \11431 , \11432 , \11433 ,
         \11434 , \11435 , \11436 , \11437 , \11438 , \11439 , \11440 , \11441 , \11442 , \11443 ,
         \11444 , \11445 , \11446 , \11447 , \11448 , \11449 , \11450 , \11451 , \11452 , \11453 ,
         \11454 , \11455 , \11456 , \11457 , \11458 , \11459 , \11460 , \11461 , \11462 , \11463 ,
         \11464 , \11465 , \11466 , \11467 , \11468 , \11469 , \11470 , \11471 , \11472 , \11473 ,
         \11474 , \11475 , \11476 , \11477 , \11478 , \11479 , \11480 , \11481 , \11482 , \11483 ,
         \11484 , \11485 , \11486 , \11487 , \11488 , \11489 , \11490 , \11491 , \11492 , \11493 ,
         \11494 , \11495 , \11496 , \11497 , \11498 , \11499 , \11500 , \11501 , \11502 , \11503 ,
         \11504 , \11505 , \11506 , \11507 , \11508 , \11509 , \11510 , \11511 , \11512 , \11513 ,
         \11514 , \11515 , \11516 , \11517 , \11518 , \11519 , \11520 , \11521 , \11522 , \11523 ,
         \11524 , \11525 , \11526 , \11527 , \11528 , \11529 , \11530 , \11531 , \11532 , \11533 ,
         \11534 , \11535 , \11536 , \11537 , \11538 , \11539 , \11540 , \11541 , \11542 , \11543 ,
         \11544 , \11545 , \11546 , \11547 , \11548 , \11549 , \11550 , \11551 , \11552 , \11553 ,
         \11554 , \11555 , \11556 , \11557 , \11558 , \11559 , \11560 , \11561 , \11562 , \11563 ,
         \11564 , \11565 , \11566 , \11567 , \11568 , \11569 , \11570 , \11571 , \11572 , \11573 ,
         \11574 , \11575 , \11576 , \11577 , \11578 , \11579 , \11580 , \11581 , \11582 , \11583 ,
         \11584 , \11585 , \11586 , \11587 , \11588 , \11589 , \11590 , \11591 , \11592 , \11593 ,
         \11594 , \11595 , \11596 , \11597 , \11598 , \11599 , \11600 , \11601 , \11602 , \11603 ,
         \11604 , \11605 , \11606 , \11607 , \11608 , \11609 , \11610 , \11611 , \11612 , \11613 ,
         \11614 , \11615 , \11616 , \11617 , \11618 , \11619 , \11620 , \11621 , \11622 , \11623 ,
         \11624 , \11625 , \11626 , \11627 , \11628 , \11629 , \11630 , \11631 , \11632 , \11633 ,
         \11634 , \11635 , \11636 , \11637 , \11638 , \11639 , \11640 , \11641 , \11642 , \11643 ,
         \11644 , \11645 , \11646 , \11647 , \11648 , \11649 , \11650 , \11651 , \11652 , \11653 ,
         \11654 , \11655 , \11656 , \11657 , \11658 , \11659 , \11660 , \11661 , \11662 , \11663 ,
         \11664 , \11665 , \11666 , \11667 , \11668 , \11669 , \11670 , \11671 , \11672 , \11673 ,
         \11674 , \11675 , \11676 , \11677 , \11678 , \11679 , \11680 , \11681 , \11682 , \11683 ,
         \11684 , \11685 , \11686 , \11687 , \11688 , \11689 , \11690 , \11691 , \11692 , \11693 ,
         \11694 , \11695 , \11696 , \11697 , \11698 , \11699 , \11700 , \11701 , \11702 , \11703 ,
         \11704 , \11705 , \11706 , \11707 , \11708 , \11709 , \11710 , \11711 , \11712 , \11713 ,
         \11714 , \11715 , \11716 , \11717 , \11718 , \11719 , \11720 , \11721 , \11722 , \11723 ,
         \11724 , \11725 , \11726 , \11727 , \11728 , \11729 , \11730 , \11731 , \11732 , \11733 ,
         \11734 , \11735 , \11736 , \11737 , \11738 , \11739 , \11740 , \11741 , \11742 , \11743 ,
         \11744 , \11745 , \11746 , \11747 , \11748 , \11749 , \11750 , \11751 , \11752 , \11753 ,
         \11754 , \11755 , \11756 , \11757 , \11758 , \11759 , \11760 , \11761 , \11762 , \11763 ,
         \11764 , \11765 , \11766 , \11767 , \11768 , \11769 , \11770 , \11771 , \11772 , \11773 ,
         \11774 , \11775 , \11776 , \11777 , \11778 , \11779 , \11780 , \11781 , \11782 , \11783 ,
         \11784 , \11785 , \11786 , \11787 , \11788 , \11789 , \11790 , \11791 , \11792 , \11793 ,
         \11794 , \11795 , \11796 , \11797 , \11798 , \11799 , \11800 , \11801 , \11802 , \11803 ,
         \11804 , \11805 , \11806 , \11807 , \11808 , \11809 , \11810 , \11811 , \11812 , \11813 ,
         \11814 , \11815 , \11816 , \11817 , \11818 , \11819 , \11820 , \11821 , \11822 , \11823 ,
         \11824 , \11825 , \11826 , \11827 , \11828 , \11829 , \11830 , \11831 , \11832 , \11833 ,
         \11834 , \11835 , \11836 , \11837 , \11838 , \11839 , \11840 , \11841 , \11842 , \11843 ,
         \11844 , \11845 , \11846 , \11847 , \11848 , \11849 , \11850 , \11851 , \11852 , \11853 ,
         \11854 , \11855 , \11856 , \11857 , \11858 , \11859 , \11860 , \11861 , \11862 , \11863 ,
         \11864 , \11865 , \11866 , \11867 , \11868 , \11869 , \11870 , \11871 , \11872 , \11873 ,
         \11874 , \11875 , \11876 , \11877 , \11878 , \11879 , \11880 , \11881 , \11882 , \11883 ,
         \11884 , \11885 , \11886 , \11887 , \11888 , \11889 , \11890 , \11891 , \11892 , \11893 ,
         \11894 , \11895 , \11896 , \11897 , \11898 , \11899 , \11900 , \11901 , \11902 , \11903 ,
         \11904 , \11905 , \11906 , \11907 , \11908 , \11909 , \11910 , \11911 , \11912 , \11913 ,
         \11914 , \11915 , \11916 , \11917 , \11918 , \11919 , \11920 , \11921 , \11922 , \11923 ,
         \11924 , \11925 , \11926 , \11927 , \11928 , \11929 , \11930 , \11931 , \11932 , \11933 ,
         \11934 , \11935 , \11936 , \11937 , \11938 , \11939 , \11940 , \11941 , \11942 , \11943 ,
         \11944 , \11945 , \11946 , \11947 , \11948 , \11949 , \11950 , \11951 , \11952 , \11953 ,
         \11954 , \11955 , \11956 , \11957 , \11958 , \11959 , \11960 , \11961 , \11962 , \11963 ,
         \11964 , \11965 , \11966 , \11967 , \11968 , \11969 , \11970 , \11971 , \11972 , \11973 ,
         \11974 , \11975 , \11976 , \11977 , \11978 , \11979 , \11980 , \11981 , \11982 , \11983 ,
         \11984 , \11985 , \11986 , \11987 , \11988 , \11989 , \11990 , \11991 , \11992 , \11993 ,
         \11994 , \11995 , \11996 , \11997 , \11998 , \11999 , \12000 , \12001 , \12002 , \12003 ,
         \12004 , \12005 , \12006 , \12007 , \12008 , \12009 , \12010 , \12011 , \12012 , \12013 ,
         \12014 , \12015 , \12016 , \12017 , \12018 , \12019 , \12020 , \12021 , \12022 , \12023 ,
         \12024 , \12025 , \12026 , \12027 , \12028 , \12029 , \12030 , \12031 , \12032 , \12033 ,
         \12034 , \12035 , \12036 , \12037 , \12038 , \12039 , \12040 , \12041 , \12042 , \12043 ,
         \12044 , \12045 , \12046 , \12047 , \12048 , \12049 , \12050 , \12051 , \12052 , \12053 ,
         \12054 , \12055 , \12056 , \12057 , \12058 , \12059 , \12060 , \12061 , \12062 , \12063 ,
         \12064 , \12065 , \12066 , \12067 , \12068 , \12069 , \12070 , \12071 , \12072 , \12073 ,
         \12074 , \12075 , \12076 , \12077 , \12078 , \12079 , \12080 , \12081 , \12082 , \12083 ,
         \12084 , \12085 , \12086 , \12087 , \12088 , \12089 , \12090 , \12091 , \12092 , \12093 ,
         \12094 , \12095 , \12096 , \12097 , \12098 , \12099 , \12100 , \12101 , \12102 , \12103 ,
         \12104 , \12105 , \12106 , \12107 , \12108 , \12109 , \12110 , \12111 , \12112 , \12113 ,
         \12114 , \12115 , \12116 , \12117 , \12118 , \12119 , \12120 , \12121 , \12122 , \12123 ,
         \12124 , \12125 , \12126 , \12127 , \12128 , \12129 , \12130 , \12131 , \12132 , \12133 ,
         \12134 , \12135 , \12136 , \12137 , \12138 , \12139 , \12140 , \12141 , \12142 , \12143 ,
         \12144 , \12145 , \12146 , \12147 , \12148 , \12149 , \12150 , \12151 , \12152 , \12153 ,
         \12154 , \12155 , \12156 , \12157 , \12158 , \12159 , \12160 , \12161 , \12162 , \12163 ,
         \12164 , \12165 , \12166 , \12167 , \12168 , \12169 , \12170 , \12171 , \12172 , \12173 ,
         \12174 , \12175 , \12176 , \12177 , \12178 , \12179 , \12180 , \12181 , \12182 , \12183 ,
         \12184 , \12185 , \12186 , \12187 , \12188 , \12189 , \12190 , \12191 , \12192 , \12193 ,
         \12194 , \12195 , \12196 , \12197 , \12198 , \12199 , \12200 , \12201 , \12202 , \12203 ,
         \12204 , \12205 , \12206 , \12207 , \12208 , \12209 , \12210 , \12211 , \12212 , \12213 ,
         \12214 , \12215 , \12216 , \12217 , \12218 , \12219 , \12220 , \12221 , \12222 , \12223 ,
         \12224 , \12225 , \12226 , \12227 , \12228 , \12229 , \12230 , \12231 , \12232 , \12233 ,
         \12234 , \12235 , \12236 , \12237 , \12238 , \12239 , \12240 , \12241 , \12242 , \12243 ,
         \12244 , \12245 , \12246 , \12247 , \12248 , \12249 , \12250 , \12251 , \12252 , \12253 ,
         \12254 , \12255 , \12256 , \12257 , \12258 , \12259 , \12260 , \12261 , \12262 , \12263 ,
         \12264 , \12265 , \12266 , \12267 , \12268 , \12269 , \12270 , \12271 , \12272 , \12273 ,
         \12274 , \12275 , \12276 , \12277 , \12278 , \12279 , \12280 , \12281 , \12282 , \12283 ,
         \12284 , \12285 , \12286 , \12287 , \12288 , \12289 , \12290 , \12291 , \12292 , \12293 ,
         \12294 , \12295 , \12296 , \12297 , \12298 , \12299 , \12300 , \12301 , \12302 , \12303 ,
         \12304 , \12305 , \12306 , \12307 , \12308 , \12309 , \12310 , \12311 , \12312 , \12313 ,
         \12314 , \12315 , \12316 , \12317 , \12318 , \12319 , \12320 , \12321 , \12322 , \12323 ,
         \12324 , \12325 , \12326 , \12327 , \12328 , \12329 , \12330 , \12331 , \12332 , \12333 ,
         \12334 , \12335 , \12336 , \12337 , \12338 , \12339 , \12340 , \12341 , \12342 , \12343 ,
         \12344 , \12345 , \12346 , \12347 , \12348 , \12349 , \12350 , \12351 , \12352 , \12353 ,
         \12354 , \12355 , \12356 , \12357 , \12358 , \12359 , \12360 , \12361 , \12362 , \12363 ,
         \12364 , \12365 , \12366 , \12367 , \12368 , \12369 , \12370 , \12371 , \12372 , \12373 ,
         \12374 , \12375 , \12376 , \12377 , \12378 , \12379 , \12380 , \12381 , \12382 , \12383 ,
         \12384 , \12385 , \12386 , \12387 , \12388 , \12389 , \12390 , \12391 , \12392 , \12393 ,
         \12394 , \12395 , \12396 , \12397 , \12398 , \12399 , \12400 , \12401 , \12402 , \12403 ,
         \12404 , \12405 , \12406 , \12407 , \12408 , \12409 , \12410 , \12411 , \12412 , \12413 ,
         \12414 , \12415 , \12416 , \12417 , \12418 , \12419 , \12420 , \12421 , \12422 , \12423 ,
         \12424 , \12425 , \12426 , \12427 , \12428 , \12429 , \12430 , \12431 , \12432 , \12433 ,
         \12434 , \12435 , \12436 , \12437 , \12438 , \12439 , \12440 , \12441 , \12442 , \12443 ,
         \12444 , \12445 , \12446 , \12447 , \12448 , \12449 , \12450 , \12451 , \12452 , \12453 ,
         \12454 , \12455 , \12456 , \12457 , \12458 , \12459 , \12460 , \12461 , \12462 , \12463 ,
         \12464 , \12465 , \12466 , \12467 , \12468 , \12469 , \12470 , \12471 , \12472 , \12473 ,
         \12474 , \12475 , \12476 , \12477 , \12478 , \12479 , \12480 , \12481 , \12482 , \12483 ,
         \12484 , \12485 , \12486 , \12487 , \12488 , \12489 , \12490 , \12491 , \12492 , \12493 ,
         \12494 , \12495 , \12496 , \12497 , \12498 , \12499 , \12500 , \12501 , \12502 , \12503 ,
         \12504 , \12505 , \12506 , \12507 , \12508 , \12509 , \12510 , \12511 , \12512 , \12513 ,
         \12514 , \12515 , \12516 , \12517 , \12518 , \12519 , \12520 , \12521 , \12522 , \12523 ,
         \12524 , \12525 , \12526 , \12527 , \12528 , \12529 , \12530 , \12531 , \12532 , \12533 ,
         \12534 , \12535 , \12536 , \12537 , \12538 , \12539 , \12540 , \12541 , \12542 , \12543 ,
         \12544 , \12545 , \12546 , \12547 , \12548 , \12549 , \12550 , \12551 , \12552 , \12553 ,
         \12554 , \12555 , \12556 , \12557 , \12558 , \12559 , \12560 , \12561 , \12562 , \12563 ,
         \12564 , \12565 , \12566 , \12567 , \12568 , \12569 , \12570 , \12571 , \12572 , \12573 ,
         \12574 , \12575 , \12576 , \12577 , \12578 , \12579 , \12580 , \12581 , \12582 , \12583 ,
         \12584 , \12585 , \12586 , \12587 , \12588 , \12589 , \12590 , \12591 , \12592 , \12593 ,
         \12594 , \12595 , \12596 , \12597 , \12598 , \12599 , \12600 , \12601 , \12602 , \12603 ,
         \12604 , \12605 , \12606 , \12607 , \12608 , \12609 , \12610 , \12611 , \12612 , \12613 ,
         \12614 , \12615 , \12616 , \12617 , \12618 , \12619 , \12620 , \12621 , \12622 , \12623 ,
         \12624 , \12625 , \12626 , \12627 , \12628 , \12629 , \12630 , \12631 , \12632 , \12633 ,
         \12634 , \12635 , \12636 , \12637 , \12638 , \12639 , \12640 , \12641 , \12642 , \12643 ,
         \12644 , \12645 , \12646 , \12647 , \12648 , \12649 , \12650 , \12651 , \12652 , \12653 ,
         \12654 , \12655 , \12656 , \12657 , \12658 , \12659 , \12660 , \12661 , \12662 , \12663 ,
         \12664 , \12665 , \12666 , \12667 , \12668 , \12669 , \12670 , \12671 , \12672 , \12673 ,
         \12674 , \12675 , \12676 , \12677 , \12678 , \12679 , \12680 , \12681 , \12682 , \12683 ,
         \12684 , \12685 , \12686 , \12687 , \12688 , \12689 , \12690 , \12691 , \12692 , \12693 ,
         \12694 , \12695 , \12696 , \12697 , \12698 , \12699 , \12700 , \12701 , \12702 , \12703 ,
         \12704 , \12705 , \12706 , \12707 , \12708 , \12709 , \12710 , \12711 , \12712 , \12713 ,
         \12714 , \12715 , \12716 , \12717 , \12718 , \12719 , \12720 , \12721 , \12722 , \12723 ,
         \12724 , \12725 , \12726 , \12727 , \12728 , \12729 , \12730 , \12731 , \12732 , \12733 ,
         \12734 , \12735 , \12736 , \12737 , \12738 , \12739 , \12740 , \12741 , \12742 , \12743 ,
         \12744 , \12745 , \12746 , \12747 , \12748 , \12749 , \12750 , \12751 , \12752 , \12753 ,
         \12754 , \12755 , \12756 , \12757 , \12758 , \12759 , \12760 , \12761 , \12762 , \12763 ,
         \12764 , \12765 , \12766 , \12767 , \12768 , \12769 , \12770 , \12771 , \12772 , \12773 ,
         \12774 , \12775 , \12776 , \12777 , \12778 , \12779 , \12780 , \12781 , \12782 , \12783 ,
         \12784 , \12785 , \12786 , \12787 , \12788 , \12789 , \12790 , \12791 , \12792 , \12793 ,
         \12794 , \12795 , \12796 , \12797 , \12798 , \12799 , \12800 , \12801 , \12802 , \12803 ,
         \12804 , \12805 , \12806 , \12807 , \12808 , \12809 , \12810 , \12811 , \12812 , \12813 ,
         \12814 , \12815 , \12816 , \12817 , \12818 , \12819 , \12820 , \12821 , \12822 , \12823 ,
         \12824 , \12825 , \12826 , \12827 , \12828 , \12829 , \12830 , \12831 , \12832 , \12833 ,
         \12834 , \12835 , \12836 , \12837 , \12838 , \12839 , \12840 , \12841 , \12842 , \12843 ,
         \12844 , \12845 , \12846 , \12847 , \12848 , \12849 , \12850 , \12851 , \12852 , \12853 ,
         \12854 , \12855 , \12856 , \12857 , \12858 , \12859 , \12860 , \12861 , \12862 , \12863 ,
         \12864 , \12865 , \12866 , \12867 , \12868 , \12869 , \12870 , \12871 , \12872 , \12873 ,
         \12874 , \12875 , \12876 , \12877 , \12878 , \12879 , \12880 , \12881 , \12882 , \12883 ,
         \12884 , \12885 , \12886 , \12887 , \12888 , \12889 , \12890 , \12891 , \12892 , \12893 ,
         \12894 , \12895 , \12896 , \12897 , \12898 , \12899 , \12900 , \12901 , \12902 , \12903 ,
         \12904 , \12905 , \12906 , \12907 , \12908 , \12909 , \12910 , \12911 , \12912 , \12913 ,
         \12914 , \12915 , \12916 , \12917 , \12918 , \12919 , \12920 , \12921 , \12922 , \12923 ,
         \12924 , \12925 , \12926 , \12927 , \12928 , \12929 , \12930 , \12931 , \12932 , \12933 ,
         \12934 , \12935 , \12936 , \12937 , \12938 , \12939 , \12940 , \12941 , \12942 , \12943 ,
         \12944 , \12945 , \12946 , \12947 , \12948 , \12949 , \12950 , \12951 , \12952 , \12953 ,
         \12954 , \12955 , \12956 , \12957 , \12958 , \12959 , \12960 , \12961 , \12962 , \12963 ,
         \12964 , \12965 , \12966 , \12967 , \12968 , \12969 , \12970 , \12971 , \12972 , \12973 ,
         \12974 , \12975 , \12976 , \12977 , \12978 , \12979 , \12980 , \12981 , \12982 , \12983 ,
         \12984 , \12985 , \12986 , \12987 , \12988 , \12989 , \12990 , \12991 , \12992 , \12993 ,
         \12994 , \12995 , \12996 , \12997 , \12998 , \12999 , \13000 , \13001 , \13002 , \13003 ,
         \13004 , \13005 , \13006 , \13007 , \13008 , \13009 , \13010 , \13011 , \13012 , \13013 ,
         \13014 , \13015 , \13016 , \13017 , \13018 , \13019 , \13020 , \13021 , \13022 , \13023 ,
         \13024 , \13025 , \13026 , \13027 , \13028 , \13029 , \13030 , \13031 , \13032 , \13033 ,
         \13034 , \13035 , \13036 , \13037 , \13038 , \13039 , \13040 , \13041 , \13042 , \13043 ,
         \13044 , \13045 , \13046 , \13047 , \13048 , \13049 , \13050 , \13051 , \13052 , \13053 ,
         \13054 , \13055 , \13056 , \13057 , \13058 , \13059 , \13060 , \13061 , \13062 , \13063 ,
         \13064 , \13065 , \13066 , \13067 , \13068 , \13069 , \13070 , \13071 , \13072 , \13073 ,
         \13074 , \13075 , \13076 , \13077 , \13078 , \13079 , \13080 , \13081 , \13082 , \13083 ,
         \13084 , \13085 , \13086 , \13087 , \13088 , \13089 , \13090 , \13091 , \13092 , \13093 ,
         \13094 , \13095 , \13096 , \13097 , \13098 , \13099 , \13100 , \13101 , \13102 , \13103 ,
         \13104 , \13105 , \13106 , \13107 , \13108 , \13109 , \13110 , \13111 , \13112 , \13113 ,
         \13114 , \13115 , \13116 , \13117 , \13118 , \13119 , \13120 , \13121 , \13122 , \13123 ,
         \13124 , \13125 , \13126 , \13127 , \13128 , \13129 , \13130 , \13131 , \13132 , \13133 ,
         \13134 , \13135 , \13136 , \13137 , \13138 , \13139 , \13140 , \13141 , \13142 , \13143 ,
         \13144 , \13145 , \13146 , \13147 , \13148 , \13149 , \13150 , \13151 , \13152 , \13153 ,
         \13154 , \13155 , \13156 , \13157 , \13158 , \13159 , \13160 , \13161 , \13162 , \13163 ,
         \13164 , \13165 , \13166 , \13167 , \13168 , \13169 , \13170 , \13171 , \13172 , \13173 ,
         \13174 , \13175 , \13176 , \13177 , \13178 , \13179 , \13180 , \13181 , \13182 , \13183 ,
         \13184 , \13185 , \13186 , \13187 , \13188 , \13189 , \13190 , \13191 , \13192 , \13193 ,
         \13194 , \13195 , \13196 , \13197 , \13198 , \13199 , \13200 , \13201 , \13202 , \13203 ,
         \13204 , \13205 , \13206 , \13207 , \13208 , \13209 , \13210 , \13211 , \13212 , \13213 ,
         \13214 , \13215 , \13216 , \13217 , \13218 , \13219 , \13220 , \13221 , \13222 , \13223 ,
         \13224 , \13225 , \13226 , \13227 , \13228 , \13229 , \13230 , \13231 , \13232 , \13233 ,
         \13234 , \13235 , \13236 , \13237 , \13238 , \13239 , \13240 , \13241 , \13242 , \13243 ,
         \13244 , \13245 , \13246 , \13247 , \13248 , \13249 , \13250 , \13251 , \13252 , \13253 ,
         \13254 , \13255 , \13256 , \13257 , \13258 , \13259 , \13260 , \13261 , \13262 , \13263 ,
         \13264 , \13265 , \13266 , \13267 , \13268 , \13269 , \13270 , \13271 , \13272 , \13273 ,
         \13274 , \13275 , \13276 , \13277 , \13278 , \13279 , \13280 , \13281 , \13282 , \13283 ,
         \13284 , \13285 , \13286 , \13287 , \13288 , \13289 , \13290 , \13291 , \13292 , \13293 ,
         \13294 , \13295 , \13296 , \13297 , \13298 , \13299 , \13300 , \13301 , \13302 , \13303 ,
         \13304 , \13305 , \13306 , \13307 , \13308 , \13309 , \13310 , \13311 , \13312 , \13313 ,
         \13314 , \13315 , \13316 , \13317 , \13318 , \13319 , \13320 , \13321 , \13322 , \13323 ,
         \13324 , \13325 , \13326 , \13327 , \13328 , \13329 , \13330 , \13331 , \13332 , \13333 ,
         \13334 , \13335 , \13336 , \13337 , \13338 , \13339 , \13340 , \13341 , \13342 , \13343 ,
         \13344 , \13345 , \13346 , \13347 , \13348 , \13349 , \13350 , \13351 , \13352 , \13353 ,
         \13354 , \13355 , \13356 , \13357 , \13358 , \13359 , \13360 , \13361 , \13362 , \13363 ,
         \13364 , \13365 , \13366 , \13367 , \13368 , \13369 , \13370 , \13371 , \13372 , \13373 ,
         \13374 , \13375 , \13376 , \13377 , \13378 , \13379 , \13380 , \13381 , \13382 , \13383 ,
         \13384 , \13385 , \13386 , \13387 , \13388 , \13389 , \13390 , \13391 , \13392 , \13393 ,
         \13394 , \13395 , \13396 , \13397 , \13398 , \13399 , \13400 , \13401 , \13402 , \13403 ,
         \13404 , \13405 , \13406 , \13407 , \13408 , \13409 , \13410 , \13411 , \13412 , \13413 ,
         \13414 , \13415 , \13416 , \13417 , \13418 , \13419 , \13420 , \13421 , \13422 , \13423 ,
         \13424 , \13425 , \13426 , \13427 , \13428 , \13429 , \13430 , \13431 , \13432 , \13433 ,
         \13434 , \13435 , \13436 , \13437 , \13438 , \13439 , \13440 , \13441 , \13442 , \13443 ,
         \13444 , \13445 , \13446 , \13447 , \13448 , \13449 , \13450 , \13451 , \13452 , \13453 ,
         \13454 , \13455 , \13456 , \13457 , \13458 , \13459 , \13460 , \13461 , \13462 , \13463 ,
         \13464 , \13465 , \13466 , \13467 , \13468 , \13469 , \13470 , \13471 , \13472 , \13473 ,
         \13474 , \13475 , \13476 , \13477 , \13478 , \13479 , \13480 , \13481 , \13482 , \13483 ,
         \13484 , \13485 , \13486 , \13487 , \13488 , \13489 , \13490 , \13491 , \13492 , \13493 ,
         \13494 , \13495 , \13496 , \13497 , \13498 , \13499 , \13500 , \13501 , \13502 , \13503 ,
         \13504 , \13505 , \13506 , \13507 , \13508 , \13509 , \13510 , \13511 , \13512 , \13513 ,
         \13514 , \13515 , \13516 , \13517 , \13518 , \13519 , \13520 , \13521 , \13522 , \13523 ,
         \13524 , \13525 , \13526 , \13527 , \13528 , \13529 , \13530 , \13531 , \13532 , \13533 ,
         \13534 , \13535 , \13536 , \13537 , \13538 , \13539 , \13540 , \13541 , \13542 , \13543 ,
         \13544 , \13545 , \13546 , \13547 , \13548 , \13549 , \13550 , \13551 , \13552 , \13553 ,
         \13554 , \13555 , \13556 , \13557 , \13558 , \13559 , \13560 , \13561 , \13562 , \13563 ,
         \13564 , \13565 , \13566 , \13567 , \13568 , \13569 , \13570 , \13571 , \13572 , \13573 ,
         \13574 , \13575 , \13576 , \13577 , \13578 , \13579 , \13580 , \13581 , \13582 , \13583 ,
         \13584 , \13585 , \13586 , \13587 , \13588 , \13589 , \13590 , \13591 , \13592 , \13593 ,
         \13594 , \13595 , \13596 , \13597 , \13598 , \13599 , \13600 , \13601 , \13602 , \13603 ,
         \13604 , \13605 , \13606 , \13607 , \13608 , \13609 , \13610 , \13611 , \13612 , \13613 ,
         \13614 , \13615 , \13616 , \13617 , \13618 , \13619 , \13620 , \13621 , \13622 , \13623 ,
         \13624 , \13625 , \13626 , \13627 , \13628 , \13629 , \13630 , \13631 , \13632 , \13633 ,
         \13634 , \13635 , \13636 , \13637 , \13638 , \13639 , \13640 , \13641 , \13642 , \13643 ,
         \13644 , \13645 , \13646 , \13647 , \13648 , \13649 , \13650 , \13651 , \13652 , \13653 ,
         \13654 , \13655 , \13656 , \13657 , \13658 , \13659 , \13660 , \13661 , \13662 , \13663 ,
         \13664 , \13665 , \13666 , \13667 , \13668 , \13669 , \13670 , \13671 , \13672 , \13673 ,
         \13674 , \13675 , \13676 , \13677 , \13678 , \13679 , \13680 , \13681 , \13682 , \13683 ,
         \13684 , \13685 , \13686 , \13687 , \13688 , \13689 , \13690 , \13691 , \13692 , \13693 ,
         \13694 , \13695 , \13696 , \13697 , \13698 , \13699 , \13700 , \13701 , \13702 , \13703 ,
         \13704 , \13705 , \13706 , \13707 , \13708 , \13709 , \13710 , \13711 , \13712 , \13713 ,
         \13714 , \13715 , \13716 , \13717 , \13718 , \13719 , \13720 , \13721 , \13722 , \13723 ,
         \13724 , \13725 , \13726 , \13727 , \13728 , \13729 , \13730 , \13731 , \13732 , \13733 ,
         \13734 , \13735 , \13736 , \13737 , \13738 , \13739 , \13740 , \13741 , \13742 , \13743 ,
         \13744 , \13745 , \13746 , \13747 , \13748 , \13749 , \13750 , \13751 , \13752 , \13753 ,
         \13754 , \13755 , \13756 , \13757 , \13758 , \13759 , \13760 , \13761 , \13762 , \13763 ,
         \13764 , \13765 , \13766 , \13767 , \13768 , \13769 , \13770 , \13771 , \13772 , \13773 ,
         \13774 , \13775 , \13776 , \13777 , \13778 , \13779 , \13780 , \13781 , \13782 , \13783 ,
         \13784 , \13785 , \13786 , \13787 , \13788 , \13789 , \13790 , \13791 , \13792 , \13793 ,
         \13794 , \13795 , \13796 , \13797 , \13798 , \13799 , \13800 , \13801 , \13802 , \13803 ,
         \13804 , \13805 , \13806 , \13807 , \13808 , \13809 , \13810 , \13811 , \13812 , \13813 ,
         \13814 , \13815 , \13816 , \13817 , \13818 , \13819 , \13820 , \13821 , \13822 , \13823 ,
         \13824 , \13825 , \13826 , \13827 , \13828 , \13829 , \13830 , \13831 , \13832 , \13833 ,
         \13834 , \13835 , \13836 , \13837 , \13838 , \13839 , \13840 , \13841 , \13842 , \13843 ,
         \13844 , \13845 , \13846 , \13847 , \13848 , \13849 , \13850 , \13851 , \13852 , \13853 ,
         \13854 , \13855 , \13856 , \13857 , \13858 , \13859 , \13860 , \13861 , \13862 , \13863 ,
         \13864 , \13865 , \13866 , \13867 , \13868 , \13869 , \13870 , \13871 , \13872 , \13873 ,
         \13874 , \13875 , \13876 , \13877 , \13878 , \13879 , \13880 , \13881 , \13882 , \13883 ,
         \13884 , \13885 , \13886 , \13887 , \13888 , \13889 , \13890 , \13891 , \13892 , \13893 ,
         \13894 , \13895 , \13896 , \13897 , \13898 , \13899 , \13900 , \13901 , \13902 , \13903 ,
         \13904 , \13905 , \13906 , \13907 , \13908 , \13909 , \13910 , \13911 , \13912 , \13913 ,
         \13914 , \13915 , \13916 , \13917 , \13918 , \13919 , \13920 , \13921 , \13922 , \13923 ,
         \13924 , \13925 , \13926 , \13927 , \13928 , \13929 , \13930 , \13931 , \13932 , \13933 ,
         \13934 , \13935 , \13936 , \13937 , \13938 , \13939 , \13940 , \13941 , \13942 , \13943 ,
         \13944 , \13945 , \13946 , \13947 , \13948 , \13949 , \13950 , \13951 , \13952 , \13953 ,
         \13954 , \13955 , \13956 , \13957 , \13958 , \13959 , \13960 , \13961 , \13962 , \13963 ,
         \13964 , \13965 , \13966 , \13967 , \13968 , \13969 , \13970 , \13971 , \13972 , \13973 ,
         \13974 , \13975 , \13976 , \13977 , \13978 , \13979 , \13980 , \13981 , \13982 , \13983 ,
         \13984 , \13985 , \13986 , \13987 , \13988 , \13989 , \13990 , \13991 , \13992 , \13993 ,
         \13994 , \13995 , \13996 , \13997 , \13998 , \13999 , \14000 , \14001 , \14002 , \14003 ,
         \14004 , \14005 , \14006 , \14007 , \14008 , \14009 , \14010 , \14011 , \14012 , \14013 ,
         \14014 , \14015 , \14016 , \14017 , \14018 , \14019 , \14020 , \14021 , \14022 , \14023 ,
         \14024 , \14025 , \14026 , \14027 , \14028 , \14029 , \14030 , \14031 , \14032 , \14033 ,
         \14034 , \14035 , \14036 , \14037 , \14038 , \14039 , \14040 , \14041 , \14042 , \14043 ,
         \14044 , \14045 , \14046 , \14047 , \14048 , \14049 , \14050 , \14051 , \14052 , \14053 ,
         \14054 , \14055 , \14056 , \14057 , \14058 , \14059 , \14060 , \14061 , \14062 , \14063 ,
         \14064 , \14065 , \14066 , \14067 , \14068 , \14069 , \14070 , \14071 , \14072 , \14073 ,
         \14074 , \14075 , \14076 , \14077 , \14078 , \14079 , \14080 , \14081 , \14082 , \14083 ,
         \14084 , \14085 , \14086 , \14087 , \14088 , \14089 , \14090 , \14091 , \14092 , \14093 ,
         \14094 , \14095 , \14096 , \14097 , \14098 , \14099 , \14100 , \14101 , \14102 , \14103 ,
         \14104 , \14105 , \14106 , \14107 , \14108 , \14109 , \14110 , \14111 , \14112 , \14113 ,
         \14114 , \14115 , \14116 , \14117 , \14118 , \14119 , \14120 , \14121 , \14122 , \14123 ,
         \14124 , \14125 , \14126 , \14127 , \14128 , \14129 , \14130 , \14131 , \14132 , \14133 ,
         \14134 , \14135 , \14136 , \14137 , \14138 , \14139 , \14140 , \14141 , \14142 , \14143 ,
         \14144 , \14145 , \14146 , \14147 , \14148 , \14149 , \14150 , \14151 , \14152 , \14153 ,
         \14154 , \14155 , \14156 , \14157 , \14158 , \14159 , \14160 , \14161 , \14162 , \14163 ,
         \14164 , \14165 , \14166 , \14167 , \14168 , \14169 , \14170 , \14171 , \14172 , \14173 ,
         \14174 , \14175 , \14176 , \14177 , \14178 , \14179 , \14180 , \14181 , \14182 , \14183 ,
         \14184 , \14185 , \14186 , \14187 , \14188 , \14189 , \14190 , \14191 , \14192 , \14193 ,
         \14194 , \14195 , \14196 , \14197 , \14198 , \14199 , \14200 , \14201 , \14202 , \14203 ,
         \14204 , \14205 , \14206 , \14207 , \14208 , \14209 , \14210 , \14211 , \14212 , \14213 ,
         \14214 , \14215 , \14216 , \14217 , \14218 , \14219 , \14220 , \14221 , \14222 , \14223 ,
         \14224 , \14225 , \14226 , \14227 , \14228 , \14229 , \14230 , \14231 , \14232 , \14233 ,
         \14234 , \14235 , \14236 , \14237 , \14238 , \14239 , \14240 , \14241 , \14242 , \14243 ,
         \14244 , \14245 , \14246 , \14247 , \14248 , \14249 , \14250 , \14251 , \14252 , \14253 ,
         \14254 , \14255 , \14256 , \14257 , \14258 , \14259 , \14260 , \14261 , \14262 , \14263 ,
         \14264 , \14265 , \14266 , \14267 , \14268 , \14269 , \14270 , \14271 , \14272 , \14273 ,
         \14274 , \14275 , \14276 , \14277 , \14278 , \14279 , \14280 , \14281 , \14282 , \14283 ,
         \14284 , \14285 , \14286 , \14287 , \14288 , \14289 , \14290 , \14291 , \14292 , \14293 ,
         \14294 , \14295 , \14296 , \14297 , \14298 , \14299 , \14300 , \14301 , \14302 , \14303 ,
         \14304 , \14305 , \14306 , \14307 , \14308 , \14309 , \14310 , \14311 , \14312 , \14313 ,
         \14314 , \14315 , \14316 , \14317 , \14318 , \14319 , \14320 , \14321 , \14322 , \14323 ,
         \14324 , \14325 , \14326 , \14327 , \14328 , \14329 , \14330 , \14331 , \14332 , \14333 ,
         \14334 , \14335 , \14336 , \14337 , \14338 , \14339 , \14340 , \14341 , \14342 , \14343 ,
         \14344 , \14345 , \14346 , \14347 , \14348 , \14349 , \14350 , \14351 , \14352 , \14353 ,
         \14354 , \14355 , \14356 , \14357 , \14358 , \14359 , \14360 , \14361 , \14362 , \14363 ,
         \14364 , \14365 , \14366 , \14367 , \14368 , \14369 , \14370 , \14371 , \14372 , \14373 ,
         \14374 , \14375 , \14376 , \14377 , \14378 , \14379 , \14380 , \14381 , \14382 , \14383 ,
         \14384 , \14385 , \14386 , \14387 , \14388 , \14389 , \14390 , \14391 , \14392 , \14393 ,
         \14394 , \14395 , \14396 , \14397 , \14398 , \14399 , \14400 , \14401 , \14402 , \14403 ,
         \14404 , \14405 , \14406 , \14407 , \14408 , \14409 , \14410 , \14411 , \14412 , \14413 ,
         \14414 , \14415 , \14416 , \14417 , \14418 , \14419 , \14420 , \14421 , \14422 , \14423 ,
         \14424 , \14425 , \14426 , \14427 , \14428 , \14429 , \14430 , \14431 , \14432 , \14433 ,
         \14434 , \14435 , \14436 , \14437 , \14438 , \14439 , \14440 , \14441 , \14442 , \14443 ,
         \14444 , \14445 , \14446 , \14447 , \14448 , \14449 , \14450 , \14451 , \14452 , \14453 ,
         \14454 , \14455 , \14456 , \14457 , \14458 , \14459 , \14460 , \14461 , \14462 , \14463 ,
         \14464 , \14465 , \14466 , \14467 , \14468 , \14469 , \14470 , \14471 , \14472 , \14473 ,
         \14474 , \14475 , \14476 , \14477 , \14478 , \14479 , \14480 , \14481 , \14482 , \14483 ,
         \14484 , \14485 , \14486 , \14487 , \14488 , \14489 , \14490 , \14491 , \14492 , \14493 ,
         \14494 , \14495 , \14496 , \14497 , \14498 , \14499 , \14500 , \14501 , \14502 , \14503 ,
         \14504 , \14505 , \14506 , \14507 , \14508 , \14509 , \14510 , \14511 , \14512 , \14513 ,
         \14514 , \14515 , \14516 , \14517 , \14518 , \14519 , \14520 , \14521 , \14522 , \14523 ,
         \14524 , \14525 , \14526 , \14527 , \14528 , \14529 , \14530 , \14531 , \14532 , \14533 ,
         \14534 , \14535 , \14536 , \14537 , \14538 , \14539 , \14540 , \14541 , \14542 , \14543 ,
         \14544 , \14545 , \14546 , \14547 , \14548 , \14549 , \14550 , \14551 , \14552 , \14553 ,
         \14554 , \14555 , \14556 , \14557 , \14558 , \14559 , \14560 , \14561 , \14562 , \14563 ,
         \14564 , \14565 , \14566 , \14567 , \14568 , \14569 , \14570 , \14571 , \14572 , \14573 ,
         \14574 , \14575 , \14576 , \14577 , \14578 , \14579 , \14580 , \14581 , \14582 , \14583 ,
         \14584 , \14585 , \14586 , \14587 , \14588 , \14589 , \14590 , \14591 , \14592 , \14593 ,
         \14594 , \14595 , \14596 , \14597 , \14598 , \14599 , \14600 , \14601 , \14602 , \14603 ,
         \14604 , \14605 , \14606 , \14607 , \14608 , \14609 , \14610 , \14611 , \14612 , \14613 ,
         \14614 , \14615 , \14616 , \14617 , \14618 , \14619 , \14620 , \14621 , \14622 , \14623 ,
         \14624 , \14625 , \14626 , \14627 , \14628 , \14629 , \14630 , \14631 , \14632 , \14633 ,
         \14634 , \14635 , \14636 , \14637 , \14638 , \14639 , \14640 , \14641 , \14642 , \14643 ,
         \14644 , \14645 , \14646 , \14647 , \14648 , \14649 , \14650 , \14651 , \14652 , \14653 ,
         \14654 , \14655 , \14656 , \14657 , \14658 , \14659 , \14660 , \14661 , \14662 , \14663 ,
         \14664 , \14665 , \14666 , \14667 , \14668 , \14669 , \14670 , \14671 , \14672 , \14673 ,
         \14674 , \14675 , \14676 , \14677 , \14678 , \14679 , \14680 , \14681 , \14682 , \14683 ,
         \14684 , \14685 , \14686 , \14687 , \14688 , \14689 , \14690 , \14691 , \14692 , \14693 ,
         \14694 , \14695 , \14696 , \14697 , \14698 , \14699 , \14700 , \14701 , \14702 , \14703 ,
         \14704 , \14705 , \14706 , \14707 , \14708 , \14709 , \14710 , \14711 , \14712 , \14713 ,
         \14714 , \14715 , \14716 , \14717 , \14718 , \14719 , \14720 , \14721 , \14722 , \14723 ,
         \14724 , \14725 , \14726 , \14727 , \14728 , \14729 , \14730 , \14731 , \14732 , \14733 ,
         \14734 , \14735 , \14736 , \14737 , \14738 , \14739 , \14740 , \14741 , \14742 , \14743 ,
         \14744 , \14745 , \14746 , \14747 , \14748 , \14749 , \14750 , \14751 , \14752 , \14753 ,
         \14754 , \14755 , \14756 , \14757 , \14758 , \14759 , \14760 , \14761 , \14762 , \14763 ,
         \14764 , \14765 , \14766 , \14767 , \14768 , \14769 , \14770 , \14771 , \14772 , \14773 ,
         \14774 , \14775 , \14776 , \14777 , \14778 , \14779 , \14780 , \14781 , \14782 , \14783 ,
         \14784 , \14785 , \14786 , \14787 , \14788 , \14789 , \14790 , \14791 , \14792 , \14793 ,
         \14794 , \14795 , \14796 , \14797 , \14798 , \14799 , \14800 , \14801 , \14802 , \14803 ,
         \14804 , \14805 , \14806 , \14807 , \14808 , \14809 , \14810 , \14811 , \14812 , \14813 ,
         \14814 , \14815 , \14816 , \14817 , \14818 , \14819 , \14820 , \14821 , \14822 , \14823 ,
         \14824 , \14825 , \14826 , \14827 , \14828 , \14829 , \14830 , \14831 , \14832 , \14833 ,
         \14834 , \14835 , \14836 , \14837 , \14838 , \14839 , \14840 , \14841 , \14842 , \14843 ,
         \14844 , \14845 , \14846 , \14847 , \14848 , \14849 , \14850 , \14851 , \14852 , \14853 ,
         \14854 , \14855 , \14856 , \14857 , \14858 , \14859 , \14860 , \14861 , \14862 , \14863 ,
         \14864 , \14865 , \14866 , \14867 , \14868 , \14869 , \14870 , \14871 , \14872 , \14873 ,
         \14874 , \14875 , \14876 , \14877 , \14878 , \14879 , \14880 , \14881 , \14882 , \14883 ,
         \14884 , \14885 , \14886 , \14887 , \14888 , \14889 , \14890 , \14891 , \14892 , \14893 ,
         \14894 , \14895 , \14896 , \14897 , \14898 , \14899 , \14900 , \14901 , \14902 , \14903 ,
         \14904 , \14905 , \14906 , \14907 , \14908 , \14909 , \14910 , \14911 , \14912 , \14913 ,
         \14914 , \14915 , \14916 , \14917 , \14918 , \14919 , \14920 , \14921 , \14922 , \14923 ,
         \14924 , \14925 , \14926 , \14927 , \14928 , \14929 , \14930 , \14931 , \14932 , \14933 ,
         \14934 , \14935 , \14936 , \14937 , \14938 , \14939 , \14940 , \14941 , \14942 , \14943 ,
         \14944 , \14945 , \14946 , \14947 , \14948 , \14949 , \14950 , \14951 , \14952 , \14953 ,
         \14954 , \14955 , \14956 , \14957 , \14958 , \14959 , \14960 , \14961 , \14962 , \14963 ,
         \14964 , \14965 , \14966 , \14967 , \14968 , \14969 , \14970 , \14971 , \14972 , \14973 ,
         \14974 , \14975 , \14976 , \14977 , \14978 , \14979 , \14980 , \14981 , \14982 , \14983 ,
         \14984 , \14985 , \14986 , \14987 , \14988 , \14989 , \14990 , \14991 , \14992 , \14993 ,
         \14994 , \14995 , \14996 , \14997 , \14998 , \14999 , \15000 , \15001 , \15002 , \15003 ,
         \15004 , \15005 , \15006 , \15007 , \15008 , \15009 , \15010 , \15011 , \15012 , \15013 ,
         \15014 , \15015 , \15016 , \15017 , \15018 , \15019 , \15020 , \15021 , \15022 , \15023 ,
         \15024 , \15025 , \15026 , \15027 , \15028 , \15029 , \15030 , \15031 ;
buf \U$labaj1525 ( R_61_85b54e8, \14014 );
buf \U$labaj1526 ( R_62_85b5590, \14196 );
buf \U$labaj1527 ( R_63_85b5638, \14286 );
buf \U$labaj1528 ( R_64_85b56e0, \14377 );
buf \U$labaj1529 ( R_65_85b5788, \14422 );
buf \U$labaj1530 ( R_66_85b5830, \14467 );
buf \U$labaj1531 ( R_67_85b58d8, \14510 );
buf \U$labaj1532 ( R_68_85b5980, \14553 );
buf \U$labaj1533 ( R_69_85b5a28, \14576 );
buf \U$labaj1534 ( R_6a_85b5ad0, \14599 );
buf \U$labaj1535 ( R_6b_85b5b78, \14621 );
buf \U$labaj1536 ( R_6c_85b5c20, \14643 );
buf \U$labaj1537 ( R_6d_85b5cc8, \14665 );
buf \U$labaj1538 ( R_6e_85b5d70, \14687 );
buf \U$labaj1539 ( R_6f_85b5e18, \14707 );
buf \U$labaj1540 ( R_70_85b5ec0, \14727 );
buf \U$labaj1541 ( R_71_85b5f68, \14739 );
buf \U$labaj1542 ( R_72_85b6010, \14751 );
buf \U$labaj1543 ( R_73_85b60b8, \14763 );
buf \U$labaj1544 ( R_74_85b6160, \14775 );
buf \U$labaj1545 ( R_75_85b6208, \14787 );
buf \U$labaj1546 ( R_76_85b62b0, \14799 );
buf \U$labaj1547 ( R_77_85b6358, \14810 );
buf \U$labaj1548 ( R_78_85b6400, \14821 );
buf \U$labaj1549 ( R_79_85b64a8, \14832 );
buf \U$labaj1550 ( R_7a_85b6550, \14843 );
buf \U$labaj1551 ( R_7b_85b65f8, \14854 );
buf \U$labaj1552 ( R_7c_85b66a0, \14865 );
buf \U$labaj1553 ( R_7d_85b6748, \14876 );
buf \U$labaj1554 ( R_7e_85b67f0, \14887 );
buf \U$labaj1555 ( R_7f_85b6898, \14894 );
buf \U$labaj1556 ( R_80_85b6940, \14901 );
buf \U$labaj1557 ( R_81_85b69e8, \14906 );
buf \U$labaj1558 ( R_82_85b6a90, \14911 );
buf \U$labaj1559 ( R_83_85b6b38, \14916 );
buf \U$labaj1560 ( R_84_85b6be0, \14921 );
buf \U$labaj1561 ( R_85_85b6c88, \14926 );
buf \U$labaj1562 ( R_86_85b6d30, \14931 );
buf \U$labaj1563 ( R_87_85b6dd8, \14936 );
buf \U$labaj1564 ( R_88_85b6e80, \14941 );
buf \U$labaj1565 ( R_89_85b6f28, \14946 );
buf \U$labaj1566 ( R_8a_85b6fd0, \14951 );
buf \U$labaj1567 ( R_8b_85b7078, \14956 );
buf \U$labaj1568 ( R_8c_85b7120, \14961 );
buf \U$labaj1569 ( R_8d_85b71c8, \14966 );
buf \U$labaj1570 ( R_8e_85b7270, \14971 );
buf \U$labaj1571 ( R_8f_85b7318, \14976 );
buf \U$labaj1572 ( R_90_85b73c0, \14981 );
buf \U$labaj1573 ( R_91_85b7468, \14986 );
buf \U$labaj1574 ( R_92_85b7510, \14991 );
buf \U$labaj1575 ( R_93_85b75b8, \14996 );
buf \U$labaj1576 ( R_94_85b7660, \15001 );
buf \U$labaj1577 ( R_95_85b7708, \15006 );
buf \U$labaj1578 ( R_96_85b77b0, \15011 );
buf \U$labaj1579 ( R_97_85b7858, \15016 );
buf \U$labaj1580 ( R_98_85b7900, \15021 );
buf \U$labaj1581 ( R_99_85b79a8, \15026 );
buf \U$labaj1582 ( R_9a_85b7a50, \15031 );
buf \U$1 ( \159 , RIb4bfa38_65);
buf \U$2 ( \160 , RIa167a08_1);
buf \U$3 ( \161 , RIb4ca3e8_33);
xor \U$4 ( \162 , \160 , \161 );
buf \U$5 ( \163 , RIa167990_2);
buf \U$6 ( \164 , RIb4c6c20_34);
xor \U$7 ( \165 , \163 , \164 );
or \U$8 ( \166 , \162 , \165 );
buf \U$9 ( \167 , RIa167918_3);
buf \U$10 ( \168 , RIb4c6ba8_35);
xor \U$11 ( \169 , \167 , \168 );
or \U$12 ( \170 , \166 , \169 );
buf \U$13 ( \171 , RIa1678a0_4);
buf \U$14 ( \172 , RIb4c6b30_36);
xor \U$15 ( \173 , \171 , \172 );
or \U$16 ( \174 , \170 , \173 );
buf \U$17 ( \175 , RIa167828_5);
buf \U$18 ( \176 , RIb4c6ab8_37);
xor \U$19 ( \177 , \175 , \176 );
or \U$20 ( \178 , \174 , \177 );
buf \U$21 ( \179 , RIa1677b0_6);
buf \U$22 ( \180 , RIb4c6a40_38);
xor \U$23 ( \181 , \179 , \180 );
or \U$24 ( \182 , \178 , \181 );
buf \U$25 ( \183 , RIa167738_7);
buf \U$26 ( \184 , RIb4c69c8_39);
xor \U$27 ( \185 , \183 , \184 );
or \U$28 ( \186 , \182 , \185 );
buf \U$29 ( \187 , RIa1676c0_8);
buf \U$30 ( \188 , RIb4c6950_40);
xor \U$31 ( \189 , \187 , \188 );
or \U$32 ( \190 , \186 , \189 );
buf \U$33 ( \191 , RIa167648_9);
buf \U$34 ( \192 , RIb4c68d8_41);
xor \U$35 ( \193 , \191 , \192 );
or \U$36 ( \194 , \190 , \193 );
buf \U$37 ( \195 , RIa1675d0_10);
buf \U$38 ( \196 , RIb4c6860_42);
xor \U$39 ( \197 , \195 , \196 );
or \U$40 ( \198 , \194 , \197 );
buf \U$41 ( \199 , RIa167558_11);
buf \U$42 ( \200 , RIb4c67e8_43);
xor \U$43 ( \201 , \199 , \200 );
or \U$44 ( \202 , \198 , \201 );
buf \U$45 ( \203 , RIa1674e0_12);
buf \U$46 ( \204 , RIb4c6770_44);
xor \U$47 ( \205 , \203 , \204 );
or \U$48 ( \206 , \202 , \205 );
buf \U$49 ( \207 , RIa167468_13);
buf \U$50 ( \208 , RIb4c3368_45);
xor \U$51 ( \209 , \207 , \208 );
or \U$52 ( \210 , \206 , \209 );
buf \U$53 ( \211 , RIa1673f0_14);
buf \U$54 ( \212 , RIb4c32f0_46);
xor \U$55 ( \213 , \211 , \212 );
or \U$56 ( \214 , \210 , \213 );
buf \U$57 ( \215 , RIa167378_15);
buf \U$58 ( \216 , RIb4c3278_47);
xor \U$59 ( \217 , \215 , \216 );
or \U$60 ( \218 , \214 , \217 );
buf \U$61 ( \219 , RIa167300_16);
buf \U$62 ( \220 , RIb4c3200_48);
xor \U$63 ( \221 , \219 , \220 );
or \U$64 ( \222 , \218 , \221 );
buf \U$65 ( \223 , RIa167288_17);
buf \U$66 ( \224 , RIb4c3188_49);
xor \U$67 ( \225 , \223 , \224 );
or \U$68 ( \226 , \222 , \225 );
buf \U$69 ( \227 , RIa167210_18);
buf \U$70 ( \228 , RIb4c3110_50);
xor \U$71 ( \229 , \227 , \228 );
or \U$72 ( \230 , \226 , \229 );
buf \U$73 ( \231 , RIa167198_19);
buf \U$74 ( \232 , RIb4c3098_51);
xor \U$75 ( \233 , \231 , \232 );
or \U$76 ( \234 , \230 , \233 );
buf \U$77 ( \235 , RIa167120_20);
buf \U$78 ( \236 , RIb4c3020_52);
xor \U$79 ( \237 , \235 , \236 );
or \U$80 ( \238 , \234 , \237 );
buf \U$81 ( \239 , RIa1670a8_21);
buf \U$82 ( \240 , RIb4c2fa8_53);
xor \U$83 ( \241 , \239 , \240 );
or \U$84 ( \242 , \238 , \241 );
buf \U$85 ( \243 , RIa167030_22);
buf \U$86 ( \244 , RIb4c2f30_54);
xor \U$87 ( \245 , \243 , \244 );
or \U$88 ( \246 , \242 , \245 );
buf \U$89 ( \247 , RIa166fb8_23);
buf \U$90 ( \248 , RIb4c2eb8_55);
xor \U$91 ( \249 , \247 , \248 );
or \U$92 ( \250 , \246 , \249 );
buf \U$93 ( \251 , RIa166f40_24);
buf \U$94 ( \252 , RIb4c2e40_56);
xor \U$95 ( \253 , \251 , \252 );
or \U$96 ( \254 , \250 , \253 );
buf \U$97 ( \255 , RIa166ec8_25);
buf \U$98 ( \256 , RIb4c2dc8_57);
xor \U$99 ( \257 , \255 , \256 );
or \U$100 ( \258 , \254 , \257 );
buf \U$101 ( \259 , RIa166e50_26);
buf \U$102 ( \260 , RIb4c2d50_58);
xor \U$103 ( \261 , \259 , \260 );
or \U$104 ( \262 , \258 , \261 );
buf \U$105 ( \263 , RIa166dd8_27);
buf \U$106 ( \264 , RIb4c2cd8_59);
xor \U$107 ( \265 , \263 , \264 );
or \U$108 ( \266 , \262 , \265 );
buf \U$109 ( \267 , RIa166d60_28);
buf \U$110 ( \268 , RIb4c2c60_60);
xor \U$111 ( \269 , \267 , \268 );
or \U$112 ( \270 , \266 , \269 );
buf \U$113 ( \271 , RIa166ce8_29);
buf \U$114 ( \272 , RIb4c2be8_61);
xor \U$115 ( \273 , \271 , \272 );
or \U$116 ( \274 , \270 , \273 );
buf \U$117 ( \275 , RIa166c70_30);
buf \U$118 ( \276 , RIb4c2b70_62);
xor \U$119 ( \277 , \275 , \276 );
or \U$120 ( \278 , \274 , \277 );
buf \U$121 ( \279 , RIb4ca4d8_31);
buf \U$122 ( \280 , RIb4c2af8_63);
xor \U$123 ( \281 , \279 , \280 );
or \U$124 ( \282 , \278 , \281 );
buf \U$125 ( \283 , RIb4ca460_32);
buf \U$126 ( \284 , RIb4bfab0_64);
xor \U$127 ( \285 , \283 , \284 );
or \U$128 ( \286 , \282 , \285 );
buf \U$129 ( \287 , \286 );
not \U$130 ( \288 , \287 );
_DC r13d ( \289_nR13d , RIb4c69c8_39 , \288 );
buf \U$131 ( \290 , \289_nR13d );
_DC r13c ( \291_nR13c , RIb4c6950_40 , \288 );
buf \U$132 ( \292 , \291_nR13c );
xor \U$133 ( \293 , \290 , \292 );
_DC r13b ( \294_nR13b , RIb4c68d8_41 , \288 );
buf \U$134 ( \295 , \294_nR13b );
xor \U$135 ( \296 , \292 , \295 );
not \U$136 ( \297 , \296 );
and \U$137 ( \298 , \293 , \297 );
and \U$138 ( \299 , \159 , \298 );
not \U$139 ( \300 , \299 );
and \U$140 ( \301 , \292 , \295 );
not \U$141 ( \302 , \301 );
and \U$142 ( \303 , \290 , \302 );
xnor \U$143 ( \304 , \300 , \303 );
buf \U$144 ( \305 , RIb4bf948_67);
_DC r13f ( \306_nR13f , RIb4c6ab8_37 , \288 );
buf \U$145 ( \307 , \306_nR13f );
_DC r13e ( \308_nR13e , RIb4c6a40_38 , \288 );
buf \U$146 ( \309 , \308_nR13e );
xor \U$147 ( \310 , \307 , \309 );
xor \U$148 ( \311 , \309 , \290 );
not \U$149 ( \312 , \311 );
and \U$150 ( \313 , \310 , \312 );
and \U$151 ( \314 , \305 , \313 );
buf \U$152 ( \315 , RIb4bf9c0_66);
and \U$153 ( \316 , \315 , \311 );
nor \U$154 ( \317 , \314 , \316 );
and \U$155 ( \318 , \309 , \290 );
not \U$156 ( \319 , \318 );
and \U$157 ( \320 , \307 , \319 );
xnor \U$158 ( \321 , \317 , \320 );
and \U$159 ( \322 , \304 , \321 );
buf \U$160 ( \323 , RIb4bf858_69);
_DC r141 ( \324_nR141 , RIb4c6ba8_35 , \288 );
buf \U$161 ( \325 , \324_nR141 );
_DC r140 ( \326_nR140 , RIb4c6b30_36 , \288 );
buf \U$162 ( \327 , \326_nR140 );
xor \U$163 ( \328 , \325 , \327 );
xor \U$164 ( \329 , \327 , \307 );
not \U$165 ( \330 , \329 );
and \U$166 ( \331 , \328 , \330 );
and \U$167 ( \332 , \323 , \331 );
buf \U$168 ( \333 , RIb4bf8d0_68);
and \U$169 ( \334 , \333 , \329 );
nor \U$170 ( \335 , \332 , \334 );
and \U$171 ( \336 , \327 , \307 );
not \U$172 ( \337 , \336 );
and \U$173 ( \338 , \325 , \337 );
xnor \U$174 ( \339 , \335 , \338 );
and \U$175 ( \340 , \321 , \339 );
and \U$176 ( \341 , \304 , \339 );
or \U$177 ( \342 , \322 , \340 , \341 );
buf \U$178 ( \343 , RIb4bf768_71);
_DC r143 ( \344_nR143 , RIb4ca3e8_33 , \288 );
buf \U$179 ( \345 , \344_nR143 );
_DC r142 ( \346_nR142 , RIb4c6c20_34 , \288 );
buf \U$180 ( \347 , \346_nR142 );
xor \U$181 ( \348 , \345 , \347 );
xor \U$182 ( \349 , \347 , \325 );
not \U$183 ( \350 , \349 );
and \U$184 ( \351 , \348 , \350 );
and \U$185 ( \352 , \343 , \351 );
buf \U$186 ( \353 , RIb4bf7e0_70);
and \U$187 ( \354 , \353 , \349 );
nor \U$188 ( \355 , \352 , \354 );
and \U$189 ( \356 , \347 , \325 );
not \U$190 ( \357 , \356 );
and \U$191 ( \358 , \345 , \357 );
xnor \U$192 ( \359 , \355 , \358 );
buf \U$193 ( \360 , RIb4bf6f0_72);
and \U$194 ( \361 , \360 , \345 );
or \U$195 ( \362 , \359 , \361 );
and \U$196 ( \363 , \342 , \362 );
and \U$197 ( \364 , \353 , \351 );
and \U$198 ( \365 , \323 , \349 );
nor \U$199 ( \366 , \364 , \365 );
xnor \U$200 ( \367 , \366 , \358 );
and \U$201 ( \368 , \362 , \367 );
and \U$202 ( \369 , \342 , \367 );
or \U$203 ( \370 , \363 , \368 , \369 );
and \U$204 ( \371 , \343 , \345 );
not \U$205 ( \372 , \303 );
and \U$206 ( \373 , \315 , \313 );
and \U$207 ( \374 , \159 , \311 );
nor \U$208 ( \375 , \373 , \374 );
xnor \U$209 ( \376 , \375 , \320 );
xor \U$210 ( \377 , \372 , \376 );
and \U$211 ( \378 , \333 , \331 );
and \U$212 ( \379 , \305 , \329 );
nor \U$213 ( \380 , \378 , \379 );
xnor \U$214 ( \381 , \380 , \338 );
xor \U$215 ( \382 , \377 , \381 );
and \U$216 ( \383 , \371 , \382 );
and \U$217 ( \384 , \370 , \383 );
and \U$218 ( \385 , \372 , \376 );
and \U$219 ( \386 , \376 , \381 );
and \U$220 ( \387 , \372 , \381 );
or \U$221 ( \388 , \385 , \386 , \387 );
and \U$222 ( \389 , \159 , \313 );
not \U$223 ( \390 , \389 );
xnor \U$224 ( \391 , \390 , \320 );
and \U$225 ( \392 , \305 , \331 );
and \U$226 ( \393 , \315 , \329 );
nor \U$227 ( \394 , \392 , \393 );
xnor \U$228 ( \395 , \394 , \338 );
xor \U$229 ( \396 , \391 , \395 );
and \U$230 ( \397 , \323 , \351 );
and \U$231 ( \398 , \333 , \349 );
nor \U$232 ( \399 , \397 , \398 );
xnor \U$233 ( \400 , \399 , \358 );
xor \U$234 ( \401 , \396 , \400 );
xor \U$235 ( \402 , \388 , \401 );
and \U$236 ( \403 , \353 , \345 );
not \U$237 ( \404 , \403 );
xor \U$238 ( \405 , \402 , \404 );
and \U$239 ( \406 , \383 , \405 );
and \U$240 ( \407 , \370 , \405 );
or \U$241 ( \408 , \384 , \406 , \407 );
and \U$242 ( \409 , \388 , \401 );
and \U$243 ( \410 , \401 , \404 );
and \U$244 ( \411 , \388 , \404 );
or \U$245 ( \412 , \409 , \410 , \411 );
not \U$246 ( \413 , \320 );
and \U$247 ( \414 , \315 , \331 );
and \U$248 ( \415 , \159 , \329 );
nor \U$249 ( \416 , \414 , \415 );
xnor \U$250 ( \417 , \416 , \338 );
xor \U$251 ( \418 , \413 , \417 );
and \U$252 ( \419 , \333 , \351 );
and \U$253 ( \420 , \305 , \349 );
nor \U$254 ( \421 , \419 , \420 );
xnor \U$255 ( \422 , \421 , \358 );
xor \U$256 ( \423 , \418 , \422 );
xor \U$257 ( \424 , \412 , \423 );
and \U$258 ( \425 , \391 , \395 );
and \U$259 ( \426 , \395 , \400 );
and \U$260 ( \427 , \391 , \400 );
or \U$261 ( \428 , \425 , \426 , \427 );
buf \U$262 ( \429 , \403 );
xor \U$263 ( \430 , \428 , \429 );
and \U$264 ( \431 , \323 , \345 );
xor \U$265 ( \432 , \430 , \431 );
xor \U$266 ( \433 , \424 , \432 );
xor \U$267 ( \434 , \408 , \433 );
and \U$268 ( \435 , \353 , \331 );
and \U$269 ( \436 , \323 , \329 );
nor \U$270 ( \437 , \435 , \436 );
xnor \U$271 ( \438 , \437 , \338 );
and \U$272 ( \439 , \360 , \351 );
and \U$273 ( \440 , \343 , \349 );
nor \U$274 ( \441 , \439 , \440 );
xnor \U$275 ( \442 , \441 , \358 );
and \U$276 ( \443 , \438 , \442 );
buf \U$277 ( \444 , RIb4bf678_73);
and \U$278 ( \445 , \444 , \345 );
and \U$279 ( \446 , \442 , \445 );
and \U$280 ( \447 , \438 , \445 );
or \U$281 ( \448 , \443 , \446 , \447 );
_DC r13a ( \449_nR13a , RIb4c6860_42 , \288 );
buf \U$282 ( \450 , \449_nR13a );
_DC r139 ( \451_nR139 , RIb4c67e8_43 , \288 );
buf \U$283 ( \452 , \451_nR139 );
and \U$284 ( \453 , \450 , \452 );
not \U$285 ( \454 , \453 );
and \U$286 ( \455 , \295 , \454 );
not \U$287 ( \456 , \455 );
and \U$288 ( \457 , \315 , \298 );
and \U$289 ( \458 , \159 , \296 );
nor \U$290 ( \459 , \457 , \458 );
xnor \U$291 ( \460 , \459 , \303 );
and \U$292 ( \461 , \456 , \460 );
and \U$293 ( \462 , \333 , \313 );
and \U$294 ( \463 , \305 , \311 );
nor \U$295 ( \464 , \462 , \463 );
xnor \U$296 ( \465 , \464 , \320 );
and \U$297 ( \466 , \460 , \465 );
and \U$298 ( \467 , \456 , \465 );
or \U$299 ( \468 , \461 , \466 , \467 );
and \U$300 ( \469 , \448 , \468 );
xnor \U$301 ( \470 , \359 , \361 );
and \U$302 ( \471 , \468 , \470 );
and \U$303 ( \472 , \448 , \470 );
or \U$304 ( \473 , \469 , \471 , \472 );
xor \U$305 ( \474 , \342 , \362 );
xor \U$306 ( \475 , \474 , \367 );
and \U$307 ( \476 , \473 , \475 );
xor \U$308 ( \477 , \371 , \382 );
and \U$309 ( \478 , \475 , \477 );
and \U$310 ( \479 , \473 , \477 );
or \U$311 ( \480 , \476 , \478 , \479 );
xor \U$312 ( \481 , \370 , \383 );
xor \U$313 ( \482 , \481 , \405 );
and \U$314 ( \483 , \480 , \482 );
xor \U$315 ( \484 , \434 , \483 );
xor \U$316 ( \485 , \480 , \482 );
and \U$317 ( \486 , \343 , \331 );
and \U$318 ( \487 , \353 , \329 );
nor \U$319 ( \488 , \486 , \487 );
xnor \U$320 ( \489 , \488 , \338 );
and \U$321 ( \490 , \444 , \351 );
and \U$322 ( \491 , \360 , \349 );
nor \U$323 ( \492 , \490 , \491 );
xnor \U$324 ( \493 , \492 , \358 );
and \U$325 ( \494 , \489 , \493 );
buf \U$326 ( \495 , RIb4bf600_74);
and \U$327 ( \496 , \495 , \345 );
and \U$328 ( \497 , \493 , \496 );
and \U$329 ( \498 , \489 , \496 );
or \U$330 ( \499 , \494 , \497 , \498 );
xor \U$331 ( \500 , \295 , \450 );
xor \U$332 ( \501 , \450 , \452 );
not \U$333 ( \502 , \501 );
and \U$334 ( \503 , \500 , \502 );
and \U$335 ( \504 , \159 , \503 );
not \U$336 ( \505 , \504 );
xnor \U$337 ( \506 , \505 , \455 );
and \U$338 ( \507 , \305 , \298 );
and \U$339 ( \508 , \315 , \296 );
nor \U$340 ( \509 , \507 , \508 );
xnor \U$341 ( \510 , \509 , \303 );
and \U$342 ( \511 , \506 , \510 );
and \U$343 ( \512 , \323 , \313 );
and \U$344 ( \513 , \333 , \311 );
nor \U$345 ( \514 , \512 , \513 );
xnor \U$346 ( \515 , \514 , \320 );
and \U$347 ( \516 , \510 , \515 );
and \U$348 ( \517 , \506 , \515 );
or \U$349 ( \518 , \511 , \516 , \517 );
and \U$350 ( \519 , \499 , \518 );
xor \U$351 ( \520 , \438 , \442 );
xor \U$352 ( \521 , \520 , \445 );
and \U$353 ( \522 , \518 , \521 );
and \U$354 ( \523 , \499 , \521 );
or \U$355 ( \524 , \519 , \522 , \523 );
xor \U$356 ( \525 , \304 , \321 );
xor \U$357 ( \526 , \525 , \339 );
and \U$358 ( \527 , \524 , \526 );
xor \U$359 ( \528 , \448 , \468 );
xor \U$360 ( \529 , \528 , \470 );
and \U$361 ( \530 , \526 , \529 );
and \U$362 ( \531 , \524 , \529 );
or \U$363 ( \532 , \527 , \530 , \531 );
xor \U$364 ( \533 , \473 , \475 );
xor \U$365 ( \534 , \533 , \477 );
and \U$366 ( \535 , \532 , \534 );
and \U$367 ( \536 , \485 , \535 );
xor \U$368 ( \537 , \485 , \535 );
xor \U$369 ( \538 , \532 , \534 );
and \U$370 ( \539 , \353 , \313 );
and \U$371 ( \540 , \323 , \311 );
nor \U$372 ( \541 , \539 , \540 );
xnor \U$373 ( \542 , \541 , \320 );
and \U$374 ( \543 , \360 , \331 );
and \U$375 ( \544 , \343 , \329 );
nor \U$376 ( \545 , \543 , \544 );
xnor \U$377 ( \546 , \545 , \338 );
and \U$378 ( \547 , \542 , \546 );
and \U$379 ( \548 , \495 , \351 );
and \U$380 ( \549 , \444 , \349 );
nor \U$381 ( \550 , \548 , \549 );
xnor \U$382 ( \551 , \550 , \358 );
and \U$383 ( \552 , \546 , \551 );
and \U$384 ( \553 , \542 , \551 );
or \U$385 ( \554 , \547 , \552 , \553 );
_DC r138 ( \555_nR138 , RIb4c6770_44 , \288 );
buf \U$386 ( \556 , \555_nR138 );
_DC r137 ( \557_nR137 , RIb4c3368_45 , \288 );
buf \U$387 ( \558 , \557_nR137 );
and \U$388 ( \559 , \556 , \558 );
not \U$389 ( \560 , \559 );
and \U$390 ( \561 , \452 , \560 );
not \U$391 ( \562 , \561 );
and \U$392 ( \563 , \315 , \503 );
and \U$393 ( \564 , \159 , \501 );
nor \U$394 ( \565 , \563 , \564 );
xnor \U$395 ( \566 , \565 , \455 );
and \U$396 ( \567 , \562 , \566 );
and \U$397 ( \568 , \333 , \298 );
and \U$398 ( \569 , \305 , \296 );
nor \U$399 ( \570 , \568 , \569 );
xnor \U$400 ( \571 , \570 , \303 );
and \U$401 ( \572 , \566 , \571 );
and \U$402 ( \573 , \562 , \571 );
or \U$403 ( \574 , \567 , \572 , \573 );
or \U$404 ( \575 , \554 , \574 );
xor \U$405 ( \576 , \456 , \460 );
xor \U$406 ( \577 , \576 , \465 );
and \U$407 ( \578 , \575 , \577 );
xor \U$408 ( \579 , \499 , \518 );
xor \U$409 ( \580 , \579 , \521 );
and \U$410 ( \581 , \577 , \580 );
and \U$411 ( \582 , \575 , \580 );
or \U$412 ( \583 , \578 , \581 , \582 );
and \U$413 ( \584 , \343 , \313 );
and \U$414 ( \585 , \353 , \311 );
nor \U$415 ( \586 , \584 , \585 );
xnor \U$416 ( \587 , \586 , \320 );
and \U$417 ( \588 , \444 , \331 );
and \U$418 ( \589 , \360 , \329 );
nor \U$419 ( \590 , \588 , \589 );
xnor \U$420 ( \591 , \590 , \338 );
and \U$421 ( \592 , \587 , \591 );
buf \U$422 ( \593 , RIb4bf588_75);
and \U$423 ( \594 , \593 , \351 );
and \U$424 ( \595 , \495 , \349 );
nor \U$425 ( \596 , \594 , \595 );
xnor \U$426 ( \597 , \596 , \358 );
and \U$427 ( \598 , \591 , \597 );
and \U$428 ( \599 , \587 , \597 );
or \U$429 ( \600 , \592 , \598 , \599 );
xor \U$430 ( \601 , \452 , \556 );
xor \U$431 ( \602 , \556 , \558 );
not \U$432 ( \603 , \602 );
and \U$433 ( \604 , \601 , \603 );
and \U$434 ( \605 , \159 , \604 );
not \U$435 ( \606 , \605 );
xnor \U$436 ( \607 , \606 , \561 );
and \U$437 ( \608 , \305 , \503 );
and \U$438 ( \609 , \315 , \501 );
nor \U$439 ( \610 , \608 , \609 );
xnor \U$440 ( \611 , \610 , \455 );
and \U$441 ( \612 , \607 , \611 );
and \U$442 ( \613 , \323 , \298 );
and \U$443 ( \614 , \333 , \296 );
nor \U$444 ( \615 , \613 , \614 );
xnor \U$445 ( \616 , \615 , \303 );
and \U$446 ( \617 , \611 , \616 );
and \U$447 ( \618 , \607 , \616 );
or \U$448 ( \619 , \612 , \617 , \618 );
and \U$449 ( \620 , \600 , \619 );
buf \U$450 ( \621 , RIb4bf510_76);
and \U$451 ( \622 , \621 , \345 );
buf \U$452 ( \623 , \622 );
and \U$453 ( \624 , \619 , \623 );
and \U$454 ( \625 , \600 , \623 );
or \U$455 ( \626 , \620 , \624 , \625 );
and \U$456 ( \627 , \593 , \345 );
xor \U$457 ( \628 , \542 , \546 );
xor \U$458 ( \629 , \628 , \551 );
and \U$459 ( \630 , \627 , \629 );
xor \U$460 ( \631 , \562 , \566 );
xor \U$461 ( \632 , \631 , \571 );
and \U$462 ( \633 , \629 , \632 );
and \U$463 ( \634 , \627 , \632 );
or \U$464 ( \635 , \630 , \633 , \634 );
and \U$465 ( \636 , \626 , \635 );
xor \U$466 ( \637 , \489 , \493 );
xor \U$467 ( \638 , \637 , \496 );
and \U$468 ( \639 , \635 , \638 );
and \U$469 ( \640 , \626 , \638 );
or \U$470 ( \641 , \636 , \639 , \640 );
xor \U$471 ( \642 , \506 , \510 );
xor \U$472 ( \643 , \642 , \515 );
xnor \U$473 ( \644 , \554 , \574 );
and \U$474 ( \645 , \643 , \644 );
and \U$475 ( \646 , \641 , \645 );
xor \U$476 ( \647 , \575 , \577 );
xor \U$477 ( \648 , \647 , \580 );
and \U$478 ( \649 , \645 , \648 );
and \U$479 ( \650 , \641 , \648 );
or \U$480 ( \651 , \646 , \649 , \650 );
and \U$481 ( \652 , \583 , \651 );
xor \U$482 ( \653 , \524 , \526 );
xor \U$483 ( \654 , \653 , \529 );
and \U$484 ( \655 , \651 , \654 );
and \U$485 ( \656 , \583 , \654 );
or \U$486 ( \657 , \652 , \655 , \656 );
and \U$487 ( \658 , \538 , \657 );
xor \U$488 ( \659 , \538 , \657 );
xor \U$489 ( \660 , \583 , \651 );
xor \U$490 ( \661 , \660 , \654 );
_DC r136 ( \662_nR136 , RIb4c32f0_46 , \288 );
buf \U$491 ( \663 , \662_nR136 );
_DC r135 ( \664_nR135 , RIb4c3278_47 , \288 );
buf \U$492 ( \665 , \664_nR135 );
and \U$493 ( \666 , \663 , \665 );
not \U$494 ( \667 , \666 );
and \U$495 ( \668 , \558 , \667 );
not \U$496 ( \669 , \668 );
and \U$497 ( \670 , \315 , \604 );
and \U$498 ( \671 , \159 , \602 );
nor \U$499 ( \672 , \670 , \671 );
xnor \U$500 ( \673 , \672 , \561 );
and \U$501 ( \674 , \669 , \673 );
and \U$502 ( \675 , \333 , \503 );
and \U$503 ( \676 , \305 , \501 );
nor \U$504 ( \677 , \675 , \676 );
xnor \U$505 ( \678 , \677 , \455 );
and \U$506 ( \679 , \673 , \678 );
and \U$507 ( \680 , \669 , \678 );
or \U$508 ( \681 , \674 , \679 , \680 );
and \U$509 ( \682 , \353 , \298 );
and \U$510 ( \683 , \323 , \296 );
nor \U$511 ( \684 , \682 , \683 );
xnor \U$512 ( \685 , \684 , \303 );
and \U$513 ( \686 , \360 , \313 );
and \U$514 ( \687 , \343 , \311 );
nor \U$515 ( \688 , \686 , \687 );
xnor \U$516 ( \689 , \688 , \320 );
and \U$517 ( \690 , \685 , \689 );
and \U$518 ( \691 , \495 , \331 );
and \U$519 ( \692 , \444 , \329 );
nor \U$520 ( \693 , \691 , \692 );
xnor \U$521 ( \694 , \693 , \338 );
and \U$522 ( \695 , \689 , \694 );
and \U$523 ( \696 , \685 , \694 );
or \U$524 ( \697 , \690 , \695 , \696 );
and \U$525 ( \698 , \681 , \697 );
and \U$526 ( \699 , \621 , \351 );
and \U$527 ( \700 , \593 , \349 );
nor \U$528 ( \701 , \699 , \700 );
xnor \U$529 ( \702 , \701 , \358 );
buf \U$530 ( \703 , RIb4bf498_77);
and \U$531 ( \704 , \703 , \345 );
and \U$532 ( \705 , \702 , \704 );
and \U$533 ( \706 , \697 , \705 );
and \U$534 ( \707 , \681 , \705 );
or \U$535 ( \708 , \698 , \706 , \707 );
xor \U$536 ( \709 , \587 , \591 );
xor \U$537 ( \710 , \709 , \597 );
xor \U$538 ( \711 , \607 , \611 );
xor \U$539 ( \712 , \711 , \616 );
and \U$540 ( \713 , \710 , \712 );
not \U$541 ( \714 , \622 );
and \U$542 ( \715 , \712 , \714 );
and \U$543 ( \716 , \710 , \714 );
or \U$544 ( \717 , \713 , \715 , \716 );
and \U$545 ( \718 , \708 , \717 );
xor \U$546 ( \719 , \627 , \629 );
xor \U$547 ( \720 , \719 , \632 );
and \U$548 ( \721 , \717 , \720 );
and \U$549 ( \722 , \708 , \720 );
or \U$550 ( \723 , \718 , \721 , \722 );
xor \U$551 ( \724 , \626 , \635 );
xor \U$552 ( \725 , \724 , \638 );
and \U$553 ( \726 , \723 , \725 );
xor \U$554 ( \727 , \643 , \644 );
and \U$555 ( \728 , \725 , \727 );
and \U$556 ( \729 , \723 , \727 );
or \U$557 ( \730 , \726 , \728 , \729 );
xor \U$558 ( \731 , \641 , \645 );
xor \U$559 ( \732 , \731 , \648 );
and \U$560 ( \733 , \730 , \732 );
and \U$561 ( \734 , \661 , \733 );
xor \U$562 ( \735 , \661 , \733 );
xor \U$563 ( \736 , \730 , \732 );
xor \U$564 ( \737 , \558 , \663 );
xor \U$565 ( \738 , \663 , \665 );
not \U$566 ( \739 , \738 );
and \U$567 ( \740 , \737 , \739 );
and \U$568 ( \741 , \159 , \740 );
not \U$569 ( \742 , \741 );
xnor \U$570 ( \743 , \742 , \668 );
and \U$571 ( \744 , \305 , \604 );
and \U$572 ( \745 , \315 , \602 );
nor \U$573 ( \746 , \744 , \745 );
xnor \U$574 ( \747 , \746 , \561 );
and \U$575 ( \748 , \743 , \747 );
and \U$576 ( \749 , \323 , \503 );
and \U$577 ( \750 , \333 , \501 );
nor \U$578 ( \751 , \749 , \750 );
xnor \U$579 ( \752 , \751 , \455 );
and \U$580 ( \753 , \747 , \752 );
and \U$581 ( \754 , \743 , \752 );
or \U$582 ( \755 , \748 , \753 , \754 );
and \U$583 ( \756 , \343 , \298 );
and \U$584 ( \757 , \353 , \296 );
nor \U$585 ( \758 , \756 , \757 );
xnor \U$586 ( \759 , \758 , \303 );
and \U$587 ( \760 , \444 , \313 );
and \U$588 ( \761 , \360 , \311 );
nor \U$589 ( \762 , \760 , \761 );
xnor \U$590 ( \763 , \762 , \320 );
and \U$591 ( \764 , \759 , \763 );
and \U$592 ( \765 , \593 , \331 );
and \U$593 ( \766 , \495 , \329 );
nor \U$594 ( \767 , \765 , \766 );
xnor \U$595 ( \768 , \767 , \338 );
and \U$596 ( \769 , \763 , \768 );
and \U$597 ( \770 , \759 , \768 );
or \U$598 ( \771 , \764 , \769 , \770 );
and \U$599 ( \772 , \755 , \771 );
and \U$600 ( \773 , \703 , \351 );
and \U$601 ( \774 , \621 , \349 );
nor \U$602 ( \775 , \773 , \774 );
xnor \U$603 ( \776 , \775 , \358 );
buf \U$604 ( \777 , RIb4bf420_78);
and \U$605 ( \778 , \777 , \345 );
or \U$606 ( \779 , \776 , \778 );
and \U$607 ( \780 , \771 , \779 );
and \U$608 ( \781 , \755 , \779 );
or \U$609 ( \782 , \772 , \780 , \781 );
xor \U$610 ( \783 , \669 , \673 );
xor \U$611 ( \784 , \783 , \678 );
xor \U$612 ( \785 , \685 , \689 );
xor \U$613 ( \786 , \785 , \694 );
and \U$614 ( \787 , \784 , \786 );
xor \U$615 ( \788 , \702 , \704 );
and \U$616 ( \789 , \786 , \788 );
and \U$617 ( \790 , \784 , \788 );
or \U$618 ( \791 , \787 , \789 , \790 );
and \U$619 ( \792 , \782 , \791 );
xor \U$620 ( \793 , \710 , \712 );
xor \U$621 ( \794 , \793 , \714 );
and \U$622 ( \795 , \791 , \794 );
and \U$623 ( \796 , \782 , \794 );
or \U$624 ( \797 , \792 , \795 , \796 );
xor \U$625 ( \798 , \600 , \619 );
xor \U$626 ( \799 , \798 , \623 );
and \U$627 ( \800 , \797 , \799 );
xor \U$628 ( \801 , \708 , \717 );
xor \U$629 ( \802 , \801 , \720 );
and \U$630 ( \803 , \799 , \802 );
and \U$631 ( \804 , \797 , \802 );
or \U$632 ( \805 , \800 , \803 , \804 );
xor \U$633 ( \806 , \723 , \725 );
xor \U$634 ( \807 , \806 , \727 );
and \U$635 ( \808 , \805 , \807 );
and \U$636 ( \809 , \736 , \808 );
xor \U$637 ( \810 , \736 , \808 );
xor \U$638 ( \811 , \805 , \807 );
_DC r134 ( \812_nR134 , RIb4c3200_48 , \288 );
buf \U$639 ( \813 , \812_nR134 );
_DC r133 ( \814_nR133 , RIb4c3188_49 , \288 );
buf \U$640 ( \815 , \814_nR133 );
and \U$641 ( \816 , \813 , \815 );
not \U$642 ( \817 , \816 );
and \U$643 ( \818 , \665 , \817 );
not \U$644 ( \819 , \818 );
and \U$645 ( \820 , \315 , \740 );
and \U$646 ( \821 , \159 , \738 );
nor \U$647 ( \822 , \820 , \821 );
xnor \U$648 ( \823 , \822 , \668 );
and \U$649 ( \824 , \819 , \823 );
and \U$650 ( \825 , \333 , \604 );
and \U$651 ( \826 , \305 , \602 );
nor \U$652 ( \827 , \825 , \826 );
xnor \U$653 ( \828 , \827 , \561 );
and \U$654 ( \829 , \823 , \828 );
and \U$655 ( \830 , \819 , \828 );
or \U$656 ( \831 , \824 , \829 , \830 );
and \U$657 ( \832 , \621 , \331 );
and \U$658 ( \833 , \593 , \329 );
nor \U$659 ( \834 , \832 , \833 );
xnor \U$660 ( \835 , \834 , \338 );
and \U$661 ( \836 , \777 , \351 );
and \U$662 ( \837 , \703 , \349 );
nor \U$663 ( \838 , \836 , \837 );
xnor \U$664 ( \839 , \838 , \358 );
and \U$665 ( \840 , \835 , \839 );
buf \U$666 ( \841 , RIb4bf3a8_79);
and \U$667 ( \842 , \841 , \345 );
and \U$668 ( \843 , \839 , \842 );
and \U$669 ( \844 , \835 , \842 );
or \U$670 ( \845 , \840 , \843 , \844 );
and \U$671 ( \846 , \831 , \845 );
and \U$672 ( \847 , \353 , \503 );
and \U$673 ( \848 , \323 , \501 );
nor \U$674 ( \849 , \847 , \848 );
xnor \U$675 ( \850 , \849 , \455 );
and \U$676 ( \851 , \360 , \298 );
and \U$677 ( \852 , \343 , \296 );
nor \U$678 ( \853 , \851 , \852 );
xnor \U$679 ( \854 , \853 , \303 );
and \U$680 ( \855 , \850 , \854 );
and \U$681 ( \856 , \495 , \313 );
and \U$682 ( \857 , \444 , \311 );
nor \U$683 ( \858 , \856 , \857 );
xnor \U$684 ( \859 , \858 , \320 );
and \U$685 ( \860 , \854 , \859 );
and \U$686 ( \861 , \850 , \859 );
or \U$687 ( \862 , \855 , \860 , \861 );
and \U$688 ( \863 , \845 , \862 );
and \U$689 ( \864 , \831 , \862 );
or \U$690 ( \865 , \846 , \863 , \864 );
xor \U$691 ( \866 , \743 , \747 );
xor \U$692 ( \867 , \866 , \752 );
xor \U$693 ( \868 , \759 , \763 );
xor \U$694 ( \869 , \868 , \768 );
and \U$695 ( \870 , \867 , \869 );
xnor \U$696 ( \871 , \776 , \778 );
and \U$697 ( \872 , \869 , \871 );
and \U$698 ( \873 , \867 , \871 );
or \U$699 ( \874 , \870 , \872 , \873 );
and \U$700 ( \875 , \865 , \874 );
xor \U$701 ( \876 , \784 , \786 );
xor \U$702 ( \877 , \876 , \788 );
and \U$703 ( \878 , \874 , \877 );
and \U$704 ( \879 , \865 , \877 );
or \U$705 ( \880 , \875 , \878 , \879 );
xor \U$706 ( \881 , \681 , \697 );
xor \U$707 ( \882 , \881 , \705 );
and \U$708 ( \883 , \880 , \882 );
xor \U$709 ( \884 , \782 , \791 );
xor \U$710 ( \885 , \884 , \794 );
and \U$711 ( \886 , \882 , \885 );
and \U$712 ( \887 , \880 , \885 );
or \U$713 ( \888 , \883 , \886 , \887 );
xor \U$714 ( \889 , \797 , \799 );
xor \U$715 ( \890 , \889 , \802 );
and \U$716 ( \891 , \888 , \890 );
and \U$717 ( \892 , \811 , \891 );
xor \U$718 ( \893 , \811 , \891 );
xor \U$719 ( \894 , \888 , \890 );
and \U$720 ( \895 , \703 , \331 );
and \U$721 ( \896 , \621 , \329 );
nor \U$722 ( \897 , \895 , \896 );
xnor \U$723 ( \898 , \897 , \338 );
and \U$724 ( \899 , \841 , \351 );
and \U$725 ( \900 , \777 , \349 );
nor \U$726 ( \901 , \899 , \900 );
xnor \U$727 ( \902 , \901 , \358 );
and \U$728 ( \903 , \898 , \902 );
buf \U$729 ( \904 , RIb4bf330_80);
and \U$730 ( \905 , \904 , \345 );
and \U$731 ( \906 , \902 , \905 );
and \U$732 ( \907 , \898 , \905 );
or \U$733 ( \908 , \903 , \906 , \907 );
xor \U$734 ( \909 , \665 , \813 );
xor \U$735 ( \910 , \813 , \815 );
not \U$736 ( \911 , \910 );
and \U$737 ( \912 , \909 , \911 );
and \U$738 ( \913 , \159 , \912 );
not \U$739 ( \914 , \913 );
xnor \U$740 ( \915 , \914 , \818 );
and \U$741 ( \916 , \305 , \740 );
and \U$742 ( \917 , \315 , \738 );
nor \U$743 ( \918 , \916 , \917 );
xnor \U$744 ( \919 , \918 , \668 );
and \U$745 ( \920 , \915 , \919 );
and \U$746 ( \921 , \323 , \604 );
and \U$747 ( \922 , \333 , \602 );
nor \U$748 ( \923 , \921 , \922 );
xnor \U$749 ( \924 , \923 , \561 );
and \U$750 ( \925 , \919 , \924 );
and \U$751 ( \926 , \915 , \924 );
or \U$752 ( \927 , \920 , \925 , \926 );
and \U$753 ( \928 , \908 , \927 );
and \U$754 ( \929 , \343 , \503 );
and \U$755 ( \930 , \353 , \501 );
nor \U$756 ( \931 , \929 , \930 );
xnor \U$757 ( \932 , \931 , \455 );
and \U$758 ( \933 , \444 , \298 );
and \U$759 ( \934 , \360 , \296 );
nor \U$760 ( \935 , \933 , \934 );
xnor \U$761 ( \936 , \935 , \303 );
and \U$762 ( \937 , \932 , \936 );
and \U$763 ( \938 , \593 , \313 );
and \U$764 ( \939 , \495 , \311 );
nor \U$765 ( \940 , \938 , \939 );
xnor \U$766 ( \941 , \940 , \320 );
and \U$767 ( \942 , \936 , \941 );
and \U$768 ( \943 , \932 , \941 );
or \U$769 ( \944 , \937 , \942 , \943 );
and \U$770 ( \945 , \927 , \944 );
and \U$771 ( \946 , \908 , \944 );
or \U$772 ( \947 , \928 , \945 , \946 );
xor \U$773 ( \948 , \819 , \823 );
xor \U$774 ( \949 , \948 , \828 );
xor \U$775 ( \950 , \835 , \839 );
xor \U$776 ( \951 , \950 , \842 );
and \U$777 ( \952 , \949 , \951 );
xor \U$778 ( \953 , \850 , \854 );
xor \U$779 ( \954 , \953 , \859 );
and \U$780 ( \955 , \951 , \954 );
and \U$781 ( \956 , \949 , \954 );
or \U$782 ( \957 , \952 , \955 , \956 );
and \U$783 ( \958 , \947 , \957 );
xor \U$784 ( \959 , \867 , \869 );
xor \U$785 ( \960 , \959 , \871 );
and \U$786 ( \961 , \957 , \960 );
and \U$787 ( \962 , \947 , \960 );
or \U$788 ( \963 , \958 , \961 , \962 );
xor \U$789 ( \964 , \755 , \771 );
xor \U$790 ( \965 , \964 , \779 );
and \U$791 ( \966 , \963 , \965 );
xor \U$792 ( \967 , \865 , \874 );
xor \U$793 ( \968 , \967 , \877 );
and \U$794 ( \969 , \965 , \968 );
and \U$795 ( \970 , \963 , \968 );
or \U$796 ( \971 , \966 , \969 , \970 );
xor \U$797 ( \972 , \880 , \882 );
xor \U$798 ( \973 , \972 , \885 );
and \U$799 ( \974 , \971 , \973 );
and \U$800 ( \975 , \894 , \974 );
xor \U$801 ( \976 , \894 , \974 );
xor \U$802 ( \977 , \971 , \973 );
_DC r132 ( \978_nR132 , RIb4c3110_50 , \288 );
buf \U$803 ( \979 , \978_nR132 );
_DC r131 ( \980_nR131 , RIb4c3098_51 , \288 );
buf \U$804 ( \981 , \980_nR131 );
and \U$805 ( \982 , \979 , \981 );
not \U$806 ( \983 , \982 );
and \U$807 ( \984 , \815 , \983 );
not \U$808 ( \985 , \984 );
and \U$809 ( \986 , \315 , \912 );
and \U$810 ( \987 , \159 , \910 );
nor \U$811 ( \988 , \986 , \987 );
xnor \U$812 ( \989 , \988 , \818 );
and \U$813 ( \990 , \985 , \989 );
and \U$814 ( \991 , \333 , \740 );
and \U$815 ( \992 , \305 , \738 );
nor \U$816 ( \993 , \991 , \992 );
xnor \U$817 ( \994 , \993 , \668 );
and \U$818 ( \995 , \989 , \994 );
and \U$819 ( \996 , \985 , \994 );
or \U$820 ( \997 , \990 , \995 , \996 );
and \U$821 ( \998 , \353 , \604 );
and \U$822 ( \999 , \323 , \602 );
nor \U$823 ( \1000 , \998 , \999 );
xnor \U$824 ( \1001 , \1000 , \561 );
and \U$825 ( \1002 , \360 , \503 );
and \U$826 ( \1003 , \343 , \501 );
nor \U$827 ( \1004 , \1002 , \1003 );
xnor \U$828 ( \1005 , \1004 , \455 );
and \U$829 ( \1006 , \1001 , \1005 );
and \U$830 ( \1007 , \495 , \298 );
and \U$831 ( \1008 , \444 , \296 );
nor \U$832 ( \1009 , \1007 , \1008 );
xnor \U$833 ( \1010 , \1009 , \303 );
and \U$834 ( \1011 , \1005 , \1010 );
and \U$835 ( \1012 , \1001 , \1010 );
or \U$836 ( \1013 , \1006 , \1011 , \1012 );
and \U$837 ( \1014 , \997 , \1013 );
and \U$838 ( \1015 , \621 , \313 );
and \U$839 ( \1016 , \593 , \311 );
nor \U$840 ( \1017 , \1015 , \1016 );
xnor \U$841 ( \1018 , \1017 , \320 );
and \U$842 ( \1019 , \777 , \331 );
and \U$843 ( \1020 , \703 , \329 );
nor \U$844 ( \1021 , \1019 , \1020 );
xnor \U$845 ( \1022 , \1021 , \338 );
and \U$846 ( \1023 , \1018 , \1022 );
and \U$847 ( \1024 , \904 , \351 );
and \U$848 ( \1025 , \841 , \349 );
nor \U$849 ( \1026 , \1024 , \1025 );
xnor \U$850 ( \1027 , \1026 , \358 );
and \U$851 ( \1028 , \1022 , \1027 );
and \U$852 ( \1029 , \1018 , \1027 );
or \U$853 ( \1030 , \1023 , \1028 , \1029 );
and \U$854 ( \1031 , \1013 , \1030 );
and \U$855 ( \1032 , \997 , \1030 );
or \U$856 ( \1033 , \1014 , \1031 , \1032 );
xor \U$857 ( \1034 , \898 , \902 );
xor \U$858 ( \1035 , \1034 , \905 );
xor \U$859 ( \1036 , \932 , \936 );
xor \U$860 ( \1037 , \1036 , \941 );
or \U$861 ( \1038 , \1035 , \1037 );
and \U$862 ( \1039 , \1033 , \1038 );
xor \U$863 ( \1040 , \949 , \951 );
xor \U$864 ( \1041 , \1040 , \954 );
and \U$865 ( \1042 , \1038 , \1041 );
and \U$866 ( \1043 , \1033 , \1041 );
or \U$867 ( \1044 , \1039 , \1042 , \1043 );
xor \U$868 ( \1045 , \831 , \845 );
xor \U$869 ( \1046 , \1045 , \862 );
and \U$870 ( \1047 , \1044 , \1046 );
xor \U$871 ( \1048 , \947 , \957 );
xor \U$872 ( \1049 , \1048 , \960 );
and \U$873 ( \1050 , \1046 , \1049 );
and \U$874 ( \1051 , \1044 , \1049 );
or \U$875 ( \1052 , \1047 , \1050 , \1051 );
xor \U$876 ( \1053 , \963 , \965 );
xor \U$877 ( \1054 , \1053 , \968 );
and \U$878 ( \1055 , \1052 , \1054 );
and \U$879 ( \1056 , \977 , \1055 );
xor \U$880 ( \1057 , \977 , \1055 );
xor \U$881 ( \1058 , \1052 , \1054 );
xor \U$882 ( \1059 , \815 , \979 );
xor \U$883 ( \1060 , \979 , \981 );
not \U$884 ( \1061 , \1060 );
and \U$885 ( \1062 , \1059 , \1061 );
and \U$886 ( \1063 , \159 , \1062 );
not \U$887 ( \1064 , \1063 );
xnor \U$888 ( \1065 , \1064 , \984 );
and \U$889 ( \1066 , \305 , \912 );
and \U$890 ( \1067 , \315 , \910 );
nor \U$891 ( \1068 , \1066 , \1067 );
xnor \U$892 ( \1069 , \1068 , \818 );
and \U$893 ( \1070 , \1065 , \1069 );
and \U$894 ( \1071 , \323 , \740 );
and \U$895 ( \1072 , \333 , \738 );
nor \U$896 ( \1073 , \1071 , \1072 );
xnor \U$897 ( \1074 , \1073 , \668 );
and \U$898 ( \1075 , \1069 , \1074 );
and \U$899 ( \1076 , \1065 , \1074 );
or \U$900 ( \1077 , \1070 , \1075 , \1076 );
and \U$901 ( \1078 , \343 , \604 );
and \U$902 ( \1079 , \353 , \602 );
nor \U$903 ( \1080 , \1078 , \1079 );
xnor \U$904 ( \1081 , \1080 , \561 );
and \U$905 ( \1082 , \444 , \503 );
and \U$906 ( \1083 , \360 , \501 );
nor \U$907 ( \1084 , \1082 , \1083 );
xnor \U$908 ( \1085 , \1084 , \455 );
and \U$909 ( \1086 , \1081 , \1085 );
and \U$910 ( \1087 , \593 , \298 );
and \U$911 ( \1088 , \495 , \296 );
nor \U$912 ( \1089 , \1087 , \1088 );
xnor \U$913 ( \1090 , \1089 , \303 );
and \U$914 ( \1091 , \1085 , \1090 );
and \U$915 ( \1092 , \1081 , \1090 );
or \U$916 ( \1093 , \1086 , \1091 , \1092 );
and \U$917 ( \1094 , \1077 , \1093 );
and \U$918 ( \1095 , \703 , \313 );
and \U$919 ( \1096 , \621 , \311 );
nor \U$920 ( \1097 , \1095 , \1096 );
xnor \U$921 ( \1098 , \1097 , \320 );
and \U$922 ( \1099 , \841 , \331 );
and \U$923 ( \1100 , \777 , \329 );
nor \U$924 ( \1101 , \1099 , \1100 );
xnor \U$925 ( \1102 , \1101 , \338 );
and \U$926 ( \1103 , \1098 , \1102 );
buf \U$927 ( \1104 , RIb4bf2b8_81);
and \U$928 ( \1105 , \1104 , \351 );
and \U$929 ( \1106 , \904 , \349 );
nor \U$930 ( \1107 , \1105 , \1106 );
xnor \U$931 ( \1108 , \1107 , \358 );
and \U$932 ( \1109 , \1102 , \1108 );
and \U$933 ( \1110 , \1098 , \1108 );
or \U$934 ( \1111 , \1103 , \1109 , \1110 );
and \U$935 ( \1112 , \1093 , \1111 );
and \U$936 ( \1113 , \1077 , \1111 );
or \U$937 ( \1114 , \1094 , \1112 , \1113 );
and \U$938 ( \1115 , \1104 , \345 );
xor \U$939 ( \1116 , \1001 , \1005 );
xor \U$940 ( \1117 , \1116 , \1010 );
and \U$941 ( \1118 , \1115 , \1117 );
xor \U$942 ( \1119 , \1018 , \1022 );
xor \U$943 ( \1120 , \1119 , \1027 );
and \U$944 ( \1121 , \1117 , \1120 );
and \U$945 ( \1122 , \1115 , \1120 );
or \U$946 ( \1123 , \1118 , \1121 , \1122 );
and \U$947 ( \1124 , \1114 , \1123 );
xor \U$948 ( \1125 , \915 , \919 );
xor \U$949 ( \1126 , \1125 , \924 );
and \U$950 ( \1127 , \1123 , \1126 );
and \U$951 ( \1128 , \1114 , \1126 );
or \U$952 ( \1129 , \1124 , \1127 , \1128 );
xor \U$953 ( \1130 , \908 , \927 );
xor \U$954 ( \1131 , \1130 , \944 );
and \U$955 ( \1132 , \1129 , \1131 );
xor \U$956 ( \1133 , \1033 , \1038 );
xor \U$957 ( \1134 , \1133 , \1041 );
and \U$958 ( \1135 , \1131 , \1134 );
and \U$959 ( \1136 , \1129 , \1134 );
or \U$960 ( \1137 , \1132 , \1135 , \1136 );
and \U$961 ( \1138 , \353 , \740 );
and \U$962 ( \1139 , \323 , \738 );
nor \U$963 ( \1140 , \1138 , \1139 );
xnor \U$964 ( \1141 , \1140 , \668 );
and \U$965 ( \1142 , \360 , \604 );
and \U$966 ( \1143 , \343 , \602 );
nor \U$967 ( \1144 , \1142 , \1143 );
xnor \U$968 ( \1145 , \1144 , \561 );
and \U$969 ( \1146 , \1141 , \1145 );
and \U$970 ( \1147 , \495 , \503 );
and \U$971 ( \1148 , \444 , \501 );
nor \U$972 ( \1149 , \1147 , \1148 );
xnor \U$973 ( \1150 , \1149 , \455 );
and \U$974 ( \1151 , \1145 , \1150 );
and \U$975 ( \1152 , \1141 , \1150 );
or \U$976 ( \1153 , \1146 , \1151 , \1152 );
and \U$977 ( \1154 , \621 , \298 );
and \U$978 ( \1155 , \593 , \296 );
nor \U$979 ( \1156 , \1154 , \1155 );
xnor \U$980 ( \1157 , \1156 , \303 );
and \U$981 ( \1158 , \777 , \313 );
and \U$982 ( \1159 , \703 , \311 );
nor \U$983 ( \1160 , \1158 , \1159 );
xnor \U$984 ( \1161 , \1160 , \320 );
and \U$985 ( \1162 , \1157 , \1161 );
and \U$986 ( \1163 , \904 , \331 );
and \U$987 ( \1164 , \841 , \329 );
nor \U$988 ( \1165 , \1163 , \1164 );
xnor \U$989 ( \1166 , \1165 , \338 );
and \U$990 ( \1167 , \1161 , \1166 );
and \U$991 ( \1168 , \1157 , \1166 );
or \U$992 ( \1169 , \1162 , \1167 , \1168 );
and \U$993 ( \1170 , \1153 , \1169 );
_DC r130 ( \1171_nR130 , RIb4c3020_52 , \288 );
buf \U$994 ( \1172 , \1171_nR130 );
_DC r12f ( \1173_nR12f , RIb4c2fa8_53 , \288 );
buf \U$995 ( \1174 , \1173_nR12f );
and \U$996 ( \1175 , \1172 , \1174 );
not \U$997 ( \1176 , \1175 );
and \U$998 ( \1177 , \981 , \1176 );
not \U$999 ( \1178 , \1177 );
and \U$1000 ( \1179 , \315 , \1062 );
and \U$1001 ( \1180 , \159 , \1060 );
nor \U$1002 ( \1181 , \1179 , \1180 );
xnor \U$1003 ( \1182 , \1181 , \984 );
and \U$1004 ( \1183 , \1178 , \1182 );
and \U$1005 ( \1184 , \333 , \912 );
and \U$1006 ( \1185 , \305 , \910 );
nor \U$1007 ( \1186 , \1184 , \1185 );
xnor \U$1008 ( \1187 , \1186 , \818 );
and \U$1009 ( \1188 , \1182 , \1187 );
and \U$1010 ( \1189 , \1178 , \1187 );
or \U$1011 ( \1190 , \1183 , \1188 , \1189 );
and \U$1012 ( \1191 , \1169 , \1190 );
and \U$1013 ( \1192 , \1153 , \1190 );
or \U$1014 ( \1193 , \1170 , \1191 , \1192 );
buf \U$1015 ( \1194 , RIb4bf240_82);
and \U$1016 ( \1195 , \1194 , \345 );
xor \U$1017 ( \1196 , \1098 , \1102 );
xor \U$1018 ( \1197 , \1196 , \1108 );
or \U$1019 ( \1198 , \1195 , \1197 );
and \U$1020 ( \1199 , \1193 , \1198 );
xor \U$1021 ( \1200 , \1065 , \1069 );
xor \U$1022 ( \1201 , \1200 , \1074 );
xor \U$1023 ( \1202 , \1081 , \1085 );
xor \U$1024 ( \1203 , \1202 , \1090 );
and \U$1025 ( \1204 , \1201 , \1203 );
and \U$1026 ( \1205 , \1198 , \1204 );
and \U$1027 ( \1206 , \1193 , \1204 );
or \U$1028 ( \1207 , \1199 , \1205 , \1206 );
xor \U$1029 ( \1208 , \985 , \989 );
xor \U$1030 ( \1209 , \1208 , \994 );
xor \U$1031 ( \1210 , \1077 , \1093 );
xor \U$1032 ( \1211 , \1210 , \1111 );
and \U$1033 ( \1212 , \1209 , \1211 );
xor \U$1034 ( \1213 , \1115 , \1117 );
xor \U$1035 ( \1214 , \1213 , \1120 );
and \U$1036 ( \1215 , \1211 , \1214 );
and \U$1037 ( \1216 , \1209 , \1214 );
or \U$1038 ( \1217 , \1212 , \1215 , \1216 );
and \U$1039 ( \1218 , \1207 , \1217 );
xnor \U$1040 ( \1219 , \1035 , \1037 );
and \U$1041 ( \1220 , \1217 , \1219 );
and \U$1042 ( \1221 , \1207 , \1219 );
or \U$1043 ( \1222 , \1218 , \1220 , \1221 );
xor \U$1044 ( \1223 , \997 , \1013 );
xor \U$1045 ( \1224 , \1223 , \1030 );
xor \U$1046 ( \1225 , \1114 , \1123 );
xor \U$1047 ( \1226 , \1225 , \1126 );
and \U$1048 ( \1227 , \1224 , \1226 );
and \U$1049 ( \1228 , \1222 , \1227 );
xor \U$1050 ( \1229 , \1129 , \1131 );
xor \U$1051 ( \1230 , \1229 , \1134 );
and \U$1052 ( \1231 , \1227 , \1230 );
and \U$1053 ( \1232 , \1222 , \1230 );
or \U$1054 ( \1233 , \1228 , \1231 , \1232 );
and \U$1055 ( \1234 , \1137 , \1233 );
xor \U$1056 ( \1235 , \1044 , \1046 );
xor \U$1057 ( \1236 , \1235 , \1049 );
and \U$1058 ( \1237 , \1233 , \1236 );
and \U$1059 ( \1238 , \1137 , \1236 );
or \U$1060 ( \1239 , \1234 , \1237 , \1238 );
and \U$1061 ( \1240 , \1058 , \1239 );
xor \U$1062 ( \1241 , \1058 , \1239 );
xor \U$1063 ( \1242 , \1137 , \1233 );
xor \U$1064 ( \1243 , \1242 , \1236 );
and \U$1065 ( \1244 , \343 , \740 );
and \U$1066 ( \1245 , \353 , \738 );
nor \U$1067 ( \1246 , \1244 , \1245 );
xnor \U$1068 ( \1247 , \1246 , \668 );
and \U$1069 ( \1248 , \444 , \604 );
and \U$1070 ( \1249 , \360 , \602 );
nor \U$1071 ( \1250 , \1248 , \1249 );
xnor \U$1072 ( \1251 , \1250 , \561 );
and \U$1073 ( \1252 , \1247 , \1251 );
and \U$1074 ( \1253 , \593 , \503 );
and \U$1075 ( \1254 , \495 , \501 );
nor \U$1076 ( \1255 , \1253 , \1254 );
xnor \U$1077 ( \1256 , \1255 , \455 );
and \U$1078 ( \1257 , \1251 , \1256 );
and \U$1079 ( \1258 , \1247 , \1256 );
or \U$1080 ( \1259 , \1252 , \1257 , \1258 );
and \U$1081 ( \1260 , \703 , \298 );
and \U$1082 ( \1261 , \621 , \296 );
nor \U$1083 ( \1262 , \1260 , \1261 );
xnor \U$1084 ( \1263 , \1262 , \303 );
and \U$1085 ( \1264 , \841 , \313 );
and \U$1086 ( \1265 , \777 , \311 );
nor \U$1087 ( \1266 , \1264 , \1265 );
xnor \U$1088 ( \1267 , \1266 , \320 );
and \U$1089 ( \1268 , \1263 , \1267 );
and \U$1090 ( \1269 , \1104 , \331 );
and \U$1091 ( \1270 , \904 , \329 );
nor \U$1092 ( \1271 , \1269 , \1270 );
xnor \U$1093 ( \1272 , \1271 , \338 );
and \U$1094 ( \1273 , \1267 , \1272 );
and \U$1095 ( \1274 , \1263 , \1272 );
or \U$1096 ( \1275 , \1268 , \1273 , \1274 );
and \U$1097 ( \1276 , \1259 , \1275 );
xor \U$1098 ( \1277 , \981 , \1172 );
xor \U$1099 ( \1278 , \1172 , \1174 );
not \U$1100 ( \1279 , \1278 );
and \U$1101 ( \1280 , \1277 , \1279 );
and \U$1102 ( \1281 , \159 , \1280 );
not \U$1103 ( \1282 , \1281 );
xnor \U$1104 ( \1283 , \1282 , \1177 );
and \U$1105 ( \1284 , \305 , \1062 );
and \U$1106 ( \1285 , \315 , \1060 );
nor \U$1107 ( \1286 , \1284 , \1285 );
xnor \U$1108 ( \1287 , \1286 , \984 );
and \U$1109 ( \1288 , \1283 , \1287 );
and \U$1110 ( \1289 , \323 , \912 );
and \U$1111 ( \1290 , \333 , \910 );
nor \U$1112 ( \1291 , \1289 , \1290 );
xnor \U$1113 ( \1292 , \1291 , \818 );
and \U$1114 ( \1293 , \1287 , \1292 );
and \U$1115 ( \1294 , \1283 , \1292 );
or \U$1116 ( \1295 , \1288 , \1293 , \1294 );
and \U$1117 ( \1296 , \1275 , \1295 );
and \U$1118 ( \1297 , \1259 , \1295 );
or \U$1119 ( \1298 , \1276 , \1296 , \1297 );
buf \U$1120 ( \1299 , RIb4bf1c8_83);
and \U$1121 ( \1300 , \1299 , \351 );
and \U$1122 ( \1301 , \1194 , \349 );
nor \U$1123 ( \1302 , \1300 , \1301 );
xnor \U$1124 ( \1303 , \1302 , \358 );
buf \U$1125 ( \1304 , RIb4bf150_84);
and \U$1126 ( \1305 , \1304 , \345 );
or \U$1127 ( \1306 , \1303 , \1305 );
and \U$1128 ( \1307 , \1194 , \351 );
and \U$1129 ( \1308 , \1104 , \349 );
nor \U$1130 ( \1309 , \1307 , \1308 );
xnor \U$1131 ( \1310 , \1309 , \358 );
and \U$1132 ( \1311 , \1306 , \1310 );
and \U$1133 ( \1312 , \1299 , \345 );
and \U$1134 ( \1313 , \1310 , \1312 );
and \U$1135 ( \1314 , \1306 , \1312 );
or \U$1136 ( \1315 , \1311 , \1313 , \1314 );
and \U$1137 ( \1316 , \1298 , \1315 );
xor \U$1138 ( \1317 , \1141 , \1145 );
xor \U$1139 ( \1318 , \1317 , \1150 );
xor \U$1140 ( \1319 , \1157 , \1161 );
xor \U$1141 ( \1320 , \1319 , \1166 );
and \U$1142 ( \1321 , \1318 , \1320 );
xor \U$1143 ( \1322 , \1178 , \1182 );
xor \U$1144 ( \1323 , \1322 , \1187 );
and \U$1145 ( \1324 , \1320 , \1323 );
and \U$1146 ( \1325 , \1318 , \1323 );
or \U$1147 ( \1326 , \1321 , \1324 , \1325 );
and \U$1148 ( \1327 , \1315 , \1326 );
and \U$1149 ( \1328 , \1298 , \1326 );
or \U$1150 ( \1329 , \1316 , \1327 , \1328 );
xor \U$1151 ( \1330 , \1153 , \1169 );
xor \U$1152 ( \1331 , \1330 , \1190 );
xnor \U$1153 ( \1332 , \1195 , \1197 );
and \U$1154 ( \1333 , \1331 , \1332 );
xor \U$1155 ( \1334 , \1201 , \1203 );
and \U$1156 ( \1335 , \1332 , \1334 );
and \U$1157 ( \1336 , \1331 , \1334 );
or \U$1158 ( \1337 , \1333 , \1335 , \1336 );
and \U$1159 ( \1338 , \1329 , \1337 );
xor \U$1160 ( \1339 , \1209 , \1211 );
xor \U$1161 ( \1340 , \1339 , \1214 );
and \U$1162 ( \1341 , \1337 , \1340 );
and \U$1163 ( \1342 , \1329 , \1340 );
or \U$1164 ( \1343 , \1338 , \1341 , \1342 );
xor \U$1165 ( \1344 , \1207 , \1217 );
xor \U$1166 ( \1345 , \1344 , \1219 );
and \U$1167 ( \1346 , \1343 , \1345 );
xor \U$1168 ( \1347 , \1224 , \1226 );
and \U$1169 ( \1348 , \1345 , \1347 );
and \U$1170 ( \1349 , \1343 , \1347 );
or \U$1171 ( \1350 , \1346 , \1348 , \1349 );
xor \U$1172 ( \1351 , \1222 , \1227 );
xor \U$1173 ( \1352 , \1351 , \1230 );
and \U$1174 ( \1353 , \1350 , \1352 );
and \U$1175 ( \1354 , \1243 , \1353 );
xor \U$1176 ( \1355 , \1243 , \1353 );
xor \U$1177 ( \1356 , \1350 , \1352 );
_DC r12e ( \1357_nR12e , RIb4c2f30_54 , \288 );
buf \U$1178 ( \1358 , \1357_nR12e );
_DC r12d ( \1359_nR12d , RIb4c2eb8_55 , \288 );
buf \U$1179 ( \1360 , \1359_nR12d );
and \U$1180 ( \1361 , \1358 , \1360 );
not \U$1181 ( \1362 , \1361 );
and \U$1182 ( \1363 , \1174 , \1362 );
not \U$1183 ( \1364 , \1363 );
and \U$1184 ( \1365 , \315 , \1280 );
and \U$1185 ( \1366 , \159 , \1278 );
nor \U$1186 ( \1367 , \1365 , \1366 );
xnor \U$1187 ( \1368 , \1367 , \1177 );
and \U$1188 ( \1369 , \1364 , \1368 );
and \U$1189 ( \1370 , \333 , \1062 );
and \U$1190 ( \1371 , \305 , \1060 );
nor \U$1191 ( \1372 , \1370 , \1371 );
xnor \U$1192 ( \1373 , \1372 , \984 );
and \U$1193 ( \1374 , \1368 , \1373 );
and \U$1194 ( \1375 , \1364 , \1373 );
or \U$1195 ( \1376 , \1369 , \1374 , \1375 );
and \U$1196 ( \1377 , \353 , \912 );
and \U$1197 ( \1378 , \323 , \910 );
nor \U$1198 ( \1379 , \1377 , \1378 );
xnor \U$1199 ( \1380 , \1379 , \818 );
and \U$1200 ( \1381 , \360 , \740 );
and \U$1201 ( \1382 , \343 , \738 );
nor \U$1202 ( \1383 , \1381 , \1382 );
xnor \U$1203 ( \1384 , \1383 , \668 );
and \U$1204 ( \1385 , \1380 , \1384 );
and \U$1205 ( \1386 , \495 , \604 );
and \U$1206 ( \1387 , \444 , \602 );
nor \U$1207 ( \1388 , \1386 , \1387 );
xnor \U$1208 ( \1389 , \1388 , \561 );
and \U$1209 ( \1390 , \1384 , \1389 );
and \U$1210 ( \1391 , \1380 , \1389 );
or \U$1211 ( \1392 , \1385 , \1390 , \1391 );
and \U$1212 ( \1393 , \1376 , \1392 );
and \U$1213 ( \1394 , \621 , \503 );
and \U$1214 ( \1395 , \593 , \501 );
nor \U$1215 ( \1396 , \1394 , \1395 );
xnor \U$1216 ( \1397 , \1396 , \455 );
and \U$1217 ( \1398 , \777 , \298 );
and \U$1218 ( \1399 , \703 , \296 );
nor \U$1219 ( \1400 , \1398 , \1399 );
xnor \U$1220 ( \1401 , \1400 , \303 );
and \U$1221 ( \1402 , \1397 , \1401 );
and \U$1222 ( \1403 , \904 , \313 );
and \U$1223 ( \1404 , \841 , \311 );
nor \U$1224 ( \1405 , \1403 , \1404 );
xnor \U$1225 ( \1406 , \1405 , \320 );
and \U$1226 ( \1407 , \1401 , \1406 );
and \U$1227 ( \1408 , \1397 , \1406 );
or \U$1228 ( \1409 , \1402 , \1407 , \1408 );
and \U$1229 ( \1410 , \1392 , \1409 );
and \U$1230 ( \1411 , \1376 , \1409 );
or \U$1231 ( \1412 , \1393 , \1410 , \1411 );
and \U$1232 ( \1413 , \1194 , \331 );
and \U$1233 ( \1414 , \1104 , \329 );
nor \U$1234 ( \1415 , \1413 , \1414 );
xnor \U$1235 ( \1416 , \1415 , \338 );
and \U$1236 ( \1417 , \1304 , \351 );
and \U$1237 ( \1418 , \1299 , \349 );
nor \U$1238 ( \1419 , \1417 , \1418 );
xnor \U$1239 ( \1420 , \1419 , \358 );
and \U$1240 ( \1421 , \1416 , \1420 );
buf \U$1241 ( \1422 , RIb4bf0d8_85);
and \U$1242 ( \1423 , \1422 , \345 );
and \U$1243 ( \1424 , \1420 , \1423 );
and \U$1244 ( \1425 , \1416 , \1423 );
or \U$1245 ( \1426 , \1421 , \1424 , \1425 );
xor \U$1246 ( \1427 , \1263 , \1267 );
xor \U$1247 ( \1428 , \1427 , \1272 );
and \U$1248 ( \1429 , \1426 , \1428 );
xnor \U$1249 ( \1430 , \1303 , \1305 );
and \U$1250 ( \1431 , \1428 , \1430 );
and \U$1251 ( \1432 , \1426 , \1430 );
or \U$1252 ( \1433 , \1429 , \1431 , \1432 );
and \U$1253 ( \1434 , \1412 , \1433 );
xor \U$1254 ( \1435 , \1247 , \1251 );
xor \U$1255 ( \1436 , \1435 , \1256 );
xor \U$1256 ( \1437 , \1283 , \1287 );
xor \U$1257 ( \1438 , \1437 , \1292 );
and \U$1258 ( \1439 , \1436 , \1438 );
and \U$1259 ( \1440 , \1433 , \1439 );
and \U$1260 ( \1441 , \1412 , \1439 );
or \U$1261 ( \1442 , \1434 , \1440 , \1441 );
xor \U$1262 ( \1443 , \1259 , \1275 );
xor \U$1263 ( \1444 , \1443 , \1295 );
xor \U$1264 ( \1445 , \1306 , \1310 );
xor \U$1265 ( \1446 , \1445 , \1312 );
and \U$1266 ( \1447 , \1444 , \1446 );
xor \U$1267 ( \1448 , \1318 , \1320 );
xor \U$1268 ( \1449 , \1448 , \1323 );
and \U$1269 ( \1450 , \1446 , \1449 );
and \U$1270 ( \1451 , \1444 , \1449 );
or \U$1271 ( \1452 , \1447 , \1450 , \1451 );
and \U$1272 ( \1453 , \1442 , \1452 );
xor \U$1273 ( \1454 , \1331 , \1332 );
xor \U$1274 ( \1455 , \1454 , \1334 );
and \U$1275 ( \1456 , \1452 , \1455 );
and \U$1276 ( \1457 , \1442 , \1455 );
or \U$1277 ( \1458 , \1453 , \1456 , \1457 );
xor \U$1278 ( \1459 , \1193 , \1198 );
xor \U$1279 ( \1460 , \1459 , \1204 );
and \U$1280 ( \1461 , \1458 , \1460 );
xor \U$1281 ( \1462 , \1329 , \1337 );
xor \U$1282 ( \1463 , \1462 , \1340 );
and \U$1283 ( \1464 , \1460 , \1463 );
and \U$1284 ( \1465 , \1458 , \1463 );
or \U$1285 ( \1466 , \1461 , \1464 , \1465 );
xor \U$1286 ( \1467 , \1343 , \1345 );
xor \U$1287 ( \1468 , \1467 , \1347 );
and \U$1288 ( \1469 , \1466 , \1468 );
and \U$1289 ( \1470 , \1356 , \1469 );
xor \U$1290 ( \1471 , \1356 , \1469 );
xor \U$1291 ( \1472 , \1466 , \1468 );
xor \U$1292 ( \1473 , \1174 , \1358 );
xor \U$1293 ( \1474 , \1358 , \1360 );
not \U$1294 ( \1475 , \1474 );
and \U$1295 ( \1476 , \1473 , \1475 );
and \U$1296 ( \1477 , \159 , \1476 );
not \U$1297 ( \1478 , \1477 );
xnor \U$1298 ( \1479 , \1478 , \1363 );
and \U$1299 ( \1480 , \305 , \1280 );
and \U$1300 ( \1481 , \315 , \1278 );
nor \U$1301 ( \1482 , \1480 , \1481 );
xnor \U$1302 ( \1483 , \1482 , \1177 );
and \U$1303 ( \1484 , \1479 , \1483 );
and \U$1304 ( \1485 , \323 , \1062 );
and \U$1305 ( \1486 , \333 , \1060 );
nor \U$1306 ( \1487 , \1485 , \1486 );
xnor \U$1307 ( \1488 , \1487 , \984 );
and \U$1308 ( \1489 , \1483 , \1488 );
and \U$1309 ( \1490 , \1479 , \1488 );
or \U$1310 ( \1491 , \1484 , \1489 , \1490 );
and \U$1311 ( \1492 , \343 , \912 );
and \U$1312 ( \1493 , \353 , \910 );
nor \U$1313 ( \1494 , \1492 , \1493 );
xnor \U$1314 ( \1495 , \1494 , \818 );
and \U$1315 ( \1496 , \444 , \740 );
and \U$1316 ( \1497 , \360 , \738 );
nor \U$1317 ( \1498 , \1496 , \1497 );
xnor \U$1318 ( \1499 , \1498 , \668 );
and \U$1319 ( \1500 , \1495 , \1499 );
and \U$1320 ( \1501 , \593 , \604 );
and \U$1321 ( \1502 , \495 , \602 );
nor \U$1322 ( \1503 , \1501 , \1502 );
xnor \U$1323 ( \1504 , \1503 , \561 );
and \U$1324 ( \1505 , \1499 , \1504 );
and \U$1325 ( \1506 , \1495 , \1504 );
or \U$1326 ( \1507 , \1500 , \1505 , \1506 );
and \U$1327 ( \1508 , \1491 , \1507 );
and \U$1328 ( \1509 , \703 , \503 );
and \U$1329 ( \1510 , \621 , \501 );
nor \U$1330 ( \1511 , \1509 , \1510 );
xnor \U$1331 ( \1512 , \1511 , \455 );
and \U$1332 ( \1513 , \841 , \298 );
and \U$1333 ( \1514 , \777 , \296 );
nor \U$1334 ( \1515 , \1513 , \1514 );
xnor \U$1335 ( \1516 , \1515 , \303 );
and \U$1336 ( \1517 , \1512 , \1516 );
and \U$1337 ( \1518 , \1104 , \313 );
and \U$1338 ( \1519 , \904 , \311 );
nor \U$1339 ( \1520 , \1518 , \1519 );
xnor \U$1340 ( \1521 , \1520 , \320 );
and \U$1341 ( \1522 , \1516 , \1521 );
and \U$1342 ( \1523 , \1512 , \1521 );
or \U$1343 ( \1524 , \1517 , \1522 , \1523 );
and \U$1344 ( \1525 , \1507 , \1524 );
and \U$1345 ( \1526 , \1491 , \1524 );
or \U$1346 ( \1527 , \1508 , \1525 , \1526 );
and \U$1347 ( \1528 , \1299 , \331 );
and \U$1348 ( \1529 , \1194 , \329 );
nor \U$1349 ( \1530 , \1528 , \1529 );
xnor \U$1350 ( \1531 , \1530 , \338 );
and \U$1351 ( \1532 , \1422 , \351 );
and \U$1352 ( \1533 , \1304 , \349 );
nor \U$1353 ( \1534 , \1532 , \1533 );
xnor \U$1354 ( \1535 , \1534 , \358 );
and \U$1355 ( \1536 , \1531 , \1535 );
buf \U$1356 ( \1537 , RIb4bf060_86);
and \U$1357 ( \1538 , \1537 , \345 );
and \U$1358 ( \1539 , \1535 , \1538 );
and \U$1359 ( \1540 , \1531 , \1538 );
or \U$1360 ( \1541 , \1536 , \1539 , \1540 );
xor \U$1361 ( \1542 , \1416 , \1420 );
xor \U$1362 ( \1543 , \1542 , \1423 );
and \U$1363 ( \1544 , \1541 , \1543 );
xor \U$1364 ( \1545 , \1397 , \1401 );
xor \U$1365 ( \1546 , \1545 , \1406 );
and \U$1366 ( \1547 , \1543 , \1546 );
and \U$1367 ( \1548 , \1541 , \1546 );
or \U$1368 ( \1549 , \1544 , \1547 , \1548 );
and \U$1369 ( \1550 , \1527 , \1549 );
xor \U$1370 ( \1551 , \1364 , \1368 );
xor \U$1371 ( \1552 , \1551 , \1373 );
xor \U$1372 ( \1553 , \1380 , \1384 );
xor \U$1373 ( \1554 , \1553 , \1389 );
and \U$1374 ( \1555 , \1552 , \1554 );
and \U$1375 ( \1556 , \1549 , \1555 );
and \U$1376 ( \1557 , \1527 , \1555 );
or \U$1377 ( \1558 , \1550 , \1556 , \1557 );
xor \U$1378 ( \1559 , \1376 , \1392 );
xor \U$1379 ( \1560 , \1559 , \1409 );
xor \U$1380 ( \1561 , \1426 , \1428 );
xor \U$1381 ( \1562 , \1561 , \1430 );
and \U$1382 ( \1563 , \1560 , \1562 );
xor \U$1383 ( \1564 , \1436 , \1438 );
and \U$1384 ( \1565 , \1562 , \1564 );
and \U$1385 ( \1566 , \1560 , \1564 );
or \U$1386 ( \1567 , \1563 , \1565 , \1566 );
and \U$1387 ( \1568 , \1558 , \1567 );
xor \U$1388 ( \1569 , \1444 , \1446 );
xor \U$1389 ( \1570 , \1569 , \1449 );
and \U$1390 ( \1571 , \1567 , \1570 );
and \U$1391 ( \1572 , \1558 , \1570 );
or \U$1392 ( \1573 , \1568 , \1571 , \1572 );
xor \U$1393 ( \1574 , \1298 , \1315 );
xor \U$1394 ( \1575 , \1574 , \1326 );
and \U$1395 ( \1576 , \1573 , \1575 );
xor \U$1396 ( \1577 , \1442 , \1452 );
xor \U$1397 ( \1578 , \1577 , \1455 );
and \U$1398 ( \1579 , \1575 , \1578 );
and \U$1399 ( \1580 , \1573 , \1578 );
or \U$1400 ( \1581 , \1576 , \1579 , \1580 );
xor \U$1401 ( \1582 , \1458 , \1460 );
xor \U$1402 ( \1583 , \1582 , \1463 );
and \U$1403 ( \1584 , \1581 , \1583 );
and \U$1404 ( \1585 , \1472 , \1584 );
xor \U$1405 ( \1586 , \1472 , \1584 );
xor \U$1406 ( \1587 , \1581 , \1583 );
and \U$1407 ( \1588 , \621 , \604 );
and \U$1408 ( \1589 , \593 , \602 );
nor \U$1409 ( \1590 , \1588 , \1589 );
xnor \U$1410 ( \1591 , \1590 , \561 );
and \U$1411 ( \1592 , \777 , \503 );
and \U$1412 ( \1593 , \703 , \501 );
nor \U$1413 ( \1594 , \1592 , \1593 );
xnor \U$1414 ( \1595 , \1594 , \455 );
and \U$1415 ( \1596 , \1591 , \1595 );
and \U$1416 ( \1597 , \904 , \298 );
and \U$1417 ( \1598 , \841 , \296 );
nor \U$1418 ( \1599 , \1597 , \1598 );
xnor \U$1419 ( \1600 , \1599 , \303 );
and \U$1420 ( \1601 , \1595 , \1600 );
and \U$1421 ( \1602 , \1591 , \1600 );
or \U$1422 ( \1603 , \1596 , \1601 , \1602 );
_DC r12c ( \1604_nR12c , RIb4c2e40_56 , \288 );
buf \U$1423 ( \1605 , \1604_nR12c );
_DC r12b ( \1606_nR12b , RIb4c2dc8_57 , \288 );
buf \U$1424 ( \1607 , \1606_nR12b );
and \U$1425 ( \1608 , \1605 , \1607 );
not \U$1426 ( \1609 , \1608 );
and \U$1427 ( \1610 , \1360 , \1609 );
not \U$1428 ( \1611 , \1610 );
and \U$1429 ( \1612 , \315 , \1476 );
and \U$1430 ( \1613 , \159 , \1474 );
nor \U$1431 ( \1614 , \1612 , \1613 );
xnor \U$1432 ( \1615 , \1614 , \1363 );
and \U$1433 ( \1616 , \1611 , \1615 );
and \U$1434 ( \1617 , \333 , \1280 );
and \U$1435 ( \1618 , \305 , \1278 );
nor \U$1436 ( \1619 , \1617 , \1618 );
xnor \U$1437 ( \1620 , \1619 , \1177 );
and \U$1438 ( \1621 , \1615 , \1620 );
and \U$1439 ( \1622 , \1611 , \1620 );
or \U$1440 ( \1623 , \1616 , \1621 , \1622 );
and \U$1441 ( \1624 , \1603 , \1623 );
and \U$1442 ( \1625 , \353 , \1062 );
and \U$1443 ( \1626 , \323 , \1060 );
nor \U$1444 ( \1627 , \1625 , \1626 );
xnor \U$1445 ( \1628 , \1627 , \984 );
and \U$1446 ( \1629 , \360 , \912 );
and \U$1447 ( \1630 , \343 , \910 );
nor \U$1448 ( \1631 , \1629 , \1630 );
xnor \U$1449 ( \1632 , \1631 , \818 );
and \U$1450 ( \1633 , \1628 , \1632 );
and \U$1451 ( \1634 , \495 , \740 );
and \U$1452 ( \1635 , \444 , \738 );
nor \U$1453 ( \1636 , \1634 , \1635 );
xnor \U$1454 ( \1637 , \1636 , \668 );
and \U$1455 ( \1638 , \1632 , \1637 );
and \U$1456 ( \1639 , \1628 , \1637 );
or \U$1457 ( \1640 , \1633 , \1638 , \1639 );
and \U$1458 ( \1641 , \1623 , \1640 );
and \U$1459 ( \1642 , \1603 , \1640 );
or \U$1460 ( \1643 , \1624 , \1641 , \1642 );
xor \U$1461 ( \1644 , \1479 , \1483 );
xor \U$1462 ( \1645 , \1644 , \1488 );
xor \U$1463 ( \1646 , \1495 , \1499 );
xor \U$1464 ( \1647 , \1646 , \1504 );
and \U$1465 ( \1648 , \1645 , \1647 );
xor \U$1466 ( \1649 , \1512 , \1516 );
xor \U$1467 ( \1650 , \1649 , \1521 );
and \U$1468 ( \1651 , \1647 , \1650 );
and \U$1469 ( \1652 , \1645 , \1650 );
or \U$1470 ( \1653 , \1648 , \1651 , \1652 );
and \U$1471 ( \1654 , \1643 , \1653 );
and \U$1472 ( \1655 , \1194 , \313 );
and \U$1473 ( \1656 , \1104 , \311 );
nor \U$1474 ( \1657 , \1655 , \1656 );
xnor \U$1475 ( \1658 , \1657 , \320 );
and \U$1476 ( \1659 , \1304 , \331 );
and \U$1477 ( \1660 , \1299 , \329 );
nor \U$1478 ( \1661 , \1659 , \1660 );
xnor \U$1479 ( \1662 , \1661 , \338 );
and \U$1480 ( \1663 , \1658 , \1662 );
and \U$1481 ( \1664 , \1537 , \351 );
and \U$1482 ( \1665 , \1422 , \349 );
nor \U$1483 ( \1666 , \1664 , \1665 );
xnor \U$1484 ( \1667 , \1666 , \358 );
and \U$1485 ( \1668 , \1662 , \1667 );
and \U$1486 ( \1669 , \1658 , \1667 );
or \U$1487 ( \1670 , \1663 , \1668 , \1669 );
xor \U$1488 ( \1671 , \1531 , \1535 );
xor \U$1489 ( \1672 , \1671 , \1538 );
or \U$1490 ( \1673 , \1670 , \1672 );
and \U$1491 ( \1674 , \1653 , \1673 );
and \U$1492 ( \1675 , \1643 , \1673 );
or \U$1493 ( \1676 , \1654 , \1674 , \1675 );
xor \U$1494 ( \1677 , \1491 , \1507 );
xor \U$1495 ( \1678 , \1677 , \1524 );
xor \U$1496 ( \1679 , \1541 , \1543 );
xor \U$1497 ( \1680 , \1679 , \1546 );
and \U$1498 ( \1681 , \1678 , \1680 );
xor \U$1499 ( \1682 , \1552 , \1554 );
and \U$1500 ( \1683 , \1680 , \1682 );
and \U$1501 ( \1684 , \1678 , \1682 );
or \U$1502 ( \1685 , \1681 , \1683 , \1684 );
and \U$1503 ( \1686 , \1676 , \1685 );
xor \U$1504 ( \1687 , \1560 , \1562 );
xor \U$1505 ( \1688 , \1687 , \1564 );
and \U$1506 ( \1689 , \1685 , \1688 );
and \U$1507 ( \1690 , \1676 , \1688 );
or \U$1508 ( \1691 , \1686 , \1689 , \1690 );
xor \U$1509 ( \1692 , \1412 , \1433 );
xor \U$1510 ( \1693 , \1692 , \1439 );
and \U$1511 ( \1694 , \1691 , \1693 );
xor \U$1512 ( \1695 , \1558 , \1567 );
xor \U$1513 ( \1696 , \1695 , \1570 );
and \U$1514 ( \1697 , \1693 , \1696 );
and \U$1515 ( \1698 , \1691 , \1696 );
or \U$1516 ( \1699 , \1694 , \1697 , \1698 );
xor \U$1517 ( \1700 , \1573 , \1575 );
xor \U$1518 ( \1701 , \1700 , \1578 );
and \U$1519 ( \1702 , \1699 , \1701 );
and \U$1520 ( \1703 , \1587 , \1702 );
xor \U$1521 ( \1704 , \1587 , \1702 );
xor \U$1522 ( \1705 , \1699 , \1701 );
and \U$1523 ( \1706 , \703 , \604 );
and \U$1524 ( \1707 , \621 , \602 );
nor \U$1525 ( \1708 , \1706 , \1707 );
xnor \U$1526 ( \1709 , \1708 , \561 );
and \U$1527 ( \1710 , \841 , \503 );
and \U$1528 ( \1711 , \777 , \501 );
nor \U$1529 ( \1712 , \1710 , \1711 );
xnor \U$1530 ( \1713 , \1712 , \455 );
and \U$1531 ( \1714 , \1709 , \1713 );
and \U$1532 ( \1715 , \1104 , \298 );
and \U$1533 ( \1716 , \904 , \296 );
nor \U$1534 ( \1717 , \1715 , \1716 );
xnor \U$1535 ( \1718 , \1717 , \303 );
and \U$1536 ( \1719 , \1713 , \1718 );
and \U$1537 ( \1720 , \1709 , \1718 );
or \U$1538 ( \1721 , \1714 , \1719 , \1720 );
and \U$1539 ( \1722 , \343 , \1062 );
and \U$1540 ( \1723 , \353 , \1060 );
nor \U$1541 ( \1724 , \1722 , \1723 );
xnor \U$1542 ( \1725 , \1724 , \984 );
and \U$1543 ( \1726 , \444 , \912 );
and \U$1544 ( \1727 , \360 , \910 );
nor \U$1545 ( \1728 , \1726 , \1727 );
xnor \U$1546 ( \1729 , \1728 , \818 );
and \U$1547 ( \1730 , \1725 , \1729 );
and \U$1548 ( \1731 , \593 , \740 );
and \U$1549 ( \1732 , \495 , \738 );
nor \U$1550 ( \1733 , \1731 , \1732 );
xnor \U$1551 ( \1734 , \1733 , \668 );
and \U$1552 ( \1735 , \1729 , \1734 );
and \U$1553 ( \1736 , \1725 , \1734 );
or \U$1554 ( \1737 , \1730 , \1735 , \1736 );
and \U$1555 ( \1738 , \1721 , \1737 );
xor \U$1556 ( \1739 , \1360 , \1605 );
xor \U$1557 ( \1740 , \1605 , \1607 );
not \U$1558 ( \1741 , \1740 );
and \U$1559 ( \1742 , \1739 , \1741 );
and \U$1560 ( \1743 , \159 , \1742 );
not \U$1561 ( \1744 , \1743 );
xnor \U$1562 ( \1745 , \1744 , \1610 );
and \U$1563 ( \1746 , \305 , \1476 );
and \U$1564 ( \1747 , \315 , \1474 );
nor \U$1565 ( \1748 , \1746 , \1747 );
xnor \U$1566 ( \1749 , \1748 , \1363 );
and \U$1567 ( \1750 , \1745 , \1749 );
and \U$1568 ( \1751 , \323 , \1280 );
and \U$1569 ( \1752 , \333 , \1278 );
nor \U$1570 ( \1753 , \1751 , \1752 );
xnor \U$1571 ( \1754 , \1753 , \1177 );
and \U$1572 ( \1755 , \1749 , \1754 );
and \U$1573 ( \1756 , \1745 , \1754 );
or \U$1574 ( \1757 , \1750 , \1755 , \1756 );
and \U$1575 ( \1758 , \1737 , \1757 );
and \U$1576 ( \1759 , \1721 , \1757 );
or \U$1577 ( \1760 , \1738 , \1758 , \1759 );
and \U$1578 ( \1761 , \1299 , \313 );
and \U$1579 ( \1762 , \1194 , \311 );
nor \U$1580 ( \1763 , \1761 , \1762 );
xnor \U$1581 ( \1764 , \1763 , \320 );
and \U$1582 ( \1765 , \1422 , \331 );
and \U$1583 ( \1766 , \1304 , \329 );
nor \U$1584 ( \1767 , \1765 , \1766 );
xnor \U$1585 ( \1768 , \1767 , \338 );
and \U$1586 ( \1769 , \1764 , \1768 );
buf \U$1587 ( \1770 , RIb4befe8_87);
and \U$1588 ( \1771 , \1770 , \351 );
and \U$1589 ( \1772 , \1537 , \349 );
nor \U$1590 ( \1773 , \1771 , \1772 );
xnor \U$1591 ( \1774 , \1773 , \358 );
and \U$1592 ( \1775 , \1768 , \1774 );
and \U$1593 ( \1776 , \1764 , \1774 );
or \U$1594 ( \1777 , \1769 , \1775 , \1776 );
buf \U$1595 ( \1778 , RIb4bef70_88);
and \U$1596 ( \1779 , \1778 , \345 );
buf \U$1597 ( \1780 , \1779 );
and \U$1598 ( \1781 , \1777 , \1780 );
and \U$1599 ( \1782 , \1770 , \345 );
and \U$1600 ( \1783 , \1780 , \1782 );
and \U$1601 ( \1784 , \1777 , \1782 );
or \U$1602 ( \1785 , \1781 , \1783 , \1784 );
and \U$1603 ( \1786 , \1760 , \1785 );
xor \U$1604 ( \1787 , \1658 , \1662 );
xor \U$1605 ( \1788 , \1787 , \1667 );
xor \U$1606 ( \1789 , \1591 , \1595 );
xor \U$1607 ( \1790 , \1789 , \1600 );
and \U$1608 ( \1791 , \1788 , \1790 );
xor \U$1609 ( \1792 , \1628 , \1632 );
xor \U$1610 ( \1793 , \1792 , \1637 );
and \U$1611 ( \1794 , \1790 , \1793 );
and \U$1612 ( \1795 , \1788 , \1793 );
or \U$1613 ( \1796 , \1791 , \1794 , \1795 );
and \U$1614 ( \1797 , \1785 , \1796 );
and \U$1615 ( \1798 , \1760 , \1796 );
or \U$1616 ( \1799 , \1786 , \1797 , \1798 );
xor \U$1617 ( \1800 , \1603 , \1623 );
xor \U$1618 ( \1801 , \1800 , \1640 );
xor \U$1619 ( \1802 , \1645 , \1647 );
xor \U$1620 ( \1803 , \1802 , \1650 );
and \U$1621 ( \1804 , \1801 , \1803 );
xnor \U$1622 ( \1805 , \1670 , \1672 );
and \U$1623 ( \1806 , \1803 , \1805 );
and \U$1624 ( \1807 , \1801 , \1805 );
or \U$1625 ( \1808 , \1804 , \1806 , \1807 );
and \U$1626 ( \1809 , \1799 , \1808 );
xor \U$1627 ( \1810 , \1678 , \1680 );
xor \U$1628 ( \1811 , \1810 , \1682 );
and \U$1629 ( \1812 , \1808 , \1811 );
and \U$1630 ( \1813 , \1799 , \1811 );
or \U$1631 ( \1814 , \1809 , \1812 , \1813 );
xor \U$1632 ( \1815 , \1527 , \1549 );
xor \U$1633 ( \1816 , \1815 , \1555 );
and \U$1634 ( \1817 , \1814 , \1816 );
xor \U$1635 ( \1818 , \1676 , \1685 );
xor \U$1636 ( \1819 , \1818 , \1688 );
and \U$1637 ( \1820 , \1816 , \1819 );
and \U$1638 ( \1821 , \1814 , \1819 );
or \U$1639 ( \1822 , \1817 , \1820 , \1821 );
xor \U$1640 ( \1823 , \1691 , \1693 );
xor \U$1641 ( \1824 , \1823 , \1696 );
and \U$1642 ( \1825 , \1822 , \1824 );
and \U$1643 ( \1826 , \1705 , \1825 );
xor \U$1644 ( \1827 , \1705 , \1825 );
xor \U$1645 ( \1828 , \1822 , \1824 );
_DC r12a ( \1829_nR12a , RIb4c2d50_58 , \288 );
buf \U$1646 ( \1830 , \1829_nR12a );
_DC r129 ( \1831_nR129 , RIb4c2cd8_59 , \288 );
buf \U$1647 ( \1832 , \1831_nR129 );
and \U$1648 ( \1833 , \1830 , \1832 );
not \U$1649 ( \1834 , \1833 );
and \U$1650 ( \1835 , \1607 , \1834 );
not \U$1651 ( \1836 , \1835 );
and \U$1652 ( \1837 , \315 , \1742 );
and \U$1653 ( \1838 , \159 , \1740 );
nor \U$1654 ( \1839 , \1837 , \1838 );
xnor \U$1655 ( \1840 , \1839 , \1610 );
and \U$1656 ( \1841 , \1836 , \1840 );
and \U$1657 ( \1842 , \333 , \1476 );
and \U$1658 ( \1843 , \305 , \1474 );
nor \U$1659 ( \1844 , \1842 , \1843 );
xnor \U$1660 ( \1845 , \1844 , \1363 );
and \U$1661 ( \1846 , \1840 , \1845 );
and \U$1662 ( \1847 , \1836 , \1845 );
or \U$1663 ( \1848 , \1841 , \1846 , \1847 );
and \U$1664 ( \1849 , \353 , \1280 );
and \U$1665 ( \1850 , \323 , \1278 );
nor \U$1666 ( \1851 , \1849 , \1850 );
xnor \U$1667 ( \1852 , \1851 , \1177 );
and \U$1668 ( \1853 , \360 , \1062 );
and \U$1669 ( \1854 , \343 , \1060 );
nor \U$1670 ( \1855 , \1853 , \1854 );
xnor \U$1671 ( \1856 , \1855 , \984 );
and \U$1672 ( \1857 , \1852 , \1856 );
and \U$1673 ( \1858 , \495 , \912 );
and \U$1674 ( \1859 , \444 , \910 );
nor \U$1675 ( \1860 , \1858 , \1859 );
xnor \U$1676 ( \1861 , \1860 , \818 );
and \U$1677 ( \1862 , \1856 , \1861 );
and \U$1678 ( \1863 , \1852 , \1861 );
or \U$1679 ( \1864 , \1857 , \1862 , \1863 );
and \U$1680 ( \1865 , \1848 , \1864 );
and \U$1681 ( \1866 , \621 , \740 );
and \U$1682 ( \1867 , \593 , \738 );
nor \U$1683 ( \1868 , \1866 , \1867 );
xnor \U$1684 ( \1869 , \1868 , \668 );
and \U$1685 ( \1870 , \777 , \604 );
and \U$1686 ( \1871 , \703 , \602 );
nor \U$1687 ( \1872 , \1870 , \1871 );
xnor \U$1688 ( \1873 , \1872 , \561 );
and \U$1689 ( \1874 , \1869 , \1873 );
and \U$1690 ( \1875 , \904 , \503 );
and \U$1691 ( \1876 , \841 , \501 );
nor \U$1692 ( \1877 , \1875 , \1876 );
xnor \U$1693 ( \1878 , \1877 , \455 );
and \U$1694 ( \1879 , \1873 , \1878 );
and \U$1695 ( \1880 , \1869 , \1878 );
or \U$1696 ( \1881 , \1874 , \1879 , \1880 );
and \U$1697 ( \1882 , \1864 , \1881 );
and \U$1698 ( \1883 , \1848 , \1881 );
or \U$1699 ( \1884 , \1865 , \1882 , \1883 );
xor \U$1700 ( \1885 , \1709 , \1713 );
xor \U$1701 ( \1886 , \1885 , \1718 );
xor \U$1702 ( \1887 , \1725 , \1729 );
xor \U$1703 ( \1888 , \1887 , \1734 );
and \U$1704 ( \1889 , \1886 , \1888 );
xor \U$1705 ( \1890 , \1745 , \1749 );
xor \U$1706 ( \1891 , \1890 , \1754 );
and \U$1707 ( \1892 , \1888 , \1891 );
and \U$1708 ( \1893 , \1886 , \1891 );
or \U$1709 ( \1894 , \1889 , \1892 , \1893 );
and \U$1710 ( \1895 , \1884 , \1894 );
and \U$1711 ( \1896 , \1194 , \298 );
and \U$1712 ( \1897 , \1104 , \296 );
nor \U$1713 ( \1898 , \1896 , \1897 );
xnor \U$1714 ( \1899 , \1898 , \303 );
and \U$1715 ( \1900 , \1304 , \313 );
and \U$1716 ( \1901 , \1299 , \311 );
nor \U$1717 ( \1902 , \1900 , \1901 );
xnor \U$1718 ( \1903 , \1902 , \320 );
and \U$1719 ( \1904 , \1899 , \1903 );
and \U$1720 ( \1905 , \1537 , \331 );
and \U$1721 ( \1906 , \1422 , \329 );
nor \U$1722 ( \1907 , \1905 , \1906 );
xnor \U$1723 ( \1908 , \1907 , \338 );
and \U$1724 ( \1909 , \1903 , \1908 );
and \U$1725 ( \1910 , \1899 , \1908 );
or \U$1726 ( \1911 , \1904 , \1909 , \1910 );
xor \U$1727 ( \1912 , \1764 , \1768 );
xor \U$1728 ( \1913 , \1912 , \1774 );
and \U$1729 ( \1914 , \1911 , \1913 );
not \U$1730 ( \1915 , \1779 );
and \U$1731 ( \1916 , \1913 , \1915 );
and \U$1732 ( \1917 , \1911 , \1915 );
or \U$1733 ( \1918 , \1914 , \1916 , \1917 );
and \U$1734 ( \1919 , \1894 , \1918 );
and \U$1735 ( \1920 , \1884 , \1918 );
or \U$1736 ( \1921 , \1895 , \1919 , \1920 );
xor \U$1737 ( \1922 , \1611 , \1615 );
xor \U$1738 ( \1923 , \1922 , \1620 );
xor \U$1739 ( \1924 , \1777 , \1780 );
xor \U$1740 ( \1925 , \1924 , \1782 );
and \U$1741 ( \1926 , \1923 , \1925 );
xor \U$1742 ( \1927 , \1788 , \1790 );
xor \U$1743 ( \1928 , \1927 , \1793 );
and \U$1744 ( \1929 , \1925 , \1928 );
and \U$1745 ( \1930 , \1923 , \1928 );
or \U$1746 ( \1931 , \1926 , \1929 , \1930 );
and \U$1747 ( \1932 , \1921 , \1931 );
xor \U$1748 ( \1933 , \1801 , \1803 );
xor \U$1749 ( \1934 , \1933 , \1805 );
and \U$1750 ( \1935 , \1931 , \1934 );
and \U$1751 ( \1936 , \1921 , \1934 );
or \U$1752 ( \1937 , \1932 , \1935 , \1936 );
xor \U$1753 ( \1938 , \1643 , \1653 );
xor \U$1754 ( \1939 , \1938 , \1673 );
and \U$1755 ( \1940 , \1937 , \1939 );
xor \U$1756 ( \1941 , \1799 , \1808 );
xor \U$1757 ( \1942 , \1941 , \1811 );
and \U$1758 ( \1943 , \1939 , \1942 );
and \U$1759 ( \1944 , \1937 , \1942 );
or \U$1760 ( \1945 , \1940 , \1943 , \1944 );
xor \U$1761 ( \1946 , \1814 , \1816 );
xor \U$1762 ( \1947 , \1946 , \1819 );
and \U$1763 ( \1948 , \1945 , \1947 );
and \U$1764 ( \1949 , \1828 , \1948 );
xor \U$1765 ( \1950 , \1828 , \1948 );
xor \U$1766 ( \1951 , \1945 , \1947 );
xor \U$1767 ( \1952 , \1607 , \1830 );
xor \U$1768 ( \1953 , \1830 , \1832 );
not \U$1769 ( \1954 , \1953 );
and \U$1770 ( \1955 , \1952 , \1954 );
and \U$1771 ( \1956 , \159 , \1955 );
not \U$1772 ( \1957 , \1956 );
xnor \U$1773 ( \1958 , \1957 , \1835 );
and \U$1774 ( \1959 , \305 , \1742 );
and \U$1775 ( \1960 , \315 , \1740 );
nor \U$1776 ( \1961 , \1959 , \1960 );
xnor \U$1777 ( \1962 , \1961 , \1610 );
and \U$1778 ( \1963 , \1958 , \1962 );
and \U$1779 ( \1964 , \323 , \1476 );
and \U$1780 ( \1965 , \333 , \1474 );
nor \U$1781 ( \1966 , \1964 , \1965 );
xnor \U$1782 ( \1967 , \1966 , \1363 );
and \U$1783 ( \1968 , \1962 , \1967 );
and \U$1784 ( \1969 , \1958 , \1967 );
or \U$1785 ( \1970 , \1963 , \1968 , \1969 );
and \U$1786 ( \1971 , \343 , \1280 );
and \U$1787 ( \1972 , \353 , \1278 );
nor \U$1788 ( \1973 , \1971 , \1972 );
xnor \U$1789 ( \1974 , \1973 , \1177 );
and \U$1790 ( \1975 , \444 , \1062 );
and \U$1791 ( \1976 , \360 , \1060 );
nor \U$1792 ( \1977 , \1975 , \1976 );
xnor \U$1793 ( \1978 , \1977 , \984 );
and \U$1794 ( \1979 , \1974 , \1978 );
and \U$1795 ( \1980 , \593 , \912 );
and \U$1796 ( \1981 , \495 , \910 );
nor \U$1797 ( \1982 , \1980 , \1981 );
xnor \U$1798 ( \1983 , \1982 , \818 );
and \U$1799 ( \1984 , \1978 , \1983 );
and \U$1800 ( \1985 , \1974 , \1983 );
or \U$1801 ( \1986 , \1979 , \1984 , \1985 );
and \U$1802 ( \1987 , \1970 , \1986 );
and \U$1803 ( \1988 , \703 , \740 );
and \U$1804 ( \1989 , \621 , \738 );
nor \U$1805 ( \1990 , \1988 , \1989 );
xnor \U$1806 ( \1991 , \1990 , \668 );
and \U$1807 ( \1992 , \841 , \604 );
and \U$1808 ( \1993 , \777 , \602 );
nor \U$1809 ( \1994 , \1992 , \1993 );
xnor \U$1810 ( \1995 , \1994 , \561 );
and \U$1811 ( \1996 , \1991 , \1995 );
and \U$1812 ( \1997 , \1104 , \503 );
and \U$1813 ( \1998 , \904 , \501 );
nor \U$1814 ( \1999 , \1997 , \1998 );
xnor \U$1815 ( \2000 , \1999 , \455 );
and \U$1816 ( \2001 , \1995 , \2000 );
and \U$1817 ( \2002 , \1991 , \2000 );
or \U$1818 ( \2003 , \1996 , \2001 , \2002 );
and \U$1819 ( \2004 , \1986 , \2003 );
and \U$1820 ( \2005 , \1970 , \2003 );
or \U$1821 ( \2006 , \1987 , \2004 , \2005 );
and \U$1822 ( \2007 , \1299 , \298 );
and \U$1823 ( \2008 , \1194 , \296 );
nor \U$1824 ( \2009 , \2007 , \2008 );
xnor \U$1825 ( \2010 , \2009 , \303 );
and \U$1826 ( \2011 , \1422 , \313 );
and \U$1827 ( \2012 , \1304 , \311 );
nor \U$1828 ( \2013 , \2011 , \2012 );
xnor \U$1829 ( \2014 , \2013 , \320 );
and \U$1830 ( \2015 , \2010 , \2014 );
and \U$1831 ( \2016 , \1770 , \331 );
and \U$1832 ( \2017 , \1537 , \329 );
nor \U$1833 ( \2018 , \2016 , \2017 );
xnor \U$1834 ( \2019 , \2018 , \338 );
and \U$1835 ( \2020 , \2014 , \2019 );
and \U$1836 ( \2021 , \2010 , \2019 );
or \U$1837 ( \2022 , \2015 , \2020 , \2021 );
buf \U$1838 ( \2023 , RIb4beef8_89);
and \U$1839 ( \2024 , \2023 , \351 );
and \U$1840 ( \2025 , \1778 , \349 );
nor \U$1841 ( \2026 , \2024 , \2025 );
xnor \U$1842 ( \2027 , \2026 , \358 );
buf \U$1843 ( \2028 , RIb4bee80_90);
and \U$1844 ( \2029 , \2028 , \345 );
or \U$1845 ( \2030 , \2027 , \2029 );
and \U$1846 ( \2031 , \2022 , \2030 );
and \U$1847 ( \2032 , \1778 , \351 );
and \U$1848 ( \2033 , \1770 , \349 );
nor \U$1849 ( \2034 , \2032 , \2033 );
xnor \U$1850 ( \2035 , \2034 , \358 );
and \U$1851 ( \2036 , \2030 , \2035 );
and \U$1852 ( \2037 , \2022 , \2035 );
or \U$1853 ( \2038 , \2031 , \2036 , \2037 );
and \U$1854 ( \2039 , \2006 , \2038 );
and \U$1855 ( \2040 , \2023 , \345 );
xor \U$1856 ( \2041 , \1899 , \1903 );
xor \U$1857 ( \2042 , \2041 , \1908 );
and \U$1858 ( \2043 , \2040 , \2042 );
xor \U$1859 ( \2044 , \1869 , \1873 );
xor \U$1860 ( \2045 , \2044 , \1878 );
and \U$1861 ( \2046 , \2042 , \2045 );
and \U$1862 ( \2047 , \2040 , \2045 );
or \U$1863 ( \2048 , \2043 , \2046 , \2047 );
and \U$1864 ( \2049 , \2038 , \2048 );
and \U$1865 ( \2050 , \2006 , \2048 );
or \U$1866 ( \2051 , \2039 , \2049 , \2050 );
xor \U$1867 ( \2052 , \1848 , \1864 );
xor \U$1868 ( \2053 , \2052 , \1881 );
xor \U$1869 ( \2054 , \1886 , \1888 );
xor \U$1870 ( \2055 , \2054 , \1891 );
and \U$1871 ( \2056 , \2053 , \2055 );
xor \U$1872 ( \2057 , \1911 , \1913 );
xor \U$1873 ( \2058 , \2057 , \1915 );
and \U$1874 ( \2059 , \2055 , \2058 );
and \U$1875 ( \2060 , \2053 , \2058 );
or \U$1876 ( \2061 , \2056 , \2059 , \2060 );
and \U$1877 ( \2062 , \2051 , \2061 );
xor \U$1878 ( \2063 , \1721 , \1737 );
xor \U$1879 ( \2064 , \2063 , \1757 );
and \U$1880 ( \2065 , \2061 , \2064 );
and \U$1881 ( \2066 , \2051 , \2064 );
or \U$1882 ( \2067 , \2062 , \2065 , \2066 );
xor \U$1883 ( \2068 , \1884 , \1894 );
xor \U$1884 ( \2069 , \2068 , \1918 );
xor \U$1885 ( \2070 , \1923 , \1925 );
xor \U$1886 ( \2071 , \2070 , \1928 );
and \U$1887 ( \2072 , \2069 , \2071 );
and \U$1888 ( \2073 , \2067 , \2072 );
xor \U$1889 ( \2074 , \1760 , \1785 );
xor \U$1890 ( \2075 , \2074 , \1796 );
and \U$1891 ( \2076 , \2072 , \2075 );
and \U$1892 ( \2077 , \2067 , \2075 );
or \U$1893 ( \2078 , \2073 , \2076 , \2077 );
xor \U$1894 ( \2079 , \1937 , \1939 );
xor \U$1895 ( \2080 , \2079 , \1942 );
and \U$1896 ( \2081 , \2078 , \2080 );
and \U$1897 ( \2082 , \1951 , \2081 );
xor \U$1898 ( \2083 , \1951 , \2081 );
xor \U$1899 ( \2084 , \2078 , \2080 );
and \U$1900 ( \2085 , \621 , \912 );
and \U$1901 ( \2086 , \593 , \910 );
nor \U$1902 ( \2087 , \2085 , \2086 );
xnor \U$1903 ( \2088 , \2087 , \818 );
and \U$1904 ( \2089 , \777 , \740 );
and \U$1905 ( \2090 , \703 , \738 );
nor \U$1906 ( \2091 , \2089 , \2090 );
xnor \U$1907 ( \2092 , \2091 , \668 );
and \U$1908 ( \2093 , \2088 , \2092 );
and \U$1909 ( \2094 , \904 , \604 );
and \U$1910 ( \2095 , \841 , \602 );
nor \U$1911 ( \2096 , \2094 , \2095 );
xnor \U$1912 ( \2097 , \2096 , \561 );
and \U$1913 ( \2098 , \2092 , \2097 );
and \U$1914 ( \2099 , \2088 , \2097 );
or \U$1915 ( \2100 , \2093 , \2098 , \2099 );
and \U$1916 ( \2101 , \353 , \1476 );
and \U$1917 ( \2102 , \323 , \1474 );
nor \U$1918 ( \2103 , \2101 , \2102 );
xnor \U$1919 ( \2104 , \2103 , \1363 );
and \U$1920 ( \2105 , \360 , \1280 );
and \U$1921 ( \2106 , \343 , \1278 );
nor \U$1922 ( \2107 , \2105 , \2106 );
xnor \U$1923 ( \2108 , \2107 , \1177 );
and \U$1924 ( \2109 , \2104 , \2108 );
and \U$1925 ( \2110 , \495 , \1062 );
and \U$1926 ( \2111 , \444 , \1060 );
nor \U$1927 ( \2112 , \2110 , \2111 );
xnor \U$1928 ( \2113 , \2112 , \984 );
and \U$1929 ( \2114 , \2108 , \2113 );
and \U$1930 ( \2115 , \2104 , \2113 );
or \U$1931 ( \2116 , \2109 , \2114 , \2115 );
and \U$1932 ( \2117 , \2100 , \2116 );
_DC r128 ( \2118_nR128 , RIb4c2c60_60 , \288 );
buf \U$1933 ( \2119 , \2118_nR128 );
_DC r127 ( \2120_nR127 , RIb4c2be8_61 , \288 );
buf \U$1934 ( \2121 , \2120_nR127 );
and \U$1935 ( \2122 , \2119 , \2121 );
not \U$1936 ( \2123 , \2122 );
and \U$1937 ( \2124 , \1832 , \2123 );
not \U$1938 ( \2125 , \2124 );
and \U$1939 ( \2126 , \315 , \1955 );
and \U$1940 ( \2127 , \159 , \1953 );
nor \U$1941 ( \2128 , \2126 , \2127 );
xnor \U$1942 ( \2129 , \2128 , \1835 );
and \U$1943 ( \2130 , \2125 , \2129 );
and \U$1944 ( \2131 , \333 , \1742 );
and \U$1945 ( \2132 , \305 , \1740 );
nor \U$1946 ( \2133 , \2131 , \2132 );
xnor \U$1947 ( \2134 , \2133 , \1610 );
and \U$1948 ( \2135 , \2129 , \2134 );
and \U$1949 ( \2136 , \2125 , \2134 );
or \U$1950 ( \2137 , \2130 , \2135 , \2136 );
and \U$1951 ( \2138 , \2116 , \2137 );
and \U$1952 ( \2139 , \2100 , \2137 );
or \U$1953 ( \2140 , \2117 , \2138 , \2139 );
xor \U$1954 ( \2141 , \2010 , \2014 );
xor \U$1955 ( \2142 , \2141 , \2019 );
xor \U$1956 ( \2143 , \1974 , \1978 );
xor \U$1957 ( \2144 , \2143 , \1983 );
and \U$1958 ( \2145 , \2142 , \2144 );
xor \U$1959 ( \2146 , \1991 , \1995 );
xor \U$1960 ( \2147 , \2146 , \2000 );
and \U$1961 ( \2148 , \2144 , \2147 );
and \U$1962 ( \2149 , \2142 , \2147 );
or \U$1963 ( \2150 , \2145 , \2148 , \2149 );
and \U$1964 ( \2151 , \2140 , \2150 );
and \U$1965 ( \2152 , \1778 , \331 );
and \U$1966 ( \2153 , \1770 , \329 );
nor \U$1967 ( \2154 , \2152 , \2153 );
xnor \U$1968 ( \2155 , \2154 , \338 );
and \U$1969 ( \2156 , \2028 , \351 );
and \U$1970 ( \2157 , \2023 , \349 );
nor \U$1971 ( \2158 , \2156 , \2157 );
xnor \U$1972 ( \2159 , \2158 , \358 );
and \U$1973 ( \2160 , \2155 , \2159 );
buf \U$1974 ( \2161 , RIb4bc1f8_91);
and \U$1975 ( \2162 , \2161 , \345 );
and \U$1976 ( \2163 , \2159 , \2162 );
and \U$1977 ( \2164 , \2155 , \2162 );
or \U$1978 ( \2165 , \2160 , \2163 , \2164 );
and \U$1979 ( \2166 , \1194 , \503 );
and \U$1980 ( \2167 , \1104 , \501 );
nor \U$1981 ( \2168 , \2166 , \2167 );
xnor \U$1982 ( \2169 , \2168 , \455 );
and \U$1983 ( \2170 , \1304 , \298 );
and \U$1984 ( \2171 , \1299 , \296 );
nor \U$1985 ( \2172 , \2170 , \2171 );
xnor \U$1986 ( \2173 , \2172 , \303 );
and \U$1987 ( \2174 , \2169 , \2173 );
and \U$1988 ( \2175 , \1537 , \313 );
and \U$1989 ( \2176 , \1422 , \311 );
nor \U$1990 ( \2177 , \2175 , \2176 );
xnor \U$1991 ( \2178 , \2177 , \320 );
and \U$1992 ( \2179 , \2173 , \2178 );
and \U$1993 ( \2180 , \2169 , \2178 );
or \U$1994 ( \2181 , \2174 , \2179 , \2180 );
and \U$1995 ( \2182 , \2165 , \2181 );
xnor \U$1996 ( \2183 , \2027 , \2029 );
and \U$1997 ( \2184 , \2181 , \2183 );
and \U$1998 ( \2185 , \2165 , \2183 );
or \U$1999 ( \2186 , \2182 , \2184 , \2185 );
and \U$2000 ( \2187 , \2150 , \2186 );
and \U$2001 ( \2188 , \2140 , \2186 );
or \U$2002 ( \2189 , \2151 , \2187 , \2188 );
xor \U$2003 ( \2190 , \1836 , \1840 );
xor \U$2004 ( \2191 , \2190 , \1845 );
xor \U$2005 ( \2192 , \1852 , \1856 );
xor \U$2006 ( \2193 , \2192 , \1861 );
and \U$2007 ( \2194 , \2191 , \2193 );
xor \U$2008 ( \2195 , \2040 , \2042 );
xor \U$2009 ( \2196 , \2195 , \2045 );
and \U$2010 ( \2197 , \2193 , \2196 );
and \U$2011 ( \2198 , \2191 , \2196 );
or \U$2012 ( \2199 , \2194 , \2197 , \2198 );
and \U$2013 ( \2200 , \2189 , \2199 );
xor \U$2014 ( \2201 , \2053 , \2055 );
xor \U$2015 ( \2202 , \2201 , \2058 );
and \U$2016 ( \2203 , \2199 , \2202 );
and \U$2017 ( \2204 , \2189 , \2202 );
or \U$2018 ( \2205 , \2200 , \2203 , \2204 );
xor \U$2019 ( \2206 , \2051 , \2061 );
xor \U$2020 ( \2207 , \2206 , \2064 );
and \U$2021 ( \2208 , \2205 , \2207 );
xor \U$2022 ( \2209 , \2069 , \2071 );
and \U$2023 ( \2210 , \2207 , \2209 );
and \U$2024 ( \2211 , \2205 , \2209 );
or \U$2025 ( \2212 , \2208 , \2210 , \2211 );
xor \U$2026 ( \2213 , \2067 , \2072 );
xor \U$2027 ( \2214 , \2213 , \2075 );
and \U$2028 ( \2215 , \2212 , \2214 );
xor \U$2029 ( \2216 , \1921 , \1931 );
xor \U$2030 ( \2217 , \2216 , \1934 );
and \U$2031 ( \2218 , \2214 , \2217 );
and \U$2032 ( \2219 , \2212 , \2217 );
or \U$2033 ( \2220 , \2215 , \2218 , \2219 );
and \U$2034 ( \2221 , \2084 , \2220 );
xor \U$2035 ( \2222 , \2084 , \2220 );
xor \U$2036 ( \2223 , \2212 , \2214 );
xor \U$2037 ( \2224 , \2223 , \2217 );
and \U$2038 ( \2225 , \703 , \912 );
and \U$2039 ( \2226 , \621 , \910 );
nor \U$2040 ( \2227 , \2225 , \2226 );
xnor \U$2041 ( \2228 , \2227 , \818 );
and \U$2042 ( \2229 , \841 , \740 );
and \U$2043 ( \2230 , \777 , \738 );
nor \U$2044 ( \2231 , \2229 , \2230 );
xnor \U$2045 ( \2232 , \2231 , \668 );
and \U$2046 ( \2233 , \2228 , \2232 );
and \U$2047 ( \2234 , \1104 , \604 );
and \U$2048 ( \2235 , \904 , \602 );
nor \U$2049 ( \2236 , \2234 , \2235 );
xnor \U$2050 ( \2237 , \2236 , \561 );
and \U$2051 ( \2238 , \2232 , \2237 );
and \U$2052 ( \2239 , \2228 , \2237 );
or \U$2053 ( \2240 , \2233 , \2238 , \2239 );
and \U$2054 ( \2241 , \343 , \1476 );
and \U$2055 ( \2242 , \353 , \1474 );
nor \U$2056 ( \2243 , \2241 , \2242 );
xnor \U$2057 ( \2244 , \2243 , \1363 );
and \U$2058 ( \2245 , \444 , \1280 );
and \U$2059 ( \2246 , \360 , \1278 );
nor \U$2060 ( \2247 , \2245 , \2246 );
xnor \U$2061 ( \2248 , \2247 , \1177 );
and \U$2062 ( \2249 , \2244 , \2248 );
and \U$2063 ( \2250 , \593 , \1062 );
and \U$2064 ( \2251 , \495 , \1060 );
nor \U$2065 ( \2252 , \2250 , \2251 );
xnor \U$2066 ( \2253 , \2252 , \984 );
and \U$2067 ( \2254 , \2248 , \2253 );
and \U$2068 ( \2255 , \2244 , \2253 );
or \U$2069 ( \2256 , \2249 , \2254 , \2255 );
and \U$2070 ( \2257 , \2240 , \2256 );
xor \U$2071 ( \2258 , \1832 , \2119 );
xor \U$2072 ( \2259 , \2119 , \2121 );
not \U$2073 ( \2260 , \2259 );
and \U$2074 ( \2261 , \2258 , \2260 );
and \U$2075 ( \2262 , \159 , \2261 );
not \U$2076 ( \2263 , \2262 );
xnor \U$2077 ( \2264 , \2263 , \2124 );
and \U$2078 ( \2265 , \305 , \1955 );
and \U$2079 ( \2266 , \315 , \1953 );
nor \U$2080 ( \2267 , \2265 , \2266 );
xnor \U$2081 ( \2268 , \2267 , \1835 );
and \U$2082 ( \2269 , \2264 , \2268 );
and \U$2083 ( \2270 , \323 , \1742 );
and \U$2084 ( \2271 , \333 , \1740 );
nor \U$2085 ( \2272 , \2270 , \2271 );
xnor \U$2086 ( \2273 , \2272 , \1610 );
and \U$2087 ( \2274 , \2268 , \2273 );
and \U$2088 ( \2275 , \2264 , \2273 );
or \U$2089 ( \2276 , \2269 , \2274 , \2275 );
and \U$2090 ( \2277 , \2256 , \2276 );
and \U$2091 ( \2278 , \2240 , \2276 );
or \U$2092 ( \2279 , \2257 , \2277 , \2278 );
and \U$2093 ( \2280 , \1299 , \503 );
and \U$2094 ( \2281 , \1194 , \501 );
nor \U$2095 ( \2282 , \2280 , \2281 );
xnor \U$2096 ( \2283 , \2282 , \455 );
and \U$2097 ( \2284 , \1422 , \298 );
and \U$2098 ( \2285 , \1304 , \296 );
nor \U$2099 ( \2286 , \2284 , \2285 );
xnor \U$2100 ( \2287 , \2286 , \303 );
and \U$2101 ( \2288 , \2283 , \2287 );
and \U$2102 ( \2289 , \1770 , \313 );
and \U$2103 ( \2290 , \1537 , \311 );
nor \U$2104 ( \2291 , \2289 , \2290 );
xnor \U$2105 ( \2292 , \2291 , \320 );
and \U$2106 ( \2293 , \2287 , \2292 );
and \U$2107 ( \2294 , \2283 , \2292 );
or \U$2108 ( \2295 , \2288 , \2293 , \2294 );
and \U$2109 ( \2296 , \2023 , \331 );
and \U$2110 ( \2297 , \1778 , \329 );
nor \U$2111 ( \2298 , \2296 , \2297 );
xnor \U$2112 ( \2299 , \2298 , \338 );
and \U$2113 ( \2300 , \2161 , \351 );
and \U$2114 ( \2301 , \2028 , \349 );
nor \U$2115 ( \2302 , \2300 , \2301 );
xnor \U$2116 ( \2303 , \2302 , \358 );
and \U$2117 ( \2304 , \2299 , \2303 );
buf \U$2118 ( \2305 , RIb4bc180_92);
and \U$2119 ( \2306 , \2305 , \345 );
and \U$2120 ( \2307 , \2303 , \2306 );
and \U$2121 ( \2308 , \2299 , \2306 );
or \U$2122 ( \2309 , \2304 , \2307 , \2308 );
and \U$2123 ( \2310 , \2295 , \2309 );
xor \U$2124 ( \2311 , \2155 , \2159 );
xor \U$2125 ( \2312 , \2311 , \2162 );
and \U$2126 ( \2313 , \2309 , \2312 );
and \U$2127 ( \2314 , \2295 , \2312 );
or \U$2128 ( \2315 , \2310 , \2313 , \2314 );
and \U$2129 ( \2316 , \2279 , \2315 );
xor \U$2130 ( \2317 , \2088 , \2092 );
xor \U$2131 ( \2318 , \2317 , \2097 );
xor \U$2132 ( \2319 , \2104 , \2108 );
xor \U$2133 ( \2320 , \2319 , \2113 );
and \U$2134 ( \2321 , \2318 , \2320 );
xor \U$2135 ( \2322 , \2169 , \2173 );
xor \U$2136 ( \2323 , \2322 , \2178 );
and \U$2137 ( \2324 , \2320 , \2323 );
and \U$2138 ( \2325 , \2318 , \2323 );
or \U$2139 ( \2326 , \2321 , \2324 , \2325 );
and \U$2140 ( \2327 , \2315 , \2326 );
and \U$2141 ( \2328 , \2279 , \2326 );
or \U$2142 ( \2329 , \2316 , \2327 , \2328 );
xor \U$2143 ( \2330 , \1958 , \1962 );
xor \U$2144 ( \2331 , \2330 , \1967 );
xor \U$2145 ( \2332 , \2142 , \2144 );
xor \U$2146 ( \2333 , \2332 , \2147 );
and \U$2147 ( \2334 , \2331 , \2333 );
xor \U$2148 ( \2335 , \2165 , \2181 );
xor \U$2149 ( \2336 , \2335 , \2183 );
and \U$2150 ( \2337 , \2333 , \2336 );
and \U$2151 ( \2338 , \2331 , \2336 );
or \U$2152 ( \2339 , \2334 , \2337 , \2338 );
and \U$2153 ( \2340 , \2329 , \2339 );
xor \U$2154 ( \2341 , \2022 , \2030 );
xor \U$2155 ( \2342 , \2341 , \2035 );
and \U$2156 ( \2343 , \2339 , \2342 );
and \U$2157 ( \2344 , \2329 , \2342 );
or \U$2158 ( \2345 , \2340 , \2343 , \2344 );
xor \U$2159 ( \2346 , \1970 , \1986 );
xor \U$2160 ( \2347 , \2346 , \2003 );
xor \U$2161 ( \2348 , \2140 , \2150 );
xor \U$2162 ( \2349 , \2348 , \2186 );
and \U$2163 ( \2350 , \2347 , \2349 );
xor \U$2164 ( \2351 , \2191 , \2193 );
xor \U$2165 ( \2352 , \2351 , \2196 );
and \U$2166 ( \2353 , \2349 , \2352 );
and \U$2167 ( \2354 , \2347 , \2352 );
or \U$2168 ( \2355 , \2350 , \2353 , \2354 );
and \U$2169 ( \2356 , \2345 , \2355 );
xor \U$2170 ( \2357 , \2006 , \2038 );
xor \U$2171 ( \2358 , \2357 , \2048 );
and \U$2172 ( \2359 , \2355 , \2358 );
and \U$2173 ( \2360 , \2345 , \2358 );
or \U$2174 ( \2361 , \2356 , \2359 , \2360 );
xor \U$2175 ( \2362 , \2205 , \2207 );
xor \U$2176 ( \2363 , \2362 , \2209 );
and \U$2177 ( \2364 , \2361 , \2363 );
and \U$2178 ( \2365 , \2224 , \2364 );
xor \U$2179 ( \2366 , \2224 , \2364 );
xor \U$2180 ( \2367 , \2361 , \2363 );
_DC r126 ( \2368_nR126 , RIb4c2b70_62 , \288 );
buf \U$2181 ( \2369 , \2368_nR126 );
_DC r125 ( \2370_nR125 , RIb4c2af8_63 , \288 );
buf \U$2182 ( \2371 , \2370_nR125 );
and \U$2183 ( \2372 , \2369 , \2371 );
not \U$2184 ( \2373 , \2372 );
and \U$2185 ( \2374 , \2121 , \2373 );
not \U$2186 ( \2375 , \2374 );
and \U$2187 ( \2376 , \315 , \2261 );
and \U$2188 ( \2377 , \159 , \2259 );
nor \U$2189 ( \2378 , \2376 , \2377 );
xnor \U$2190 ( \2379 , \2378 , \2124 );
and \U$2191 ( \2380 , \2375 , \2379 );
and \U$2192 ( \2381 , \333 , \1955 );
and \U$2193 ( \2382 , \305 , \1953 );
nor \U$2194 ( \2383 , \2381 , \2382 );
xnor \U$2195 ( \2384 , \2383 , \1835 );
and \U$2196 ( \2385 , \2379 , \2384 );
and \U$2197 ( \2386 , \2375 , \2384 );
or \U$2198 ( \2387 , \2380 , \2385 , \2386 );
and \U$2199 ( \2388 , \353 , \1742 );
and \U$2200 ( \2389 , \323 , \1740 );
nor \U$2201 ( \2390 , \2388 , \2389 );
xnor \U$2202 ( \2391 , \2390 , \1610 );
and \U$2203 ( \2392 , \360 , \1476 );
and \U$2204 ( \2393 , \343 , \1474 );
nor \U$2205 ( \2394 , \2392 , \2393 );
xnor \U$2206 ( \2395 , \2394 , \1363 );
and \U$2207 ( \2396 , \2391 , \2395 );
and \U$2208 ( \2397 , \495 , \1280 );
and \U$2209 ( \2398 , \444 , \1278 );
nor \U$2210 ( \2399 , \2397 , \2398 );
xnor \U$2211 ( \2400 , \2399 , \1177 );
and \U$2212 ( \2401 , \2395 , \2400 );
and \U$2213 ( \2402 , \2391 , \2400 );
or \U$2214 ( \2403 , \2396 , \2401 , \2402 );
and \U$2215 ( \2404 , \2387 , \2403 );
and \U$2216 ( \2405 , \621 , \1062 );
and \U$2217 ( \2406 , \593 , \1060 );
nor \U$2218 ( \2407 , \2405 , \2406 );
xnor \U$2219 ( \2408 , \2407 , \984 );
and \U$2220 ( \2409 , \777 , \912 );
and \U$2221 ( \2410 , \703 , \910 );
nor \U$2222 ( \2411 , \2409 , \2410 );
xnor \U$2223 ( \2412 , \2411 , \818 );
and \U$2224 ( \2413 , \2408 , \2412 );
and \U$2225 ( \2414 , \904 , \740 );
and \U$2226 ( \2415 , \841 , \738 );
nor \U$2227 ( \2416 , \2414 , \2415 );
xnor \U$2228 ( \2417 , \2416 , \668 );
and \U$2229 ( \2418 , \2412 , \2417 );
and \U$2230 ( \2419 , \2408 , \2417 );
or \U$2231 ( \2420 , \2413 , \2418 , \2419 );
and \U$2232 ( \2421 , \2403 , \2420 );
and \U$2233 ( \2422 , \2387 , \2420 );
or \U$2234 ( \2423 , \2404 , \2421 , \2422 );
xor \U$2235 ( \2424 , \2228 , \2232 );
xor \U$2236 ( \2425 , \2424 , \2237 );
xor \U$2237 ( \2426 , \2283 , \2287 );
xor \U$2238 ( \2427 , \2426 , \2292 );
and \U$2239 ( \2428 , \2425 , \2427 );
xor \U$2240 ( \2429 , \2299 , \2303 );
xor \U$2241 ( \2430 , \2429 , \2306 );
and \U$2242 ( \2431 , \2427 , \2430 );
and \U$2243 ( \2432 , \2425 , \2430 );
or \U$2244 ( \2433 , \2428 , \2431 , \2432 );
and \U$2245 ( \2434 , \2423 , \2433 );
and \U$2246 ( \2435 , \1778 , \313 );
and \U$2247 ( \2436 , \1770 , \311 );
nor \U$2248 ( \2437 , \2435 , \2436 );
xnor \U$2249 ( \2438 , \2437 , \320 );
and \U$2250 ( \2439 , \2028 , \331 );
and \U$2251 ( \2440 , \2023 , \329 );
nor \U$2252 ( \2441 , \2439 , \2440 );
xnor \U$2253 ( \2442 , \2441 , \338 );
and \U$2254 ( \2443 , \2438 , \2442 );
and \U$2255 ( \2444 , \2305 , \351 );
and \U$2256 ( \2445 , \2161 , \349 );
nor \U$2257 ( \2446 , \2444 , \2445 );
xnor \U$2258 ( \2447 , \2446 , \358 );
and \U$2259 ( \2448 , \2442 , \2447 );
and \U$2260 ( \2449 , \2438 , \2447 );
or \U$2261 ( \2450 , \2443 , \2448 , \2449 );
and \U$2262 ( \2451 , \1194 , \604 );
and \U$2263 ( \2452 , \1104 , \602 );
nor \U$2264 ( \2453 , \2451 , \2452 );
xnor \U$2265 ( \2454 , \2453 , \561 );
and \U$2266 ( \2455 , \1304 , \503 );
and \U$2267 ( \2456 , \1299 , \501 );
nor \U$2268 ( \2457 , \2455 , \2456 );
xnor \U$2269 ( \2458 , \2457 , \455 );
and \U$2270 ( \2459 , \2454 , \2458 );
and \U$2271 ( \2460 , \1537 , \298 );
and \U$2272 ( \2461 , \1422 , \296 );
nor \U$2273 ( \2462 , \2460 , \2461 );
xnor \U$2274 ( \2463 , \2462 , \303 );
and \U$2275 ( \2464 , \2458 , \2463 );
and \U$2276 ( \2465 , \2454 , \2463 );
or \U$2277 ( \2466 , \2459 , \2464 , \2465 );
or \U$2278 ( \2467 , \2450 , \2466 );
and \U$2279 ( \2468 , \2433 , \2467 );
and \U$2280 ( \2469 , \2423 , \2467 );
or \U$2281 ( \2470 , \2434 , \2468 , \2469 );
xor \U$2282 ( \2471 , \2125 , \2129 );
xor \U$2283 ( \2472 , \2471 , \2134 );
xor \U$2284 ( \2473 , \2295 , \2309 );
xor \U$2285 ( \2474 , \2473 , \2312 );
and \U$2286 ( \2475 , \2472 , \2474 );
xor \U$2287 ( \2476 , \2318 , \2320 );
xor \U$2288 ( \2477 , \2476 , \2323 );
and \U$2289 ( \2478 , \2474 , \2477 );
and \U$2290 ( \2479 , \2472 , \2477 );
or \U$2291 ( \2480 , \2475 , \2478 , \2479 );
and \U$2292 ( \2481 , \2470 , \2480 );
xor \U$2293 ( \2482 , \2100 , \2116 );
xor \U$2294 ( \2483 , \2482 , \2137 );
and \U$2295 ( \2484 , \2480 , \2483 );
and \U$2296 ( \2485 , \2470 , \2483 );
or \U$2297 ( \2486 , \2481 , \2484 , \2485 );
xor \U$2298 ( \2487 , \2329 , \2339 );
xor \U$2299 ( \2488 , \2487 , \2342 );
and \U$2300 ( \2489 , \2486 , \2488 );
xor \U$2301 ( \2490 , \2347 , \2349 );
xor \U$2302 ( \2491 , \2490 , \2352 );
and \U$2303 ( \2492 , \2488 , \2491 );
and \U$2304 ( \2493 , \2486 , \2491 );
or \U$2305 ( \2494 , \2489 , \2492 , \2493 );
xor \U$2306 ( \2495 , \2345 , \2355 );
xor \U$2307 ( \2496 , \2495 , \2358 );
and \U$2308 ( \2497 , \2494 , \2496 );
xor \U$2309 ( \2498 , \2189 , \2199 );
xor \U$2310 ( \2499 , \2498 , \2202 );
and \U$2311 ( \2500 , \2496 , \2499 );
and \U$2312 ( \2501 , \2494 , \2499 );
or \U$2313 ( \2502 , \2497 , \2500 , \2501 );
and \U$2314 ( \2503 , \2367 , \2502 );
xor \U$2315 ( \2504 , \2367 , \2502 );
xor \U$2316 ( \2505 , \2494 , \2496 );
xor \U$2317 ( \2506 , \2505 , \2499 );
and \U$2318 ( \2507 , \1299 , \604 );
and \U$2319 ( \2508 , \1194 , \602 );
nor \U$2320 ( \2509 , \2507 , \2508 );
xnor \U$2321 ( \2510 , \2509 , \561 );
and \U$2322 ( \2511 , \1422 , \503 );
and \U$2323 ( \2512 , \1304 , \501 );
nor \U$2324 ( \2513 , \2511 , \2512 );
xnor \U$2325 ( \2514 , \2513 , \455 );
and \U$2326 ( \2515 , \2510 , \2514 );
and \U$2327 ( \2516 , \1770 , \298 );
and \U$2328 ( \2517 , \1537 , \296 );
nor \U$2329 ( \2518 , \2516 , \2517 );
xnor \U$2330 ( \2519 , \2518 , \303 );
and \U$2331 ( \2520 , \2514 , \2519 );
and \U$2332 ( \2521 , \2510 , \2519 );
or \U$2333 ( \2522 , \2515 , \2520 , \2521 );
and \U$2334 ( \2523 , \2023 , \313 );
and \U$2335 ( \2524 , \1778 , \311 );
nor \U$2336 ( \2525 , \2523 , \2524 );
xnor \U$2337 ( \2526 , \2525 , \320 );
and \U$2338 ( \2527 , \2161 , \331 );
and \U$2339 ( \2528 , \2028 , \329 );
nor \U$2340 ( \2529 , \2527 , \2528 );
xnor \U$2341 ( \2530 , \2529 , \338 );
and \U$2342 ( \2531 , \2526 , \2530 );
buf \U$2343 ( \2532 , RIb4bc108_93);
and \U$2344 ( \2533 , \2532 , \351 );
and \U$2345 ( \2534 , \2305 , \349 );
nor \U$2346 ( \2535 , \2533 , \2534 );
xnor \U$2347 ( \2536 , \2535 , \358 );
and \U$2348 ( \2537 , \2530 , \2536 );
and \U$2349 ( \2538 , \2526 , \2536 );
or \U$2350 ( \2539 , \2531 , \2537 , \2538 );
and \U$2351 ( \2540 , \2522 , \2539 );
buf \U$2352 ( \2541 , RIb4bc090_94);
and \U$2353 ( \2542 , \2541 , \345 );
buf \U$2354 ( \2543 , \2542 );
and \U$2355 ( \2544 , \2539 , \2543 );
and \U$2356 ( \2545 , \2522 , \2543 );
or \U$2357 ( \2546 , \2540 , \2544 , \2545 );
xor \U$2358 ( \2547 , \2121 , \2369 );
xor \U$2359 ( \2548 , \2369 , \2371 );
not \U$2360 ( \2549 , \2548 );
and \U$2361 ( \2550 , \2547 , \2549 );
and \U$2362 ( \2551 , \159 , \2550 );
not \U$2363 ( \2552 , \2551 );
xnor \U$2364 ( \2553 , \2552 , \2374 );
and \U$2365 ( \2554 , \305 , \2261 );
and \U$2366 ( \2555 , \315 , \2259 );
nor \U$2367 ( \2556 , \2554 , \2555 );
xnor \U$2368 ( \2557 , \2556 , \2124 );
and \U$2369 ( \2558 , \2553 , \2557 );
and \U$2370 ( \2559 , \323 , \1955 );
and \U$2371 ( \2560 , \333 , \1953 );
nor \U$2372 ( \2561 , \2559 , \2560 );
xnor \U$2373 ( \2562 , \2561 , \1835 );
and \U$2374 ( \2563 , \2557 , \2562 );
and \U$2375 ( \2564 , \2553 , \2562 );
or \U$2376 ( \2565 , \2558 , \2563 , \2564 );
and \U$2377 ( \2566 , \343 , \1742 );
and \U$2378 ( \2567 , \353 , \1740 );
nor \U$2379 ( \2568 , \2566 , \2567 );
xnor \U$2380 ( \2569 , \2568 , \1610 );
and \U$2381 ( \2570 , \444 , \1476 );
and \U$2382 ( \2571 , \360 , \1474 );
nor \U$2383 ( \2572 , \2570 , \2571 );
xnor \U$2384 ( \2573 , \2572 , \1363 );
and \U$2385 ( \2574 , \2569 , \2573 );
and \U$2386 ( \2575 , \593 , \1280 );
and \U$2387 ( \2576 , \495 , \1278 );
nor \U$2388 ( \2577 , \2575 , \2576 );
xnor \U$2389 ( \2578 , \2577 , \1177 );
and \U$2390 ( \2579 , \2573 , \2578 );
and \U$2391 ( \2580 , \2569 , \2578 );
or \U$2392 ( \2581 , \2574 , \2579 , \2580 );
and \U$2393 ( \2582 , \2565 , \2581 );
and \U$2394 ( \2583 , \703 , \1062 );
and \U$2395 ( \2584 , \621 , \1060 );
nor \U$2396 ( \2585 , \2583 , \2584 );
xnor \U$2397 ( \2586 , \2585 , \984 );
and \U$2398 ( \2587 , \841 , \912 );
and \U$2399 ( \2588 , \777 , \910 );
nor \U$2400 ( \2589 , \2587 , \2588 );
xnor \U$2401 ( \2590 , \2589 , \818 );
and \U$2402 ( \2591 , \2586 , \2590 );
and \U$2403 ( \2592 , \1104 , \740 );
and \U$2404 ( \2593 , \904 , \738 );
nor \U$2405 ( \2594 , \2592 , \2593 );
xnor \U$2406 ( \2595 , \2594 , \668 );
and \U$2407 ( \2596 , \2590 , \2595 );
and \U$2408 ( \2597 , \2586 , \2595 );
or \U$2409 ( \2598 , \2591 , \2596 , \2597 );
and \U$2410 ( \2599 , \2581 , \2598 );
and \U$2411 ( \2600 , \2565 , \2598 );
or \U$2412 ( \2601 , \2582 , \2599 , \2600 );
and \U$2413 ( \2602 , \2546 , \2601 );
and \U$2414 ( \2603 , \2532 , \345 );
xor \U$2415 ( \2604 , \2438 , \2442 );
xor \U$2416 ( \2605 , \2604 , \2447 );
and \U$2417 ( \2606 , \2603 , \2605 );
xor \U$2418 ( \2607 , \2454 , \2458 );
xor \U$2419 ( \2608 , \2607 , \2463 );
and \U$2420 ( \2609 , \2605 , \2608 );
and \U$2421 ( \2610 , \2603 , \2608 );
or \U$2422 ( \2611 , \2606 , \2609 , \2610 );
and \U$2423 ( \2612 , \2601 , \2611 );
and \U$2424 ( \2613 , \2546 , \2611 );
or \U$2425 ( \2614 , \2602 , \2612 , \2613 );
xor \U$2426 ( \2615 , \2375 , \2379 );
xor \U$2427 ( \2616 , \2615 , \2384 );
xor \U$2428 ( \2617 , \2391 , \2395 );
xor \U$2429 ( \2618 , \2617 , \2400 );
and \U$2430 ( \2619 , \2616 , \2618 );
xor \U$2431 ( \2620 , \2408 , \2412 );
xor \U$2432 ( \2621 , \2620 , \2417 );
and \U$2433 ( \2622 , \2618 , \2621 );
and \U$2434 ( \2623 , \2616 , \2621 );
or \U$2435 ( \2624 , \2619 , \2622 , \2623 );
xor \U$2436 ( \2625 , \2244 , \2248 );
xor \U$2437 ( \2626 , \2625 , \2253 );
and \U$2438 ( \2627 , \2624 , \2626 );
xor \U$2439 ( \2628 , \2264 , \2268 );
xor \U$2440 ( \2629 , \2628 , \2273 );
and \U$2441 ( \2630 , \2626 , \2629 );
and \U$2442 ( \2631 , \2624 , \2629 );
or \U$2443 ( \2632 , \2627 , \2630 , \2631 );
and \U$2444 ( \2633 , \2614 , \2632 );
xor \U$2445 ( \2634 , \2387 , \2403 );
xor \U$2446 ( \2635 , \2634 , \2420 );
xor \U$2447 ( \2636 , \2425 , \2427 );
xor \U$2448 ( \2637 , \2636 , \2430 );
and \U$2449 ( \2638 , \2635 , \2637 );
xnor \U$2450 ( \2639 , \2450 , \2466 );
and \U$2451 ( \2640 , \2637 , \2639 );
and \U$2452 ( \2641 , \2635 , \2639 );
or \U$2453 ( \2642 , \2638 , \2640 , \2641 );
and \U$2454 ( \2643 , \2632 , \2642 );
and \U$2455 ( \2644 , \2614 , \2642 );
or \U$2456 ( \2645 , \2633 , \2643 , \2644 );
xor \U$2457 ( \2646 , \2240 , \2256 );
xor \U$2458 ( \2647 , \2646 , \2276 );
xor \U$2459 ( \2648 , \2423 , \2433 );
xor \U$2460 ( \2649 , \2648 , \2467 );
and \U$2461 ( \2650 , \2647 , \2649 );
xor \U$2462 ( \2651 , \2472 , \2474 );
xor \U$2463 ( \2652 , \2651 , \2477 );
and \U$2464 ( \2653 , \2649 , \2652 );
and \U$2465 ( \2654 , \2647 , \2652 );
or \U$2466 ( \2655 , \2650 , \2653 , \2654 );
and \U$2467 ( \2656 , \2645 , \2655 );
xor \U$2468 ( \2657 , \2331 , \2333 );
xor \U$2469 ( \2658 , \2657 , \2336 );
and \U$2470 ( \2659 , \2655 , \2658 );
and \U$2471 ( \2660 , \2645 , \2658 );
or \U$2472 ( \2661 , \2656 , \2659 , \2660 );
xor \U$2473 ( \2662 , \2279 , \2315 );
xor \U$2474 ( \2663 , \2662 , \2326 );
xor \U$2475 ( \2664 , \2470 , \2480 );
xor \U$2476 ( \2665 , \2664 , \2483 );
and \U$2477 ( \2666 , \2663 , \2665 );
and \U$2478 ( \2667 , \2661 , \2666 );
xor \U$2479 ( \2668 , \2486 , \2488 );
xor \U$2480 ( \2669 , \2668 , \2491 );
and \U$2481 ( \2670 , \2666 , \2669 );
and \U$2482 ( \2671 , \2661 , \2669 );
or \U$2483 ( \2672 , \2667 , \2670 , \2671 );
and \U$2484 ( \2673 , \2506 , \2672 );
xor \U$2485 ( \2674 , \2506 , \2672 );
xor \U$2486 ( \2675 , \2661 , \2666 );
xor \U$2487 ( \2676 , \2675 , \2669 );
and \U$2488 ( \2677 , \621 , \1280 );
and \U$2489 ( \2678 , \593 , \1278 );
nor \U$2490 ( \2679 , \2677 , \2678 );
xnor \U$2491 ( \2680 , \2679 , \1177 );
and \U$2492 ( \2681 , \777 , \1062 );
and \U$2493 ( \2682 , \703 , \1060 );
nor \U$2494 ( \2683 , \2681 , \2682 );
xnor \U$2495 ( \2684 , \2683 , \984 );
and \U$2496 ( \2685 , \2680 , \2684 );
and \U$2497 ( \2686 , \904 , \912 );
and \U$2498 ( \2687 , \841 , \910 );
nor \U$2499 ( \2688 , \2686 , \2687 );
xnor \U$2500 ( \2689 , \2688 , \818 );
and \U$2501 ( \2690 , \2684 , \2689 );
and \U$2502 ( \2691 , \2680 , \2689 );
or \U$2503 ( \2692 , \2685 , \2690 , \2691 );
not \U$2504 ( \2693 , \2371 );
and \U$2505 ( \2694 , \315 , \2550 );
and \U$2506 ( \2695 , \159 , \2548 );
nor \U$2507 ( \2696 , \2694 , \2695 );
xnor \U$2508 ( \2697 , \2696 , \2374 );
and \U$2509 ( \2698 , \2693 , \2697 );
and \U$2510 ( \2699 , \333 , \2261 );
and \U$2511 ( \2700 , \305 , \2259 );
nor \U$2512 ( \2701 , \2699 , \2700 );
xnor \U$2513 ( \2702 , \2701 , \2124 );
and \U$2514 ( \2703 , \2697 , \2702 );
and \U$2515 ( \2704 , \2693 , \2702 );
or \U$2516 ( \2705 , \2698 , \2703 , \2704 );
and \U$2517 ( \2706 , \2692 , \2705 );
and \U$2518 ( \2707 , \353 , \1955 );
and \U$2519 ( \2708 , \323 , \1953 );
nor \U$2520 ( \2709 , \2707 , \2708 );
xnor \U$2521 ( \2710 , \2709 , \1835 );
and \U$2522 ( \2711 , \360 , \1742 );
and \U$2523 ( \2712 , \343 , \1740 );
nor \U$2524 ( \2713 , \2711 , \2712 );
xnor \U$2525 ( \2714 , \2713 , \1610 );
and \U$2526 ( \2715 , \2710 , \2714 );
and \U$2527 ( \2716 , \495 , \1476 );
and \U$2528 ( \2717 , \444 , \1474 );
nor \U$2529 ( \2718 , \2716 , \2717 );
xnor \U$2530 ( \2719 , \2718 , \1363 );
and \U$2531 ( \2720 , \2714 , \2719 );
and \U$2532 ( \2721 , \2710 , \2719 );
or \U$2533 ( \2722 , \2715 , \2720 , \2721 );
and \U$2534 ( \2723 , \2705 , \2722 );
and \U$2535 ( \2724 , \2692 , \2722 );
or \U$2536 ( \2725 , \2706 , \2723 , \2724 );
and \U$2537 ( \2726 , \1778 , \298 );
and \U$2538 ( \2727 , \1770 , \296 );
nor \U$2539 ( \2728 , \2726 , \2727 );
xnor \U$2540 ( \2729 , \2728 , \303 );
and \U$2541 ( \2730 , \2028 , \313 );
and \U$2542 ( \2731 , \2023 , \311 );
nor \U$2543 ( \2732 , \2730 , \2731 );
xnor \U$2544 ( \2733 , \2732 , \320 );
and \U$2545 ( \2734 , \2729 , \2733 );
and \U$2546 ( \2735 , \2305 , \331 );
and \U$2547 ( \2736 , \2161 , \329 );
nor \U$2548 ( \2737 , \2735 , \2736 );
xnor \U$2549 ( \2738 , \2737 , \338 );
and \U$2550 ( \2739 , \2733 , \2738 );
and \U$2551 ( \2740 , \2729 , \2738 );
or \U$2552 ( \2741 , \2734 , \2739 , \2740 );
and \U$2553 ( \2742 , \1194 , \740 );
and \U$2554 ( \2743 , \1104 , \738 );
nor \U$2555 ( \2744 , \2742 , \2743 );
xnor \U$2556 ( \2745 , \2744 , \668 );
and \U$2557 ( \2746 , \1304 , \604 );
and \U$2558 ( \2747 , \1299 , \602 );
nor \U$2559 ( \2748 , \2746 , \2747 );
xnor \U$2560 ( \2749 , \2748 , \561 );
and \U$2561 ( \2750 , \2745 , \2749 );
and \U$2562 ( \2751 , \1537 , \503 );
and \U$2563 ( \2752 , \1422 , \501 );
nor \U$2564 ( \2753 , \2751 , \2752 );
xnor \U$2565 ( \2754 , \2753 , \455 );
and \U$2566 ( \2755 , \2749 , \2754 );
and \U$2567 ( \2756 , \2745 , \2754 );
or \U$2568 ( \2757 , \2750 , \2755 , \2756 );
and \U$2569 ( \2758 , \2741 , \2757 );
and \U$2570 ( \2759 , \2541 , \351 );
and \U$2571 ( \2760 , \2532 , \349 );
nor \U$2572 ( \2761 , \2759 , \2760 );
xnor \U$2573 ( \2762 , \2761 , \358 );
buf \U$2574 ( \2763 , RIb4bc018_95);
and \U$2575 ( \2764 , \2763 , \345 );
or \U$2576 ( \2765 , \2762 , \2764 );
and \U$2577 ( \2766 , \2757 , \2765 );
and \U$2578 ( \2767 , \2741 , \2765 );
or \U$2579 ( \2768 , \2758 , \2766 , \2767 );
and \U$2580 ( \2769 , \2725 , \2768 );
xor \U$2581 ( \2770 , \2510 , \2514 );
xor \U$2582 ( \2771 , \2770 , \2519 );
xor \U$2583 ( \2772 , \2526 , \2530 );
xor \U$2584 ( \2773 , \2772 , \2536 );
and \U$2585 ( \2774 , \2771 , \2773 );
not \U$2586 ( \2775 , \2542 );
and \U$2587 ( \2776 , \2773 , \2775 );
and \U$2588 ( \2777 , \2771 , \2775 );
or \U$2589 ( \2778 , \2774 , \2776 , \2777 );
and \U$2590 ( \2779 , \2768 , \2778 );
and \U$2591 ( \2780 , \2725 , \2778 );
or \U$2592 ( \2781 , \2769 , \2779 , \2780 );
xor \U$2593 ( \2782 , \2553 , \2557 );
xor \U$2594 ( \2783 , \2782 , \2562 );
xor \U$2595 ( \2784 , \2569 , \2573 );
xor \U$2596 ( \2785 , \2784 , \2578 );
and \U$2597 ( \2786 , \2783 , \2785 );
xor \U$2598 ( \2787 , \2586 , \2590 );
xor \U$2599 ( \2788 , \2787 , \2595 );
and \U$2600 ( \2789 , \2785 , \2788 );
and \U$2601 ( \2790 , \2783 , \2788 );
or \U$2602 ( \2791 , \2786 , \2789 , \2790 );
xor \U$2603 ( \2792 , \2603 , \2605 );
xor \U$2604 ( \2793 , \2792 , \2608 );
and \U$2605 ( \2794 , \2791 , \2793 );
xor \U$2606 ( \2795 , \2616 , \2618 );
xor \U$2607 ( \2796 , \2795 , \2621 );
and \U$2608 ( \2797 , \2793 , \2796 );
and \U$2609 ( \2798 , \2791 , \2796 );
or \U$2610 ( \2799 , \2794 , \2797 , \2798 );
and \U$2611 ( \2800 , \2781 , \2799 );
xor \U$2612 ( \2801 , \2635 , \2637 );
xor \U$2613 ( \2802 , \2801 , \2639 );
and \U$2614 ( \2803 , \2799 , \2802 );
and \U$2615 ( \2804 , \2781 , \2802 );
or \U$2616 ( \2805 , \2800 , \2803 , \2804 );
xor \U$2617 ( \2806 , \2614 , \2632 );
xor \U$2618 ( \2807 , \2806 , \2642 );
and \U$2619 ( \2808 , \2805 , \2807 );
xor \U$2620 ( \2809 , \2647 , \2649 );
xor \U$2621 ( \2810 , \2809 , \2652 );
and \U$2622 ( \2811 , \2807 , \2810 );
and \U$2623 ( \2812 , \2805 , \2810 );
or \U$2624 ( \2813 , \2808 , \2811 , \2812 );
xor \U$2625 ( \2814 , \2645 , \2655 );
xor \U$2626 ( \2815 , \2814 , \2658 );
and \U$2627 ( \2816 , \2813 , \2815 );
xor \U$2628 ( \2817 , \2663 , \2665 );
and \U$2629 ( \2818 , \2815 , \2817 );
and \U$2630 ( \2819 , \2813 , \2817 );
or \U$2631 ( \2820 , \2816 , \2818 , \2819 );
and \U$2632 ( \2821 , \2676 , \2820 );
xor \U$2633 ( \2822 , \2676 , \2820 );
xor \U$2634 ( \2823 , \2813 , \2815 );
xor \U$2635 ( \2824 , \2823 , \2817 );
and \U$2636 ( \2825 , \1770 , \503 );
and \U$2637 ( \2826 , \1537 , \501 );
nor \U$2638 ( \2827 , \2825 , \2826 );
xnor \U$2639 ( \2828 , \2827 , \455 );
and \U$2640 ( \2829 , \2023 , \298 );
and \U$2641 ( \2830 , \1778 , \296 );
nor \U$2642 ( \2831 , \2829 , \2830 );
xnor \U$2643 ( \2832 , \2831 , \303 );
and \U$2644 ( \2833 , \2828 , \2832 );
and \U$2645 ( \2834 , \2161 , \313 );
and \U$2646 ( \2835 , \2028 , \311 );
nor \U$2647 ( \2836 , \2834 , \2835 );
xnor \U$2648 ( \2837 , \2836 , \320 );
and \U$2649 ( \2838 , \2832 , \2837 );
and \U$2650 ( \2839 , \2828 , \2837 );
or \U$2651 ( \2840 , \2833 , \2838 , \2839 );
and \U$2652 ( \2841 , \2532 , \331 );
and \U$2653 ( \2842 , \2305 , \329 );
nor \U$2654 ( \2843 , \2841 , \2842 );
xnor \U$2655 ( \2844 , \2843 , \338 );
and \U$2656 ( \2845 , \2763 , \351 );
and \U$2657 ( \2846 , \2541 , \349 );
nor \U$2658 ( \2847 , \2845 , \2846 );
xnor \U$2659 ( \2848 , \2847 , \358 );
and \U$2660 ( \2849 , \2844 , \2848 );
buf \U$2661 ( \2850 , RIb4bbfa0_96);
nand \U$2662 ( \2851 , \2850 , \345 );
not \U$2663 ( \2852 , \2851 );
and \U$2664 ( \2853 , \2848 , \2852 );
and \U$2665 ( \2854 , \2844 , \2852 );
or \U$2666 ( \2855 , \2849 , \2853 , \2854 );
and \U$2667 ( \2856 , \2840 , \2855 );
and \U$2668 ( \2857 , \1104 , \912 );
and \U$2669 ( \2858 , \904 , \910 );
nor \U$2670 ( \2859 , \2857 , \2858 );
xnor \U$2671 ( \2860 , \2859 , \818 );
and \U$2672 ( \2861 , \1299 , \740 );
and \U$2673 ( \2862 , \1194 , \738 );
nor \U$2674 ( \2863 , \2861 , \2862 );
xnor \U$2675 ( \2864 , \2863 , \668 );
and \U$2676 ( \2865 , \2860 , \2864 );
and \U$2677 ( \2866 , \1422 , \604 );
and \U$2678 ( \2867 , \1304 , \602 );
nor \U$2679 ( \2868 , \2866 , \2867 );
xnor \U$2680 ( \2869 , \2868 , \561 );
and \U$2681 ( \2870 , \2864 , \2869 );
and \U$2682 ( \2871 , \2860 , \2869 );
or \U$2683 ( \2872 , \2865 , \2870 , \2871 );
and \U$2684 ( \2873 , \2855 , \2872 );
and \U$2685 ( \2874 , \2840 , \2872 );
or \U$2686 ( \2875 , \2856 , \2873 , \2874 );
and \U$2687 ( \2876 , \593 , \1476 );
and \U$2688 ( \2877 , \495 , \1474 );
nor \U$2689 ( \2878 , \2876 , \2877 );
xnor \U$2690 ( \2879 , \2878 , \1363 );
and \U$2691 ( \2880 , \703 , \1280 );
and \U$2692 ( \2881 , \621 , \1278 );
nor \U$2693 ( \2882 , \2880 , \2881 );
xnor \U$2694 ( \2883 , \2882 , \1177 );
and \U$2695 ( \2884 , \2879 , \2883 );
and \U$2696 ( \2885 , \841 , \1062 );
and \U$2697 ( \2886 , \777 , \1060 );
nor \U$2698 ( \2887 , \2885 , \2886 );
xnor \U$2699 ( \2888 , \2887 , \984 );
and \U$2700 ( \2889 , \2883 , \2888 );
and \U$2701 ( \2890 , \2879 , \2888 );
or \U$2702 ( \2891 , \2884 , \2889 , \2890 );
and \U$2703 ( \2892 , \323 , \2261 );
and \U$2704 ( \2893 , \333 , \2259 );
nor \U$2705 ( \2894 , \2892 , \2893 );
xnor \U$2706 ( \2895 , \2894 , \2124 );
and \U$2707 ( \2896 , \343 , \1955 );
and \U$2708 ( \2897 , \353 , \1953 );
nor \U$2709 ( \2898 , \2896 , \2897 );
xnor \U$2710 ( \2899 , \2898 , \1835 );
and \U$2711 ( \2900 , \2895 , \2899 );
and \U$2712 ( \2901 , \444 , \1742 );
and \U$2713 ( \2902 , \360 , \1740 );
nor \U$2714 ( \2903 , \2901 , \2902 );
xnor \U$2715 ( \2904 , \2903 , \1610 );
and \U$2716 ( \2905 , \2899 , \2904 );
and \U$2717 ( \2906 , \2895 , \2904 );
or \U$2718 ( \2907 , \2900 , \2905 , \2906 );
and \U$2719 ( \2908 , \2891 , \2907 );
_HMUX r123 ( \2909_nR123 , 1'b0 , RIb4bfab0_64 , \287 );
buf \U$2721 ( \2910 , \2909_nR123 );
xor \U$2722 ( \2911 , \2371 , \2910 );
not \U$2723 ( \2912 , \2910 );
and \U$2724 ( \2913 , \2911 , \2912 );
and \U$2725 ( \2914 , \159 , \2913 );
not \U$2726 ( \2915 , \2914 );
xnor \U$2727 ( \2916 , \2915 , \2371 );
and \U$2728 ( \2917 , \305 , \2550 );
and \U$2729 ( \2918 , \315 , \2548 );
nor \U$2730 ( \2919 , \2917 , \2918 );
xnor \U$2731 ( \2920 , \2919 , \2374 );
and \U$2732 ( \2921 , \2916 , \2920 );
and \U$2733 ( \2922 , \2907 , \2921 );
and \U$2734 ( \2923 , \2891 , \2921 );
or \U$2735 ( \2924 , \2908 , \2922 , \2923 );
and \U$2736 ( \2925 , \2875 , \2924 );
xor \U$2737 ( \2926 , \2729 , \2733 );
xor \U$2738 ( \2927 , \2926 , \2738 );
xor \U$2739 ( \2928 , \2745 , \2749 );
xor \U$2740 ( \2929 , \2928 , \2754 );
and \U$2741 ( \2930 , \2927 , \2929 );
xnor \U$2742 ( \2931 , \2762 , \2764 );
and \U$2743 ( \2932 , \2929 , \2931 );
and \U$2744 ( \2933 , \2927 , \2931 );
or \U$2745 ( \2934 , \2930 , \2932 , \2933 );
and \U$2746 ( \2935 , \2924 , \2934 );
and \U$2747 ( \2936 , \2875 , \2934 );
or \U$2748 ( \2937 , \2925 , \2935 , \2936 );
xor \U$2749 ( \2938 , \2680 , \2684 );
xor \U$2750 ( \2939 , \2938 , \2689 );
xor \U$2751 ( \2940 , \2693 , \2697 );
xor \U$2752 ( \2941 , \2940 , \2702 );
and \U$2753 ( \2942 , \2939 , \2941 );
xor \U$2754 ( \2943 , \2710 , \2714 );
xor \U$2755 ( \2944 , \2943 , \2719 );
and \U$2756 ( \2945 , \2941 , \2944 );
and \U$2757 ( \2946 , \2939 , \2944 );
or \U$2758 ( \2947 , \2942 , \2945 , \2946 );
xor \U$2759 ( \2948 , \2783 , \2785 );
xor \U$2760 ( \2949 , \2948 , \2788 );
and \U$2761 ( \2950 , \2947 , \2949 );
xor \U$2762 ( \2951 , \2771 , \2773 );
xor \U$2763 ( \2952 , \2951 , \2775 );
and \U$2764 ( \2953 , \2949 , \2952 );
and \U$2765 ( \2954 , \2947 , \2952 );
or \U$2766 ( \2955 , \2950 , \2953 , \2954 );
and \U$2767 ( \2956 , \2937 , \2955 );
xor \U$2768 ( \2957 , \2522 , \2539 );
xor \U$2769 ( \2958 , \2957 , \2543 );
and \U$2770 ( \2959 , \2955 , \2958 );
and \U$2771 ( \2960 , \2937 , \2958 );
or \U$2772 ( \2961 , \2956 , \2959 , \2960 );
xor \U$2773 ( \2962 , \2565 , \2581 );
xor \U$2774 ( \2963 , \2962 , \2598 );
xor \U$2775 ( \2964 , \2725 , \2768 );
xor \U$2776 ( \2965 , \2964 , \2778 );
and \U$2777 ( \2966 , \2963 , \2965 );
xor \U$2778 ( \2967 , \2791 , \2793 );
xor \U$2779 ( \2968 , \2967 , \2796 );
and \U$2780 ( \2969 , \2965 , \2968 );
and \U$2781 ( \2970 , \2963 , \2968 );
or \U$2782 ( \2971 , \2966 , \2969 , \2970 );
and \U$2783 ( \2972 , \2961 , \2971 );
xor \U$2784 ( \2973 , \2624 , \2626 );
xor \U$2785 ( \2974 , \2973 , \2629 );
and \U$2786 ( \2975 , \2971 , \2974 );
and \U$2787 ( \2976 , \2961 , \2974 );
or \U$2788 ( \2977 , \2972 , \2975 , \2976 );
xor \U$2789 ( \2978 , \2546 , \2601 );
xor \U$2790 ( \2979 , \2978 , \2611 );
xor \U$2791 ( \2980 , \2781 , \2799 );
xor \U$2792 ( \2981 , \2980 , \2802 );
and \U$2793 ( \2982 , \2979 , \2981 );
and \U$2794 ( \2983 , \2977 , \2982 );
xor \U$2795 ( \2984 , \2805 , \2807 );
xor \U$2796 ( \2985 , \2984 , \2810 );
and \U$2797 ( \2986 , \2982 , \2985 );
and \U$2798 ( \2987 , \2977 , \2985 );
or \U$2799 ( \2988 , \2983 , \2986 , \2987 );
and \U$2800 ( \2989 , \2824 , \2988 );
xor \U$2801 ( \2990 , \2824 , \2988 );
xor \U$2802 ( \2991 , \2977 , \2982 );
xor \U$2803 ( \2992 , \2991 , \2985 );
and \U$2804 ( \2993 , \360 , \1955 );
and \U$2805 ( \2994 , \343 , \1953 );
nor \U$2806 ( \2995 , \2993 , \2994 );
xnor \U$2807 ( \2996 , \2995 , \1835 );
and \U$2808 ( \2997 , \495 , \1742 );
and \U$2809 ( \2998 , \444 , \1740 );
nor \U$2810 ( \2999 , \2997 , \2998 );
xnor \U$2811 ( \3000 , \2999 , \1610 );
and \U$2812 ( \3001 , \2996 , \3000 );
and \U$2813 ( \3002 , \621 , \1476 );
and \U$2814 ( \3003 , \593 , \1474 );
nor \U$2815 ( \3004 , \3002 , \3003 );
xnor \U$2816 ( \3005 , \3004 , \1363 );
and \U$2817 ( \3006 , \3000 , \3005 );
and \U$2818 ( \3007 , \2996 , \3005 );
or \U$2819 ( \3008 , \3001 , \3006 , \3007 );
and \U$2820 ( \3009 , \315 , \2913 );
and \U$2821 ( \3010 , \159 , \2910 );
nor \U$2822 ( \3011 , \3009 , \3010 );
xnor \U$2823 ( \3012 , \3011 , \2371 );
and \U$2824 ( \3013 , \333 , \2550 );
and \U$2825 ( \3014 , \305 , \2548 );
nor \U$2826 ( \3015 , \3013 , \3014 );
xnor \U$2827 ( \3016 , \3015 , \2374 );
and \U$2828 ( \3017 , \3012 , \3016 );
and \U$2829 ( \3018 , \353 , \2261 );
and \U$2830 ( \3019 , \323 , \2259 );
nor \U$2831 ( \3020 , \3018 , \3019 );
xnor \U$2832 ( \3021 , \3020 , \2124 );
and \U$2833 ( \3022 , \3016 , \3021 );
and \U$2834 ( \3023 , \3012 , \3021 );
or \U$2835 ( \3024 , \3017 , \3022 , \3023 );
and \U$2836 ( \3025 , \3008 , \3024 );
and \U$2837 ( \3026 , \777 , \1280 );
and \U$2838 ( \3027 , \703 , \1278 );
nor \U$2839 ( \3028 , \3026 , \3027 );
xnor \U$2840 ( \3029 , \3028 , \1177 );
and \U$2841 ( \3030 , \904 , \1062 );
and \U$2842 ( \3031 , \841 , \1060 );
nor \U$2843 ( \3032 , \3030 , \3031 );
xnor \U$2844 ( \3033 , \3032 , \984 );
and \U$2845 ( \3034 , \3029 , \3033 );
and \U$2846 ( \3035 , \1194 , \912 );
and \U$2847 ( \3036 , \1104 , \910 );
nor \U$2848 ( \3037 , \3035 , \3036 );
xnor \U$2849 ( \3038 , \3037 , \818 );
and \U$2850 ( \3039 , \3033 , \3038 );
and \U$2851 ( \3040 , \3029 , \3038 );
or \U$2852 ( \3041 , \3034 , \3039 , \3040 );
and \U$2853 ( \3042 , \3024 , \3041 );
and \U$2854 ( \3043 , \3008 , \3041 );
or \U$2855 ( \3044 , \3025 , \3042 , \3043 );
xor \U$2856 ( \3045 , \2828 , \2832 );
xor \U$2857 ( \3046 , \3045 , \2837 );
xor \U$2858 ( \3047 , \2879 , \2883 );
xor \U$2859 ( \3048 , \3047 , \2888 );
and \U$2860 ( \3049 , \3046 , \3048 );
xor \U$2861 ( \3050 , \2860 , \2864 );
xor \U$2862 ( \3051 , \3050 , \2869 );
and \U$2863 ( \3052 , \3048 , \3051 );
and \U$2864 ( \3053 , \3046 , \3051 );
or \U$2865 ( \3054 , \3049 , \3052 , \3053 );
and \U$2866 ( \3055 , \3044 , \3054 );
and \U$2867 ( \3056 , \1304 , \740 );
and \U$2868 ( \3057 , \1299 , \738 );
nor \U$2869 ( \3058 , \3056 , \3057 );
xnor \U$2870 ( \3059 , \3058 , \668 );
and \U$2871 ( \3060 , \1537 , \604 );
and \U$2872 ( \3061 , \1422 , \602 );
nor \U$2873 ( \3062 , \3060 , \3061 );
xnor \U$2874 ( \3063 , \3062 , \561 );
and \U$2875 ( \3064 , \3059 , \3063 );
and \U$2876 ( \3065 , \1778 , \503 );
and \U$2877 ( \3066 , \1770 , \501 );
nor \U$2878 ( \3067 , \3065 , \3066 );
xnor \U$2879 ( \3068 , \3067 , \455 );
and \U$2880 ( \3069 , \3063 , \3068 );
and \U$2881 ( \3070 , \3059 , \3068 );
or \U$2882 ( \3071 , \3064 , \3069 , \3070 );
and \U$2883 ( \3072 , \2028 , \298 );
and \U$2884 ( \3073 , \2023 , \296 );
nor \U$2885 ( \3074 , \3072 , \3073 );
xnor \U$2886 ( \3075 , \3074 , \303 );
and \U$2887 ( \3076 , \2305 , \313 );
and \U$2888 ( \3077 , \2161 , \311 );
nor \U$2889 ( \3078 , \3076 , \3077 );
xnor \U$2890 ( \3079 , \3078 , \320 );
and \U$2891 ( \3080 , \3075 , \3079 );
and \U$2892 ( \3081 , \2541 , \331 );
and \U$2893 ( \3082 , \2532 , \329 );
nor \U$2894 ( \3083 , \3081 , \3082 );
xnor \U$2895 ( \3084 , \3083 , \338 );
and \U$2896 ( \3085 , \3079 , \3084 );
and \U$2897 ( \3086 , \3075 , \3084 );
or \U$2898 ( \3087 , \3080 , \3085 , \3086 );
and \U$2899 ( \3088 , \3071 , \3087 );
xor \U$2900 ( \3089 , \2844 , \2848 );
xor \U$2901 ( \3090 , \3089 , \2852 );
and \U$2902 ( \3091 , \3087 , \3090 );
and \U$2903 ( \3092 , \3071 , \3090 );
or \U$2904 ( \3093 , \3088 , \3091 , \3092 );
and \U$2905 ( \3094 , \3054 , \3093 );
and \U$2906 ( \3095 , \3044 , \3093 );
or \U$2907 ( \3096 , \3055 , \3094 , \3095 );
xor \U$2908 ( \3097 , \2840 , \2855 );
xor \U$2909 ( \3098 , \3097 , \2872 );
xor \U$2910 ( \3099 , \2939 , \2941 );
xor \U$2911 ( \3100 , \3099 , \2944 );
and \U$2912 ( \3101 , \3098 , \3100 );
xor \U$2913 ( \3102 , \2927 , \2929 );
xor \U$2914 ( \3103 , \3102 , \2931 );
and \U$2915 ( \3104 , \3100 , \3103 );
and \U$2916 ( \3105 , \3098 , \3103 );
or \U$2917 ( \3106 , \3101 , \3104 , \3105 );
and \U$2918 ( \3107 , \3096 , \3106 );
xor \U$2919 ( \3108 , \2741 , \2757 );
xor \U$2920 ( \3109 , \3108 , \2765 );
and \U$2921 ( \3110 , \3106 , \3109 );
and \U$2922 ( \3111 , \3096 , \3109 );
or \U$2923 ( \3112 , \3107 , \3110 , \3111 );
xor \U$2924 ( \3113 , \2692 , \2705 );
xor \U$2925 ( \3114 , \3113 , \2722 );
xor \U$2926 ( \3115 , \2875 , \2924 );
xor \U$2927 ( \3116 , \3115 , \2934 );
and \U$2928 ( \3117 , \3114 , \3116 );
xor \U$2929 ( \3118 , \2947 , \2949 );
xor \U$2930 ( \3119 , \3118 , \2952 );
and \U$2931 ( \3120 , \3116 , \3119 );
and \U$2932 ( \3121 , \3114 , \3119 );
or \U$2933 ( \3122 , \3117 , \3120 , \3121 );
and \U$2934 ( \3123 , \3112 , \3122 );
xor \U$2935 ( \3124 , \2963 , \2965 );
xor \U$2936 ( \3125 , \3124 , \2968 );
and \U$2937 ( \3126 , \3122 , \3125 );
and \U$2938 ( \3127 , \3112 , \3125 );
or \U$2939 ( \3128 , \3123 , \3126 , \3127 );
xor \U$2940 ( \3129 , \2961 , \2971 );
xor \U$2941 ( \3130 , \3129 , \2974 );
and \U$2942 ( \3131 , \3128 , \3130 );
xor \U$2943 ( \3132 , \2979 , \2981 );
and \U$2944 ( \3133 , \3130 , \3132 );
and \U$2945 ( \3134 , \3128 , \3132 );
or \U$2946 ( \3135 , \3131 , \3133 , \3134 );
and \U$2947 ( \3136 , \2992 , \3135 );
xor \U$2948 ( \3137 , \2992 , \3135 );
xor \U$2949 ( \3138 , \3128 , \3130 );
xor \U$2950 ( \3139 , \3138 , \3132 );
and \U$2951 ( \3140 , \343 , \2261 );
and \U$2952 ( \3141 , \353 , \2259 );
nor \U$2953 ( \3142 , \3140 , \3141 );
xnor \U$2954 ( \3143 , \3142 , \2124 );
and \U$2955 ( \3144 , \444 , \1955 );
and \U$2956 ( \3145 , \360 , \1953 );
nor \U$2957 ( \3146 , \3144 , \3145 );
xnor \U$2958 ( \3147 , \3146 , \1835 );
and \U$2959 ( \3148 , \3143 , \3147 );
and \U$2960 ( \3149 , \593 , \1742 );
and \U$2961 ( \3150 , \495 , \1740 );
nor \U$2962 ( \3151 , \3149 , \3150 );
xnor \U$2963 ( \3152 , \3151 , \1610 );
and \U$2964 ( \3153 , \3147 , \3152 );
and \U$2965 ( \3154 , \3143 , \3152 );
or \U$2966 ( \3155 , \3148 , \3153 , \3154 );
and \U$2967 ( \3156 , \703 , \1476 );
and \U$2968 ( \3157 , \621 , \1474 );
nor \U$2969 ( \3158 , \3156 , \3157 );
xnor \U$2970 ( \3159 , \3158 , \1363 );
and \U$2971 ( \3160 , \841 , \1280 );
and \U$2972 ( \3161 , \777 , \1278 );
nor \U$2973 ( \3162 , \3160 , \3161 );
xnor \U$2974 ( \3163 , \3162 , \1177 );
and \U$2975 ( \3164 , \3159 , \3163 );
and \U$2976 ( \3165 , \1104 , \1062 );
and \U$2977 ( \3166 , \904 , \1060 );
nor \U$2978 ( \3167 , \3165 , \3166 );
xnor \U$2979 ( \3168 , \3167 , \984 );
and \U$2980 ( \3169 , \3163 , \3168 );
and \U$2981 ( \3170 , \3159 , \3168 );
or \U$2982 ( \3171 , \3164 , \3169 , \3170 );
and \U$2983 ( \3172 , \3155 , \3171 );
and \U$2984 ( \3173 , \305 , \2913 );
and \U$2985 ( \3174 , \315 , \2910 );
nor \U$2986 ( \3175 , \3173 , \3174 );
xnor \U$2987 ( \3176 , \3175 , \2371 );
and \U$2988 ( \3177 , \323 , \2550 );
and \U$2989 ( \3178 , \333 , \2548 );
nor \U$2990 ( \3179 , \3177 , \3178 );
xnor \U$2991 ( \3180 , \3179 , \2374 );
and \U$2992 ( \3181 , \3176 , \3180 );
and \U$2993 ( \3182 , \3180 , \358 );
and \U$2994 ( \3183 , \3176 , \358 );
or \U$2995 ( \3184 , \3181 , \3182 , \3183 );
and \U$2996 ( \3185 , \3171 , \3184 );
and \U$2997 ( \3186 , \3155 , \3184 );
or \U$2998 ( \3187 , \3172 , \3185 , \3186 );
and \U$2999 ( \3188 , \2023 , \503 );
and \U$3000 ( \3189 , \1778 , \501 );
nor \U$3001 ( \3190 , \3188 , \3189 );
xnor \U$3002 ( \3191 , \3190 , \455 );
and \U$3003 ( \3192 , \2161 , \298 );
and \U$3004 ( \3193 , \2028 , \296 );
nor \U$3005 ( \3194 , \3192 , \3193 );
xnor \U$3006 ( \3195 , \3194 , \303 );
and \U$3007 ( \3196 , \3191 , \3195 );
and \U$3008 ( \3197 , \2532 , \313 );
and \U$3009 ( \3198 , \2305 , \311 );
nor \U$3010 ( \3199 , \3197 , \3198 );
xnor \U$3011 ( \3200 , \3199 , \320 );
and \U$3012 ( \3201 , \3195 , \3200 );
and \U$3013 ( \3202 , \3191 , \3200 );
or \U$3014 ( \3203 , \3196 , \3201 , \3202 );
and \U$3015 ( \3204 , \1299 , \912 );
and \U$3016 ( \3205 , \1194 , \910 );
nor \U$3017 ( \3206 , \3204 , \3205 );
xnor \U$3018 ( \3207 , \3206 , \818 );
and \U$3019 ( \3208 , \1422 , \740 );
and \U$3020 ( \3209 , \1304 , \738 );
nor \U$3021 ( \3210 , \3208 , \3209 );
xnor \U$3022 ( \3211 , \3210 , \668 );
and \U$3023 ( \3212 , \3207 , \3211 );
and \U$3024 ( \3213 , \1770 , \604 );
and \U$3025 ( \3214 , \1537 , \602 );
nor \U$3026 ( \3215 , \3213 , \3214 );
xnor \U$3027 ( \3216 , \3215 , \561 );
and \U$3028 ( \3217 , \3211 , \3216 );
and \U$3029 ( \3218 , \3207 , \3216 );
or \U$3030 ( \3219 , \3212 , \3217 , \3218 );
and \U$3031 ( \3220 , \3203 , \3219 );
and \U$3032 ( \3221 , \2850 , \351 );
and \U$3033 ( \3222 , \2763 , \349 );
nor \U$3034 ( \3223 , \3221 , \3222 );
xnor \U$3035 ( \3224 , \3223 , \358 );
and \U$3036 ( \3225 , \3219 , \3224 );
and \U$3037 ( \3226 , \3203 , \3224 );
or \U$3038 ( \3227 , \3220 , \3225 , \3226 );
and \U$3039 ( \3228 , \3187 , \3227 );
xor \U$3040 ( \3229 , \3059 , \3063 );
xor \U$3041 ( \3230 , \3229 , \3068 );
xor \U$3042 ( \3231 , \3075 , \3079 );
xor \U$3043 ( \3232 , \3231 , \3084 );
and \U$3044 ( \3233 , \3230 , \3232 );
xor \U$3045 ( \3234 , \3029 , \3033 );
xor \U$3046 ( \3235 , \3234 , \3038 );
and \U$3047 ( \3236 , \3232 , \3235 );
and \U$3048 ( \3237 , \3230 , \3235 );
or \U$3049 ( \3238 , \3233 , \3236 , \3237 );
and \U$3050 ( \3239 , \3227 , \3238 );
and \U$3051 ( \3240 , \3187 , \3238 );
or \U$3052 ( \3241 , \3228 , \3239 , \3240 );
xor \U$3053 ( \3242 , \2895 , \2899 );
xor \U$3054 ( \3243 , \3242 , \2904 );
xor \U$3055 ( \3244 , \3046 , \3048 );
xor \U$3056 ( \3245 , \3244 , \3051 );
and \U$3057 ( \3246 , \3243 , \3245 );
xor \U$3058 ( \3247 , \2916 , \2920 );
and \U$3059 ( \3248 , \3245 , \3247 );
and \U$3060 ( \3249 , \3243 , \3247 );
or \U$3061 ( \3250 , \3246 , \3248 , \3249 );
and \U$3062 ( \3251 , \3241 , \3250 );
xor \U$3063 ( \3252 , \3008 , \3024 );
xor \U$3064 ( \3253 , \3252 , \3041 );
xor \U$3065 ( \3254 , \3071 , \3087 );
xor \U$3066 ( \3255 , \3254 , \3090 );
and \U$3067 ( \3256 , \3253 , \3255 );
and \U$3068 ( \3257 , \3250 , \3256 );
and \U$3069 ( \3258 , \3241 , \3256 );
or \U$3070 ( \3259 , \3251 , \3257 , \3258 );
xor \U$3071 ( \3260 , \2891 , \2907 );
xor \U$3072 ( \3261 , \3260 , \2921 );
xor \U$3073 ( \3262 , \3044 , \3054 );
xor \U$3074 ( \3263 , \3262 , \3093 );
and \U$3075 ( \3264 , \3261 , \3263 );
xor \U$3076 ( \3265 , \3098 , \3100 );
xor \U$3077 ( \3266 , \3265 , \3103 );
and \U$3078 ( \3267 , \3263 , \3266 );
and \U$3079 ( \3268 , \3261 , \3266 );
or \U$3080 ( \3269 , \3264 , \3267 , \3268 );
and \U$3081 ( \3270 , \3259 , \3269 );
xor \U$3082 ( \3271 , \3114 , \3116 );
xor \U$3083 ( \3272 , \3271 , \3119 );
and \U$3084 ( \3273 , \3269 , \3272 );
and \U$3085 ( \3274 , \3259 , \3272 );
or \U$3086 ( \3275 , \3270 , \3273 , \3274 );
xor \U$3087 ( \3276 , \2937 , \2955 );
xor \U$3088 ( \3277 , \3276 , \2958 );
and \U$3089 ( \3278 , \3275 , \3277 );
xor \U$3090 ( \3279 , \3112 , \3122 );
xor \U$3091 ( \3280 , \3279 , \3125 );
and \U$3092 ( \3281 , \3277 , \3280 );
and \U$3093 ( \3282 , \3275 , \3280 );
or \U$3094 ( \3283 , \3278 , \3281 , \3282 );
and \U$3095 ( \3284 , \3139 , \3283 );
xor \U$3096 ( \3285 , \3139 , \3283 );
xor \U$3097 ( \3286 , \3275 , \3277 );
xor \U$3098 ( \3287 , \3286 , \3280 );
and \U$3099 ( \3288 , \904 , \1280 );
and \U$3100 ( \3289 , \841 , \1278 );
nor \U$3101 ( \3290 , \3288 , \3289 );
xnor \U$3102 ( \3291 , \3290 , \1177 );
and \U$3103 ( \3292 , \1194 , \1062 );
and \U$3104 ( \3293 , \1104 , \1060 );
nor \U$3105 ( \3294 , \3292 , \3293 );
xnor \U$3106 ( \3295 , \3294 , \984 );
and \U$3107 ( \3296 , \3291 , \3295 );
and \U$3108 ( \3297 , \1304 , \912 );
and \U$3109 ( \3298 , \1299 , \910 );
nor \U$3110 ( \3299 , \3297 , \3298 );
xnor \U$3111 ( \3300 , \3299 , \818 );
and \U$3112 ( \3301 , \3295 , \3300 );
and \U$3113 ( \3302 , \3291 , \3300 );
or \U$3114 ( \3303 , \3296 , \3301 , \3302 );
and \U$3115 ( \3304 , \495 , \1955 );
and \U$3116 ( \3305 , \444 , \1953 );
nor \U$3117 ( \3306 , \3304 , \3305 );
xnor \U$3118 ( \3307 , \3306 , \1835 );
and \U$3119 ( \3308 , \621 , \1742 );
and \U$3120 ( \3309 , \593 , \1740 );
nor \U$3121 ( \3310 , \3308 , \3309 );
xnor \U$3122 ( \3311 , \3310 , \1610 );
and \U$3123 ( \3312 , \3307 , \3311 );
and \U$3124 ( \3313 , \777 , \1476 );
and \U$3125 ( \3314 , \703 , \1474 );
nor \U$3126 ( \3315 , \3313 , \3314 );
xnor \U$3127 ( \3316 , \3315 , \1363 );
and \U$3128 ( \3317 , \3311 , \3316 );
and \U$3129 ( \3318 , \3307 , \3316 );
or \U$3130 ( \3319 , \3312 , \3317 , \3318 );
and \U$3131 ( \3320 , \3303 , \3319 );
and \U$3132 ( \3321 , \333 , \2913 );
and \U$3133 ( \3322 , \305 , \2910 );
nor \U$3134 ( \3323 , \3321 , \3322 );
xnor \U$3135 ( \3324 , \3323 , \2371 );
and \U$3136 ( \3325 , \353 , \2550 );
and \U$3137 ( \3326 , \323 , \2548 );
nor \U$3138 ( \3327 , \3325 , \3326 );
xnor \U$3139 ( \3328 , \3327 , \2374 );
and \U$3140 ( \3329 , \3324 , \3328 );
and \U$3141 ( \3330 , \360 , \2261 );
and \U$3142 ( \3331 , \343 , \2259 );
nor \U$3143 ( \3332 , \3330 , \3331 );
xnor \U$3144 ( \3333 , \3332 , \2124 );
and \U$3145 ( \3334 , \3328 , \3333 );
and \U$3146 ( \3335 , \3324 , \3333 );
or \U$3147 ( \3336 , \3329 , \3334 , \3335 );
and \U$3148 ( \3337 , \3319 , \3336 );
and \U$3149 ( \3338 , \3303 , \3336 );
or \U$3150 ( \3339 , \3320 , \3337 , \3338 );
and \U$3151 ( \3340 , \2305 , \298 );
and \U$3152 ( \3341 , \2161 , \296 );
nor \U$3153 ( \3342 , \3340 , \3341 );
xnor \U$3154 ( \3343 , \3342 , \303 );
and \U$3155 ( \3344 , \2541 , \313 );
and \U$3156 ( \3345 , \2532 , \311 );
nor \U$3157 ( \3346 , \3344 , \3345 );
xnor \U$3158 ( \3347 , \3346 , \320 );
and \U$3159 ( \3348 , \3343 , \3347 );
and \U$3160 ( \3349 , \2850 , \331 );
and \U$3161 ( \3350 , \2763 , \329 );
nor \U$3162 ( \3351 , \3349 , \3350 );
xnor \U$3163 ( \3352 , \3351 , \338 );
and \U$3164 ( \3353 , \3347 , \3352 );
and \U$3165 ( \3354 , \3343 , \3352 );
or \U$3166 ( \3355 , \3348 , \3353 , \3354 );
and \U$3167 ( \3356 , \1537 , \740 );
and \U$3168 ( \3357 , \1422 , \738 );
nor \U$3169 ( \3358 , \3356 , \3357 );
xnor \U$3170 ( \3359 , \3358 , \668 );
and \U$3171 ( \3360 , \1778 , \604 );
and \U$3172 ( \3361 , \1770 , \602 );
nor \U$3173 ( \3362 , \3360 , \3361 );
xnor \U$3174 ( \3363 , \3362 , \561 );
and \U$3175 ( \3364 , \3359 , \3363 );
and \U$3176 ( \3365 , \2028 , \503 );
and \U$3177 ( \3366 , \2023 , \501 );
nor \U$3178 ( \3367 , \3365 , \3366 );
xnor \U$3179 ( \3368 , \3367 , \455 );
and \U$3180 ( \3369 , \3363 , \3368 );
and \U$3181 ( \3370 , \3359 , \3368 );
or \U$3182 ( \3371 , \3364 , \3369 , \3370 );
and \U$3183 ( \3372 , \3355 , \3371 );
and \U$3184 ( \3373 , \2763 , \331 );
and \U$3185 ( \3374 , \2541 , \329 );
nor \U$3186 ( \3375 , \3373 , \3374 );
xnor \U$3187 ( \3376 , \3375 , \338 );
and \U$3188 ( \3377 , \3371 , \3376 );
and \U$3189 ( \3378 , \3355 , \3376 );
or \U$3190 ( \3379 , \3372 , \3377 , \3378 );
and \U$3191 ( \3380 , \3339 , \3379 );
nand \U$3192 ( \3381 , \2850 , \349 );
xnor \U$3193 ( \3382 , \3381 , \358 );
xor \U$3194 ( \3383 , \3191 , \3195 );
xor \U$3195 ( \3384 , \3383 , \3200 );
and \U$3196 ( \3385 , \3382 , \3384 );
xor \U$3197 ( \3386 , \3207 , \3211 );
xor \U$3198 ( \3387 , \3386 , \3216 );
and \U$3199 ( \3388 , \3384 , \3387 );
and \U$3200 ( \3389 , \3382 , \3387 );
or \U$3201 ( \3390 , \3385 , \3388 , \3389 );
and \U$3202 ( \3391 , \3379 , \3390 );
and \U$3203 ( \3392 , \3339 , \3390 );
or \U$3204 ( \3393 , \3380 , \3391 , \3392 );
xor \U$3205 ( \3394 , \3143 , \3147 );
xor \U$3206 ( \3395 , \3394 , \3152 );
xor \U$3207 ( \3396 , \3159 , \3163 );
xor \U$3208 ( \3397 , \3396 , \3168 );
and \U$3209 ( \3398 , \3395 , \3397 );
xor \U$3210 ( \3399 , \3176 , \3180 );
xor \U$3211 ( \3400 , \3399 , \358 );
and \U$3212 ( \3401 , \3397 , \3400 );
and \U$3213 ( \3402 , \3395 , \3400 );
or \U$3214 ( \3403 , \3398 , \3401 , \3402 );
xor \U$3215 ( \3404 , \2996 , \3000 );
xor \U$3216 ( \3405 , \3404 , \3005 );
and \U$3217 ( \3406 , \3403 , \3405 );
xor \U$3218 ( \3407 , \3012 , \3016 );
xor \U$3219 ( \3408 , \3407 , \3021 );
and \U$3220 ( \3409 , \3405 , \3408 );
and \U$3221 ( \3410 , \3403 , \3408 );
or \U$3222 ( \3411 , \3406 , \3409 , \3410 );
and \U$3223 ( \3412 , \3393 , \3411 );
xor \U$3224 ( \3413 , \3155 , \3171 );
xor \U$3225 ( \3414 , \3413 , \3184 );
xor \U$3226 ( \3415 , \3203 , \3219 );
xor \U$3227 ( \3416 , \3415 , \3224 );
and \U$3228 ( \3417 , \3414 , \3416 );
xor \U$3229 ( \3418 , \3230 , \3232 );
xor \U$3230 ( \3419 , \3418 , \3235 );
and \U$3231 ( \3420 , \3416 , \3419 );
and \U$3232 ( \3421 , \3414 , \3419 );
or \U$3233 ( \3422 , \3417 , \3420 , \3421 );
and \U$3234 ( \3423 , \3411 , \3422 );
and \U$3235 ( \3424 , \3393 , \3422 );
or \U$3236 ( \3425 , \3412 , \3423 , \3424 );
xor \U$3237 ( \3426 , \3187 , \3227 );
xor \U$3238 ( \3427 , \3426 , \3238 );
xor \U$3239 ( \3428 , \3243 , \3245 );
xor \U$3240 ( \3429 , \3428 , \3247 );
and \U$3241 ( \3430 , \3427 , \3429 );
xor \U$3242 ( \3431 , \3253 , \3255 );
and \U$3243 ( \3432 , \3429 , \3431 );
and \U$3244 ( \3433 , \3427 , \3431 );
or \U$3245 ( \3434 , \3430 , \3432 , \3433 );
and \U$3246 ( \3435 , \3425 , \3434 );
xor \U$3247 ( \3436 , \3261 , \3263 );
xor \U$3248 ( \3437 , \3436 , \3266 );
and \U$3249 ( \3438 , \3434 , \3437 );
and \U$3250 ( \3439 , \3425 , \3437 );
or \U$3251 ( \3440 , \3435 , \3438 , \3439 );
xor \U$3252 ( \3441 , \3096 , \3106 );
xor \U$3253 ( \3442 , \3441 , \3109 );
and \U$3254 ( \3443 , \3440 , \3442 );
xor \U$3255 ( \3444 , \3259 , \3269 );
xor \U$3256 ( \3445 , \3444 , \3272 );
and \U$3257 ( \3446 , \3442 , \3445 );
and \U$3258 ( \3447 , \3440 , \3445 );
or \U$3259 ( \3448 , \3443 , \3446 , \3447 );
and \U$3260 ( \3449 , \3287 , \3448 );
xor \U$3261 ( \3450 , \3287 , \3448 );
xor \U$3262 ( \3451 , \3440 , \3442 );
xor \U$3263 ( \3452 , \3451 , \3445 );
and \U$3264 ( \3453 , \841 , \1476 );
and \U$3265 ( \3454 , \777 , \1474 );
nor \U$3266 ( \3455 , \3453 , \3454 );
xnor \U$3267 ( \3456 , \3455 , \1363 );
and \U$3268 ( \3457 , \1104 , \1280 );
and \U$3269 ( \3458 , \904 , \1278 );
nor \U$3270 ( \3459 , \3457 , \3458 );
xnor \U$3271 ( \3460 , \3459 , \1177 );
and \U$3272 ( \3461 , \3456 , \3460 );
and \U$3273 ( \3462 , \1299 , \1062 );
and \U$3274 ( \3463 , \1194 , \1060 );
nor \U$3275 ( \3464 , \3462 , \3463 );
xnor \U$3276 ( \3465 , \3464 , \984 );
and \U$3277 ( \3466 , \3460 , \3465 );
and \U$3278 ( \3467 , \3456 , \3465 );
or \U$3279 ( \3468 , \3461 , \3466 , \3467 );
and \U$3280 ( \3469 , \444 , \2261 );
and \U$3281 ( \3470 , \360 , \2259 );
nor \U$3282 ( \3471 , \3469 , \3470 );
xnor \U$3283 ( \3472 , \3471 , \2124 );
and \U$3284 ( \3473 , \593 , \1955 );
and \U$3285 ( \3474 , \495 , \1953 );
nor \U$3286 ( \3475 , \3473 , \3474 );
xnor \U$3287 ( \3476 , \3475 , \1835 );
and \U$3288 ( \3477 , \3472 , \3476 );
and \U$3289 ( \3478 , \703 , \1742 );
and \U$3290 ( \3479 , \621 , \1740 );
nor \U$3291 ( \3480 , \3478 , \3479 );
xnor \U$3292 ( \3481 , \3480 , \1610 );
and \U$3293 ( \3482 , \3476 , \3481 );
and \U$3294 ( \3483 , \3472 , \3481 );
or \U$3295 ( \3484 , \3477 , \3482 , \3483 );
and \U$3296 ( \3485 , \3468 , \3484 );
and \U$3297 ( \3486 , \323 , \2913 );
and \U$3298 ( \3487 , \333 , \2910 );
nor \U$3299 ( \3488 , \3486 , \3487 );
xnor \U$3300 ( \3489 , \3488 , \2371 );
and \U$3301 ( \3490 , \343 , \2550 );
and \U$3302 ( \3491 , \353 , \2548 );
nor \U$3303 ( \3492 , \3490 , \3491 );
xnor \U$3304 ( \3493 , \3492 , \2374 );
and \U$3305 ( \3494 , \3489 , \3493 );
and \U$3306 ( \3495 , \3493 , \338 );
and \U$3307 ( \3496 , \3489 , \338 );
or \U$3308 ( \3497 , \3494 , \3495 , \3496 );
and \U$3309 ( \3498 , \3484 , \3497 );
and \U$3310 ( \3499 , \3468 , \3497 );
or \U$3311 ( \3500 , \3485 , \3498 , \3499 );
and \U$3312 ( \3501 , \1422 , \912 );
and \U$3313 ( \3502 , \1304 , \910 );
nor \U$3314 ( \3503 , \3501 , \3502 );
xnor \U$3315 ( \3504 , \3503 , \818 );
and \U$3316 ( \3505 , \1770 , \740 );
and \U$3317 ( \3506 , \1537 , \738 );
nor \U$3318 ( \3507 , \3505 , \3506 );
xnor \U$3319 ( \3508 , \3507 , \668 );
and \U$3320 ( \3509 , \3504 , \3508 );
and \U$3321 ( \3510 , \2023 , \604 );
and \U$3322 ( \3511 , \1778 , \602 );
nor \U$3323 ( \3512 , \3510 , \3511 );
xnor \U$3324 ( \3513 , \3512 , \561 );
and \U$3325 ( \3514 , \3508 , \3513 );
and \U$3326 ( \3515 , \3504 , \3513 );
or \U$3327 ( \3516 , \3509 , \3514 , \3515 );
and \U$3328 ( \3517 , \2161 , \503 );
and \U$3329 ( \3518 , \2028 , \501 );
nor \U$3330 ( \3519 , \3517 , \3518 );
xnor \U$3331 ( \3520 , \3519 , \455 );
and \U$3332 ( \3521 , \2532 , \298 );
and \U$3333 ( \3522 , \2305 , \296 );
nor \U$3334 ( \3523 , \3521 , \3522 );
xnor \U$3335 ( \3524 , \3523 , \303 );
and \U$3336 ( \3525 , \3520 , \3524 );
and \U$3337 ( \3526 , \2763 , \313 );
and \U$3338 ( \3527 , \2541 , \311 );
nor \U$3339 ( \3528 , \3526 , \3527 );
xnor \U$3340 ( \3529 , \3528 , \320 );
and \U$3341 ( \3530 , \3524 , \3529 );
and \U$3342 ( \3531 , \3520 , \3529 );
or \U$3343 ( \3532 , \3525 , \3530 , \3531 );
and \U$3344 ( \3533 , \3516 , \3532 );
xor \U$3345 ( \3534 , \3343 , \3347 );
xor \U$3346 ( \3535 , \3534 , \3352 );
and \U$3347 ( \3536 , \3532 , \3535 );
and \U$3348 ( \3537 , \3516 , \3535 );
or \U$3349 ( \3538 , \3533 , \3536 , \3537 );
and \U$3350 ( \3539 , \3500 , \3538 );
xor \U$3351 ( \3540 , \3291 , \3295 );
xor \U$3352 ( \3541 , \3540 , \3300 );
xor \U$3353 ( \3542 , \3307 , \3311 );
xor \U$3354 ( \3543 , \3542 , \3316 );
and \U$3355 ( \3544 , \3541 , \3543 );
xor \U$3356 ( \3545 , \3359 , \3363 );
xor \U$3357 ( \3546 , \3545 , \3368 );
and \U$3358 ( \3547 , \3543 , \3546 );
and \U$3359 ( \3548 , \3541 , \3546 );
or \U$3360 ( \3549 , \3544 , \3547 , \3548 );
and \U$3361 ( \3550 , \3538 , \3549 );
and \U$3362 ( \3551 , \3500 , \3549 );
or \U$3363 ( \3552 , \3539 , \3550 , \3551 );
xor \U$3364 ( \3553 , \3355 , \3371 );
xor \U$3365 ( \3554 , \3553 , \3376 );
xor \U$3366 ( \3555 , \3395 , \3397 );
xor \U$3367 ( \3556 , \3555 , \3400 );
and \U$3368 ( \3557 , \3554 , \3556 );
xor \U$3369 ( \3558 , \3382 , \3384 );
xor \U$3370 ( \3559 , \3558 , \3387 );
and \U$3371 ( \3560 , \3556 , \3559 );
and \U$3372 ( \3561 , \3554 , \3559 );
or \U$3373 ( \3562 , \3557 , \3560 , \3561 );
and \U$3374 ( \3563 , \3552 , \3562 );
xor \U$3375 ( \3564 , \3414 , \3416 );
xor \U$3376 ( \3565 , \3564 , \3419 );
and \U$3377 ( \3566 , \3562 , \3565 );
and \U$3378 ( \3567 , \3552 , \3565 );
or \U$3379 ( \3568 , \3563 , \3566 , \3567 );
xor \U$3380 ( \3569 , \3339 , \3379 );
xor \U$3381 ( \3570 , \3569 , \3390 );
xor \U$3382 ( \3571 , \3403 , \3405 );
xor \U$3383 ( \3572 , \3571 , \3408 );
and \U$3384 ( \3573 , \3570 , \3572 );
and \U$3385 ( \3574 , \3568 , \3573 );
xor \U$3386 ( \3575 , \3427 , \3429 );
xor \U$3387 ( \3576 , \3575 , \3431 );
and \U$3388 ( \3577 , \3573 , \3576 );
and \U$3389 ( \3578 , \3568 , \3576 );
or \U$3390 ( \3579 , \3574 , \3577 , \3578 );
xor \U$3391 ( \3580 , \3241 , \3250 );
xor \U$3392 ( \3581 , \3580 , \3256 );
and \U$3393 ( \3582 , \3579 , \3581 );
xor \U$3394 ( \3583 , \3425 , \3434 );
xor \U$3395 ( \3584 , \3583 , \3437 );
and \U$3396 ( \3585 , \3581 , \3584 );
and \U$3397 ( \3586 , \3579 , \3584 );
or \U$3398 ( \3587 , \3582 , \3585 , \3586 );
and \U$3399 ( \3588 , \3452 , \3587 );
xor \U$3400 ( \3589 , \3452 , \3587 );
xor \U$3401 ( \3590 , \3579 , \3581 );
xor \U$3402 ( \3591 , \3590 , \3584 );
and \U$3403 ( \3592 , \353 , \2913 );
and \U$3404 ( \3593 , \323 , \2910 );
nor \U$3405 ( \3594 , \3592 , \3593 );
xnor \U$3406 ( \3595 , \3594 , \2371 );
and \U$3407 ( \3596 , \360 , \2550 );
and \U$3408 ( \3597 , \343 , \2548 );
nor \U$3409 ( \3598 , \3596 , \3597 );
xnor \U$3410 ( \3599 , \3598 , \2374 );
and \U$3411 ( \3600 , \3595 , \3599 );
and \U$3412 ( \3601 , \495 , \2261 );
and \U$3413 ( \3602 , \444 , \2259 );
nor \U$3414 ( \3603 , \3601 , \3602 );
xnor \U$3415 ( \3604 , \3603 , \2124 );
and \U$3416 ( \3605 , \3599 , \3604 );
and \U$3417 ( \3606 , \3595 , \3604 );
or \U$3418 ( \3607 , \3600 , \3605 , \3606 );
and \U$3419 ( \3608 , \1194 , \1280 );
and \U$3420 ( \3609 , \1104 , \1278 );
nor \U$3421 ( \3610 , \3608 , \3609 );
xnor \U$3422 ( \3611 , \3610 , \1177 );
and \U$3423 ( \3612 , \1304 , \1062 );
and \U$3424 ( \3613 , \1299 , \1060 );
nor \U$3425 ( \3614 , \3612 , \3613 );
xnor \U$3426 ( \3615 , \3614 , \984 );
and \U$3427 ( \3616 , \3611 , \3615 );
and \U$3428 ( \3617 , \1537 , \912 );
and \U$3429 ( \3618 , \1422 , \910 );
nor \U$3430 ( \3619 , \3617 , \3618 );
xnor \U$3431 ( \3620 , \3619 , \818 );
and \U$3432 ( \3621 , \3615 , \3620 );
and \U$3433 ( \3622 , \3611 , \3620 );
or \U$3434 ( \3623 , \3616 , \3621 , \3622 );
and \U$3435 ( \3624 , \3607 , \3623 );
and \U$3436 ( \3625 , \621 , \1955 );
and \U$3437 ( \3626 , \593 , \1953 );
nor \U$3438 ( \3627 , \3625 , \3626 );
xnor \U$3439 ( \3628 , \3627 , \1835 );
and \U$3440 ( \3629 , \777 , \1742 );
and \U$3441 ( \3630 , \703 , \1740 );
nor \U$3442 ( \3631 , \3629 , \3630 );
xnor \U$3443 ( \3632 , \3631 , \1610 );
and \U$3444 ( \3633 , \3628 , \3632 );
and \U$3445 ( \3634 , \904 , \1476 );
and \U$3446 ( \3635 , \841 , \1474 );
nor \U$3447 ( \3636 , \3634 , \3635 );
xnor \U$3448 ( \3637 , \3636 , \1363 );
and \U$3449 ( \3638 , \3632 , \3637 );
and \U$3450 ( \3639 , \3628 , \3637 );
or \U$3451 ( \3640 , \3633 , \3638 , \3639 );
and \U$3452 ( \3641 , \3623 , \3640 );
and \U$3453 ( \3642 , \3607 , \3640 );
or \U$3454 ( \3643 , \3624 , \3641 , \3642 );
xor \U$3455 ( \3644 , \3456 , \3460 );
xor \U$3456 ( \3645 , \3644 , \3465 );
xor \U$3457 ( \3646 , \3472 , \3476 );
xor \U$3458 ( \3647 , \3646 , \3481 );
and \U$3459 ( \3648 , \3645 , \3647 );
xor \U$3460 ( \3649 , \3504 , \3508 );
xor \U$3461 ( \3650 , \3649 , \3513 );
and \U$3462 ( \3651 , \3647 , \3650 );
and \U$3463 ( \3652 , \3645 , \3650 );
or \U$3464 ( \3653 , \3648 , \3651 , \3652 );
and \U$3465 ( \3654 , \3643 , \3653 );
and \U$3466 ( \3655 , \1778 , \740 );
and \U$3467 ( \3656 , \1770 , \738 );
nor \U$3468 ( \3657 , \3655 , \3656 );
xnor \U$3469 ( \3658 , \3657 , \668 );
and \U$3470 ( \3659 , \2028 , \604 );
and \U$3471 ( \3660 , \2023 , \602 );
nor \U$3472 ( \3661 , \3659 , \3660 );
xnor \U$3473 ( \3662 , \3661 , \561 );
and \U$3474 ( \3663 , \3658 , \3662 );
and \U$3475 ( \3664 , \2305 , \503 );
and \U$3476 ( \3665 , \2161 , \501 );
nor \U$3477 ( \3666 , \3664 , \3665 );
xnor \U$3478 ( \3667 , \3666 , \455 );
and \U$3479 ( \3668 , \3662 , \3667 );
and \U$3480 ( \3669 , \3658 , \3667 );
or \U$3481 ( \3670 , \3663 , \3668 , \3669 );
nand \U$3482 ( \3671 , \2850 , \329 );
xnor \U$3483 ( \3672 , \3671 , \338 );
and \U$3484 ( \3673 , \3670 , \3672 );
xor \U$3485 ( \3674 , \3520 , \3524 );
xor \U$3486 ( \3675 , \3674 , \3529 );
and \U$3487 ( \3676 , \3672 , \3675 );
and \U$3488 ( \3677 , \3670 , \3675 );
or \U$3489 ( \3678 , \3673 , \3676 , \3677 );
and \U$3490 ( \3679 , \3653 , \3678 );
and \U$3491 ( \3680 , \3643 , \3678 );
or \U$3492 ( \3681 , \3654 , \3679 , \3680 );
xor \U$3493 ( \3682 , \3324 , \3328 );
xor \U$3494 ( \3683 , \3682 , \3333 );
xor \U$3495 ( \3684 , \3516 , \3532 );
xor \U$3496 ( \3685 , \3684 , \3535 );
and \U$3497 ( \3686 , \3683 , \3685 );
xor \U$3498 ( \3687 , \3541 , \3543 );
xor \U$3499 ( \3688 , \3687 , \3546 );
and \U$3500 ( \3689 , \3685 , \3688 );
and \U$3501 ( \3690 , \3683 , \3688 );
or \U$3502 ( \3691 , \3686 , \3689 , \3690 );
and \U$3503 ( \3692 , \3681 , \3691 );
xor \U$3504 ( \3693 , \3303 , \3319 );
xor \U$3505 ( \3694 , \3693 , \3336 );
and \U$3506 ( \3695 , \3691 , \3694 );
and \U$3507 ( \3696 , \3681 , \3694 );
or \U$3508 ( \3697 , \3692 , \3695 , \3696 );
xor \U$3509 ( \3698 , \3552 , \3562 );
xor \U$3510 ( \3699 , \3698 , \3565 );
and \U$3511 ( \3700 , \3697 , \3699 );
xor \U$3512 ( \3701 , \3570 , \3572 );
and \U$3513 ( \3702 , \3699 , \3701 );
and \U$3514 ( \3703 , \3697 , \3701 );
or \U$3515 ( \3704 , \3700 , \3702 , \3703 );
xor \U$3516 ( \3705 , \3393 , \3411 );
xor \U$3517 ( \3706 , \3705 , \3422 );
and \U$3518 ( \3707 , \3704 , \3706 );
xor \U$3519 ( \3708 , \3568 , \3573 );
xor \U$3520 ( \3709 , \3708 , \3576 );
and \U$3521 ( \3710 , \3706 , \3709 );
and \U$3522 ( \3711 , \3704 , \3709 );
or \U$3523 ( \3712 , \3707 , \3710 , \3711 );
and \U$3524 ( \3713 , \3591 , \3712 );
xor \U$3525 ( \3714 , \3591 , \3712 );
xor \U$3526 ( \3715 , \3704 , \3706 );
xor \U$3527 ( \3716 , \3715 , \3709 );
and \U$3528 ( \3717 , \1770 , \912 );
and \U$3529 ( \3718 , \1537 , \910 );
nor \U$3530 ( \3719 , \3717 , \3718 );
xnor \U$3531 ( \3720 , \3719 , \818 );
and \U$3532 ( \3721 , \2023 , \740 );
and \U$3533 ( \3722 , \1778 , \738 );
nor \U$3534 ( \3723 , \3721 , \3722 );
xnor \U$3535 ( \3724 , \3723 , \668 );
and \U$3536 ( \3725 , \3720 , \3724 );
and \U$3537 ( \3726 , \2161 , \604 );
and \U$3538 ( \3727 , \2028 , \602 );
nor \U$3539 ( \3728 , \3726 , \3727 );
xnor \U$3540 ( \3729 , \3728 , \561 );
and \U$3541 ( \3730 , \3724 , \3729 );
and \U$3542 ( \3731 , \3720 , \3729 );
or \U$3543 ( \3732 , \3725 , \3730 , \3731 );
and \U$3544 ( \3733 , \2532 , \503 );
and \U$3545 ( \3734 , \2305 , \501 );
nor \U$3546 ( \3735 , \3733 , \3734 );
xnor \U$3547 ( \3736 , \3735 , \455 );
and \U$3548 ( \3737 , \2763 , \298 );
and \U$3549 ( \3738 , \2541 , \296 );
nor \U$3550 ( \3739 , \3737 , \3738 );
xnor \U$3551 ( \3740 , \3739 , \303 );
and \U$3552 ( \3741 , \3736 , \3740 );
nand \U$3553 ( \3742 , \2850 , \311 );
xnor \U$3554 ( \3743 , \3742 , \320 );
and \U$3555 ( \3744 , \3740 , \3743 );
and \U$3556 ( \3745 , \3736 , \3743 );
or \U$3557 ( \3746 , \3741 , \3744 , \3745 );
and \U$3558 ( \3747 , \3732 , \3746 );
and \U$3559 ( \3748 , \2541 , \298 );
and \U$3560 ( \3749 , \2532 , \296 );
nor \U$3561 ( \3750 , \3748 , \3749 );
xnor \U$3562 ( \3751 , \3750 , \303 );
and \U$3563 ( \3752 , \3746 , \3751 );
and \U$3564 ( \3753 , \3732 , \3751 );
or \U$3565 ( \3754 , \3747 , \3752 , \3753 );
and \U$3566 ( \3755 , \1104 , \1476 );
and \U$3567 ( \3756 , \904 , \1474 );
nor \U$3568 ( \3757 , \3755 , \3756 );
xnor \U$3569 ( \3758 , \3757 , \1363 );
and \U$3570 ( \3759 , \1299 , \1280 );
and \U$3571 ( \3760 , \1194 , \1278 );
nor \U$3572 ( \3761 , \3759 , \3760 );
xnor \U$3573 ( \3762 , \3761 , \1177 );
and \U$3574 ( \3763 , \3758 , \3762 );
and \U$3575 ( \3764 , \1422 , \1062 );
and \U$3576 ( \3765 , \1304 , \1060 );
nor \U$3577 ( \3766 , \3764 , \3765 );
xnor \U$3578 ( \3767 , \3766 , \984 );
and \U$3579 ( \3768 , \3762 , \3767 );
and \U$3580 ( \3769 , \3758 , \3767 );
or \U$3581 ( \3770 , \3763 , \3768 , \3769 );
and \U$3582 ( \3771 , \343 , \2913 );
and \U$3583 ( \3772 , \353 , \2910 );
nor \U$3584 ( \3773 , \3771 , \3772 );
xnor \U$3585 ( \3774 , \3773 , \2371 );
and \U$3586 ( \3775 , \444 , \2550 );
and \U$3587 ( \3776 , \360 , \2548 );
nor \U$3588 ( \3777 , \3775 , \3776 );
xnor \U$3589 ( \3778 , \3777 , \2374 );
and \U$3590 ( \3779 , \3774 , \3778 );
and \U$3591 ( \3780 , \3778 , \320 );
and \U$3592 ( \3781 , \3774 , \320 );
or \U$3593 ( \3782 , \3779 , \3780 , \3781 );
and \U$3594 ( \3783 , \3770 , \3782 );
and \U$3595 ( \3784 , \593 , \2261 );
and \U$3596 ( \3785 , \495 , \2259 );
nor \U$3597 ( \3786 , \3784 , \3785 );
xnor \U$3598 ( \3787 , \3786 , \2124 );
and \U$3599 ( \3788 , \703 , \1955 );
and \U$3600 ( \3789 , \621 , \1953 );
nor \U$3601 ( \3790 , \3788 , \3789 );
xnor \U$3602 ( \3791 , \3790 , \1835 );
and \U$3603 ( \3792 , \3787 , \3791 );
and \U$3604 ( \3793 , \841 , \1742 );
and \U$3605 ( \3794 , \777 , \1740 );
nor \U$3606 ( \3795 , \3793 , \3794 );
xnor \U$3607 ( \3796 , \3795 , \1610 );
and \U$3608 ( \3797 , \3791 , \3796 );
and \U$3609 ( \3798 , \3787 , \3796 );
or \U$3610 ( \3799 , \3792 , \3797 , \3798 );
and \U$3611 ( \3800 , \3782 , \3799 );
and \U$3612 ( \3801 , \3770 , \3799 );
or \U$3613 ( \3802 , \3783 , \3800 , \3801 );
and \U$3614 ( \3803 , \3754 , \3802 );
and \U$3615 ( \3804 , \2850 , \313 );
and \U$3616 ( \3805 , \2763 , \311 );
nor \U$3617 ( \3806 , \3804 , \3805 );
xnor \U$3618 ( \3807 , \3806 , \320 );
xor \U$3619 ( \3808 , \3658 , \3662 );
xor \U$3620 ( \3809 , \3808 , \3667 );
and \U$3621 ( \3810 , \3807 , \3809 );
xor \U$3622 ( \3811 , \3611 , \3615 );
xor \U$3623 ( \3812 , \3811 , \3620 );
and \U$3624 ( \3813 , \3809 , \3812 );
and \U$3625 ( \3814 , \3807 , \3812 );
or \U$3626 ( \3815 , \3810 , \3813 , \3814 );
and \U$3627 ( \3816 , \3802 , \3815 );
and \U$3628 ( \3817 , \3754 , \3815 );
or \U$3629 ( \3818 , \3803 , \3816 , \3817 );
xor \U$3630 ( \3819 , \3489 , \3493 );
xor \U$3631 ( \3820 , \3819 , \338 );
xor \U$3632 ( \3821 , \3645 , \3647 );
xor \U$3633 ( \3822 , \3821 , \3650 );
and \U$3634 ( \3823 , \3820 , \3822 );
xor \U$3635 ( \3824 , \3670 , \3672 );
xor \U$3636 ( \3825 , \3824 , \3675 );
and \U$3637 ( \3826 , \3822 , \3825 );
and \U$3638 ( \3827 , \3820 , \3825 );
or \U$3639 ( \3828 , \3823 , \3826 , \3827 );
and \U$3640 ( \3829 , \3818 , \3828 );
xor \U$3641 ( \3830 , \3468 , \3484 );
xor \U$3642 ( \3831 , \3830 , \3497 );
and \U$3643 ( \3832 , \3828 , \3831 );
and \U$3644 ( \3833 , \3818 , \3831 );
or \U$3645 ( \3834 , \3829 , \3832 , \3833 );
xor \U$3646 ( \3835 , \3643 , \3653 );
xor \U$3647 ( \3836 , \3835 , \3678 );
xor \U$3648 ( \3837 , \3683 , \3685 );
xor \U$3649 ( \3838 , \3837 , \3688 );
and \U$3650 ( \3839 , \3836 , \3838 );
and \U$3651 ( \3840 , \3834 , \3839 );
xor \U$3652 ( \3841 , \3554 , \3556 );
xor \U$3653 ( \3842 , \3841 , \3559 );
and \U$3654 ( \3843 , \3839 , \3842 );
and \U$3655 ( \3844 , \3834 , \3842 );
or \U$3656 ( \3845 , \3840 , \3843 , \3844 );
xor \U$3657 ( \3846 , \3500 , \3538 );
xor \U$3658 ( \3847 , \3846 , \3549 );
xor \U$3659 ( \3848 , \3681 , \3691 );
xor \U$3660 ( \3849 , \3848 , \3694 );
and \U$3661 ( \3850 , \3847 , \3849 );
and \U$3662 ( \3851 , \3845 , \3850 );
xor \U$3663 ( \3852 , \3697 , \3699 );
xor \U$3664 ( \3853 , \3852 , \3701 );
and \U$3665 ( \3854 , \3850 , \3853 );
and \U$3666 ( \3855 , \3845 , \3853 );
or \U$3667 ( \3856 , \3851 , \3854 , \3855 );
and \U$3668 ( \3857 , \3716 , \3856 );
xor \U$3669 ( \3858 , \3716 , \3856 );
xor \U$3670 ( \3859 , \3845 , \3850 );
xor \U$3671 ( \3860 , \3859 , \3853 );
and \U$3672 ( \3861 , \777 , \1955 );
and \U$3673 ( \3862 , \703 , \1953 );
nor \U$3674 ( \3863 , \3861 , \3862 );
xnor \U$3675 ( \3864 , \3863 , \1835 );
and \U$3676 ( \3865 , \904 , \1742 );
and \U$3677 ( \3866 , \841 , \1740 );
nor \U$3678 ( \3867 , \3865 , \3866 );
xnor \U$3679 ( \3868 , \3867 , \1610 );
and \U$3680 ( \3869 , \3864 , \3868 );
and \U$3681 ( \3870 , \1194 , \1476 );
and \U$3682 ( \3871 , \1104 , \1474 );
nor \U$3683 ( \3872 , \3870 , \3871 );
xnor \U$3684 ( \3873 , \3872 , \1363 );
and \U$3685 ( \3874 , \3868 , \3873 );
and \U$3686 ( \3875 , \3864 , \3873 );
or \U$3687 ( \3876 , \3869 , \3874 , \3875 );
and \U$3688 ( \3877 , \360 , \2913 );
and \U$3689 ( \3878 , \343 , \2910 );
nor \U$3690 ( \3879 , \3877 , \3878 );
xnor \U$3691 ( \3880 , \3879 , \2371 );
and \U$3692 ( \3881 , \495 , \2550 );
and \U$3693 ( \3882 , \444 , \2548 );
nor \U$3694 ( \3883 , \3881 , \3882 );
xnor \U$3695 ( \3884 , \3883 , \2374 );
and \U$3696 ( \3885 , \3880 , \3884 );
and \U$3697 ( \3886 , \621 , \2261 );
and \U$3698 ( \3887 , \593 , \2259 );
nor \U$3699 ( \3888 , \3886 , \3887 );
xnor \U$3700 ( \3889 , \3888 , \2124 );
and \U$3701 ( \3890 , \3884 , \3889 );
and \U$3702 ( \3891 , \3880 , \3889 );
or \U$3703 ( \3892 , \3885 , \3890 , \3891 );
and \U$3704 ( \3893 , \3876 , \3892 );
and \U$3705 ( \3894 , \1304 , \1280 );
and \U$3706 ( \3895 , \1299 , \1278 );
nor \U$3707 ( \3896 , \3894 , \3895 );
xnor \U$3708 ( \3897 , \3896 , \1177 );
and \U$3709 ( \3898 , \1537 , \1062 );
and \U$3710 ( \3899 , \1422 , \1060 );
nor \U$3711 ( \3900 , \3898 , \3899 );
xnor \U$3712 ( \3901 , \3900 , \984 );
and \U$3713 ( \3902 , \3897 , \3901 );
and \U$3714 ( \3903 , \1778 , \912 );
and \U$3715 ( \3904 , \1770 , \910 );
nor \U$3716 ( \3905 , \3903 , \3904 );
xnor \U$3717 ( \3906 , \3905 , \818 );
and \U$3718 ( \3907 , \3901 , \3906 );
and \U$3719 ( \3908 , \3897 , \3906 );
or \U$3720 ( \3909 , \3902 , \3907 , \3908 );
and \U$3721 ( \3910 , \3892 , \3909 );
and \U$3722 ( \3911 , \3876 , \3909 );
or \U$3723 ( \3912 , \3893 , \3910 , \3911 );
xor \U$3724 ( \3913 , \3758 , \3762 );
xor \U$3725 ( \3914 , \3913 , \3767 );
xor \U$3726 ( \3915 , \3774 , \3778 );
xor \U$3727 ( \3916 , \3915 , \320 );
and \U$3728 ( \3917 , \3914 , \3916 );
xor \U$3729 ( \3918 , \3787 , \3791 );
xor \U$3730 ( \3919 , \3918 , \3796 );
and \U$3731 ( \3920 , \3916 , \3919 );
and \U$3732 ( \3921 , \3914 , \3919 );
or \U$3733 ( \3922 , \3917 , \3920 , \3921 );
and \U$3734 ( \3923 , \3912 , \3922 );
and \U$3735 ( \3924 , \2028 , \740 );
and \U$3736 ( \3925 , \2023 , \738 );
nor \U$3737 ( \3926 , \3924 , \3925 );
xnor \U$3738 ( \3927 , \3926 , \668 );
and \U$3739 ( \3928 , \2305 , \604 );
and \U$3740 ( \3929 , \2161 , \602 );
nor \U$3741 ( \3930 , \3928 , \3929 );
xnor \U$3742 ( \3931 , \3930 , \561 );
and \U$3743 ( \3932 , \3927 , \3931 );
and \U$3744 ( \3933 , \2541 , \503 );
and \U$3745 ( \3934 , \2532 , \501 );
nor \U$3746 ( \3935 , \3933 , \3934 );
xnor \U$3747 ( \3936 , \3935 , \455 );
and \U$3748 ( \3937 , \3931 , \3936 );
and \U$3749 ( \3938 , \3927 , \3936 );
or \U$3750 ( \3939 , \3932 , \3937 , \3938 );
xor \U$3751 ( \3940 , \3720 , \3724 );
xor \U$3752 ( \3941 , \3940 , \3729 );
and \U$3753 ( \3942 , \3939 , \3941 );
xor \U$3754 ( \3943 , \3736 , \3740 );
xor \U$3755 ( \3944 , \3943 , \3743 );
and \U$3756 ( \3945 , \3941 , \3944 );
and \U$3757 ( \3946 , \3939 , \3944 );
or \U$3758 ( \3947 , \3942 , \3945 , \3946 );
and \U$3759 ( \3948 , \3922 , \3947 );
and \U$3760 ( \3949 , \3912 , \3947 );
or \U$3761 ( \3950 , \3923 , \3948 , \3949 );
xor \U$3762 ( \3951 , \3595 , \3599 );
xor \U$3763 ( \3952 , \3951 , \3604 );
xor \U$3764 ( \3953 , \3628 , \3632 );
xor \U$3765 ( \3954 , \3953 , \3637 );
and \U$3766 ( \3955 , \3952 , \3954 );
xor \U$3767 ( \3956 , \3807 , \3809 );
xor \U$3768 ( \3957 , \3956 , \3812 );
and \U$3769 ( \3958 , \3954 , \3957 );
and \U$3770 ( \3959 , \3952 , \3957 );
or \U$3771 ( \3960 , \3955 , \3958 , \3959 );
and \U$3772 ( \3961 , \3950 , \3960 );
xor \U$3773 ( \3962 , \3607 , \3623 );
xor \U$3774 ( \3963 , \3962 , \3640 );
and \U$3775 ( \3964 , \3960 , \3963 );
and \U$3776 ( \3965 , \3950 , \3963 );
or \U$3777 ( \3966 , \3961 , \3964 , \3965 );
xor \U$3778 ( \3967 , \3818 , \3828 );
xor \U$3779 ( \3968 , \3967 , \3831 );
and \U$3780 ( \3969 , \3966 , \3968 );
xor \U$3781 ( \3970 , \3836 , \3838 );
and \U$3782 ( \3971 , \3968 , \3970 );
and \U$3783 ( \3972 , \3966 , \3970 );
or \U$3784 ( \3973 , \3969 , \3971 , \3972 );
xor \U$3785 ( \3974 , \3834 , \3839 );
xor \U$3786 ( \3975 , \3974 , \3842 );
and \U$3787 ( \3976 , \3973 , \3975 );
xor \U$3788 ( \3977 , \3847 , \3849 );
and \U$3789 ( \3978 , \3975 , \3977 );
and \U$3790 ( \3979 , \3973 , \3977 );
or \U$3791 ( \3980 , \3976 , \3978 , \3979 );
and \U$3792 ( \3981 , \3860 , \3980 );
xor \U$3793 ( \3982 , \3860 , \3980 );
xor \U$3794 ( \3983 , \3973 , \3975 );
xor \U$3795 ( \3984 , \3983 , \3977 );
and \U$3796 ( \3985 , \703 , \2261 );
and \U$3797 ( \3986 , \621 , \2259 );
nor \U$3798 ( \3987 , \3985 , \3986 );
xnor \U$3799 ( \3988 , \3987 , \2124 );
and \U$3800 ( \3989 , \841 , \1955 );
and \U$3801 ( \3990 , \777 , \1953 );
nor \U$3802 ( \3991 , \3989 , \3990 );
xnor \U$3803 ( \3992 , \3991 , \1835 );
and \U$3804 ( \3993 , \3988 , \3992 );
and \U$3805 ( \3994 , \1104 , \1742 );
and \U$3806 ( \3995 , \904 , \1740 );
nor \U$3807 ( \3996 , \3994 , \3995 );
xnor \U$3808 ( \3997 , \3996 , \1610 );
and \U$3809 ( \3998 , \3992 , \3997 );
and \U$3810 ( \3999 , \3988 , \3997 );
or \U$3811 ( \4000 , \3993 , \3998 , \3999 );
and \U$3812 ( \4001 , \444 , \2913 );
and \U$3813 ( \4002 , \360 , \2910 );
nor \U$3814 ( \4003 , \4001 , \4002 );
xnor \U$3815 ( \4004 , \4003 , \2371 );
and \U$3816 ( \4005 , \593 , \2550 );
and \U$3817 ( \4006 , \495 , \2548 );
nor \U$3818 ( \4007 , \4005 , \4006 );
xnor \U$3819 ( \4008 , \4007 , \2374 );
and \U$3820 ( \4009 , \4004 , \4008 );
and \U$3821 ( \4010 , \4008 , \303 );
and \U$3822 ( \4011 , \4004 , \303 );
or \U$3823 ( \4012 , \4009 , \4010 , \4011 );
and \U$3824 ( \4013 , \4000 , \4012 );
and \U$3825 ( \4014 , \1299 , \1476 );
and \U$3826 ( \4015 , \1194 , \1474 );
nor \U$3827 ( \4016 , \4014 , \4015 );
xnor \U$3828 ( \4017 , \4016 , \1363 );
and \U$3829 ( \4018 , \1422 , \1280 );
and \U$3830 ( \4019 , \1304 , \1278 );
nor \U$3831 ( \4020 , \4018 , \4019 );
xnor \U$3832 ( \4021 , \4020 , \1177 );
and \U$3833 ( \4022 , \4017 , \4021 );
and \U$3834 ( \4023 , \1770 , \1062 );
and \U$3835 ( \4024 , \1537 , \1060 );
nor \U$3836 ( \4025 , \4023 , \4024 );
xnor \U$3837 ( \4026 , \4025 , \984 );
and \U$3838 ( \4027 , \4021 , \4026 );
and \U$3839 ( \4028 , \4017 , \4026 );
or \U$3840 ( \4029 , \4022 , \4027 , \4028 );
and \U$3841 ( \4030 , \4012 , \4029 );
and \U$3842 ( \4031 , \4000 , \4029 );
or \U$3843 ( \4032 , \4013 , \4030 , \4031 );
and \U$3844 ( \4033 , \2023 , \912 );
and \U$3845 ( \4034 , \1778 , \910 );
nor \U$3846 ( \4035 , \4033 , \4034 );
xnor \U$3847 ( \4036 , \4035 , \818 );
and \U$3848 ( \4037 , \2161 , \740 );
and \U$3849 ( \4038 , \2028 , \738 );
nor \U$3850 ( \4039 , \4037 , \4038 );
xnor \U$3851 ( \4040 , \4039 , \668 );
and \U$3852 ( \4041 , \4036 , \4040 );
and \U$3853 ( \4042 , \2532 , \604 );
and \U$3854 ( \4043 , \2305 , \602 );
nor \U$3855 ( \4044 , \4042 , \4043 );
xnor \U$3856 ( \4045 , \4044 , \561 );
and \U$3857 ( \4046 , \4040 , \4045 );
and \U$3858 ( \4047 , \4036 , \4045 );
or \U$3859 ( \4048 , \4041 , \4046 , \4047 );
and \U$3860 ( \4049 , \2763 , \503 );
and \U$3861 ( \4050 , \2541 , \501 );
nor \U$3862 ( \4051 , \4049 , \4050 );
xnor \U$3863 ( \4052 , \4051 , \455 );
nand \U$3864 ( \4053 , \2850 , \296 );
xnor \U$3865 ( \4054 , \4053 , \303 );
and \U$3866 ( \4055 , \4052 , \4054 );
and \U$3867 ( \4056 , \4048 , \4055 );
and \U$3868 ( \4057 , \2850 , \298 );
and \U$3869 ( \4058 , \2763 , \296 );
nor \U$3870 ( \4059 , \4057 , \4058 );
xnor \U$3871 ( \4060 , \4059 , \303 );
and \U$3872 ( \4061 , \4055 , \4060 );
and \U$3873 ( \4062 , \4048 , \4060 );
or \U$3874 ( \4063 , \4056 , \4061 , \4062 );
and \U$3875 ( \4064 , \4032 , \4063 );
xor \U$3876 ( \4065 , \3864 , \3868 );
xor \U$3877 ( \4066 , \4065 , \3873 );
xor \U$3878 ( \4067 , \3927 , \3931 );
xor \U$3879 ( \4068 , \4067 , \3936 );
and \U$3880 ( \4069 , \4066 , \4068 );
xor \U$3881 ( \4070 , \3897 , \3901 );
xor \U$3882 ( \4071 , \4070 , \3906 );
and \U$3883 ( \4072 , \4068 , \4071 );
and \U$3884 ( \4073 , \4066 , \4071 );
or \U$3885 ( \4074 , \4069 , \4072 , \4073 );
and \U$3886 ( \4075 , \4063 , \4074 );
and \U$3887 ( \4076 , \4032 , \4074 );
or \U$3888 ( \4077 , \4064 , \4075 , \4076 );
xor \U$3889 ( \4078 , \3876 , \3892 );
xor \U$3890 ( \4079 , \4078 , \3909 );
xor \U$3891 ( \4080 , \3914 , \3916 );
xor \U$3892 ( \4081 , \4080 , \3919 );
and \U$3893 ( \4082 , \4079 , \4081 );
xor \U$3894 ( \4083 , \3939 , \3941 );
xor \U$3895 ( \4084 , \4083 , \3944 );
and \U$3896 ( \4085 , \4081 , \4084 );
and \U$3897 ( \4086 , \4079 , \4084 );
or \U$3898 ( \4087 , \4082 , \4085 , \4086 );
and \U$3899 ( \4088 , \4077 , \4087 );
xor \U$3900 ( \4089 , \3732 , \3746 );
xor \U$3901 ( \4090 , \4089 , \3751 );
and \U$3902 ( \4091 , \4087 , \4090 );
and \U$3903 ( \4092 , \4077 , \4090 );
or \U$3904 ( \4093 , \4088 , \4091 , \4092 );
xor \U$3905 ( \4094 , \3770 , \3782 );
xor \U$3906 ( \4095 , \4094 , \3799 );
xor \U$3907 ( \4096 , \3912 , \3922 );
xor \U$3908 ( \4097 , \4096 , \3947 );
and \U$3909 ( \4098 , \4095 , \4097 );
xor \U$3910 ( \4099 , \3952 , \3954 );
xor \U$3911 ( \4100 , \4099 , \3957 );
and \U$3912 ( \4101 , \4097 , \4100 );
and \U$3913 ( \4102 , \4095 , \4100 );
or \U$3914 ( \4103 , \4098 , \4101 , \4102 );
and \U$3915 ( \4104 , \4093 , \4103 );
xor \U$3916 ( \4105 , \3820 , \3822 );
xor \U$3917 ( \4106 , \4105 , \3825 );
and \U$3918 ( \4107 , \4103 , \4106 );
and \U$3919 ( \4108 , \4093 , \4106 );
or \U$3920 ( \4109 , \4104 , \4107 , \4108 );
xor \U$3921 ( \4110 , \3754 , \3802 );
xor \U$3922 ( \4111 , \4110 , \3815 );
xor \U$3923 ( \4112 , \3950 , \3960 );
xor \U$3924 ( \4113 , \4112 , \3963 );
and \U$3925 ( \4114 , \4111 , \4113 );
and \U$3926 ( \4115 , \4109 , \4114 );
xor \U$3927 ( \4116 , \3966 , \3968 );
xor \U$3928 ( \4117 , \4116 , \3970 );
and \U$3929 ( \4118 , \4114 , \4117 );
and \U$3930 ( \4119 , \4109 , \4117 );
or \U$3931 ( \4120 , \4115 , \4118 , \4119 );
and \U$3932 ( \4121 , \3984 , \4120 );
xor \U$3933 ( \4122 , \3984 , \4120 );
xor \U$3934 ( \4123 , \4109 , \4114 );
xor \U$3935 ( \4124 , \4123 , \4117 );
and \U$3936 ( \4125 , \904 , \1955 );
and \U$3937 ( \4126 , \841 , \1953 );
nor \U$3938 ( \4127 , \4125 , \4126 );
xnor \U$3939 ( \4128 , \4127 , \1835 );
and \U$3940 ( \4129 , \1194 , \1742 );
and \U$3941 ( \4130 , \1104 , \1740 );
nor \U$3942 ( \4131 , \4129 , \4130 );
xnor \U$3943 ( \4132 , \4131 , \1610 );
and \U$3944 ( \4133 , \4128 , \4132 );
and \U$3945 ( \4134 , \1304 , \1476 );
and \U$3946 ( \4135 , \1299 , \1474 );
nor \U$3947 ( \4136 , \4134 , \4135 );
xnor \U$3948 ( \4137 , \4136 , \1363 );
and \U$3949 ( \4138 , \4132 , \4137 );
and \U$3950 ( \4139 , \4128 , \4137 );
or \U$3951 ( \4140 , \4133 , \4138 , \4139 );
and \U$3952 ( \4141 , \1537 , \1280 );
and \U$3953 ( \4142 , \1422 , \1278 );
nor \U$3954 ( \4143 , \4141 , \4142 );
xnor \U$3955 ( \4144 , \4143 , \1177 );
and \U$3956 ( \4145 , \1778 , \1062 );
and \U$3957 ( \4146 , \1770 , \1060 );
nor \U$3958 ( \4147 , \4145 , \4146 );
xnor \U$3959 ( \4148 , \4147 , \984 );
and \U$3960 ( \4149 , \4144 , \4148 );
and \U$3961 ( \4150 , \2028 , \912 );
and \U$3962 ( \4151 , \2023 , \910 );
nor \U$3963 ( \4152 , \4150 , \4151 );
xnor \U$3964 ( \4153 , \4152 , \818 );
and \U$3965 ( \4154 , \4148 , \4153 );
and \U$3966 ( \4155 , \4144 , \4153 );
or \U$3967 ( \4156 , \4149 , \4154 , \4155 );
and \U$3968 ( \4157 , \4140 , \4156 );
and \U$3969 ( \4158 , \495 , \2913 );
and \U$3970 ( \4159 , \444 , \2910 );
nor \U$3971 ( \4160 , \4158 , \4159 );
xnor \U$3972 ( \4161 , \4160 , \2371 );
and \U$3973 ( \4162 , \621 , \2550 );
and \U$3974 ( \4163 , \593 , \2548 );
nor \U$3975 ( \4164 , \4162 , \4163 );
xnor \U$3976 ( \4165 , \4164 , \2374 );
and \U$3977 ( \4166 , \4161 , \4165 );
and \U$3978 ( \4167 , \777 , \2261 );
and \U$3979 ( \4168 , \703 , \2259 );
nor \U$3980 ( \4169 , \4167 , \4168 );
xnor \U$3981 ( \4170 , \4169 , \2124 );
and \U$3982 ( \4171 , \4165 , \4170 );
and \U$3983 ( \4172 , \4161 , \4170 );
or \U$3984 ( \4173 , \4166 , \4171 , \4172 );
and \U$3985 ( \4174 , \4156 , \4173 );
and \U$3986 ( \4175 , \4140 , \4173 );
or \U$3987 ( \4176 , \4157 , \4174 , \4175 );
xor \U$3988 ( \4177 , \3988 , \3992 );
xor \U$3989 ( \4178 , \4177 , \3997 );
xor \U$3990 ( \4179 , \4004 , \4008 );
xor \U$3991 ( \4180 , \4179 , \303 );
and \U$3992 ( \4181 , \4178 , \4180 );
xor \U$3993 ( \4182 , \4017 , \4021 );
xor \U$3994 ( \4183 , \4182 , \4026 );
and \U$3995 ( \4184 , \4180 , \4183 );
and \U$3996 ( \4185 , \4178 , \4183 );
or \U$3997 ( \4186 , \4181 , \4184 , \4185 );
and \U$3998 ( \4187 , \4176 , \4186 );
and \U$3999 ( \4188 , \2305 , \740 );
and \U$4000 ( \4189 , \2161 , \738 );
nor \U$4001 ( \4190 , \4188 , \4189 );
xnor \U$4002 ( \4191 , \4190 , \668 );
and \U$4003 ( \4192 , \2541 , \604 );
and \U$4004 ( \4193 , \2532 , \602 );
nor \U$4005 ( \4194 , \4192 , \4193 );
xnor \U$4006 ( \4195 , \4194 , \561 );
and \U$4007 ( \4196 , \4191 , \4195 );
and \U$4008 ( \4197 , \2850 , \503 );
and \U$4009 ( \4198 , \2763 , \501 );
nor \U$4010 ( \4199 , \4197 , \4198 );
xnor \U$4011 ( \4200 , \4199 , \455 );
and \U$4012 ( \4201 , \4195 , \4200 );
and \U$4013 ( \4202 , \4191 , \4200 );
or \U$4014 ( \4203 , \4196 , \4201 , \4202 );
xor \U$4015 ( \4204 , \4036 , \4040 );
xor \U$4016 ( \4205 , \4204 , \4045 );
and \U$4017 ( \4206 , \4203 , \4205 );
xor \U$4018 ( \4207 , \4052 , \4054 );
and \U$4019 ( \4208 , \4205 , \4207 );
and \U$4020 ( \4209 , \4203 , \4207 );
or \U$4021 ( \4210 , \4206 , \4208 , \4209 );
and \U$4022 ( \4211 , \4186 , \4210 );
and \U$4023 ( \4212 , \4176 , \4210 );
or \U$4024 ( \4213 , \4187 , \4211 , \4212 );
xor \U$4025 ( \4214 , \3880 , \3884 );
xor \U$4026 ( \4215 , \4214 , \3889 );
xor \U$4027 ( \4216 , \4048 , \4055 );
xor \U$4028 ( \4217 , \4216 , \4060 );
and \U$4029 ( \4218 , \4215 , \4217 );
xor \U$4030 ( \4219 , \4066 , \4068 );
xor \U$4031 ( \4220 , \4219 , \4071 );
and \U$4032 ( \4221 , \4217 , \4220 );
and \U$4033 ( \4222 , \4215 , \4220 );
or \U$4034 ( \4223 , \4218 , \4221 , \4222 );
and \U$4035 ( \4224 , \4213 , \4223 );
xor \U$4036 ( \4225 , \4079 , \4081 );
xor \U$4037 ( \4226 , \4225 , \4084 );
and \U$4038 ( \4227 , \4223 , \4226 );
and \U$4039 ( \4228 , \4213 , \4226 );
or \U$4040 ( \4229 , \4224 , \4227 , \4228 );
xor \U$4041 ( \4230 , \4077 , \4087 );
xor \U$4042 ( \4231 , \4230 , \4090 );
and \U$4043 ( \4232 , \4229 , \4231 );
xor \U$4044 ( \4233 , \4095 , \4097 );
xor \U$4045 ( \4234 , \4233 , \4100 );
and \U$4046 ( \4235 , \4231 , \4234 );
and \U$4047 ( \4236 , \4229 , \4234 );
or \U$4048 ( \4237 , \4232 , \4235 , \4236 );
xor \U$4049 ( \4238 , \4093 , \4103 );
xor \U$4050 ( \4239 , \4238 , \4106 );
and \U$4051 ( \4240 , \4237 , \4239 );
xor \U$4052 ( \4241 , \4111 , \4113 );
and \U$4053 ( \4242 , \4239 , \4241 );
and \U$4054 ( \4243 , \4237 , \4241 );
or \U$4055 ( \4244 , \4240 , \4242 , \4243 );
and \U$4056 ( \4245 , \4124 , \4244 );
xor \U$4057 ( \4246 , \4124 , \4244 );
xor \U$4058 ( \4247 , \4237 , \4239 );
xor \U$4059 ( \4248 , \4247 , \4241 );
and \U$4060 ( \4249 , \841 , \2261 );
and \U$4061 ( \4250 , \777 , \2259 );
nor \U$4062 ( \4251 , \4249 , \4250 );
xnor \U$4063 ( \4252 , \4251 , \2124 );
and \U$4064 ( \4253 , \1104 , \1955 );
and \U$4065 ( \4254 , \904 , \1953 );
nor \U$4066 ( \4255 , \4253 , \4254 );
xnor \U$4067 ( \4256 , \4255 , \1835 );
and \U$4068 ( \4257 , \4252 , \4256 );
and \U$4069 ( \4258 , \1299 , \1742 );
and \U$4070 ( \4259 , \1194 , \1740 );
nor \U$4071 ( \4260 , \4258 , \4259 );
xnor \U$4072 ( \4261 , \4260 , \1610 );
and \U$4073 ( \4262 , \4256 , \4261 );
and \U$4074 ( \4263 , \4252 , \4261 );
or \U$4075 ( \4264 , \4257 , \4262 , \4263 );
and \U$4076 ( \4265 , \1422 , \1476 );
and \U$4077 ( \4266 , \1304 , \1474 );
nor \U$4078 ( \4267 , \4265 , \4266 );
xnor \U$4079 ( \4268 , \4267 , \1363 );
and \U$4080 ( \4269 , \1770 , \1280 );
and \U$4081 ( \4270 , \1537 , \1278 );
nor \U$4082 ( \4271 , \4269 , \4270 );
xnor \U$4083 ( \4272 , \4271 , \1177 );
and \U$4084 ( \4273 , \4268 , \4272 );
and \U$4085 ( \4274 , \2023 , \1062 );
and \U$4086 ( \4275 , \1778 , \1060 );
nor \U$4087 ( \4276 , \4274 , \4275 );
xnor \U$4088 ( \4277 , \4276 , \984 );
and \U$4089 ( \4278 , \4272 , \4277 );
and \U$4090 ( \4279 , \4268 , \4277 );
or \U$4091 ( \4280 , \4273 , \4278 , \4279 );
and \U$4092 ( \4281 , \4264 , \4280 );
and \U$4093 ( \4282 , \593 , \2913 );
and \U$4094 ( \4283 , \495 , \2910 );
nor \U$4095 ( \4284 , \4282 , \4283 );
xnor \U$4096 ( \4285 , \4284 , \2371 );
and \U$4097 ( \4286 , \703 , \2550 );
and \U$4098 ( \4287 , \621 , \2548 );
nor \U$4099 ( \4288 , \4286 , \4287 );
xnor \U$4100 ( \4289 , \4288 , \2374 );
and \U$4101 ( \4290 , \4285 , \4289 );
and \U$4102 ( \4291 , \4289 , \455 );
and \U$4103 ( \4292 , \4285 , \455 );
or \U$4104 ( \4293 , \4290 , \4291 , \4292 );
and \U$4105 ( \4294 , \4280 , \4293 );
and \U$4106 ( \4295 , \4264 , \4293 );
or \U$4107 ( \4296 , \4281 , \4294 , \4295 );
and \U$4108 ( \4297 , \2161 , \912 );
and \U$4109 ( \4298 , \2028 , \910 );
nor \U$4110 ( \4299 , \4297 , \4298 );
xnor \U$4111 ( \4300 , \4299 , \818 );
and \U$4112 ( \4301 , \2532 , \740 );
and \U$4113 ( \4302 , \2305 , \738 );
nor \U$4114 ( \4303 , \4301 , \4302 );
xnor \U$4115 ( \4304 , \4303 , \668 );
and \U$4116 ( \4305 , \4300 , \4304 );
and \U$4117 ( \4306 , \2763 , \604 );
and \U$4118 ( \4307 , \2541 , \602 );
nor \U$4119 ( \4308 , \4306 , \4307 );
xnor \U$4120 ( \4309 , \4308 , \561 );
and \U$4121 ( \4310 , \4304 , \4309 );
and \U$4122 ( \4311 , \4300 , \4309 );
or \U$4123 ( \4312 , \4305 , \4310 , \4311 );
xor \U$4124 ( \4313 , \4144 , \4148 );
xor \U$4125 ( \4314 , \4313 , \4153 );
and \U$4126 ( \4315 , \4312 , \4314 );
xor \U$4127 ( \4316 , \4191 , \4195 );
xor \U$4128 ( \4317 , \4316 , \4200 );
and \U$4129 ( \4318 , \4314 , \4317 );
and \U$4130 ( \4319 , \4312 , \4317 );
or \U$4131 ( \4320 , \4315 , \4318 , \4319 );
and \U$4132 ( \4321 , \4296 , \4320 );
xor \U$4133 ( \4322 , \4128 , \4132 );
xor \U$4134 ( \4323 , \4322 , \4137 );
xor \U$4135 ( \4324 , \4161 , \4165 );
xor \U$4136 ( \4325 , \4324 , \4170 );
and \U$4137 ( \4326 , \4323 , \4325 );
and \U$4138 ( \4327 , \4320 , \4326 );
and \U$4139 ( \4328 , \4296 , \4326 );
or \U$4140 ( \4329 , \4321 , \4327 , \4328 );
xor \U$4141 ( \4330 , \4140 , \4156 );
xor \U$4142 ( \4331 , \4330 , \4173 );
xor \U$4143 ( \4332 , \4178 , \4180 );
xor \U$4144 ( \4333 , \4332 , \4183 );
and \U$4145 ( \4334 , \4331 , \4333 );
xor \U$4146 ( \4335 , \4203 , \4205 );
xor \U$4147 ( \4336 , \4335 , \4207 );
and \U$4148 ( \4337 , \4333 , \4336 );
and \U$4149 ( \4338 , \4331 , \4336 );
or \U$4150 ( \4339 , \4334 , \4337 , \4338 );
and \U$4151 ( \4340 , \4329 , \4339 );
xor \U$4152 ( \4341 , \4000 , \4012 );
xor \U$4153 ( \4342 , \4341 , \4029 );
and \U$4154 ( \4343 , \4339 , \4342 );
and \U$4155 ( \4344 , \4329 , \4342 );
or \U$4156 ( \4345 , \4340 , \4343 , \4344 );
xor \U$4157 ( \4346 , \4176 , \4186 );
xor \U$4158 ( \4347 , \4346 , \4210 );
xor \U$4159 ( \4348 , \4215 , \4217 );
xor \U$4160 ( \4349 , \4348 , \4220 );
and \U$4161 ( \4350 , \4347 , \4349 );
and \U$4162 ( \4351 , \4345 , \4350 );
xor \U$4163 ( \4352 , \4032 , \4063 );
xor \U$4164 ( \4353 , \4352 , \4074 );
and \U$4165 ( \4354 , \4350 , \4353 );
and \U$4166 ( \4355 , \4345 , \4353 );
or \U$4167 ( \4356 , \4351 , \4354 , \4355 );
xor \U$4168 ( \4357 , \4229 , \4231 );
xor \U$4169 ( \4358 , \4357 , \4234 );
and \U$4170 ( \4359 , \4356 , \4358 );
and \U$4171 ( \4360 , \4248 , \4359 );
xor \U$4172 ( \4361 , \4248 , \4359 );
xor \U$4173 ( \4362 , \4356 , \4358 );
xor \U$4174 ( \4363 , \4345 , \4350 );
xor \U$4175 ( \4364 , \4363 , \4353 );
xor \U$4176 ( \4365 , \4213 , \4223 );
xor \U$4177 ( \4366 , \4365 , \4226 );
and \U$4178 ( \4367 , \4364 , \4366 );
and \U$4179 ( \4368 , \4362 , \4367 );
xor \U$4180 ( \4369 , \4362 , \4367 );
xor \U$4181 ( \4370 , \4364 , \4366 );
and \U$4182 ( \4371 , \621 , \2913 );
and \U$4183 ( \4372 , \593 , \2910 );
nor \U$4184 ( \4373 , \4371 , \4372 );
xnor \U$4185 ( \4374 , \4373 , \2371 );
and \U$4186 ( \4375 , \777 , \2550 );
and \U$4187 ( \4376 , \703 , \2548 );
nor \U$4188 ( \4377 , \4375 , \4376 );
xnor \U$4189 ( \4378 , \4377 , \2374 );
and \U$4190 ( \4379 , \4374 , \4378 );
and \U$4191 ( \4380 , \904 , \2261 );
and \U$4192 ( \4381 , \841 , \2259 );
nor \U$4193 ( \4382 , \4380 , \4381 );
xnor \U$4194 ( \4383 , \4382 , \2124 );
and \U$4195 ( \4384 , \4378 , \4383 );
and \U$4196 ( \4385 , \4374 , \4383 );
or \U$4197 ( \4386 , \4379 , \4384 , \4385 );
and \U$4198 ( \4387 , \1778 , \1280 );
and \U$4199 ( \4388 , \1770 , \1278 );
nor \U$4200 ( \4389 , \4387 , \4388 );
xnor \U$4201 ( \4390 , \4389 , \1177 );
and \U$4202 ( \4391 , \2028 , \1062 );
and \U$4203 ( \4392 , \2023 , \1060 );
nor \U$4204 ( \4393 , \4391 , \4392 );
xnor \U$4205 ( \4394 , \4393 , \984 );
and \U$4206 ( \4395 , \4390 , \4394 );
and \U$4207 ( \4396 , \2305 , \912 );
and \U$4208 ( \4397 , \2161 , \910 );
nor \U$4209 ( \4398 , \4396 , \4397 );
xnor \U$4210 ( \4399 , \4398 , \818 );
and \U$4211 ( \4400 , \4394 , \4399 );
and \U$4212 ( \4401 , \4390 , \4399 );
or \U$4213 ( \4402 , \4395 , \4400 , \4401 );
and \U$4214 ( \4403 , \4386 , \4402 );
and \U$4215 ( \4404 , \1194 , \1955 );
and \U$4216 ( \4405 , \1104 , \1953 );
nor \U$4217 ( \4406 , \4404 , \4405 );
xnor \U$4218 ( \4407 , \4406 , \1835 );
and \U$4219 ( \4408 , \1304 , \1742 );
and \U$4220 ( \4409 , \1299 , \1740 );
nor \U$4221 ( \4410 , \4408 , \4409 );
xnor \U$4222 ( \4411 , \4410 , \1610 );
and \U$4223 ( \4412 , \4407 , \4411 );
and \U$4224 ( \4413 , \1537 , \1476 );
and \U$4225 ( \4414 , \1422 , \1474 );
nor \U$4226 ( \4415 , \4413 , \4414 );
xnor \U$4227 ( \4416 , \4415 , \1363 );
and \U$4228 ( \4417 , \4411 , \4416 );
and \U$4229 ( \4418 , \4407 , \4416 );
or \U$4230 ( \4419 , \4412 , \4417 , \4418 );
and \U$4231 ( \4420 , \4402 , \4419 );
and \U$4232 ( \4421 , \4386 , \4419 );
or \U$4233 ( \4422 , \4403 , \4420 , \4421 );
nand \U$4234 ( \4423 , \2850 , \501 );
xnor \U$4235 ( \4424 , \4423 , \455 );
xor \U$4236 ( \4425 , \4268 , \4272 );
xor \U$4237 ( \4426 , \4425 , \4277 );
and \U$4238 ( \4427 , \4424 , \4426 );
xor \U$4239 ( \4428 , \4300 , \4304 );
xor \U$4240 ( \4429 , \4428 , \4309 );
and \U$4241 ( \4430 , \4426 , \4429 );
and \U$4242 ( \4431 , \4424 , \4429 );
or \U$4243 ( \4432 , \4427 , \4430 , \4431 );
and \U$4244 ( \4433 , \4422 , \4432 );
xor \U$4245 ( \4434 , \4252 , \4256 );
xor \U$4246 ( \4435 , \4434 , \4261 );
xor \U$4247 ( \4436 , \4285 , \4289 );
xor \U$4248 ( \4437 , \4436 , \455 );
and \U$4249 ( \4438 , \4435 , \4437 );
and \U$4250 ( \4439 , \4432 , \4438 );
and \U$4251 ( \4440 , \4422 , \4438 );
or \U$4252 ( \4441 , \4433 , \4439 , \4440 );
xor \U$4253 ( \4442 , \4264 , \4280 );
xor \U$4254 ( \4443 , \4442 , \4293 );
xor \U$4255 ( \4444 , \4312 , \4314 );
xor \U$4256 ( \4445 , \4444 , \4317 );
and \U$4257 ( \4446 , \4443 , \4445 );
xor \U$4258 ( \4447 , \4323 , \4325 );
and \U$4259 ( \4448 , \4445 , \4447 );
and \U$4260 ( \4449 , \4443 , \4447 );
or \U$4261 ( \4450 , \4446 , \4448 , \4449 );
and \U$4262 ( \4451 , \4441 , \4450 );
xor \U$4263 ( \4452 , \4331 , \4333 );
xor \U$4264 ( \4453 , \4452 , \4336 );
and \U$4265 ( \4454 , \4450 , \4453 );
and \U$4266 ( \4455 , \4441 , \4453 );
or \U$4267 ( \4456 , \4451 , \4454 , \4455 );
xor \U$4268 ( \4457 , \4329 , \4339 );
xor \U$4269 ( \4458 , \4457 , \4342 );
and \U$4270 ( \4459 , \4456 , \4458 );
xor \U$4271 ( \4460 , \4347 , \4349 );
and \U$4272 ( \4461 , \4458 , \4460 );
and \U$4273 ( \4462 , \4456 , \4460 );
or \U$4274 ( \4463 , \4459 , \4461 , \4462 );
and \U$4275 ( \4464 , \4370 , \4463 );
xor \U$4276 ( \4465 , \4370 , \4463 );
xor \U$4277 ( \4466 , \4456 , \4458 );
xor \U$4278 ( \4467 , \4466 , \4460 );
and \U$4279 ( \4468 , \2532 , \912 );
and \U$4280 ( \4469 , \2305 , \910 );
nor \U$4281 ( \4470 , \4468 , \4469 );
xnor \U$4282 ( \4471 , \4470 , \818 );
and \U$4283 ( \4472 , \2763 , \740 );
and \U$4284 ( \4473 , \2541 , \738 );
nor \U$4285 ( \4474 , \4472 , \4473 );
xnor \U$4286 ( \4475 , \4474 , \668 );
and \U$4287 ( \4476 , \4471 , \4475 );
nand \U$4288 ( \4477 , \2850 , \602 );
xnor \U$4289 ( \4478 , \4477 , \561 );
and \U$4290 ( \4479 , \4475 , \4478 );
and \U$4291 ( \4480 , \4471 , \4478 );
or \U$4292 ( \4481 , \4476 , \4479 , \4480 );
and \U$4293 ( \4482 , \2541 , \740 );
and \U$4294 ( \4483 , \2532 , \738 );
nor \U$4295 ( \4484 , \4482 , \4483 );
xnor \U$4296 ( \4485 , \4484 , \668 );
and \U$4297 ( \4486 , \4481 , \4485 );
and \U$4298 ( \4487 , \2850 , \604 );
and \U$4299 ( \4488 , \2763 , \602 );
nor \U$4300 ( \4489 , \4487 , \4488 );
xnor \U$4301 ( \4490 , \4489 , \561 );
and \U$4302 ( \4491 , \4485 , \4490 );
and \U$4303 ( \4492 , \4481 , \4490 );
or \U$4304 ( \4493 , \4486 , \4491 , \4492 );
and \U$4305 ( \4494 , \703 , \2913 );
and \U$4306 ( \4495 , \621 , \2910 );
nor \U$4307 ( \4496 , \4494 , \4495 );
xnor \U$4308 ( \4497 , \4496 , \2371 );
and \U$4309 ( \4498 , \841 , \2550 );
and \U$4310 ( \4499 , \777 , \2548 );
nor \U$4311 ( \4500 , \4498 , \4499 );
xnor \U$4312 ( \4501 , \4500 , \2374 );
and \U$4313 ( \4502 , \4497 , \4501 );
and \U$4314 ( \4503 , \4501 , \561 );
and \U$4315 ( \4504 , \4497 , \561 );
or \U$4316 ( \4505 , \4502 , \4503 , \4504 );
and \U$4317 ( \4506 , \1104 , \2261 );
and \U$4318 ( \4507 , \904 , \2259 );
nor \U$4319 ( \4508 , \4506 , \4507 );
xnor \U$4320 ( \4509 , \4508 , \2124 );
and \U$4321 ( \4510 , \1299 , \1955 );
and \U$4322 ( \4511 , \1194 , \1953 );
nor \U$4323 ( \4512 , \4510 , \4511 );
xnor \U$4324 ( \4513 , \4512 , \1835 );
and \U$4325 ( \4514 , \4509 , \4513 );
and \U$4326 ( \4515 , \1422 , \1742 );
and \U$4327 ( \4516 , \1304 , \1740 );
nor \U$4328 ( \4517 , \4515 , \4516 );
xnor \U$4329 ( \4518 , \4517 , \1610 );
and \U$4330 ( \4519 , \4513 , \4518 );
and \U$4331 ( \4520 , \4509 , \4518 );
or \U$4332 ( \4521 , \4514 , \4519 , \4520 );
and \U$4333 ( \4522 , \4505 , \4521 );
and \U$4334 ( \4523 , \1770 , \1476 );
and \U$4335 ( \4524 , \1537 , \1474 );
nor \U$4336 ( \4525 , \4523 , \4524 );
xnor \U$4337 ( \4526 , \4525 , \1363 );
and \U$4338 ( \4527 , \2023 , \1280 );
and \U$4339 ( \4528 , \1778 , \1278 );
nor \U$4340 ( \4529 , \4527 , \4528 );
xnor \U$4341 ( \4530 , \4529 , \1177 );
and \U$4342 ( \4531 , \4526 , \4530 );
and \U$4343 ( \4532 , \2161 , \1062 );
and \U$4344 ( \4533 , \2028 , \1060 );
nor \U$4345 ( \4534 , \4532 , \4533 );
xnor \U$4346 ( \4535 , \4534 , \984 );
and \U$4347 ( \4536 , \4530 , \4535 );
and \U$4348 ( \4537 , \4526 , \4535 );
or \U$4349 ( \4538 , \4531 , \4536 , \4537 );
and \U$4350 ( \4539 , \4521 , \4538 );
and \U$4351 ( \4540 , \4505 , \4538 );
or \U$4352 ( \4541 , \4522 , \4539 , \4540 );
and \U$4353 ( \4542 , \4493 , \4541 );
xor \U$4354 ( \4543 , \4374 , \4378 );
xor \U$4355 ( \4544 , \4543 , \4383 );
xor \U$4356 ( \4545 , \4390 , \4394 );
xor \U$4357 ( \4546 , \4545 , \4399 );
and \U$4358 ( \4547 , \4544 , \4546 );
xor \U$4359 ( \4548 , \4407 , \4411 );
xor \U$4360 ( \4549 , \4548 , \4416 );
and \U$4361 ( \4550 , \4546 , \4549 );
and \U$4362 ( \4551 , \4544 , \4549 );
or \U$4363 ( \4552 , \4547 , \4550 , \4551 );
and \U$4364 ( \4553 , \4541 , \4552 );
and \U$4365 ( \4554 , \4493 , \4552 );
or \U$4366 ( \4555 , \4542 , \4553 , \4554 );
xor \U$4367 ( \4556 , \4386 , \4402 );
xor \U$4368 ( \4557 , \4556 , \4419 );
xor \U$4369 ( \4558 , \4424 , \4426 );
xor \U$4370 ( \4559 , \4558 , \4429 );
and \U$4371 ( \4560 , \4557 , \4559 );
xor \U$4372 ( \4561 , \4435 , \4437 );
and \U$4373 ( \4562 , \4559 , \4561 );
and \U$4374 ( \4563 , \4557 , \4561 );
or \U$4375 ( \4564 , \4560 , \4562 , \4563 );
and \U$4376 ( \4565 , \4555 , \4564 );
xor \U$4377 ( \4566 , \4443 , \4445 );
xor \U$4378 ( \4567 , \4566 , \4447 );
and \U$4379 ( \4568 , \4564 , \4567 );
and \U$4380 ( \4569 , \4555 , \4567 );
or \U$4381 ( \4570 , \4565 , \4568 , \4569 );
xor \U$4382 ( \4571 , \4296 , \4320 );
xor \U$4383 ( \4572 , \4571 , \4326 );
and \U$4384 ( \4573 , \4570 , \4572 );
xor \U$4385 ( \4574 , \4441 , \4450 );
xor \U$4386 ( \4575 , \4574 , \4453 );
and \U$4387 ( \4576 , \4572 , \4575 );
and \U$4388 ( \4577 , \4570 , \4575 );
or \U$4389 ( \4578 , \4573 , \4576 , \4577 );
and \U$4390 ( \4579 , \4467 , \4578 );
xor \U$4391 ( \4580 , \4467 , \4578 );
xor \U$4392 ( \4581 , \4570 , \4572 );
xor \U$4393 ( \4582 , \4581 , \4575 );
and \U$4394 ( \4583 , \2028 , \1280 );
and \U$4395 ( \4584 , \2023 , \1278 );
nor \U$4396 ( \4585 , \4583 , \4584 );
xnor \U$4397 ( \4586 , \4585 , \1177 );
and \U$4398 ( \4587 , \2305 , \1062 );
and \U$4399 ( \4588 , \2161 , \1060 );
nor \U$4400 ( \4589 , \4587 , \4588 );
xnor \U$4401 ( \4590 , \4589 , \984 );
and \U$4402 ( \4591 , \4586 , \4590 );
and \U$4403 ( \4592 , \2541 , \912 );
and \U$4404 ( \4593 , \2532 , \910 );
nor \U$4405 ( \4594 , \4592 , \4593 );
xnor \U$4406 ( \4595 , \4594 , \818 );
and \U$4407 ( \4596 , \4590 , \4595 );
and \U$4408 ( \4597 , \4586 , \4595 );
or \U$4409 ( \4598 , \4591 , \4596 , \4597 );
and \U$4410 ( \4599 , \777 , \2913 );
and \U$4411 ( \4600 , \703 , \2910 );
nor \U$4412 ( \4601 , \4599 , \4600 );
xnor \U$4413 ( \4602 , \4601 , \2371 );
and \U$4414 ( \4603 , \904 , \2550 );
and \U$4415 ( \4604 , \841 , \2548 );
nor \U$4416 ( \4605 , \4603 , \4604 );
xnor \U$4417 ( \4606 , \4605 , \2374 );
and \U$4418 ( \4607 , \4602 , \4606 );
and \U$4419 ( \4608 , \1194 , \2261 );
and \U$4420 ( \4609 , \1104 , \2259 );
nor \U$4421 ( \4610 , \4608 , \4609 );
xnor \U$4422 ( \4611 , \4610 , \2124 );
and \U$4423 ( \4612 , \4606 , \4611 );
and \U$4424 ( \4613 , \4602 , \4611 );
or \U$4425 ( \4614 , \4607 , \4612 , \4613 );
and \U$4426 ( \4615 , \4598 , \4614 );
and \U$4427 ( \4616 , \1304 , \1955 );
and \U$4428 ( \4617 , \1299 , \1953 );
nor \U$4429 ( \4618 , \4616 , \4617 );
xnor \U$4430 ( \4619 , \4618 , \1835 );
and \U$4431 ( \4620 , \1537 , \1742 );
and \U$4432 ( \4621 , \1422 , \1740 );
nor \U$4433 ( \4622 , \4620 , \4621 );
xnor \U$4434 ( \4623 , \4622 , \1610 );
and \U$4435 ( \4624 , \4619 , \4623 );
and \U$4436 ( \4625 , \1778 , \1476 );
and \U$4437 ( \4626 , \1770 , \1474 );
nor \U$4438 ( \4627 , \4625 , \4626 );
xnor \U$4439 ( \4628 , \4627 , \1363 );
and \U$4440 ( \4629 , \4623 , \4628 );
and \U$4441 ( \4630 , \4619 , \4628 );
or \U$4442 ( \4631 , \4624 , \4629 , \4630 );
and \U$4443 ( \4632 , \4614 , \4631 );
and \U$4444 ( \4633 , \4598 , \4631 );
or \U$4445 ( \4634 , \4615 , \4632 , \4633 );
xor \U$4446 ( \4635 , \4509 , \4513 );
xor \U$4447 ( \4636 , \4635 , \4518 );
xor \U$4448 ( \4637 , \4471 , \4475 );
xor \U$4449 ( \4638 , \4637 , \4478 );
and \U$4450 ( \4639 , \4636 , \4638 );
xor \U$4451 ( \4640 , \4526 , \4530 );
xor \U$4452 ( \4641 , \4640 , \4535 );
and \U$4453 ( \4642 , \4638 , \4641 );
and \U$4454 ( \4643 , \4636 , \4641 );
or \U$4455 ( \4644 , \4639 , \4642 , \4643 );
and \U$4456 ( \4645 , \4634 , \4644 );
xor \U$4457 ( \4646 , \4544 , \4546 );
xor \U$4458 ( \4647 , \4646 , \4549 );
and \U$4459 ( \4648 , \4644 , \4647 );
and \U$4460 ( \4649 , \4634 , \4647 );
or \U$4461 ( \4650 , \4645 , \4648 , \4649 );
xor \U$4462 ( \4651 , \4493 , \4541 );
xor \U$4463 ( \4652 , \4651 , \4552 );
and \U$4464 ( \4653 , \4650 , \4652 );
xor \U$4465 ( \4654 , \4557 , \4559 );
xor \U$4466 ( \4655 , \4654 , \4561 );
and \U$4467 ( \4656 , \4652 , \4655 );
and \U$4468 ( \4657 , \4650 , \4655 );
or \U$4469 ( \4658 , \4653 , \4656 , \4657 );
xor \U$4470 ( \4659 , \4422 , \4432 );
xor \U$4471 ( \4660 , \4659 , \4438 );
and \U$4472 ( \4661 , \4658 , \4660 );
xor \U$4473 ( \4662 , \4555 , \4564 );
xor \U$4474 ( \4663 , \4662 , \4567 );
and \U$4475 ( \4664 , \4660 , \4663 );
and \U$4476 ( \4665 , \4658 , \4663 );
or \U$4477 ( \4666 , \4661 , \4664 , \4665 );
and \U$4478 ( \4667 , \4582 , \4666 );
xor \U$4479 ( \4668 , \4582 , \4666 );
xor \U$4480 ( \4669 , \4658 , \4660 );
xor \U$4481 ( \4670 , \4669 , \4663 );
and \U$4482 ( \4671 , \841 , \2913 );
and \U$4483 ( \4672 , \777 , \2910 );
nor \U$4484 ( \4673 , \4671 , \4672 );
xnor \U$4485 ( \4674 , \4673 , \2371 );
and \U$4486 ( \4675 , \1104 , \2550 );
and \U$4487 ( \4676 , \904 , \2548 );
nor \U$4488 ( \4677 , \4675 , \4676 );
xnor \U$4489 ( \4678 , \4677 , \2374 );
and \U$4490 ( \4679 , \4674 , \4678 );
and \U$4491 ( \4680 , \4678 , \668 );
and \U$4492 ( \4681 , \4674 , \668 );
or \U$4493 ( \4682 , \4679 , \4680 , \4681 );
and \U$4494 ( \4683 , \2023 , \1476 );
and \U$4495 ( \4684 , \1778 , \1474 );
nor \U$4496 ( \4685 , \4683 , \4684 );
xnor \U$4497 ( \4686 , \4685 , \1363 );
and \U$4498 ( \4687 , \2161 , \1280 );
and \U$4499 ( \4688 , \2028 , \1278 );
nor \U$4500 ( \4689 , \4687 , \4688 );
xnor \U$4501 ( \4690 , \4689 , \1177 );
and \U$4502 ( \4691 , \4686 , \4690 );
and \U$4503 ( \4692 , \2532 , \1062 );
and \U$4504 ( \4693 , \2305 , \1060 );
nor \U$4505 ( \4694 , \4692 , \4693 );
xnor \U$4506 ( \4695 , \4694 , \984 );
and \U$4507 ( \4696 , \4690 , \4695 );
and \U$4508 ( \4697 , \4686 , \4695 );
or \U$4509 ( \4698 , \4691 , \4696 , \4697 );
and \U$4510 ( \4699 , \4682 , \4698 );
and \U$4511 ( \4700 , \1299 , \2261 );
and \U$4512 ( \4701 , \1194 , \2259 );
nor \U$4513 ( \4702 , \4700 , \4701 );
xnor \U$4514 ( \4703 , \4702 , \2124 );
and \U$4515 ( \4704 , \1422 , \1955 );
and \U$4516 ( \4705 , \1304 , \1953 );
nor \U$4517 ( \4706 , \4704 , \4705 );
xnor \U$4518 ( \4707 , \4706 , \1835 );
and \U$4519 ( \4708 , \4703 , \4707 );
and \U$4520 ( \4709 , \1770 , \1742 );
and \U$4521 ( \4710 , \1537 , \1740 );
nor \U$4522 ( \4711 , \4709 , \4710 );
xnor \U$4523 ( \4712 , \4711 , \1610 );
and \U$4524 ( \4713 , \4707 , \4712 );
and \U$4525 ( \4714 , \4703 , \4712 );
or \U$4526 ( \4715 , \4708 , \4713 , \4714 );
and \U$4527 ( \4716 , \4698 , \4715 );
and \U$4528 ( \4717 , \4682 , \4715 );
or \U$4529 ( \4718 , \4699 , \4716 , \4717 );
and \U$4530 ( \4719 , \2850 , \740 );
and \U$4531 ( \4720 , \2763 , \738 );
nor \U$4532 ( \4721 , \4719 , \4720 );
xnor \U$4533 ( \4722 , \4721 , \668 );
xor \U$4534 ( \4723 , \4586 , \4590 );
xor \U$4535 ( \4724 , \4723 , \4595 );
and \U$4536 ( \4725 , \4722 , \4724 );
xor \U$4537 ( \4726 , \4619 , \4623 );
xor \U$4538 ( \4727 , \4726 , \4628 );
and \U$4539 ( \4728 , \4724 , \4727 );
and \U$4540 ( \4729 , \4722 , \4727 );
or \U$4541 ( \4730 , \4725 , \4728 , \4729 );
and \U$4542 ( \4731 , \4718 , \4730 );
xor \U$4543 ( \4732 , \4497 , \4501 );
xor \U$4544 ( \4733 , \4732 , \561 );
and \U$4545 ( \4734 , \4730 , \4733 );
and \U$4546 ( \4735 , \4718 , \4733 );
or \U$4547 ( \4736 , \4731 , \4734 , \4735 );
xor \U$4548 ( \4737 , \4598 , \4614 );
xor \U$4549 ( \4738 , \4737 , \4631 );
xor \U$4550 ( \4739 , \4636 , \4638 );
xor \U$4551 ( \4740 , \4739 , \4641 );
and \U$4552 ( \4741 , \4738 , \4740 );
and \U$4553 ( \4742 , \4736 , \4741 );
xor \U$4554 ( \4743 , \4481 , \4485 );
xor \U$4555 ( \4744 , \4743 , \4490 );
and \U$4556 ( \4745 , \4741 , \4744 );
and \U$4557 ( \4746 , \4736 , \4744 );
or \U$4558 ( \4747 , \4742 , \4745 , \4746 );
xor \U$4559 ( \4748 , \4505 , \4521 );
xor \U$4560 ( \4749 , \4748 , \4538 );
xor \U$4561 ( \4750 , \4634 , \4644 );
xor \U$4562 ( \4751 , \4750 , \4647 );
and \U$4563 ( \4752 , \4749 , \4751 );
and \U$4564 ( \4753 , \4747 , \4752 );
xor \U$4565 ( \4754 , \4650 , \4652 );
xor \U$4566 ( \4755 , \4754 , \4655 );
and \U$4567 ( \4756 , \4752 , \4755 );
and \U$4568 ( \4757 , \4747 , \4755 );
or \U$4569 ( \4758 , \4753 , \4756 , \4757 );
and \U$4570 ( \4759 , \4670 , \4758 );
xor \U$4571 ( \4760 , \4670 , \4758 );
xor \U$4572 ( \4761 , \4747 , \4752 );
xor \U$4573 ( \4762 , \4761 , \4755 );
and \U$4574 ( \4763 , \1537 , \1955 );
and \U$4575 ( \4764 , \1422 , \1953 );
nor \U$4576 ( \4765 , \4763 , \4764 );
xnor \U$4577 ( \4766 , \4765 , \1835 );
and \U$4578 ( \4767 , \1778 , \1742 );
and \U$4579 ( \4768 , \1770 , \1740 );
nor \U$4580 ( \4769 , \4767 , \4768 );
xnor \U$4581 ( \4770 , \4769 , \1610 );
and \U$4582 ( \4771 , \4766 , \4770 );
and \U$4583 ( \4772 , \2028 , \1476 );
and \U$4584 ( \4773 , \2023 , \1474 );
nor \U$4585 ( \4774 , \4772 , \4773 );
xnor \U$4586 ( \4775 , \4774 , \1363 );
and \U$4587 ( \4776 , \4770 , \4775 );
and \U$4588 ( \4777 , \4766 , \4775 );
or \U$4589 ( \4778 , \4771 , \4776 , \4777 );
and \U$4590 ( \4779 , \904 , \2913 );
and \U$4591 ( \4780 , \841 , \2910 );
nor \U$4592 ( \4781 , \4779 , \4780 );
xnor \U$4593 ( \4782 , \4781 , \2371 );
and \U$4594 ( \4783 , \1194 , \2550 );
and \U$4595 ( \4784 , \1104 , \2548 );
nor \U$4596 ( \4785 , \4783 , \4784 );
xnor \U$4597 ( \4786 , \4785 , \2374 );
and \U$4598 ( \4787 , \4782 , \4786 );
and \U$4599 ( \4788 , \1304 , \2261 );
and \U$4600 ( \4789 , \1299 , \2259 );
nor \U$4601 ( \4790 , \4788 , \4789 );
xnor \U$4602 ( \4791 , \4790 , \2124 );
and \U$4603 ( \4792 , \4786 , \4791 );
and \U$4604 ( \4793 , \4782 , \4791 );
or \U$4605 ( \4794 , \4787 , \4792 , \4793 );
and \U$4606 ( \4795 , \4778 , \4794 );
and \U$4607 ( \4796 , \2305 , \1280 );
and \U$4608 ( \4797 , \2161 , \1278 );
nor \U$4609 ( \4798 , \4796 , \4797 );
xnor \U$4610 ( \4799 , \4798 , \1177 );
and \U$4611 ( \4800 , \2541 , \1062 );
and \U$4612 ( \4801 , \2532 , \1060 );
nor \U$4613 ( \4802 , \4800 , \4801 );
xnor \U$4614 ( \4803 , \4802 , \984 );
and \U$4615 ( \4804 , \4799 , \4803 );
and \U$4616 ( \4805 , \2850 , \912 );
and \U$4617 ( \4806 , \2763 , \910 );
nor \U$4618 ( \4807 , \4805 , \4806 );
xnor \U$4619 ( \4808 , \4807 , \818 );
and \U$4620 ( \4809 , \4803 , \4808 );
and \U$4621 ( \4810 , \4799 , \4808 );
or \U$4622 ( \4811 , \4804 , \4809 , \4810 );
and \U$4623 ( \4812 , \4794 , \4811 );
and \U$4624 ( \4813 , \4778 , \4811 );
or \U$4625 ( \4814 , \4795 , \4812 , \4813 );
and \U$4626 ( \4815 , \2763 , \912 );
and \U$4627 ( \4816 , \2541 , \910 );
nor \U$4628 ( \4817 , \4815 , \4816 );
xnor \U$4629 ( \4818 , \4817 , \818 );
nand \U$4630 ( \4819 , \2850 , \738 );
xnor \U$4631 ( \4820 , \4819 , \668 );
and \U$4632 ( \4821 , \4818 , \4820 );
xor \U$4633 ( \4822 , \4686 , \4690 );
xor \U$4634 ( \4823 , \4822 , \4695 );
and \U$4635 ( \4824 , \4820 , \4823 );
and \U$4636 ( \4825 , \4818 , \4823 );
or \U$4637 ( \4826 , \4821 , \4824 , \4825 );
and \U$4638 ( \4827 , \4814 , \4826 );
xor \U$4639 ( \4828 , \4602 , \4606 );
xor \U$4640 ( \4829 , \4828 , \4611 );
and \U$4641 ( \4830 , \4826 , \4829 );
and \U$4642 ( \4831 , \4814 , \4829 );
or \U$4643 ( \4832 , \4827 , \4830 , \4831 );
xor \U$4644 ( \4833 , \4718 , \4730 );
xor \U$4645 ( \4834 , \4833 , \4733 );
and \U$4646 ( \4835 , \4832 , \4834 );
xor \U$4647 ( \4836 , \4738 , \4740 );
and \U$4648 ( \4837 , \4834 , \4836 );
and \U$4649 ( \4838 , \4832 , \4836 );
or \U$4650 ( \4839 , \4835 , \4837 , \4838 );
xor \U$4651 ( \4840 , \4736 , \4741 );
xor \U$4652 ( \4841 , \4840 , \4744 );
and \U$4653 ( \4842 , \4839 , \4841 );
xor \U$4654 ( \4843 , \4749 , \4751 );
and \U$4655 ( \4844 , \4841 , \4843 );
and \U$4656 ( \4845 , \4839 , \4843 );
or \U$4657 ( \4846 , \4842 , \4844 , \4845 );
and \U$4658 ( \4847 , \4762 , \4846 );
xor \U$4659 ( \4848 , \4762 , \4846 );
xor \U$4660 ( \4849 , \4839 , \4841 );
xor \U$4661 ( \4850 , \4849 , \4843 );
and \U$4662 ( \4851 , \1422 , \2261 );
and \U$4663 ( \4852 , \1304 , \2259 );
nor \U$4664 ( \4853 , \4851 , \4852 );
xnor \U$4665 ( \4854 , \4853 , \2124 );
and \U$4666 ( \4855 , \1770 , \1955 );
and \U$4667 ( \4856 , \1537 , \1953 );
nor \U$4668 ( \4857 , \4855 , \4856 );
xnor \U$4669 ( \4858 , \4857 , \1835 );
and \U$4670 ( \4859 , \4854 , \4858 );
and \U$4671 ( \4860 , \2023 , \1742 );
and \U$4672 ( \4861 , \1778 , \1740 );
nor \U$4673 ( \4862 , \4860 , \4861 );
xnor \U$4674 ( \4863 , \4862 , \1610 );
and \U$4675 ( \4864 , \4858 , \4863 );
and \U$4676 ( \4865 , \4854 , \4863 );
or \U$4677 ( \4866 , \4859 , \4864 , \4865 );
and \U$4678 ( \4867 , \1104 , \2913 );
and \U$4679 ( \4868 , \904 , \2910 );
nor \U$4680 ( \4869 , \4867 , \4868 );
xnor \U$4681 ( \4870 , \4869 , \2371 );
and \U$4682 ( \4871 , \1299 , \2550 );
and \U$4683 ( \4872 , \1194 , \2548 );
nor \U$4684 ( \4873 , \4871 , \4872 );
xnor \U$4685 ( \4874 , \4873 , \2374 );
and \U$4686 ( \4875 , \4870 , \4874 );
and \U$4687 ( \4876 , \4874 , \818 );
and \U$4688 ( \4877 , \4870 , \818 );
or \U$4689 ( \4878 , \4875 , \4876 , \4877 );
and \U$4690 ( \4879 , \4866 , \4878 );
and \U$4691 ( \4880 , \2161 , \1476 );
and \U$4692 ( \4881 , \2028 , \1474 );
nor \U$4693 ( \4882 , \4880 , \4881 );
xnor \U$4694 ( \4883 , \4882 , \1363 );
and \U$4695 ( \4884 , \2532 , \1280 );
and \U$4696 ( \4885 , \2305 , \1278 );
nor \U$4697 ( \4886 , \4884 , \4885 );
xnor \U$4698 ( \4887 , \4886 , \1177 );
and \U$4699 ( \4888 , \4883 , \4887 );
and \U$4700 ( \4889 , \2763 , \1062 );
and \U$4701 ( \4890 , \2541 , \1060 );
nor \U$4702 ( \4891 , \4889 , \4890 );
xnor \U$4703 ( \4892 , \4891 , \984 );
and \U$4704 ( \4893 , \4887 , \4892 );
and \U$4705 ( \4894 , \4883 , \4892 );
or \U$4706 ( \4895 , \4888 , \4893 , \4894 );
and \U$4707 ( \4896 , \4878 , \4895 );
and \U$4708 ( \4897 , \4866 , \4895 );
or \U$4709 ( \4898 , \4879 , \4896 , \4897 );
xor \U$4710 ( \4899 , \4766 , \4770 );
xor \U$4711 ( \4900 , \4899 , \4775 );
xor \U$4712 ( \4901 , \4782 , \4786 );
xor \U$4713 ( \4902 , \4901 , \4791 );
and \U$4714 ( \4903 , \4900 , \4902 );
xor \U$4715 ( \4904 , \4799 , \4803 );
xor \U$4716 ( \4905 , \4904 , \4808 );
and \U$4717 ( \4906 , \4902 , \4905 );
and \U$4718 ( \4907 , \4900 , \4905 );
or \U$4719 ( \4908 , \4903 , \4906 , \4907 );
and \U$4720 ( \4909 , \4898 , \4908 );
xor \U$4721 ( \4910 , \4703 , \4707 );
xor \U$4722 ( \4911 , \4910 , \4712 );
and \U$4723 ( \4912 , \4908 , \4911 );
and \U$4724 ( \4913 , \4898 , \4911 );
or \U$4725 ( \4914 , \4909 , \4912 , \4913 );
xor \U$4726 ( \4915 , \4674 , \4678 );
xor \U$4727 ( \4916 , \4915 , \668 );
xor \U$4728 ( \4917 , \4778 , \4794 );
xor \U$4729 ( \4918 , \4917 , \4811 );
and \U$4730 ( \4919 , \4916 , \4918 );
xor \U$4731 ( \4920 , \4818 , \4820 );
xor \U$4732 ( \4921 , \4920 , \4823 );
and \U$4733 ( \4922 , \4918 , \4921 );
and \U$4734 ( \4923 , \4916 , \4921 );
or \U$4735 ( \4924 , \4919 , \4922 , \4923 );
and \U$4736 ( \4925 , \4914 , \4924 );
xor \U$4737 ( \4926 , \4722 , \4724 );
xor \U$4738 ( \4927 , \4926 , \4727 );
and \U$4739 ( \4928 , \4924 , \4927 );
and \U$4740 ( \4929 , \4914 , \4927 );
or \U$4741 ( \4930 , \4925 , \4928 , \4929 );
xor \U$4742 ( \4931 , \4682 , \4698 );
xor \U$4743 ( \4932 , \4931 , \4715 );
xor \U$4744 ( \4933 , \4814 , \4826 );
xor \U$4745 ( \4934 , \4933 , \4829 );
and \U$4746 ( \4935 , \4932 , \4934 );
and \U$4747 ( \4936 , \4930 , \4935 );
xor \U$4748 ( \4937 , \4832 , \4834 );
xor \U$4749 ( \4938 , \4937 , \4836 );
and \U$4750 ( \4939 , \4935 , \4938 );
and \U$4751 ( \4940 , \4930 , \4938 );
or \U$4752 ( \4941 , \4936 , \4939 , \4940 );
and \U$4753 ( \4942 , \4850 , \4941 );
xor \U$4754 ( \4943 , \4850 , \4941 );
xor \U$4755 ( \4944 , \4930 , \4935 );
xor \U$4756 ( \4945 , \4944 , \4938 );
and \U$4757 ( \4946 , \1194 , \2913 );
and \U$4758 ( \4947 , \1104 , \2910 );
nor \U$4759 ( \4948 , \4946 , \4947 );
xnor \U$4760 ( \4949 , \4948 , \2371 );
and \U$4761 ( \4950 , \1304 , \2550 );
and \U$4762 ( \4951 , \1299 , \2548 );
nor \U$4763 ( \4952 , \4950 , \4951 );
xnor \U$4764 ( \4953 , \4952 , \2374 );
and \U$4765 ( \4954 , \4949 , \4953 );
and \U$4766 ( \4955 , \1537 , \2261 );
and \U$4767 ( \4956 , \1422 , \2259 );
nor \U$4768 ( \4957 , \4955 , \4956 );
xnor \U$4769 ( \4958 , \4957 , \2124 );
and \U$4770 ( \4959 , \4953 , \4958 );
and \U$4771 ( \4960 , \4949 , \4958 );
or \U$4772 ( \4961 , \4954 , \4959 , \4960 );
and \U$4773 ( \4962 , \1778 , \1955 );
and \U$4774 ( \4963 , \1770 , \1953 );
nor \U$4775 ( \4964 , \4962 , \4963 );
xnor \U$4776 ( \4965 , \4964 , \1835 );
and \U$4777 ( \4966 , \2028 , \1742 );
and \U$4778 ( \4967 , \2023 , \1740 );
nor \U$4779 ( \4968 , \4966 , \4967 );
xnor \U$4780 ( \4969 , \4968 , \1610 );
and \U$4781 ( \4970 , \4965 , \4969 );
and \U$4782 ( \4971 , \2305 , \1476 );
and \U$4783 ( \4972 , \2161 , \1474 );
nor \U$4784 ( \4973 , \4971 , \4972 );
xnor \U$4785 ( \4974 , \4973 , \1363 );
and \U$4786 ( \4975 , \4969 , \4974 );
and \U$4787 ( \4976 , \4965 , \4974 );
or \U$4788 ( \4977 , \4970 , \4975 , \4976 );
and \U$4789 ( \4978 , \4961 , \4977 );
and \U$4790 ( \4979 , \2541 , \1280 );
and \U$4791 ( \4980 , \2532 , \1278 );
nor \U$4792 ( \4981 , \4979 , \4980 );
xnor \U$4793 ( \4982 , \4981 , \1177 );
and \U$4794 ( \4983 , \2850 , \1062 );
and \U$4795 ( \4984 , \2763 , \1060 );
nor \U$4796 ( \4985 , \4983 , \4984 );
xnor \U$4797 ( \4986 , \4985 , \984 );
and \U$4798 ( \4987 , \4982 , \4986 );
and \U$4799 ( \4988 , \4977 , \4987 );
and \U$4800 ( \4989 , \4961 , \4987 );
or \U$4801 ( \4990 , \4978 , \4988 , \4989 );
nand \U$4802 ( \4991 , \2850 , \910 );
xnor \U$4803 ( \4992 , \4991 , \818 );
xor \U$4804 ( \4993 , \4854 , \4858 );
xor \U$4805 ( \4994 , \4993 , \4863 );
and \U$4806 ( \4995 , \4992 , \4994 );
xor \U$4807 ( \4996 , \4883 , \4887 );
xor \U$4808 ( \4997 , \4996 , \4892 );
and \U$4809 ( \4998 , \4994 , \4997 );
and \U$4810 ( \4999 , \4992 , \4997 );
or \U$4811 ( \5000 , \4995 , \4998 , \4999 );
and \U$4812 ( \5001 , \4990 , \5000 );
xor \U$4813 ( \5002 , \4900 , \4902 );
xor \U$4814 ( \5003 , \5002 , \4905 );
and \U$4815 ( \5004 , \5000 , \5003 );
and \U$4816 ( \5005 , \4990 , \5003 );
or \U$4817 ( \5006 , \5001 , \5004 , \5005 );
xor \U$4818 ( \5007 , \4898 , \4908 );
xor \U$4819 ( \5008 , \5007 , \4911 );
and \U$4820 ( \5009 , \5006 , \5008 );
xor \U$4821 ( \5010 , \4916 , \4918 );
xor \U$4822 ( \5011 , \5010 , \4921 );
and \U$4823 ( \5012 , \5008 , \5011 );
and \U$4824 ( \5013 , \5006 , \5011 );
or \U$4825 ( \5014 , \5009 , \5012 , \5013 );
xor \U$4826 ( \5015 , \4914 , \4924 );
xor \U$4827 ( \5016 , \5015 , \4927 );
and \U$4828 ( \5017 , \5014 , \5016 );
xor \U$4829 ( \5018 , \4932 , \4934 );
and \U$4830 ( \5019 , \5016 , \5018 );
and \U$4831 ( \5020 , \5014 , \5018 );
or \U$4832 ( \5021 , \5017 , \5019 , \5020 );
and \U$4833 ( \5022 , \4945 , \5021 );
xor \U$4834 ( \5023 , \4945 , \5021 );
xor \U$4835 ( \5024 , \5014 , \5016 );
xor \U$4836 ( \5025 , \5024 , \5018 );
and \U$4837 ( \5026 , \2532 , \1476 );
and \U$4838 ( \5027 , \2305 , \1474 );
nor \U$4839 ( \5028 , \5026 , \5027 );
xnor \U$4840 ( \5029 , \5028 , \1363 );
and \U$4841 ( \5030 , \2763 , \1280 );
and \U$4842 ( \5031 , \2541 , \1278 );
nor \U$4843 ( \5032 , \5030 , \5031 );
xnor \U$4844 ( \5033 , \5032 , \1177 );
and \U$4845 ( \5034 , \5029 , \5033 );
nand \U$4846 ( \5035 , \2850 , \1060 );
xnor \U$4847 ( \5036 , \5035 , \984 );
and \U$4848 ( \5037 , \5033 , \5036 );
and \U$4849 ( \5038 , \5029 , \5036 );
or \U$4850 ( \5039 , \5034 , \5037 , \5038 );
and \U$4851 ( \5040 , \1299 , \2913 );
and \U$4852 ( \5041 , \1194 , \2910 );
nor \U$4853 ( \5042 , \5040 , \5041 );
xnor \U$4854 ( \5043 , \5042 , \2371 );
and \U$4855 ( \5044 , \1422 , \2550 );
and \U$4856 ( \5045 , \1304 , \2548 );
nor \U$4857 ( \5046 , \5044 , \5045 );
xnor \U$4858 ( \5047 , \5046 , \2374 );
and \U$4859 ( \5048 , \5043 , \5047 );
and \U$4860 ( \5049 , \5047 , \984 );
and \U$4861 ( \5050 , \5043 , \984 );
or \U$4862 ( \5051 , \5048 , \5049 , \5050 );
and \U$4863 ( \5052 , \5039 , \5051 );
and \U$4864 ( \5053 , \1770 , \2261 );
and \U$4865 ( \5054 , \1537 , \2259 );
nor \U$4866 ( \5055 , \5053 , \5054 );
xnor \U$4867 ( \5056 , \5055 , \2124 );
and \U$4868 ( \5057 , \2023 , \1955 );
and \U$4869 ( \5058 , \1778 , \1953 );
nor \U$4870 ( \5059 , \5057 , \5058 );
xnor \U$4871 ( \5060 , \5059 , \1835 );
and \U$4872 ( \5061 , \5056 , \5060 );
and \U$4873 ( \5062 , \2161 , \1742 );
and \U$4874 ( \5063 , \2028 , \1740 );
nor \U$4875 ( \5064 , \5062 , \5063 );
xnor \U$4876 ( \5065 , \5064 , \1610 );
and \U$4877 ( \5066 , \5060 , \5065 );
and \U$4878 ( \5067 , \5056 , \5065 );
or \U$4879 ( \5068 , \5061 , \5066 , \5067 );
and \U$4880 ( \5069 , \5051 , \5068 );
and \U$4881 ( \5070 , \5039 , \5068 );
or \U$4882 ( \5071 , \5052 , \5069 , \5070 );
xor \U$4883 ( \5072 , \4949 , \4953 );
xor \U$4884 ( \5073 , \5072 , \4958 );
xor \U$4885 ( \5074 , \4965 , \4969 );
xor \U$4886 ( \5075 , \5074 , \4974 );
and \U$4887 ( \5076 , \5073 , \5075 );
xor \U$4888 ( \5077 , \4982 , \4986 );
and \U$4889 ( \5078 , \5075 , \5077 );
and \U$4890 ( \5079 , \5073 , \5077 );
or \U$4891 ( \5080 , \5076 , \5078 , \5079 );
and \U$4892 ( \5081 , \5071 , \5080 );
xor \U$4893 ( \5082 , \4870 , \4874 );
xor \U$4894 ( \5083 , \5082 , \818 );
and \U$4895 ( \5084 , \5080 , \5083 );
and \U$4896 ( \5085 , \5071 , \5083 );
or \U$4897 ( \5086 , \5081 , \5084 , \5085 );
xor \U$4898 ( \5087 , \4961 , \4977 );
xor \U$4899 ( \5088 , \5087 , \4987 );
xor \U$4900 ( \5089 , \4992 , \4994 );
xor \U$4901 ( \5090 , \5089 , \4997 );
and \U$4902 ( \5091 , \5088 , \5090 );
and \U$4903 ( \5092 , \5086 , \5091 );
xor \U$4904 ( \5093 , \4866 , \4878 );
xor \U$4905 ( \5094 , \5093 , \4895 );
and \U$4906 ( \5095 , \5091 , \5094 );
and \U$4907 ( \5096 , \5086 , \5094 );
or \U$4908 ( \5097 , \5092 , \5095 , \5096 );
xor \U$4909 ( \5098 , \5006 , \5008 );
xor \U$4910 ( \5099 , \5098 , \5011 );
and \U$4911 ( \5100 , \5097 , \5099 );
and \U$4912 ( \5101 , \5025 , \5100 );
xor \U$4913 ( \5102 , \5025 , \5100 );
xor \U$4914 ( \5103 , \5097 , \5099 );
xor \U$4915 ( \5104 , \5086 , \5091 );
xor \U$4916 ( \5105 , \5104 , \5094 );
xor \U$4917 ( \5106 , \4990 , \5000 );
xor \U$4918 ( \5107 , \5106 , \5003 );
and \U$4919 ( \5108 , \5105 , \5107 );
and \U$4920 ( \5109 , \5103 , \5108 );
xor \U$4921 ( \5110 , \5103 , \5108 );
xor \U$4922 ( \5111 , \5105 , \5107 );
and \U$4923 ( \5112 , \1304 , \2913 );
and \U$4924 ( \5113 , \1299 , \2910 );
nor \U$4925 ( \5114 , \5112 , \5113 );
xnor \U$4926 ( \5115 , \5114 , \2371 );
and \U$4927 ( \5116 , \1537 , \2550 );
and \U$4928 ( \5117 , \1422 , \2548 );
nor \U$4929 ( \5118 , \5116 , \5117 );
xnor \U$4930 ( \5119 , \5118 , \2374 );
and \U$4931 ( \5120 , \5115 , \5119 );
and \U$4932 ( \5121 , \1778 , \2261 );
and \U$4933 ( \5122 , \1770 , \2259 );
nor \U$4934 ( \5123 , \5121 , \5122 );
xnor \U$4935 ( \5124 , \5123 , \2124 );
and \U$4936 ( \5125 , \5119 , \5124 );
and \U$4937 ( \5126 , \5115 , \5124 );
or \U$4938 ( \5127 , \5120 , \5125 , \5126 );
and \U$4939 ( \5128 , \2028 , \1955 );
and \U$4940 ( \5129 , \2023 , \1953 );
nor \U$4941 ( \5130 , \5128 , \5129 );
xnor \U$4942 ( \5131 , \5130 , \1835 );
and \U$4943 ( \5132 , \2305 , \1742 );
and \U$4944 ( \5133 , \2161 , \1740 );
nor \U$4945 ( \5134 , \5132 , \5133 );
xnor \U$4946 ( \5135 , \5134 , \1610 );
and \U$4947 ( \5136 , \5131 , \5135 );
and \U$4948 ( \5137 , \2541 , \1476 );
and \U$4949 ( \5138 , \2532 , \1474 );
nor \U$4950 ( \5139 , \5137 , \5138 );
xnor \U$4951 ( \5140 , \5139 , \1363 );
and \U$4952 ( \5141 , \5135 , \5140 );
and \U$4953 ( \5142 , \5131 , \5140 );
or \U$4954 ( \5143 , \5136 , \5141 , \5142 );
and \U$4955 ( \5144 , \5127 , \5143 );
xor \U$4956 ( \5145 , \5029 , \5033 );
xor \U$4957 ( \5146 , \5145 , \5036 );
and \U$4958 ( \5147 , \5143 , \5146 );
and \U$4959 ( \5148 , \5127 , \5146 );
or \U$4960 ( \5149 , \5144 , \5147 , \5148 );
xor \U$4961 ( \5150 , \5043 , \5047 );
xor \U$4962 ( \5151 , \5150 , \984 );
xor \U$4963 ( \5152 , \5056 , \5060 );
xor \U$4964 ( \5153 , \5152 , \5065 );
and \U$4965 ( \5154 , \5151 , \5153 );
and \U$4966 ( \5155 , \5149 , \5154 );
xor \U$4967 ( \5156 , \5073 , \5075 );
xor \U$4968 ( \5157 , \5156 , \5077 );
and \U$4969 ( \5158 , \5154 , \5157 );
and \U$4970 ( \5159 , \5149 , \5157 );
or \U$4971 ( \5160 , \5155 , \5158 , \5159 );
xor \U$4972 ( \5161 , \5071 , \5080 );
xor \U$4973 ( \5162 , \5161 , \5083 );
and \U$4974 ( \5163 , \5160 , \5162 );
xor \U$4975 ( \5164 , \5088 , \5090 );
and \U$4976 ( \5165 , \5162 , \5164 );
and \U$4977 ( \5166 , \5160 , \5164 );
or \U$4978 ( \5167 , \5163 , \5165 , \5166 );
and \U$4979 ( \5168 , \5111 , \5167 );
xor \U$4980 ( \5169 , \5111 , \5167 );
xor \U$4981 ( \5170 , \5160 , \5162 );
xor \U$4982 ( \5171 , \5170 , \5164 );
and \U$4983 ( \5172 , \1422 , \2913 );
and \U$4984 ( \5173 , \1304 , \2910 );
nor \U$4985 ( \5174 , \5172 , \5173 );
xnor \U$4986 ( \5175 , \5174 , \2371 );
and \U$4987 ( \5176 , \1770 , \2550 );
and \U$4988 ( \5177 , \1537 , \2548 );
nor \U$4989 ( \5178 , \5176 , \5177 );
xnor \U$4990 ( \5179 , \5178 , \2374 );
and \U$4991 ( \5180 , \5175 , \5179 );
and \U$4992 ( \5181 , \5179 , \1177 );
and \U$4993 ( \5182 , \5175 , \1177 );
or \U$4994 ( \5183 , \5180 , \5181 , \5182 );
and \U$4995 ( \5184 , \2023 , \2261 );
and \U$4996 ( \5185 , \1778 , \2259 );
nor \U$4997 ( \5186 , \5184 , \5185 );
xnor \U$4998 ( \5187 , \5186 , \2124 );
and \U$4999 ( \5188 , \2161 , \1955 );
and \U$5000 ( \5189 , \2028 , \1953 );
nor \U$5001 ( \5190 , \5188 , \5189 );
xnor \U$5002 ( \5191 , \5190 , \1835 );
and \U$5003 ( \5192 , \5187 , \5191 );
and \U$5004 ( \5193 , \2532 , \1742 );
and \U$5005 ( \5194 , \2305 , \1740 );
nor \U$5006 ( \5195 , \5193 , \5194 );
xnor \U$5007 ( \5196 , \5195 , \1610 );
and \U$5008 ( \5197 , \5191 , \5196 );
and \U$5009 ( \5198 , \5187 , \5196 );
or \U$5010 ( \5199 , \5192 , \5197 , \5198 );
and \U$5011 ( \5200 , \5183 , \5199 );
and \U$5012 ( \5201 , \2850 , \1280 );
and \U$5013 ( \5202 , \2763 , \1278 );
nor \U$5014 ( \5203 , \5201 , \5202 );
xnor \U$5015 ( \5204 , \5203 , \1177 );
and \U$5016 ( \5205 , \5199 , \5204 );
and \U$5017 ( \5206 , \5183 , \5204 );
or \U$5018 ( \5207 , \5200 , \5205 , \5206 );
xor \U$5019 ( \5208 , \5127 , \5143 );
xor \U$5020 ( \5209 , \5208 , \5146 );
and \U$5021 ( \5210 , \5207 , \5209 );
xor \U$5022 ( \5211 , \5151 , \5153 );
and \U$5023 ( \5212 , \5209 , \5211 );
and \U$5024 ( \5213 , \5207 , \5211 );
or \U$5025 ( \5214 , \5210 , \5212 , \5213 );
xor \U$5026 ( \5215 , \5039 , \5051 );
xor \U$5027 ( \5216 , \5215 , \5068 );
and \U$5028 ( \5217 , \5214 , \5216 );
xor \U$5029 ( \5218 , \5149 , \5154 );
xor \U$5030 ( \5219 , \5218 , \5157 );
and \U$5031 ( \5220 , \5216 , \5219 );
and \U$5032 ( \5221 , \5214 , \5219 );
or \U$5033 ( \5222 , \5217 , \5220 , \5221 );
and \U$5034 ( \5223 , \5171 , \5222 );
xor \U$5035 ( \5224 , \5171 , \5222 );
xor \U$5036 ( \5225 , \5214 , \5216 );
xor \U$5037 ( \5226 , \5225 , \5219 );
and \U$5038 ( \5227 , \2305 , \1955 );
and \U$5039 ( \5228 , \2161 , \1953 );
nor \U$5040 ( \5229 , \5227 , \5228 );
xnor \U$5041 ( \5230 , \5229 , \1835 );
and \U$5042 ( \5231 , \2541 , \1742 );
and \U$5043 ( \5232 , \2532 , \1740 );
nor \U$5044 ( \5233 , \5231 , \5232 );
xnor \U$5045 ( \5234 , \5233 , \1610 );
and \U$5046 ( \5235 , \5230 , \5234 );
and \U$5047 ( \5236 , \2850 , \1476 );
and \U$5048 ( \5237 , \2763 , \1474 );
nor \U$5049 ( \5238 , \5236 , \5237 );
xnor \U$5050 ( \5239 , \5238 , \1363 );
and \U$5051 ( \5240 , \5234 , \5239 );
and \U$5052 ( \5241 , \5230 , \5239 );
or \U$5053 ( \5242 , \5235 , \5240 , \5241 );
and \U$5054 ( \5243 , \1537 , \2913 );
and \U$5055 ( \5244 , \1422 , \2910 );
nor \U$5056 ( \5245 , \5243 , \5244 );
xnor \U$5057 ( \5246 , \5245 , \2371 );
and \U$5058 ( \5247 , \1778 , \2550 );
and \U$5059 ( \5248 , \1770 , \2548 );
nor \U$5060 ( \5249 , \5247 , \5248 );
xnor \U$5061 ( \5250 , \5249 , \2374 );
and \U$5062 ( \5251 , \5246 , \5250 );
and \U$5063 ( \5252 , \2028 , \2261 );
and \U$5064 ( \5253 , \2023 , \2259 );
nor \U$5065 ( \5254 , \5252 , \5253 );
xnor \U$5066 ( \5255 , \5254 , \2124 );
and \U$5067 ( \5256 , \5250 , \5255 );
and \U$5068 ( \5257 , \5246 , \5255 );
or \U$5069 ( \5258 , \5251 , \5256 , \5257 );
and \U$5070 ( \5259 , \5242 , \5258 );
and \U$5071 ( \5260 , \2763 , \1476 );
and \U$5072 ( \5261 , \2541 , \1474 );
nor \U$5073 ( \5262 , \5260 , \5261 );
xnor \U$5074 ( \5263 , \5262 , \1363 );
and \U$5075 ( \5264 , \5258 , \5263 );
and \U$5076 ( \5265 , \5242 , \5263 );
or \U$5077 ( \5266 , \5259 , \5264 , \5265 );
nand \U$5078 ( \5267 , \2850 , \1278 );
xnor \U$5079 ( \5268 , \5267 , \1177 );
xor \U$5080 ( \5269 , \5175 , \5179 );
xor \U$5081 ( \5270 , \5269 , \1177 );
and \U$5082 ( \5271 , \5268 , \5270 );
xor \U$5083 ( \5272 , \5187 , \5191 );
xor \U$5084 ( \5273 , \5272 , \5196 );
and \U$5085 ( \5274 , \5270 , \5273 );
and \U$5086 ( \5275 , \5268 , \5273 );
or \U$5087 ( \5276 , \5271 , \5274 , \5275 );
and \U$5088 ( \5277 , \5266 , \5276 );
xor \U$5089 ( \5278 , \5131 , \5135 );
xor \U$5090 ( \5279 , \5278 , \5140 );
and \U$5091 ( \5280 , \5276 , \5279 );
and \U$5092 ( \5281 , \5266 , \5279 );
or \U$5093 ( \5282 , \5277 , \5280 , \5281 );
xor \U$5094 ( \5283 , \5115 , \5119 );
xor \U$5095 ( \5284 , \5283 , \5124 );
xor \U$5096 ( \5285 , \5183 , \5199 );
xor \U$5097 ( \5286 , \5285 , \5204 );
and \U$5098 ( \5287 , \5284 , \5286 );
and \U$5099 ( \5288 , \5282 , \5287 );
xor \U$5100 ( \5289 , \5207 , \5209 );
xor \U$5101 ( \5290 , \5289 , \5211 );
and \U$5102 ( \5291 , \5287 , \5290 );
and \U$5103 ( \5292 , \5282 , \5290 );
or \U$5104 ( \5293 , \5288 , \5291 , \5292 );
and \U$5105 ( \5294 , \5226 , \5293 );
xor \U$5106 ( \5295 , \5226 , \5293 );
xor \U$5107 ( \5296 , \5282 , \5287 );
xor \U$5108 ( \5297 , \5296 , \5290 );
and \U$5109 ( \5298 , \2161 , \2261 );
and \U$5110 ( \5299 , \2028 , \2259 );
nor \U$5111 ( \5300 , \5298 , \5299 );
xnor \U$5112 ( \5301 , \5300 , \2124 );
and \U$5113 ( \5302 , \2532 , \1955 );
and \U$5114 ( \5303 , \2305 , \1953 );
nor \U$5115 ( \5304 , \5302 , \5303 );
xnor \U$5116 ( \5305 , \5304 , \1835 );
and \U$5117 ( \5306 , \5301 , \5305 );
and \U$5118 ( \5307 , \2763 , \1742 );
and \U$5119 ( \5308 , \2541 , \1740 );
nor \U$5120 ( \5309 , \5307 , \5308 );
xnor \U$5121 ( \5310 , \5309 , \1610 );
and \U$5122 ( \5311 , \5305 , \5310 );
and \U$5123 ( \5312 , \5301 , \5310 );
or \U$5124 ( \5313 , \5306 , \5311 , \5312 );
and \U$5125 ( \5314 , \1770 , \2913 );
and \U$5126 ( \5315 , \1537 , \2910 );
nor \U$5127 ( \5316 , \5314 , \5315 );
xnor \U$5128 ( \5317 , \5316 , \2371 );
and \U$5129 ( \5318 , \2023 , \2550 );
and \U$5130 ( \5319 , \1778 , \2548 );
nor \U$5131 ( \5320 , \5318 , \5319 );
xnor \U$5132 ( \5321 , \5320 , \2374 );
and \U$5133 ( \5322 , \5317 , \5321 );
and \U$5134 ( \5323 , \5321 , \1363 );
and \U$5135 ( \5324 , \5317 , \1363 );
or \U$5136 ( \5325 , \5322 , \5323 , \5324 );
and \U$5137 ( \5326 , \5313 , \5325 );
xor \U$5138 ( \5327 , \5230 , \5234 );
xor \U$5139 ( \5328 , \5327 , \5239 );
and \U$5140 ( \5329 , \5325 , \5328 );
and \U$5141 ( \5330 , \5313 , \5328 );
or \U$5142 ( \5331 , \5326 , \5329 , \5330 );
xor \U$5143 ( \5332 , \5242 , \5258 );
xor \U$5144 ( \5333 , \5332 , \5263 );
and \U$5145 ( \5334 , \5331 , \5333 );
xor \U$5146 ( \5335 , \5268 , \5270 );
xor \U$5147 ( \5336 , \5335 , \5273 );
and \U$5148 ( \5337 , \5333 , \5336 );
and \U$5149 ( \5338 , \5331 , \5336 );
or \U$5150 ( \5339 , \5334 , \5337 , \5338 );
xor \U$5151 ( \5340 , \5266 , \5276 );
xor \U$5152 ( \5341 , \5340 , \5279 );
and \U$5153 ( \5342 , \5339 , \5341 );
xor \U$5154 ( \5343 , \5284 , \5286 );
and \U$5155 ( \5344 , \5341 , \5343 );
and \U$5156 ( \5345 , \5339 , \5343 );
or \U$5157 ( \5346 , \5342 , \5344 , \5345 );
and \U$5158 ( \5347 , \5297 , \5346 );
xor \U$5159 ( \5348 , \5297 , \5346 );
xor \U$5160 ( \5349 , \5339 , \5341 );
xor \U$5161 ( \5350 , \5349 , \5343 );
and \U$5162 ( \5351 , \1778 , \2913 );
and \U$5163 ( \5352 , \1770 , \2910 );
nor \U$5164 ( \5353 , \5351 , \5352 );
xnor \U$5165 ( \5354 , \5353 , \2371 );
and \U$5166 ( \5355 , \2028 , \2550 );
and \U$5167 ( \5356 , \2023 , \2548 );
nor \U$5168 ( \5357 , \5355 , \5356 );
xnor \U$5169 ( \5358 , \5357 , \2374 );
and \U$5170 ( \5359 , \5354 , \5358 );
and \U$5171 ( \5360 , \2305 , \2261 );
and \U$5172 ( \5361 , \2161 , \2259 );
nor \U$5173 ( \5362 , \5360 , \5361 );
xnor \U$5174 ( \5363 , \5362 , \2124 );
and \U$5175 ( \5364 , \5358 , \5363 );
and \U$5176 ( \5365 , \5354 , \5363 );
or \U$5177 ( \5366 , \5359 , \5364 , \5365 );
nand \U$5178 ( \5367 , \2850 , \1474 );
xnor \U$5179 ( \5368 , \5367 , \1363 );
and \U$5180 ( \5369 , \5366 , \5368 );
xor \U$5181 ( \5370 , \5301 , \5305 );
xor \U$5182 ( \5371 , \5370 , \5310 );
and \U$5183 ( \5372 , \5368 , \5371 );
and \U$5184 ( \5373 , \5366 , \5371 );
or \U$5185 ( \5374 , \5369 , \5372 , \5373 );
xor \U$5186 ( \5375 , \5246 , \5250 );
xor \U$5187 ( \5376 , \5375 , \5255 );
and \U$5188 ( \5377 , \5374 , \5376 );
xor \U$5189 ( \5378 , \5313 , \5325 );
xor \U$5190 ( \5379 , \5378 , \5328 );
and \U$5191 ( \5380 , \5376 , \5379 );
and \U$5192 ( \5381 , \5374 , \5379 );
or \U$5193 ( \5382 , \5377 , \5380 , \5381 );
xor \U$5194 ( \5383 , \5331 , \5333 );
xor \U$5195 ( \5384 , \5383 , \5336 );
and \U$5196 ( \5385 , \5382 , \5384 );
and \U$5197 ( \5386 , \5350 , \5385 );
xor \U$5198 ( \5387 , \5350 , \5385 );
xor \U$5199 ( \5388 , \5382 , \5384 );
and \U$5200 ( \5389 , \2532 , \2261 );
and \U$5201 ( \5390 , \2305 , \2259 );
nor \U$5202 ( \5391 , \5389 , \5390 );
xnor \U$5203 ( \5392 , \5391 , \2124 );
and \U$5204 ( \5393 , \2763 , \1955 );
and \U$5205 ( \5394 , \2541 , \1953 );
nor \U$5206 ( \5395 , \5393 , \5394 );
xnor \U$5207 ( \5396 , \5395 , \1835 );
and \U$5208 ( \5397 , \5392 , \5396 );
nand \U$5209 ( \5398 , \2850 , \1740 );
xnor \U$5210 ( \5399 , \5398 , \1610 );
and \U$5211 ( \5400 , \5396 , \5399 );
and \U$5212 ( \5401 , \5392 , \5399 );
or \U$5213 ( \5402 , \5397 , \5400 , \5401 );
and \U$5214 ( \5403 , \2023 , \2913 );
and \U$5215 ( \5404 , \1778 , \2910 );
nor \U$5216 ( \5405 , \5403 , \5404 );
xnor \U$5217 ( \5406 , \5405 , \2371 );
and \U$5218 ( \5407 , \2161 , \2550 );
and \U$5219 ( \5408 , \2028 , \2548 );
nor \U$5220 ( \5409 , \5407 , \5408 );
xnor \U$5221 ( \5410 , \5409 , \2374 );
and \U$5222 ( \5411 , \5406 , \5410 );
and \U$5223 ( \5412 , \5410 , \1610 );
and \U$5224 ( \5413 , \5406 , \1610 );
or \U$5225 ( \5414 , \5411 , \5412 , \5413 );
and \U$5226 ( \5415 , \5402 , \5414 );
and \U$5227 ( \5416 , \2541 , \1955 );
and \U$5228 ( \5417 , \2532 , \1953 );
nor \U$5229 ( \5418 , \5416 , \5417 );
xnor \U$5230 ( \5419 , \5418 , \1835 );
and \U$5231 ( \5420 , \5414 , \5419 );
and \U$5232 ( \5421 , \5402 , \5419 );
or \U$5233 ( \5422 , \5415 , \5420 , \5421 );
and \U$5234 ( \5423 , \2850 , \1742 );
and \U$5235 ( \5424 , \2763 , \1740 );
nor \U$5236 ( \5425 , \5423 , \5424 );
xnor \U$5237 ( \5426 , \5425 , \1610 );
xor \U$5238 ( \5427 , \5354 , \5358 );
xor \U$5239 ( \5428 , \5427 , \5363 );
and \U$5240 ( \5429 , \5426 , \5428 );
and \U$5241 ( \5430 , \5422 , \5429 );
xor \U$5242 ( \5431 , \5317 , \5321 );
xor \U$5243 ( \5432 , \5431 , \1363 );
and \U$5244 ( \5433 , \5429 , \5432 );
and \U$5245 ( \5434 , \5422 , \5432 );
or \U$5246 ( \5435 , \5430 , \5433 , \5434 );
xor \U$5247 ( \5436 , \5374 , \5376 );
xor \U$5248 ( \5437 , \5436 , \5379 );
and \U$5249 ( \5438 , \5435 , \5437 );
and \U$5250 ( \5439 , \5388 , \5438 );
xor \U$5251 ( \5440 , \5388 , \5438 );
xor \U$5252 ( \5441 , \5435 , \5437 );
xor \U$5253 ( \5442 , \5366 , \5368 );
xor \U$5254 ( \5443 , \5442 , \5371 );
xor \U$5255 ( \5444 , \5422 , \5429 );
xor \U$5256 ( \5445 , \5444 , \5432 );
and \U$5257 ( \5446 , \5443 , \5445 );
and \U$5258 ( \5447 , \5441 , \5446 );
xor \U$5259 ( \5448 , \5441 , \5446 );
xor \U$5260 ( \5449 , \5443 , \5445 );
and \U$5261 ( \5450 , \2028 , \2913 );
and \U$5262 ( \5451 , \2023 , \2910 );
nor \U$5263 ( \5452 , \5450 , \5451 );
xnor \U$5264 ( \5453 , \5452 , \2371 );
and \U$5265 ( \5454 , \2305 , \2550 );
and \U$5266 ( \5455 , \2161 , \2548 );
nor \U$5267 ( \5456 , \5454 , \5455 );
xnor \U$5268 ( \5457 , \5456 , \2374 );
and \U$5269 ( \5458 , \5453 , \5457 );
and \U$5270 ( \5459 , \2541 , \2261 );
and \U$5271 ( \5460 , \2532 , \2259 );
nor \U$5272 ( \5461 , \5459 , \5460 );
xnor \U$5273 ( \5462 , \5461 , \2124 );
and \U$5274 ( \5463 , \5457 , \5462 );
and \U$5275 ( \5464 , \5453 , \5462 );
or \U$5276 ( \5465 , \5458 , \5463 , \5464 );
xor \U$5277 ( \5466 , \5392 , \5396 );
xor \U$5278 ( \5467 , \5466 , \5399 );
and \U$5279 ( \5468 , \5465 , \5467 );
xor \U$5280 ( \5469 , \5406 , \5410 );
xor \U$5281 ( \5470 , \5469 , \1610 );
and \U$5282 ( \5471 , \5467 , \5470 );
and \U$5283 ( \5472 , \5465 , \5470 );
or \U$5284 ( \5473 , \5468 , \5471 , \5472 );
xor \U$5285 ( \5474 , \5402 , \5414 );
xor \U$5286 ( \5475 , \5474 , \5419 );
and \U$5287 ( \5476 , \5473 , \5475 );
xor \U$5288 ( \5477 , \5426 , \5428 );
and \U$5289 ( \5478 , \5475 , \5477 );
and \U$5290 ( \5479 , \5473 , \5477 );
or \U$5291 ( \5480 , \5476 , \5478 , \5479 );
and \U$5292 ( \5481 , \5449 , \5480 );
xor \U$5293 ( \5482 , \5449 , \5480 );
xor \U$5294 ( \5483 , \5473 , \5475 );
xor \U$5295 ( \5484 , \5483 , \5477 );
and \U$5296 ( \5485 , \2161 , \2913 );
and \U$5297 ( \5486 , \2028 , \2910 );
nor \U$5298 ( \5487 , \5485 , \5486 );
xnor \U$5299 ( \5488 , \5487 , \2371 );
and \U$5300 ( \5489 , \2532 , \2550 );
and \U$5301 ( \5490 , \2305 , \2548 );
nor \U$5302 ( \5491 , \5489 , \5490 );
xnor \U$5303 ( \5492 , \5491 , \2374 );
and \U$5304 ( \5493 , \5488 , \5492 );
and \U$5305 ( \5494 , \5492 , \1835 );
and \U$5306 ( \5495 , \5488 , \1835 );
or \U$5307 ( \5496 , \5493 , \5494 , \5495 );
and \U$5308 ( \5497 , \2763 , \2261 );
and \U$5309 ( \5498 , \2541 , \2259 );
nor \U$5310 ( \5499 , \5497 , \5498 );
xnor \U$5311 ( \5500 , \5499 , \2124 );
nand \U$5312 ( \5501 , \2850 , \1953 );
xnor \U$5313 ( \5502 , \5501 , \1835 );
and \U$5314 ( \5503 , \5500 , \5502 );
and \U$5315 ( \5504 , \5496 , \5503 );
and \U$5316 ( \5505 , \2850 , \1955 );
and \U$5317 ( \5506 , \2763 , \1953 );
nor \U$5318 ( \5507 , \5505 , \5506 );
xnor \U$5319 ( \5508 , \5507 , \1835 );
and \U$5320 ( \5509 , \5503 , \5508 );
and \U$5321 ( \5510 , \5496 , \5508 );
or \U$5322 ( \5511 , \5504 , \5509 , \5510 );
xor \U$5323 ( \5512 , \5465 , \5467 );
xor \U$5324 ( \5513 , \5512 , \5470 );
and \U$5325 ( \5514 , \5511 , \5513 );
and \U$5326 ( \5515 , \5484 , \5514 );
xor \U$5327 ( \5516 , \5484 , \5514 );
xor \U$5328 ( \5517 , \5511 , \5513 );
xor \U$5329 ( \5518 , \5453 , \5457 );
xor \U$5330 ( \5519 , \5518 , \5462 );
xor \U$5331 ( \5520 , \5496 , \5503 );
xor \U$5332 ( \5521 , \5520 , \5508 );
and \U$5333 ( \5522 , \5519 , \5521 );
and \U$5334 ( \5523 , \5517 , \5522 );
xor \U$5335 ( \5524 , \5517 , \5522 );
xor \U$5336 ( \5525 , \5519 , \5521 );
and \U$5337 ( \5526 , \2305 , \2913 );
and \U$5338 ( \5527 , \2161 , \2910 );
nor \U$5339 ( \5528 , \5526 , \5527 );
xnor \U$5340 ( \5529 , \5528 , \2371 );
and \U$5341 ( \5530 , \2541 , \2550 );
and \U$5342 ( \5531 , \2532 , \2548 );
nor \U$5343 ( \5532 , \5530 , \5531 );
xnor \U$5344 ( \5533 , \5532 , \2374 );
and \U$5345 ( \5534 , \5529 , \5533 );
and \U$5346 ( \5535 , \2850 , \2261 );
and \U$5347 ( \5536 , \2763 , \2259 );
nor \U$5348 ( \5537 , \5535 , \5536 );
xnor \U$5349 ( \5538 , \5537 , \2124 );
and \U$5350 ( \5539 , \5533 , \5538 );
and \U$5351 ( \5540 , \5529 , \5538 );
or \U$5352 ( \5541 , \5534 , \5539 , \5540 );
xor \U$5353 ( \5542 , \5488 , \5492 );
xor \U$5354 ( \5543 , \5542 , \1835 );
and \U$5355 ( \5544 , \5541 , \5543 );
xor \U$5356 ( \5545 , \5500 , \5502 );
and \U$5357 ( \5546 , \5543 , \5545 );
and \U$5358 ( \5547 , \5541 , \5545 );
or \U$5359 ( \5548 , \5544 , \5546 , \5547 );
and \U$5360 ( \5549 , \5525 , \5548 );
xor \U$5361 ( \5550 , \5525 , \5548 );
xor \U$5362 ( \5551 , \5541 , \5543 );
xor \U$5363 ( \5552 , \5551 , \5545 );
and \U$5364 ( \5553 , \2532 , \2913 );
and \U$5365 ( \5554 , \2305 , \2910 );
nor \U$5366 ( \5555 , \5553 , \5554 );
xnor \U$5367 ( \5556 , \5555 , \2371 );
and \U$5368 ( \5557 , \2763 , \2550 );
and \U$5369 ( \5558 , \2541 , \2548 );
nor \U$5370 ( \5559 , \5557 , \5558 );
xnor \U$5371 ( \5560 , \5559 , \2374 );
and \U$5372 ( \5561 , \5556 , \5560 );
and \U$5373 ( \5562 , \5560 , \2124 );
and \U$5374 ( \5563 , \5556 , \2124 );
or \U$5375 ( \5564 , \5561 , \5562 , \5563 );
xor \U$5376 ( \5565 , \5529 , \5533 );
xor \U$5377 ( \5566 , \5565 , \5538 );
and \U$5378 ( \5567 , \5564 , \5566 );
and \U$5379 ( \5568 , \5552 , \5567 );
xor \U$5380 ( \5569 , \5552 , \5567 );
xor \U$5381 ( \5570 , \5564 , \5566 );
nand \U$5382 ( \5571 , \2850 , \2259 );
xnor \U$5383 ( \5572 , \5571 , \2124 );
xor \U$5384 ( \5573 , \5556 , \5560 );
xor \U$5385 ( \5574 , \5573 , \2124 );
and \U$5386 ( \5575 , \5572 , \5574 );
and \U$5387 ( \5576 , \5570 , \5575 );
xor \U$5388 ( \5577 , \5570 , \5575 );
xor \U$5389 ( \5578 , \5572 , \5574 );
and \U$5390 ( \5579 , \2541 , \2913 );
and \U$5391 ( \5580 , \2532 , \2910 );
nor \U$5392 ( \5581 , \5579 , \5580 );
xnor \U$5393 ( \5582 , \5581 , \2371 );
and \U$5394 ( \5583 , \2850 , \2550 );
and \U$5395 ( \5584 , \2763 , \2548 );
nor \U$5396 ( \5585 , \5583 , \5584 );
xnor \U$5397 ( \5586 , \5585 , \2374 );
and \U$5398 ( \5587 , \5582 , \5586 );
and \U$5399 ( \5588 , \5578 , \5587 );
xor \U$5400 ( \5589 , \5578 , \5587 );
xor \U$5401 ( \5590 , \5582 , \5586 );
and \U$5402 ( \5591 , \2763 , \2913 );
and \U$5403 ( \5592 , \2541 , \2910 );
nor \U$5404 ( \5593 , \5591 , \5592 );
xnor \U$5405 ( \5594 , \5593 , \2371 );
and \U$5406 ( \5595 , \5594 , \2374 );
and \U$5407 ( \5596 , \5590 , \5595 );
xor \U$5408 ( \5597 , \5590 , \5595 );
nand \U$5409 ( \5598 , \2850 , \2548 );
xnor \U$5410 ( \5599 , \5598 , \2374 );
xor \U$5411 ( \5600 , \5594 , \2374 );
and \U$5412 ( \5601 , \5599 , \5600 );
xor \U$5413 ( \5602 , \5599 , \5600 );
and \U$5414 ( \5603 , \2850 , \2913 );
and \U$5415 ( \5604 , \2763 , \2910 );
nor \U$5416 ( \5605 , \5603 , \5604 );
xnor \U$5417 ( \5606 , \5605 , \2371 );
nand \U$5418 ( \5607 , \2850 , \2910 );
xnor \U$5419 ( \5608 , \5607 , \2371 );
and \U$5420 ( \5609 , \5608 , \2371 );
and \U$5421 ( \5610 , \5606 , \5609 );
and \U$5422 ( \5611 , \5602 , \5610 );
or \U$5423 ( \5612 , \5601 , \5611 );
and \U$5424 ( \5613 , \5597 , \5612 );
or \U$5425 ( \5614 , \5596 , \5613 );
and \U$5426 ( \5615 , \5589 , \5614 );
or \U$5427 ( \5616 , \5588 , \5615 );
and \U$5428 ( \5617 , \5577 , \5616 );
or \U$5429 ( \5618 , \5576 , \5617 );
and \U$5430 ( \5619 , \5569 , \5618 );
or \U$5431 ( \5620 , \5568 , \5619 );
and \U$5432 ( \5621 , \5550 , \5620 );
or \U$5433 ( \5622 , \5549 , \5621 );
and \U$5434 ( \5623 , \5524 , \5622 );
or \U$5435 ( \5624 , \5523 , \5623 );
and \U$5436 ( \5625 , \5516 , \5624 );
or \U$5437 ( \5626 , \5515 , \5625 );
and \U$5438 ( \5627 , \5482 , \5626 );
or \U$5439 ( \5628 , \5481 , \5627 );
and \U$5440 ( \5629 , \5448 , \5628 );
or \U$5441 ( \5630 , \5447 , \5629 );
and \U$5442 ( \5631 , \5440 , \5630 );
or \U$5443 ( \5632 , \5439 , \5631 );
and \U$5444 ( \5633 , \5387 , \5632 );
or \U$5445 ( \5634 , \5386 , \5633 );
and \U$5446 ( \5635 , \5348 , \5634 );
or \U$5447 ( \5636 , \5347 , \5635 );
and \U$5448 ( \5637 , \5295 , \5636 );
or \U$5449 ( \5638 , \5294 , \5637 );
and \U$5450 ( \5639 , \5224 , \5638 );
or \U$5451 ( \5640 , \5223 , \5639 );
and \U$5452 ( \5641 , \5169 , \5640 );
or \U$5453 ( \5642 , \5168 , \5641 );
and \U$5454 ( \5643 , \5110 , \5642 );
or \U$5455 ( \5644 , \5109 , \5643 );
and \U$5456 ( \5645 , \5102 , \5644 );
or \U$5457 ( \5646 , \5101 , \5645 );
and \U$5458 ( \5647 , \5023 , \5646 );
or \U$5459 ( \5648 , \5022 , \5647 );
and \U$5460 ( \5649 , \4943 , \5648 );
or \U$5461 ( \5650 , \4942 , \5649 );
and \U$5462 ( \5651 , \4848 , \5650 );
or \U$5463 ( \5652 , \4847 , \5651 );
and \U$5464 ( \5653 , \4760 , \5652 );
or \U$5465 ( \5654 , \4759 , \5653 );
and \U$5466 ( \5655 , \4668 , \5654 );
or \U$5467 ( \5656 , \4667 , \5655 );
and \U$5468 ( \5657 , \4580 , \5656 );
or \U$5469 ( \5658 , \4579 , \5657 );
and \U$5470 ( \5659 , \4465 , \5658 );
or \U$5471 ( \5660 , \4464 , \5659 );
and \U$5472 ( \5661 , \4369 , \5660 );
or \U$5473 ( \5662 , \4368 , \5661 );
and \U$5474 ( \5663 , \4361 , \5662 );
or \U$5475 ( \5664 , \4360 , \5663 );
and \U$5476 ( \5665 , \4246 , \5664 );
or \U$5477 ( \5666 , \4245 , \5665 );
and \U$5478 ( \5667 , \4122 , \5666 );
or \U$5479 ( \5668 , \4121 , \5667 );
and \U$5480 ( \5669 , \3982 , \5668 );
or \U$5481 ( \5670 , \3981 , \5669 );
and \U$5482 ( \5671 , \3858 , \5670 );
or \U$5483 ( \5672 , \3857 , \5671 );
and \U$5484 ( \5673 , \3714 , \5672 );
or \U$5485 ( \5674 , \3713 , \5673 );
and \U$5486 ( \5675 , \3589 , \5674 );
or \U$5487 ( \5676 , \3588 , \5675 );
and \U$5488 ( \5677 , \3450 , \5676 );
or \U$5489 ( \5678 , \3449 , \5677 );
and \U$5490 ( \5679 , \3285 , \5678 );
or \U$5491 ( \5680 , \3284 , \5679 );
and \U$5492 ( \5681 , \3137 , \5680 );
or \U$5493 ( \5682 , \3136 , \5681 );
and \U$5494 ( \5683 , \2990 , \5682 );
or \U$5495 ( \5684 , \2989 , \5683 );
and \U$5496 ( \5685 , \2822 , \5684 );
or \U$5497 ( \5686 , \2821 , \5685 );
and \U$5498 ( \5687 , \2674 , \5686 );
or \U$5499 ( \5688 , \2673 , \5687 );
and \U$5500 ( \5689 , \2504 , \5688 );
or \U$5501 ( \5690 , \2503 , \5689 );
and \U$5502 ( \5691 , \2366 , \5690 );
or \U$5503 ( \5692 , \2365 , \5691 );
and \U$5504 ( \5693 , \2222 , \5692 );
or \U$5505 ( \5694 , \2221 , \5693 );
and \U$5506 ( \5695 , \2083 , \5694 );
or \U$5507 ( \5696 , \2082 , \5695 );
and \U$5508 ( \5697 , \1950 , \5696 );
or \U$5509 ( \5698 , \1949 , \5697 );
and \U$5510 ( \5699 , \1827 , \5698 );
or \U$5511 ( \5700 , \1826 , \5699 );
and \U$5512 ( \5701 , \1704 , \5700 );
or \U$5513 ( \5702 , \1703 , \5701 );
and \U$5514 ( \5703 , \1586 , \5702 );
or \U$5515 ( \5704 , \1585 , \5703 );
and \U$5516 ( \5705 , \1471 , \5704 );
or \U$5517 ( \5706 , \1470 , \5705 );
and \U$5518 ( \5707 , \1355 , \5706 );
or \U$5519 ( \5708 , \1354 , \5707 );
and \U$5520 ( \5709 , \1241 , \5708 );
or \U$5521 ( \5710 , \1240 , \5709 );
and \U$5522 ( \5711 , \1057 , \5710 );
or \U$5523 ( \5712 , \1056 , \5711 );
and \U$5524 ( \5713 , \976 , \5712 );
or \U$5525 ( \5714 , \975 , \5713 );
and \U$5526 ( \5715 , \893 , \5714 );
or \U$5527 ( \5716 , \892 , \5715 );
and \U$5528 ( \5717 , \810 , \5716 );
or \U$5529 ( \5718 , \809 , \5717 );
and \U$5530 ( \5719 , \735 , \5718 );
or \U$5531 ( \5720 , \734 , \5719 );
and \U$5532 ( \5721 , \659 , \5720 );
or \U$5533 ( \5722 , \658 , \5721 );
and \U$5534 ( \5723 , \537 , \5722 );
or \U$5535 ( \5724 , \536 , \5723 );
xor \U$5536 ( \5725 , \484 , \5724 );
buf \U$5537 ( \5726 , \5725 );
buf \U$5538 ( \5727 , \5726 );
xor \U$5539 ( \5728 , \537 , \5722 );
buf \U$5540 ( \5729 , \5728 );
buf \U$5541 ( \5730 , \5729 );
xor \U$5542 ( \5731 , \659 , \5720 );
buf \U$5543 ( \5732 , \5731 );
buf \U$5544 ( \5733 , \5732 );
and \U$5545 ( \5734 , \5730 , \5733 );
not \U$5546 ( \5735 , \5734 );
and \U$5547 ( \5736 , \5727 , \5735 );
buf \U$5548 ( \5737 , RIa167a08_1);
xor \U$5549 ( \5738 , \4369 , \5660 );
buf \U$5550 ( \5739 , \5738 );
buf \U$5551 ( \5740 , \5739 );
xor \U$5552 ( \5741 , \4465 , \5658 );
buf \U$5553 ( \5742 , \5741 );
buf \U$5554 ( \5743 , \5742 );
xor \U$5555 ( \5744 , \5740 , \5743 );
xor \U$5556 ( \5745 , \4580 , \5656 );
buf \U$5557 ( \5746 , \5745 );
buf \U$5558 ( \5747 , \5746 );
xor \U$5559 ( \5748 , \5743 , \5747 );
not \U$5560 ( \5749 , \5748 );
and \U$5561 ( \5750 , \5744 , \5749 );
and \U$5562 ( \5751 , \5737 , \5750 );
not \U$5563 ( \5752 , \5751 );
and \U$5564 ( \5753 , \5743 , \5747 );
not \U$5565 ( \5754 , \5753 );
and \U$5566 ( \5755 , \5740 , \5754 );
xnor \U$5567 ( \5756 , \5752 , \5755 );
and \U$5568 ( \5757 , \5736 , \5756 );
buf \U$5569 ( \5758 , RIa167918_3);
xor \U$5570 ( \5759 , \4246 , \5664 );
buf \U$5571 ( \5760 , \5759 );
buf \U$5572 ( \5761 , \5760 );
xor \U$5573 ( \5762 , \4361 , \5662 );
buf \U$5574 ( \5763 , \5762 );
buf \U$5575 ( \5764 , \5763 );
xor \U$5576 ( \5765 , \5761 , \5764 );
xor \U$5577 ( \5766 , \5764 , \5740 );
not \U$5578 ( \5767 , \5766 );
and \U$5579 ( \5768 , \5765 , \5767 );
and \U$5580 ( \5769 , \5758 , \5768 );
buf \U$5581 ( \5770 , RIa167990_2);
and \U$5582 ( \5771 , \5770 , \5766 );
nor \U$5583 ( \5772 , \5769 , \5771 );
and \U$5584 ( \5773 , \5764 , \5740 );
not \U$5585 ( \5774 , \5773 );
and \U$5586 ( \5775 , \5761 , \5774 );
xnor \U$5587 ( \5776 , \5772 , \5775 );
and \U$5588 ( \5777 , \5756 , \5776 );
and \U$5589 ( \5778 , \5736 , \5776 );
or \U$5590 ( \5779 , \5757 , \5777 , \5778 );
buf \U$5591 ( \5780 , RIa167828_5);
xor \U$5592 ( \5781 , \3982 , \5668 );
buf \U$5593 ( \5782 , \5781 );
buf \U$5594 ( \5783 , \5782 );
xor \U$5595 ( \5784 , \4122 , \5666 );
buf \U$5596 ( \5785 , \5784 );
buf \U$5597 ( \5786 , \5785 );
xor \U$5598 ( \5787 , \5783 , \5786 );
xor \U$5599 ( \5788 , \5786 , \5761 );
not \U$5600 ( \5789 , \5788 );
and \U$5601 ( \5790 , \5787 , \5789 );
and \U$5602 ( \5791 , \5780 , \5790 );
buf \U$5603 ( \5792 , RIa1678a0_4);
and \U$5604 ( \5793 , \5792 , \5788 );
nor \U$5605 ( \5794 , \5791 , \5793 );
and \U$5606 ( \5795 , \5786 , \5761 );
not \U$5607 ( \5796 , \5795 );
and \U$5608 ( \5797 , \5783 , \5796 );
xnor \U$5609 ( \5798 , \5794 , \5797 );
buf \U$5610 ( \5799 , RIa167738_7);
xor \U$5611 ( \5800 , \3714 , \5672 );
buf \U$5612 ( \5801 , \5800 );
buf \U$5613 ( \5802 , \5801 );
xor \U$5614 ( \5803 , \3858 , \5670 );
buf \U$5615 ( \5804 , \5803 );
buf \U$5616 ( \5805 , \5804 );
xor \U$5617 ( \5806 , \5802 , \5805 );
xor \U$5618 ( \5807 , \5805 , \5783 );
not \U$5619 ( \5808 , \5807 );
and \U$5620 ( \5809 , \5806 , \5808 );
and \U$5621 ( \5810 , \5799 , \5809 );
buf \U$5622 ( \5811 , RIa1677b0_6);
and \U$5623 ( \5812 , \5811 , \5807 );
nor \U$5624 ( \5813 , \5810 , \5812 );
and \U$5625 ( \5814 , \5805 , \5783 );
not \U$5626 ( \5815 , \5814 );
and \U$5627 ( \5816 , \5802 , \5815 );
xnor \U$5628 ( \5817 , \5813 , \5816 );
and \U$5629 ( \5818 , \5798 , \5817 );
buf \U$5630 ( \5819 , RIa167648_9);
xor \U$5631 ( \5820 , \3450 , \5676 );
buf \U$5632 ( \5821 , \5820 );
buf \U$5633 ( \5822 , \5821 );
xor \U$5634 ( \5823 , \3589 , \5674 );
buf \U$5635 ( \5824 , \5823 );
buf \U$5636 ( \5825 , \5824 );
xor \U$5637 ( \5826 , \5822 , \5825 );
xor \U$5638 ( \5827 , \5825 , \5802 );
not \U$5639 ( \5828 , \5827 );
and \U$5640 ( \5829 , \5826 , \5828 );
and \U$5641 ( \5830 , \5819 , \5829 );
buf \U$5642 ( \5831 , RIa1676c0_8);
and \U$5643 ( \5832 , \5831 , \5827 );
nor \U$5644 ( \5833 , \5830 , \5832 );
and \U$5645 ( \5834 , \5825 , \5802 );
not \U$5646 ( \5835 , \5834 );
and \U$5647 ( \5836 , \5822 , \5835 );
xnor \U$5648 ( \5837 , \5833 , \5836 );
and \U$5649 ( \5838 , \5817 , \5837 );
and \U$5650 ( \5839 , \5798 , \5837 );
or \U$5651 ( \5840 , \5818 , \5838 , \5839 );
and \U$5652 ( \5841 , \5779 , \5840 );
buf \U$5653 ( \5842 , RIa167558_11);
xor \U$5654 ( \5843 , \3137 , \5680 );
buf \U$5655 ( \5844 , \5843 );
buf \U$5656 ( \5845 , \5844 );
xor \U$5657 ( \5846 , \3285 , \5678 );
buf \U$5658 ( \5847 , \5846 );
buf \U$5659 ( \5848 , \5847 );
xor \U$5660 ( \5849 , \5845 , \5848 );
xor \U$5661 ( \5850 , \5848 , \5822 );
not \U$5662 ( \5851 , \5850 );
and \U$5663 ( \5852 , \5849 , \5851 );
and \U$5664 ( \5853 , \5842 , \5852 );
buf \U$5665 ( \5854 , RIa1675d0_10);
and \U$5666 ( \5855 , \5854 , \5850 );
nor \U$5667 ( \5856 , \5853 , \5855 );
and \U$5668 ( \5857 , \5848 , \5822 );
not \U$5669 ( \5858 , \5857 );
and \U$5670 ( \5859 , \5845 , \5858 );
xnor \U$5671 ( \5860 , \5856 , \5859 );
buf \U$5672 ( \5861 , RIa167468_13);
xor \U$5673 ( \5862 , \2822 , \5684 );
buf \U$5674 ( \5863 , \5862 );
buf \U$5675 ( \5864 , \5863 );
xor \U$5676 ( \5865 , \2990 , \5682 );
buf \U$5677 ( \5866 , \5865 );
buf \U$5678 ( \5867 , \5866 );
xor \U$5679 ( \5868 , \5864 , \5867 );
xor \U$5680 ( \5869 , \5867 , \5845 );
not \U$5681 ( \5870 , \5869 );
and \U$5682 ( \5871 , \5868 , \5870 );
and \U$5683 ( \5872 , \5861 , \5871 );
buf \U$5684 ( \5873 , RIa1674e0_12);
and \U$5685 ( \5874 , \5873 , \5869 );
nor \U$5686 ( \5875 , \5872 , \5874 );
and \U$5687 ( \5876 , \5867 , \5845 );
not \U$5688 ( \5877 , \5876 );
and \U$5689 ( \5878 , \5864 , \5877 );
xnor \U$5690 ( \5879 , \5875 , \5878 );
and \U$5691 ( \5880 , \5860 , \5879 );
buf \U$5692 ( \5881 , RIa167378_15);
xor \U$5693 ( \5882 , \2504 , \5688 );
buf \U$5694 ( \5883 , \5882 );
buf \U$5695 ( \5884 , \5883 );
xor \U$5696 ( \5885 , \2674 , \5686 );
buf \U$5697 ( \5886 , \5885 );
buf \U$5698 ( \5887 , \5886 );
xor \U$5699 ( \5888 , \5884 , \5887 );
xor \U$5700 ( \5889 , \5887 , \5864 );
not \U$5701 ( \5890 , \5889 );
and \U$5702 ( \5891 , \5888 , \5890 );
and \U$5703 ( \5892 , \5881 , \5891 );
buf \U$5704 ( \5893 , RIa1673f0_14);
and \U$5705 ( \5894 , \5893 , \5889 );
nor \U$5706 ( \5895 , \5892 , \5894 );
and \U$5707 ( \5896 , \5887 , \5864 );
not \U$5708 ( \5897 , \5896 );
and \U$5709 ( \5898 , \5884 , \5897 );
xnor \U$5710 ( \5899 , \5895 , \5898 );
and \U$5711 ( \5900 , \5879 , \5899 );
and \U$5712 ( \5901 , \5860 , \5899 );
or \U$5713 ( \5902 , \5880 , \5900 , \5901 );
and \U$5714 ( \5903 , \5840 , \5902 );
and \U$5715 ( \5904 , \5779 , \5902 );
or \U$5716 ( \5905 , \5841 , \5903 , \5904 );
buf \U$5717 ( \5906 , RIa167288_17);
xor \U$5718 ( \5907 , \2222 , \5692 );
buf \U$5719 ( \5908 , \5907 );
buf \U$5720 ( \5909 , \5908 );
xor \U$5721 ( \5910 , \2366 , \5690 );
buf \U$5722 ( \5911 , \5910 );
buf \U$5723 ( \5912 , \5911 );
xor \U$5724 ( \5913 , \5909 , \5912 );
xor \U$5725 ( \5914 , \5912 , \5884 );
not \U$5726 ( \5915 , \5914 );
and \U$5727 ( \5916 , \5913 , \5915 );
and \U$5728 ( \5917 , \5906 , \5916 );
buf \U$5729 ( \5918 , RIa167300_16);
and \U$5730 ( \5919 , \5918 , \5914 );
nor \U$5731 ( \5920 , \5917 , \5919 );
and \U$5732 ( \5921 , \5912 , \5884 );
not \U$5733 ( \5922 , \5921 );
and \U$5734 ( \5923 , \5909 , \5922 );
xnor \U$5735 ( \5924 , \5920 , \5923 );
buf \U$5736 ( \5925 , RIa167198_19);
xor \U$5737 ( \5926 , \1950 , \5696 );
buf \U$5738 ( \5927 , \5926 );
buf \U$5739 ( \5928 , \5927 );
xor \U$5740 ( \5929 , \2083 , \5694 );
buf \U$5741 ( \5930 , \5929 );
buf \U$5742 ( \5931 , \5930 );
xor \U$5743 ( \5932 , \5928 , \5931 );
xor \U$5744 ( \5933 , \5931 , \5909 );
not \U$5745 ( \5934 , \5933 );
and \U$5746 ( \5935 , \5932 , \5934 );
and \U$5747 ( \5936 , \5925 , \5935 );
buf \U$5748 ( \5937 , RIa167210_18);
and \U$5749 ( \5938 , \5937 , \5933 );
nor \U$5750 ( \5939 , \5936 , \5938 );
and \U$5751 ( \5940 , \5931 , \5909 );
not \U$5752 ( \5941 , \5940 );
and \U$5753 ( \5942 , \5928 , \5941 );
xnor \U$5754 ( \5943 , \5939 , \5942 );
and \U$5755 ( \5944 , \5924 , \5943 );
buf \U$5756 ( \5945 , RIa1670a8_21);
xor \U$5757 ( \5946 , \1704 , \5700 );
buf \U$5758 ( \5947 , \5946 );
buf \U$5759 ( \5948 , \5947 );
xor \U$5760 ( \5949 , \1827 , \5698 );
buf \U$5761 ( \5950 , \5949 );
buf \U$5762 ( \5951 , \5950 );
xor \U$5763 ( \5952 , \5948 , \5951 );
xor \U$5764 ( \5953 , \5951 , \5928 );
not \U$5765 ( \5954 , \5953 );
and \U$5766 ( \5955 , \5952 , \5954 );
and \U$5767 ( \5956 , \5945 , \5955 );
buf \U$5768 ( \5957 , RIa167120_20);
and \U$5769 ( \5958 , \5957 , \5953 );
nor \U$5770 ( \5959 , \5956 , \5958 );
and \U$5771 ( \5960 , \5951 , \5928 );
not \U$5772 ( \5961 , \5960 );
and \U$5773 ( \5962 , \5948 , \5961 );
xnor \U$5774 ( \5963 , \5959 , \5962 );
and \U$5775 ( \5964 , \5943 , \5963 );
and \U$5776 ( \5965 , \5924 , \5963 );
or \U$5777 ( \5966 , \5944 , \5964 , \5965 );
buf \U$5778 ( \5967 , RIa166fb8_23);
xor \U$5779 ( \5968 , \1471 , \5704 );
buf \U$5780 ( \5969 , \5968 );
buf \U$5781 ( \5970 , \5969 );
xor \U$5782 ( \5971 , \1586 , \5702 );
buf \U$5783 ( \5972 , \5971 );
buf \U$5784 ( \5973 , \5972 );
xor \U$5785 ( \5974 , \5970 , \5973 );
xor \U$5786 ( \5975 , \5973 , \5948 );
not \U$5787 ( \5976 , \5975 );
and \U$5788 ( \5977 , \5974 , \5976 );
and \U$5789 ( \5978 , \5967 , \5977 );
buf \U$5790 ( \5979 , RIa167030_22);
and \U$5791 ( \5980 , \5979 , \5975 );
nor \U$5792 ( \5981 , \5978 , \5980 );
and \U$5793 ( \5982 , \5973 , \5948 );
not \U$5794 ( \5983 , \5982 );
and \U$5795 ( \5984 , \5970 , \5983 );
xnor \U$5796 ( \5985 , \5981 , \5984 );
buf \U$5797 ( \5986 , RIa166ec8_25);
xor \U$5798 ( \5987 , \1241 , \5708 );
buf \U$5799 ( \5988 , \5987 );
buf \U$5800 ( \5989 , \5988 );
xor \U$5801 ( \5990 , \1355 , \5706 );
buf \U$5802 ( \5991 , \5990 );
buf \U$5803 ( \5992 , \5991 );
xor \U$5804 ( \5993 , \5989 , \5992 );
xor \U$5805 ( \5994 , \5992 , \5970 );
not \U$5806 ( \5995 , \5994 );
and \U$5807 ( \5996 , \5993 , \5995 );
and \U$5808 ( \5997 , \5986 , \5996 );
buf \U$5809 ( \5998 , RIa166f40_24);
and \U$5810 ( \5999 , \5998 , \5994 );
nor \U$5811 ( \6000 , \5997 , \5999 );
and \U$5812 ( \6001 , \5992 , \5970 );
not \U$5813 ( \6002 , \6001 );
and \U$5814 ( \6003 , \5989 , \6002 );
xnor \U$5815 ( \6004 , \6000 , \6003 );
and \U$5816 ( \6005 , \5985 , \6004 );
buf \U$5817 ( \6006 , RIa166dd8_27);
xor \U$5818 ( \6007 , \976 , \5712 );
buf \U$5819 ( \6008 , \6007 );
buf \U$5820 ( \6009 , \6008 );
xor \U$5821 ( \6010 , \1057 , \5710 );
buf \U$5822 ( \6011 , \6010 );
buf \U$5823 ( \6012 , \6011 );
xor \U$5824 ( \6013 , \6009 , \6012 );
xor \U$5825 ( \6014 , \6012 , \5989 );
not \U$5826 ( \6015 , \6014 );
and \U$5827 ( \6016 , \6013 , \6015 );
and \U$5828 ( \6017 , \6006 , \6016 );
buf \U$5829 ( \6018 , RIa166e50_26);
and \U$5830 ( \6019 , \6018 , \6014 );
nor \U$5831 ( \6020 , \6017 , \6019 );
and \U$5832 ( \6021 , \6012 , \5989 );
not \U$5833 ( \6022 , \6021 );
and \U$5834 ( \6023 , \6009 , \6022 );
xnor \U$5835 ( \6024 , \6020 , \6023 );
and \U$5836 ( \6025 , \6004 , \6024 );
and \U$5837 ( \6026 , \5985 , \6024 );
or \U$5838 ( \6027 , \6005 , \6025 , \6026 );
and \U$5839 ( \6028 , \5966 , \6027 );
buf \U$5840 ( \6029 , RIa166ce8_29);
xor \U$5841 ( \6030 , \810 , \5716 );
buf \U$5842 ( \6031 , \6030 );
buf \U$5843 ( \6032 , \6031 );
xor \U$5844 ( \6033 , \893 , \5714 );
buf \U$5845 ( \6034 , \6033 );
buf \U$5846 ( \6035 , \6034 );
xor \U$5847 ( \6036 , \6032 , \6035 );
xor \U$5848 ( \6037 , \6035 , \6009 );
not \U$5849 ( \6038 , \6037 );
and \U$5850 ( \6039 , \6036 , \6038 );
and \U$5851 ( \6040 , \6029 , \6039 );
buf \U$5852 ( \6041 , RIa166d60_28);
and \U$5853 ( \6042 , \6041 , \6037 );
nor \U$5854 ( \6043 , \6040 , \6042 );
and \U$5855 ( \6044 , \6035 , \6009 );
not \U$5856 ( \6045 , \6044 );
and \U$5857 ( \6046 , \6032 , \6045 );
xnor \U$5858 ( \6047 , \6043 , \6046 );
buf \U$5859 ( \6048 , RIb4ca4d8_31);
xor \U$5860 ( \6049 , \735 , \5718 );
buf \U$5861 ( \6050 , \6049 );
buf \U$5862 ( \6051 , \6050 );
xor \U$5863 ( \6052 , \5733 , \6051 );
xor \U$5864 ( \6053 , \6051 , \6032 );
not \U$5865 ( \6054 , \6053 );
and \U$5866 ( \6055 , \6052 , \6054 );
and \U$5867 ( \6056 , \6048 , \6055 );
buf \U$5868 ( \6057 , RIa166c70_30);
and \U$5869 ( \6058 , \6057 , \6053 );
nor \U$5870 ( \6059 , \6056 , \6058 );
and \U$5871 ( \6060 , \6051 , \6032 );
not \U$5872 ( \6061 , \6060 );
and \U$5873 ( \6062 , \5733 , \6061 );
xnor \U$5874 ( \6063 , \6059 , \6062 );
and \U$5875 ( \6064 , \6047 , \6063 );
buf \U$5876 ( \6065 , RIb4ca460_32);
xor \U$5877 ( \6066 , \5730 , \5733 );
nand \U$5878 ( \6067 , \6065 , \6066 );
xnor \U$5879 ( \6068 , \6067 , \5736 );
and \U$5880 ( \6069 , \6063 , \6068 );
and \U$5881 ( \6070 , \6047 , \6068 );
or \U$5882 ( \6071 , \6064 , \6069 , \6070 );
and \U$5883 ( \6072 , \6027 , \6071 );
and \U$5884 ( \6073 , \5966 , \6071 );
or \U$5885 ( \6074 , \6028 , \6072 , \6073 );
and \U$5886 ( \6075 , \5905 , \6074 );
and \U$5887 ( \6076 , \6057 , \6055 );
and \U$5888 ( \6077 , \6029 , \6053 );
nor \U$5889 ( \6078 , \6076 , \6077 );
xnor \U$5890 ( \6079 , \6078 , \6062 );
xor \U$5891 ( \6080 , \5727 , \5730 );
not \U$5892 ( \6081 , \6066 );
and \U$5893 ( \6082 , \6080 , \6081 );
and \U$5894 ( \6083 , \6065 , \6082 );
and \U$5895 ( \6084 , \6048 , \6066 );
nor \U$5896 ( \6085 , \6083 , \6084 );
xnor \U$5897 ( \6086 , \6085 , \5736 );
xor \U$5898 ( \6087 , \6079 , \6086 );
and \U$5899 ( \6088 , \5998 , \5996 );
and \U$5900 ( \6089 , \5967 , \5994 );
nor \U$5901 ( \6090 , \6088 , \6089 );
xnor \U$5902 ( \6091 , \6090 , \6003 );
and \U$5903 ( \6092 , \6018 , \6016 );
and \U$5904 ( \6093 , \5986 , \6014 );
nor \U$5905 ( \6094 , \6092 , \6093 );
xnor \U$5906 ( \6095 , \6094 , \6023 );
xor \U$5907 ( \6096 , \6091 , \6095 );
and \U$5908 ( \6097 , \6041 , \6039 );
and \U$5909 ( \6098 , \6006 , \6037 );
nor \U$5910 ( \6099 , \6097 , \6098 );
xnor \U$5911 ( \6100 , \6099 , \6046 );
xor \U$5912 ( \6101 , \6096 , \6100 );
and \U$5913 ( \6102 , \6087 , \6101 );
and \U$5914 ( \6103 , \5937 , \5935 );
and \U$5915 ( \6104 , \5906 , \5933 );
nor \U$5916 ( \6105 , \6103 , \6104 );
xnor \U$5917 ( \6106 , \6105 , \5942 );
and \U$5918 ( \6107 , \5957 , \5955 );
and \U$5919 ( \6108 , \5925 , \5953 );
nor \U$5920 ( \6109 , \6107 , \6108 );
xnor \U$5921 ( \6110 , \6109 , \5962 );
xor \U$5922 ( \6111 , \6106 , \6110 );
and \U$5923 ( \6112 , \5979 , \5977 );
and \U$5924 ( \6113 , \5945 , \5975 );
nor \U$5925 ( \6114 , \6112 , \6113 );
xnor \U$5926 ( \6115 , \6114 , \5984 );
xor \U$5927 ( \6116 , \6111 , \6115 );
and \U$5928 ( \6117 , \6101 , \6116 );
and \U$5929 ( \6118 , \6087 , \6116 );
or \U$5930 ( \6119 , \6102 , \6117 , \6118 );
and \U$5931 ( \6120 , \6074 , \6119 );
and \U$5932 ( \6121 , \5905 , \6119 );
or \U$5933 ( \6122 , \6075 , \6120 , \6121 );
and \U$5934 ( \6123 , \5873 , \5871 );
and \U$5935 ( \6124 , \5842 , \5869 );
nor \U$5936 ( \6125 , \6123 , \6124 );
xnor \U$5937 ( \6126 , \6125 , \5878 );
and \U$5938 ( \6127 , \5893 , \5891 );
and \U$5939 ( \6128 , \5861 , \5889 );
nor \U$5940 ( \6129 , \6127 , \6128 );
xnor \U$5941 ( \6130 , \6129 , \5898 );
xor \U$5942 ( \6131 , \6126 , \6130 );
and \U$5943 ( \6132 , \5918 , \5916 );
and \U$5944 ( \6133 , \5881 , \5914 );
nor \U$5945 ( \6134 , \6132 , \6133 );
xnor \U$5946 ( \6135 , \6134 , \5923 );
xor \U$5947 ( \6136 , \6131 , \6135 );
and \U$5948 ( \6137 , \5811 , \5809 );
and \U$5949 ( \6138 , \5780 , \5807 );
nor \U$5950 ( \6139 , \6137 , \6138 );
xnor \U$5951 ( \6140 , \6139 , \5816 );
and \U$5952 ( \6141 , \5831 , \5829 );
and \U$5953 ( \6142 , \5799 , \5827 );
nor \U$5954 ( \6143 , \6141 , \6142 );
xnor \U$5955 ( \6144 , \6143 , \5836 );
xor \U$5956 ( \6145 , \6140 , \6144 );
and \U$5957 ( \6146 , \5854 , \5852 );
and \U$5958 ( \6147 , \5819 , \5850 );
nor \U$5959 ( \6148 , \6146 , \6147 );
xnor \U$5960 ( \6149 , \6148 , \5859 );
xor \U$5961 ( \6150 , \6145 , \6149 );
and \U$5962 ( \6151 , \6136 , \6150 );
not \U$5963 ( \6152 , \5755 );
and \U$5964 ( \6153 , \5770 , \5768 );
and \U$5965 ( \6154 , \5737 , \5766 );
nor \U$5966 ( \6155 , \6153 , \6154 );
xnor \U$5967 ( \6156 , \6155 , \5775 );
xor \U$5968 ( \6157 , \6152 , \6156 );
and \U$5969 ( \6158 , \5792 , \5790 );
and \U$5970 ( \6159 , \5758 , \5788 );
nor \U$5971 ( \6160 , \6158 , \6159 );
xnor \U$5972 ( \6161 , \6160 , \5797 );
xor \U$5973 ( \6162 , \6157 , \6161 );
and \U$5974 ( \6163 , \6150 , \6162 );
and \U$5975 ( \6164 , \6136 , \6162 );
or \U$5976 ( \6165 , \6151 , \6163 , \6164 );
and \U$5977 ( \6166 , \159 , \331 );
not \U$5978 ( \6167 , \6166 );
xnor \U$5979 ( \6168 , \6167 , \338 );
and \U$5980 ( \6169 , \305 , \351 );
and \U$5981 ( \6170 , \315 , \349 );
nor \U$5982 ( \6171 , \6169 , \6170 );
xnor \U$5983 ( \6172 , \6171 , \358 );
and \U$5984 ( \6173 , \6168 , \6172 );
and \U$5985 ( \6174 , \333 , \345 );
and \U$5986 ( \6175 , \6172 , \6174 );
and \U$5987 ( \6176 , \6168 , \6174 );
or \U$5988 ( \6177 , \6173 , \6175 , \6176 );
and \U$5989 ( \6178 , \413 , \417 );
and \U$5990 ( \6179 , \417 , \422 );
and \U$5991 ( \6180 , \413 , \422 );
or \U$5992 ( \6181 , \6178 , \6179 , \6180 );
xor \U$5993 ( \6182 , \6168 , \6172 );
xor \U$5994 ( \6183 , \6182 , \6174 );
or \U$5995 ( \6184 , \6181 , \6183 );
xor \U$5996 ( \6185 , \6177 , \6184 );
not \U$5997 ( \6186 , \338 );
and \U$5998 ( \6187 , \315 , \351 );
and \U$5999 ( \6188 , \159 , \349 );
nor \U$6000 ( \6189 , \6187 , \6188 );
xnor \U$6001 ( \6190 , \6189 , \358 );
xor \U$6002 ( \6191 , \6186 , \6190 );
and \U$6003 ( \6192 , \305 , \345 );
xor \U$6004 ( \6193 , \6191 , \6192 );
xor \U$6005 ( \6194 , \6185 , \6193 );
and \U$6006 ( \6195 , \428 , \429 );
and \U$6007 ( \6196 , \429 , \431 );
and \U$6008 ( \6197 , \428 , \431 );
or \U$6009 ( \6198 , \6195 , \6196 , \6197 );
and \U$6010 ( \6199 , \412 , \423 );
and \U$6011 ( \6200 , \423 , \432 );
and \U$6012 ( \6201 , \412 , \432 );
or \U$6013 ( \6202 , \6199 , \6200 , \6201 );
and \U$6014 ( \6203 , \6198 , \6202 );
xnor \U$6015 ( \6204 , \6181 , \6183 );
and \U$6016 ( \6205 , \6202 , \6204 );
and \U$6017 ( \6206 , \6198 , \6204 );
or \U$6018 ( \6207 , \6203 , \6205 , \6206 );
xor \U$6019 ( \6208 , \6194 , \6207 );
xor \U$6020 ( \6209 , \6198 , \6202 );
xor \U$6021 ( \6210 , \6209 , \6204 );
and \U$6022 ( \6211 , \408 , \433 );
and \U$6023 ( \6212 , \6210 , \6211 );
xor \U$6024 ( \6213 , \6210 , \6211 );
and \U$6025 ( \6214 , \434 , \483 );
and \U$6026 ( \6215 , \484 , \5724 );
or \U$6027 ( \6216 , \6214 , \6215 );
and \U$6028 ( \6217 , \6213 , \6216 );
or \U$6029 ( \6218 , \6212 , \6217 );
xor \U$6030 ( \6219 , \6208 , \6218 );
buf \U$6031 ( \6220 , \6219 );
buf \U$6032 ( \6221 , \6220 );
xor \U$6033 ( \6222 , \6213 , \6216 );
buf \U$6034 ( \6223 , \6222 );
buf \U$6035 ( \6224 , \6223 );
and \U$6036 ( \6225 , \6224 , \5727 );
not \U$6037 ( \6226 , \6225 );
and \U$6038 ( \6227 , \6221 , \6226 );
and \U$6039 ( \6228 , \5737 , \5768 );
not \U$6040 ( \6229 , \6228 );
xnor \U$6041 ( \6230 , \6229 , \5775 );
xor \U$6042 ( \6231 , \6227 , \6230 );
and \U$6043 ( \6232 , \5758 , \5790 );
and \U$6044 ( \6233 , \5770 , \5788 );
nor \U$6045 ( \6234 , \6232 , \6233 );
xnor \U$6046 ( \6235 , \6234 , \5797 );
xor \U$6047 ( \6236 , \6231 , \6235 );
and \U$6048 ( \6237 , \6165 , \6236 );
and \U$6049 ( \6238 , \5906 , \5935 );
and \U$6050 ( \6239 , \5918 , \5933 );
nor \U$6051 ( \6240 , \6238 , \6239 );
xnor \U$6052 ( \6241 , \6240 , \5942 );
and \U$6053 ( \6242 , \5925 , \5955 );
and \U$6054 ( \6243 , \5937 , \5953 );
nor \U$6055 ( \6244 , \6242 , \6243 );
xnor \U$6056 ( \6245 , \6244 , \5962 );
xor \U$6057 ( \6246 , \6241 , \6245 );
and \U$6058 ( \6247 , \5945 , \5977 );
and \U$6059 ( \6248 , \5957 , \5975 );
nor \U$6060 ( \6249 , \6247 , \6248 );
xnor \U$6061 ( \6250 , \6249 , \5984 );
xor \U$6062 ( \6251 , \6246 , \6250 );
and \U$6063 ( \6252 , \5842 , \5871 );
and \U$6064 ( \6253 , \5854 , \5869 );
nor \U$6065 ( \6254 , \6252 , \6253 );
xnor \U$6066 ( \6255 , \6254 , \5878 );
and \U$6067 ( \6256 , \5861 , \5891 );
and \U$6068 ( \6257 , \5873 , \5889 );
nor \U$6069 ( \6258 , \6256 , \6257 );
xnor \U$6070 ( \6259 , \6258 , \5898 );
xor \U$6071 ( \6260 , \6255 , \6259 );
and \U$6072 ( \6261 , \5881 , \5916 );
and \U$6073 ( \6262 , \5893 , \5914 );
nor \U$6074 ( \6263 , \6261 , \6262 );
xnor \U$6075 ( \6264 , \6263 , \5923 );
xor \U$6076 ( \6265 , \6260 , \6264 );
xor \U$6077 ( \6266 , \6251 , \6265 );
and \U$6078 ( \6267 , \5780 , \5809 );
and \U$6079 ( \6268 , \5792 , \5807 );
nor \U$6080 ( \6269 , \6267 , \6268 );
xnor \U$6081 ( \6270 , \6269 , \5816 );
and \U$6082 ( \6271 , \5799 , \5829 );
and \U$6083 ( \6272 , \5811 , \5827 );
nor \U$6084 ( \6273 , \6271 , \6272 );
xnor \U$6085 ( \6274 , \6273 , \5836 );
xor \U$6086 ( \6275 , \6270 , \6274 );
and \U$6087 ( \6276 , \5819 , \5852 );
and \U$6088 ( \6277 , \5831 , \5850 );
nor \U$6089 ( \6278 , \6276 , \6277 );
xnor \U$6090 ( \6279 , \6278 , \5859 );
xor \U$6091 ( \6280 , \6275 , \6279 );
xor \U$6092 ( \6281 , \6266 , \6280 );
and \U$6093 ( \6282 , \6236 , \6281 );
and \U$6094 ( \6283 , \6165 , \6281 );
or \U$6095 ( \6284 , \6237 , \6282 , \6283 );
and \U$6096 ( \6285 , \6122 , \6284 );
and \U$6097 ( \6286 , \6029 , \6055 );
and \U$6098 ( \6287 , \6041 , \6053 );
nor \U$6099 ( \6288 , \6286 , \6287 );
xnor \U$6100 ( \6289 , \6288 , \6062 );
and \U$6101 ( \6290 , \6048 , \6082 );
and \U$6102 ( \6291 , \6057 , \6066 );
nor \U$6103 ( \6292 , \6290 , \6291 );
xnor \U$6104 ( \6293 , \6292 , \5736 );
xor \U$6105 ( \6294 , \6289 , \6293 );
xor \U$6106 ( \6295 , \6224 , \5727 );
nand \U$6107 ( \6296 , \6065 , \6295 );
xnor \U$6108 ( \6297 , \6296 , \6227 );
xor \U$6109 ( \6298 , \6294 , \6297 );
and \U$6110 ( \6299 , \5967 , \5996 );
and \U$6111 ( \6300 , \5979 , \5994 );
nor \U$6112 ( \6301 , \6299 , \6300 );
xnor \U$6113 ( \6302 , \6301 , \6003 );
and \U$6114 ( \6303 , \5986 , \6016 );
and \U$6115 ( \6304 , \5998 , \6014 );
nor \U$6116 ( \6305 , \6303 , \6304 );
xnor \U$6117 ( \6306 , \6305 , \6023 );
xor \U$6118 ( \6307 , \6302 , \6306 );
and \U$6119 ( \6308 , \6006 , \6039 );
and \U$6120 ( \6309 , \6018 , \6037 );
nor \U$6121 ( \6310 , \6308 , \6309 );
xnor \U$6122 ( \6311 , \6310 , \6046 );
xor \U$6123 ( \6312 , \6307 , \6311 );
xnor \U$6124 ( \6313 , \6298 , \6312 );
and \U$6125 ( \6314 , \6106 , \6110 );
and \U$6126 ( \6315 , \6110 , \6115 );
and \U$6127 ( \6316 , \6106 , \6115 );
or \U$6128 ( \6317 , \6314 , \6315 , \6316 );
and \U$6129 ( \6318 , \6091 , \6095 );
and \U$6130 ( \6319 , \6095 , \6100 );
and \U$6131 ( \6320 , \6091 , \6100 );
or \U$6132 ( \6321 , \6318 , \6319 , \6320 );
xor \U$6133 ( \6322 , \6317 , \6321 );
and \U$6134 ( \6323 , \6079 , \6086 );
xor \U$6135 ( \6324 , \6322 , \6323 );
and \U$6136 ( \6325 , \6313 , \6324 );
and \U$6137 ( \6326 , \6152 , \6156 );
and \U$6138 ( \6327 , \6156 , \6161 );
and \U$6139 ( \6328 , \6152 , \6161 );
or \U$6140 ( \6329 , \6326 , \6327 , \6328 );
and \U$6141 ( \6330 , \6140 , \6144 );
and \U$6142 ( \6331 , \6144 , \6149 );
and \U$6143 ( \6332 , \6140 , \6149 );
or \U$6144 ( \6333 , \6330 , \6331 , \6332 );
xor \U$6145 ( \6334 , \6329 , \6333 );
and \U$6146 ( \6335 , \6126 , \6130 );
and \U$6147 ( \6336 , \6130 , \6135 );
and \U$6148 ( \6337 , \6126 , \6135 );
or \U$6149 ( \6338 , \6335 , \6336 , \6337 );
xor \U$6150 ( \6339 , \6334 , \6338 );
and \U$6151 ( \6340 , \6324 , \6339 );
and \U$6152 ( \6341 , \6313 , \6339 );
or \U$6153 ( \6342 , \6325 , \6340 , \6341 );
and \U$6154 ( \6343 , \6284 , \6342 );
and \U$6155 ( \6344 , \6122 , \6342 );
or \U$6156 ( \6345 , \6285 , \6343 , \6344 );
and \U$6157 ( \6346 , \6241 , \6245 );
and \U$6158 ( \6347 , \6245 , \6250 );
and \U$6159 ( \6348 , \6241 , \6250 );
or \U$6160 ( \6349 , \6346 , \6347 , \6348 );
and \U$6161 ( \6350 , \6302 , \6306 );
and \U$6162 ( \6351 , \6306 , \6311 );
and \U$6163 ( \6352 , \6302 , \6311 );
or \U$6164 ( \6353 , \6350 , \6351 , \6352 );
xor \U$6165 ( \6354 , \6349 , \6353 );
and \U$6166 ( \6355 , \6289 , \6293 );
and \U$6167 ( \6356 , \6293 , \6297 );
and \U$6168 ( \6357 , \6289 , \6297 );
or \U$6169 ( \6358 , \6355 , \6356 , \6357 );
xor \U$6170 ( \6359 , \6354 , \6358 );
and \U$6171 ( \6360 , \6227 , \6230 );
and \U$6172 ( \6361 , \6230 , \6235 );
and \U$6173 ( \6362 , \6227 , \6235 );
or \U$6174 ( \6363 , \6360 , \6361 , \6362 );
and \U$6175 ( \6364 , \6270 , \6274 );
and \U$6176 ( \6365 , \6274 , \6279 );
and \U$6177 ( \6366 , \6270 , \6279 );
or \U$6178 ( \6367 , \6364 , \6365 , \6366 );
xor \U$6179 ( \6368 , \6363 , \6367 );
and \U$6180 ( \6369 , \6255 , \6259 );
and \U$6181 ( \6370 , \6259 , \6264 );
and \U$6182 ( \6371 , \6255 , \6264 );
or \U$6183 ( \6372 , \6369 , \6370 , \6371 );
xor \U$6184 ( \6373 , \6368 , \6372 );
xor \U$6185 ( \6374 , \6359 , \6373 );
and \U$6186 ( \6375 , \6251 , \6265 );
and \U$6187 ( \6376 , \6265 , \6280 );
and \U$6188 ( \6377 , \6251 , \6280 );
or \U$6189 ( \6378 , \6375 , \6376 , \6377 );
and \U$6190 ( \6379 , \5873 , \5891 );
and \U$6191 ( \6380 , \5842 , \5889 );
nor \U$6192 ( \6381 , \6379 , \6380 );
xnor \U$6193 ( \6382 , \6381 , \5898 );
and \U$6194 ( \6383 , \5893 , \5916 );
and \U$6195 ( \6384 , \5861 , \5914 );
nor \U$6196 ( \6385 , \6383 , \6384 );
xnor \U$6197 ( \6386 , \6385 , \5923 );
xor \U$6198 ( \6387 , \6382 , \6386 );
and \U$6199 ( \6388 , \5918 , \5935 );
and \U$6200 ( \6389 , \5881 , \5933 );
nor \U$6201 ( \6390 , \6388 , \6389 );
xnor \U$6202 ( \6391 , \6390 , \5942 );
xor \U$6203 ( \6392 , \6387 , \6391 );
and \U$6204 ( \6393 , \5811 , \5829 );
and \U$6205 ( \6394 , \5780 , \5827 );
nor \U$6206 ( \6395 , \6393 , \6394 );
xnor \U$6207 ( \6396 , \6395 , \5836 );
and \U$6208 ( \6397 , \5831 , \5852 );
and \U$6209 ( \6398 , \5799 , \5850 );
nor \U$6210 ( \6399 , \6397 , \6398 );
xnor \U$6211 ( \6400 , \6399 , \5859 );
xor \U$6212 ( \6401 , \6396 , \6400 );
and \U$6213 ( \6402 , \5854 , \5871 );
and \U$6214 ( \6403 , \5819 , \5869 );
nor \U$6215 ( \6404 , \6402 , \6403 );
xnor \U$6216 ( \6405 , \6404 , \5878 );
xor \U$6217 ( \6406 , \6401 , \6405 );
xor \U$6218 ( \6407 , \6392 , \6406 );
not \U$6219 ( \6408 , \5775 );
and \U$6220 ( \6409 , \5770 , \5790 );
and \U$6221 ( \6410 , \5737 , \5788 );
nor \U$6222 ( \6411 , \6409 , \6410 );
xnor \U$6223 ( \6412 , \6411 , \5797 );
xor \U$6224 ( \6413 , \6408 , \6412 );
and \U$6225 ( \6414 , \5792 , \5809 );
and \U$6226 ( \6415 , \5758 , \5807 );
nor \U$6227 ( \6416 , \6414 , \6415 );
xnor \U$6228 ( \6417 , \6416 , \5816 );
xor \U$6229 ( \6418 , \6413 , \6417 );
xor \U$6230 ( \6419 , \6407 , \6418 );
xor \U$6231 ( \6420 , \6378 , \6419 );
and \U$6232 ( \6421 , \6057 , \6082 );
and \U$6233 ( \6422 , \6029 , \6066 );
nor \U$6234 ( \6423 , \6421 , \6422 );
xnor \U$6235 ( \6424 , \6423 , \5736 );
xor \U$6236 ( \6425 , \6221 , \6224 );
not \U$6237 ( \6426 , \6295 );
and \U$6238 ( \6427 , \6425 , \6426 );
and \U$6239 ( \6428 , \6065 , \6427 );
and \U$6240 ( \6429 , \6048 , \6295 );
nor \U$6241 ( \6430 , \6428 , \6429 );
xnor \U$6242 ( \6431 , \6430 , \6227 );
xor \U$6243 ( \6432 , \6424 , \6431 );
and \U$6244 ( \6433 , \5998 , \6016 );
and \U$6245 ( \6434 , \5967 , \6014 );
nor \U$6246 ( \6435 , \6433 , \6434 );
xnor \U$6247 ( \6436 , \6435 , \6023 );
and \U$6248 ( \6437 , \6018 , \6039 );
and \U$6249 ( \6438 , \5986 , \6037 );
nor \U$6250 ( \6439 , \6437 , \6438 );
xnor \U$6251 ( \6440 , \6439 , \6046 );
xor \U$6252 ( \6441 , \6436 , \6440 );
and \U$6253 ( \6442 , \6041 , \6055 );
and \U$6254 ( \6443 , \6006 , \6053 );
nor \U$6255 ( \6444 , \6442 , \6443 );
xnor \U$6256 ( \6445 , \6444 , \6062 );
xor \U$6257 ( \6446 , \6441 , \6445 );
xor \U$6258 ( \6447 , \6432 , \6446 );
and \U$6259 ( \6448 , \5937 , \5955 );
and \U$6260 ( \6449 , \5906 , \5953 );
nor \U$6261 ( \6450 , \6448 , \6449 );
xnor \U$6262 ( \6451 , \6450 , \5962 );
and \U$6263 ( \6452 , \5957 , \5977 );
and \U$6264 ( \6453 , \5925 , \5975 );
nor \U$6265 ( \6454 , \6452 , \6453 );
xnor \U$6266 ( \6455 , \6454 , \5984 );
xor \U$6267 ( \6456 , \6451 , \6455 );
and \U$6268 ( \6457 , \5979 , \5996 );
and \U$6269 ( \6458 , \5945 , \5994 );
nor \U$6270 ( \6459 , \6457 , \6458 );
xnor \U$6271 ( \6460 , \6459 , \6003 );
xor \U$6272 ( \6461 , \6456 , \6460 );
xor \U$6273 ( \6462 , \6447 , \6461 );
xor \U$6274 ( \6463 , \6420 , \6462 );
and \U$6275 ( \6464 , \6374 , \6463 );
and \U$6276 ( \6465 , \6329 , \6333 );
and \U$6277 ( \6466 , \6333 , \6338 );
and \U$6278 ( \6467 , \6329 , \6338 );
or \U$6279 ( \6468 , \6465 , \6466 , \6467 );
and \U$6280 ( \6469 , \6317 , \6321 );
and \U$6281 ( \6470 , \6321 , \6323 );
and \U$6282 ( \6471 , \6317 , \6323 );
or \U$6283 ( \6472 , \6469 , \6470 , \6471 );
xor \U$6284 ( \6473 , \6468 , \6472 );
or \U$6285 ( \6474 , \6298 , \6312 );
xor \U$6286 ( \6475 , \6473 , \6474 );
and \U$6287 ( \6476 , \6463 , \6475 );
and \U$6288 ( \6477 , \6374 , \6475 );
or \U$6289 ( \6478 , \6464 , \6476 , \6477 );
and \U$6290 ( \6479 , \6345 , \6478 );
and \U$6291 ( \6480 , \6029 , \6082 );
and \U$6292 ( \6481 , \6041 , \6066 );
nor \U$6293 ( \6482 , \6480 , \6481 );
xnor \U$6294 ( \6483 , \6482 , \5736 );
and \U$6295 ( \6484 , \6048 , \6427 );
and \U$6296 ( \6485 , \6057 , \6295 );
nor \U$6297 ( \6486 , \6484 , \6485 );
xnor \U$6298 ( \6487 , \6486 , \6227 );
xor \U$6299 ( \6488 , \6483 , \6487 );
and \U$6300 ( \6489 , \6186 , \6190 );
and \U$6301 ( \6490 , \6190 , \6192 );
and \U$6302 ( \6491 , \6186 , \6192 );
or \U$6303 ( \6492 , \6489 , \6490 , \6491 );
and \U$6304 ( \6493 , \159 , \351 );
not \U$6305 ( \6494 , \6493 );
xnor \U$6306 ( \6495 , \6494 , \358 );
and \U$6307 ( \6496 , \315 , \345 );
xnor \U$6308 ( \6497 , \6495 , \6496 );
xor \U$6309 ( \6498 , \6492 , \6497 );
and \U$6310 ( \6499 , \6177 , \6184 );
and \U$6311 ( \6500 , \6184 , \6193 );
and \U$6312 ( \6501 , \6177 , \6193 );
or \U$6313 ( \6502 , \6499 , \6500 , \6501 );
xor \U$6314 ( \6503 , \6498 , \6502 );
and \U$6315 ( \6504 , \6194 , \6207 );
and \U$6316 ( \6505 , \6208 , \6218 );
or \U$6317 ( \6506 , \6504 , \6505 );
xor \U$6318 ( \6507 , \6503 , \6506 );
buf \U$6319 ( \6508 , \6507 );
buf \U$6320 ( \6509 , \6508 );
xor \U$6321 ( \6510 , \6509 , \6221 );
nand \U$6322 ( \6511 , \6065 , \6510 );
or \U$6323 ( \6512 , \6495 , \6496 );
not \U$6324 ( \6513 , \358 );
xor \U$6325 ( \6514 , \6512 , \6513 );
and \U$6326 ( \6515 , \159 , \345 );
xor \U$6327 ( \6516 , \6514 , \6515 );
and \U$6328 ( \6517 , \6492 , \6497 );
xor \U$6329 ( \6518 , \6516 , \6517 );
and \U$6330 ( \6519 , \6498 , \6502 );
and \U$6331 ( \6520 , \6503 , \6506 );
or \U$6332 ( \6521 , \6519 , \6520 );
xor \U$6333 ( \6522 , \6518 , \6521 );
buf \U$6334 ( \6523 , \6522 );
buf \U$6335 ( \6524 , \6523 );
and \U$6336 ( \6525 , \6509 , \6221 );
not \U$6337 ( \6526 , \6525 );
and \U$6338 ( \6527 , \6524 , \6526 );
xnor \U$6339 ( \6528 , \6511 , \6527 );
xor \U$6340 ( \6529 , \6488 , \6528 );
and \U$6341 ( \6530 , \5967 , \6016 );
and \U$6342 ( \6531 , \5979 , \6014 );
nor \U$6343 ( \6532 , \6530 , \6531 );
xnor \U$6344 ( \6533 , \6532 , \6023 );
and \U$6345 ( \6534 , \5986 , \6039 );
and \U$6346 ( \6535 , \5998 , \6037 );
nor \U$6347 ( \6536 , \6534 , \6535 );
xnor \U$6348 ( \6537 , \6536 , \6046 );
xor \U$6349 ( \6538 , \6533 , \6537 );
and \U$6350 ( \6539 , \6006 , \6055 );
and \U$6351 ( \6540 , \6018 , \6053 );
nor \U$6352 ( \6541 , \6539 , \6540 );
xnor \U$6353 ( \6542 , \6541 , \6062 );
xor \U$6354 ( \6543 , \6538 , \6542 );
xnor \U$6355 ( \6544 , \6529 , \6543 );
and \U$6356 ( \6545 , \6451 , \6455 );
and \U$6357 ( \6546 , \6455 , \6460 );
and \U$6358 ( \6547 , \6451 , \6460 );
or \U$6359 ( \6548 , \6545 , \6546 , \6547 );
and \U$6360 ( \6549 , \6436 , \6440 );
and \U$6361 ( \6550 , \6440 , \6445 );
and \U$6362 ( \6551 , \6436 , \6445 );
or \U$6363 ( \6552 , \6549 , \6550 , \6551 );
xor \U$6364 ( \6553 , \6548 , \6552 );
and \U$6365 ( \6554 , \6424 , \6431 );
xor \U$6366 ( \6555 , \6553 , \6554 );
xor \U$6367 ( \6556 , \6544 , \6555 );
and \U$6368 ( \6557 , \6408 , \6412 );
and \U$6369 ( \6558 , \6412 , \6417 );
and \U$6370 ( \6559 , \6408 , \6417 );
or \U$6371 ( \6560 , \6557 , \6558 , \6559 );
and \U$6372 ( \6561 , \6396 , \6400 );
and \U$6373 ( \6562 , \6400 , \6405 );
and \U$6374 ( \6563 , \6396 , \6405 );
or \U$6375 ( \6564 , \6561 , \6562 , \6563 );
xor \U$6376 ( \6565 , \6560 , \6564 );
and \U$6377 ( \6566 , \6382 , \6386 );
and \U$6378 ( \6567 , \6386 , \6391 );
and \U$6379 ( \6568 , \6382 , \6391 );
or \U$6380 ( \6569 , \6566 , \6567 , \6568 );
xor \U$6381 ( \6570 , \6565 , \6569 );
xor \U$6382 ( \6571 , \6556 , \6570 );
and \U$6383 ( \6572 , \6392 , \6406 );
and \U$6384 ( \6573 , \6406 , \6418 );
and \U$6385 ( \6574 , \6392 , \6418 );
or \U$6386 ( \6575 , \6572 , \6573 , \6574 );
and \U$6387 ( \6576 , \5737 , \5790 );
not \U$6388 ( \6577 , \6576 );
xnor \U$6389 ( \6578 , \6577 , \5797 );
xor \U$6390 ( \6579 , \6527 , \6578 );
and \U$6391 ( \6580 , \5758 , \5809 );
and \U$6392 ( \6581 , \5770 , \5807 );
nor \U$6393 ( \6582 , \6580 , \6581 );
xnor \U$6394 ( \6583 , \6582 , \5816 );
xor \U$6395 ( \6584 , \6579 , \6583 );
xor \U$6396 ( \6585 , \6575 , \6584 );
and \U$6397 ( \6586 , \5906 , \5955 );
and \U$6398 ( \6587 , \5918 , \5953 );
nor \U$6399 ( \6588 , \6586 , \6587 );
xnor \U$6400 ( \6589 , \6588 , \5962 );
and \U$6401 ( \6590 , \5925 , \5977 );
and \U$6402 ( \6591 , \5937 , \5975 );
nor \U$6403 ( \6592 , \6590 , \6591 );
xnor \U$6404 ( \6593 , \6592 , \5984 );
xor \U$6405 ( \6594 , \6589 , \6593 );
and \U$6406 ( \6595 , \5945 , \5996 );
and \U$6407 ( \6596 , \5957 , \5994 );
nor \U$6408 ( \6597 , \6595 , \6596 );
xnor \U$6409 ( \6598 , \6597 , \6003 );
xor \U$6410 ( \6599 , \6594 , \6598 );
and \U$6411 ( \6600 , \5842 , \5891 );
and \U$6412 ( \6601 , \5854 , \5889 );
nor \U$6413 ( \6602 , \6600 , \6601 );
xnor \U$6414 ( \6603 , \6602 , \5898 );
and \U$6415 ( \6604 , \5861 , \5916 );
and \U$6416 ( \6605 , \5873 , \5914 );
nor \U$6417 ( \6606 , \6604 , \6605 );
xnor \U$6418 ( \6607 , \6606 , \5923 );
xor \U$6419 ( \6608 , \6603 , \6607 );
and \U$6420 ( \6609 , \5881 , \5935 );
and \U$6421 ( \6610 , \5893 , \5933 );
nor \U$6422 ( \6611 , \6609 , \6610 );
xnor \U$6423 ( \6612 , \6611 , \5942 );
xor \U$6424 ( \6613 , \6608 , \6612 );
xor \U$6425 ( \6614 , \6599 , \6613 );
and \U$6426 ( \6615 , \5780 , \5829 );
and \U$6427 ( \6616 , \5792 , \5827 );
nor \U$6428 ( \6617 , \6615 , \6616 );
xnor \U$6429 ( \6618 , \6617 , \5836 );
and \U$6430 ( \6619 , \5799 , \5852 );
and \U$6431 ( \6620 , \5811 , \5850 );
nor \U$6432 ( \6621 , \6619 , \6620 );
xnor \U$6433 ( \6622 , \6621 , \5859 );
xor \U$6434 ( \6623 , \6618 , \6622 );
and \U$6435 ( \6624 , \5819 , \5871 );
and \U$6436 ( \6625 , \5831 , \5869 );
nor \U$6437 ( \6626 , \6624 , \6625 );
xnor \U$6438 ( \6627 , \6626 , \5878 );
xor \U$6439 ( \6628 , \6623 , \6627 );
xor \U$6440 ( \6629 , \6614 , \6628 );
xor \U$6441 ( \6630 , \6585 , \6629 );
xor \U$6442 ( \6631 , \6571 , \6630 );
and \U$6443 ( \6632 , \6363 , \6367 );
and \U$6444 ( \6633 , \6367 , \6372 );
and \U$6445 ( \6634 , \6363 , \6372 );
or \U$6446 ( \6635 , \6632 , \6633 , \6634 );
and \U$6447 ( \6636 , \6349 , \6353 );
and \U$6448 ( \6637 , \6353 , \6358 );
and \U$6449 ( \6638 , \6349 , \6358 );
or \U$6450 ( \6639 , \6636 , \6637 , \6638 );
xor \U$6451 ( \6640 , \6635 , \6639 );
and \U$6452 ( \6641 , \6432 , \6446 );
and \U$6453 ( \6642 , \6446 , \6461 );
and \U$6454 ( \6643 , \6432 , \6461 );
or \U$6455 ( \6644 , \6641 , \6642 , \6643 );
xor \U$6456 ( \6645 , \6640 , \6644 );
xor \U$6457 ( \6646 , \6631 , \6645 );
and \U$6458 ( \6647 , \6478 , \6646 );
and \U$6459 ( \6648 , \6345 , \6646 );
or \U$6460 ( \6649 , \6479 , \6647 , \6648 );
and \U$6461 ( \6650 , \6635 , \6639 );
and \U$6462 ( \6651 , \6639 , \6644 );
and \U$6463 ( \6652 , \6635 , \6644 );
or \U$6464 ( \6653 , \6650 , \6651 , \6652 );
and \U$6465 ( \6654 , \6575 , \6584 );
and \U$6466 ( \6655 , \6584 , \6629 );
and \U$6467 ( \6656 , \6575 , \6629 );
or \U$6468 ( \6657 , \6654 , \6655 , \6656 );
xor \U$6469 ( \6658 , \6653 , \6657 );
and \U$6470 ( \6659 , \6544 , \6555 );
and \U$6471 ( \6660 , \6555 , \6570 );
and \U$6472 ( \6661 , \6544 , \6570 );
or \U$6473 ( \6662 , \6659 , \6660 , \6661 );
xor \U$6474 ( \6663 , \6658 , \6662 );
xor \U$6475 ( \6664 , \6649 , \6663 );
and \U$6476 ( \6665 , \6468 , \6472 );
and \U$6477 ( \6666 , \6472 , \6474 );
and \U$6478 ( \6667 , \6468 , \6474 );
or \U$6479 ( \6668 , \6665 , \6666 , \6667 );
and \U$6480 ( \6669 , \6378 , \6419 );
and \U$6481 ( \6670 , \6419 , \6462 );
and \U$6482 ( \6671 , \6378 , \6462 );
or \U$6483 ( \6672 , \6669 , \6670 , \6671 );
and \U$6484 ( \6673 , \6668 , \6672 );
and \U$6485 ( \6674 , \6359 , \6373 );
and \U$6486 ( \6675 , \6672 , \6674 );
and \U$6487 ( \6676 , \6668 , \6674 );
or \U$6488 ( \6677 , \6673 , \6675 , \6676 );
and \U$6489 ( \6678 , \6571 , \6630 );
and \U$6490 ( \6679 , \6630 , \6645 );
and \U$6491 ( \6680 , \6571 , \6645 );
or \U$6492 ( \6681 , \6678 , \6679 , \6680 );
xor \U$6493 ( \6682 , \6677 , \6681 );
and \U$6494 ( \6683 , \6589 , \6593 );
and \U$6495 ( \6684 , \6593 , \6598 );
and \U$6496 ( \6685 , \6589 , \6598 );
or \U$6497 ( \6686 , \6683 , \6684 , \6685 );
and \U$6498 ( \6687 , \6533 , \6537 );
and \U$6499 ( \6688 , \6537 , \6542 );
and \U$6500 ( \6689 , \6533 , \6542 );
or \U$6501 ( \6690 , \6687 , \6688 , \6689 );
xor \U$6502 ( \6691 , \6686 , \6690 );
and \U$6503 ( \6692 , \6483 , \6487 );
and \U$6504 ( \6693 , \6487 , \6528 );
and \U$6505 ( \6694 , \6483 , \6528 );
or \U$6506 ( \6695 , \6692 , \6693 , \6694 );
xor \U$6507 ( \6696 , \6691 , \6695 );
and \U$6508 ( \6697 , \6527 , \6578 );
and \U$6509 ( \6698 , \6578 , \6583 );
and \U$6510 ( \6699 , \6527 , \6583 );
or \U$6511 ( \6700 , \6697 , \6698 , \6699 );
and \U$6512 ( \6701 , \6618 , \6622 );
and \U$6513 ( \6702 , \6622 , \6627 );
and \U$6514 ( \6703 , \6618 , \6627 );
or \U$6515 ( \6704 , \6701 , \6702 , \6703 );
xor \U$6516 ( \6705 , \6700 , \6704 );
and \U$6517 ( \6706 , \6603 , \6607 );
and \U$6518 ( \6707 , \6607 , \6612 );
and \U$6519 ( \6708 , \6603 , \6612 );
or \U$6520 ( \6709 , \6706 , \6707 , \6708 );
xor \U$6521 ( \6710 , \6705 , \6709 );
xor \U$6522 ( \6711 , \6696 , \6710 );
and \U$6523 ( \6712 , \6599 , \6613 );
and \U$6524 ( \6713 , \6613 , \6628 );
and \U$6525 ( \6714 , \6599 , \6628 );
or \U$6526 ( \6715 , \6712 , \6713 , \6714 );
and \U$6527 ( \6716 , \5873 , \5916 );
and \U$6528 ( \6717 , \5842 , \5914 );
nor \U$6529 ( \6718 , \6716 , \6717 );
xnor \U$6530 ( \6719 , \6718 , \5923 );
and \U$6531 ( \6720 , \5893 , \5935 );
and \U$6532 ( \6721 , \5861 , \5933 );
nor \U$6533 ( \6722 , \6720 , \6721 );
xnor \U$6534 ( \6723 , \6722 , \5942 );
xor \U$6535 ( \6724 , \6719 , \6723 );
and \U$6536 ( \6725 , \5918 , \5955 );
and \U$6537 ( \6726 , \5881 , \5953 );
nor \U$6538 ( \6727 , \6725 , \6726 );
xnor \U$6539 ( \6728 , \6727 , \5962 );
xor \U$6540 ( \6729 , \6724 , \6728 );
and \U$6541 ( \6730 , \5811 , \5852 );
and \U$6542 ( \6731 , \5780 , \5850 );
nor \U$6543 ( \6732 , \6730 , \6731 );
xnor \U$6544 ( \6733 , \6732 , \5859 );
and \U$6545 ( \6734 , \5831 , \5871 );
and \U$6546 ( \6735 , \5799 , \5869 );
nor \U$6547 ( \6736 , \6734 , \6735 );
xnor \U$6548 ( \6737 , \6736 , \5878 );
xor \U$6549 ( \6738 , \6733 , \6737 );
and \U$6550 ( \6739 , \5854 , \5891 );
and \U$6551 ( \6740 , \5819 , \5889 );
nor \U$6552 ( \6741 , \6739 , \6740 );
xnor \U$6553 ( \6742 , \6741 , \5898 );
xor \U$6554 ( \6743 , \6738 , \6742 );
xor \U$6555 ( \6744 , \6729 , \6743 );
not \U$6556 ( \6745 , \5797 );
and \U$6557 ( \6746 , \5770 , \5809 );
and \U$6558 ( \6747 , \5737 , \5807 );
nor \U$6559 ( \6748 , \6746 , \6747 );
xnor \U$6560 ( \6749 , \6748 , \5816 );
xor \U$6561 ( \6750 , \6745 , \6749 );
and \U$6562 ( \6751 , \5792 , \5829 );
and \U$6563 ( \6752 , \5758 , \5827 );
nor \U$6564 ( \6753 , \6751 , \6752 );
xnor \U$6565 ( \6754 , \6753 , \5836 );
xor \U$6566 ( \6755 , \6750 , \6754 );
xor \U$6567 ( \6756 , \6744 , \6755 );
xor \U$6568 ( \6757 , \6715 , \6756 );
and \U$6569 ( \6758 , \6057 , \6427 );
and \U$6570 ( \6759 , \6029 , \6295 );
nor \U$6571 ( \6760 , \6758 , \6759 );
xnor \U$6572 ( \6761 , \6760 , \6227 );
xor \U$6573 ( \6762 , \6524 , \6509 );
not \U$6574 ( \6763 , \6510 );
and \U$6575 ( \6764 , \6762 , \6763 );
and \U$6576 ( \6765 , \6065 , \6764 );
and \U$6577 ( \6766 , \6048 , \6510 );
nor \U$6578 ( \6767 , \6765 , \6766 );
xnor \U$6579 ( \6768 , \6767 , \6527 );
xor \U$6580 ( \6769 , \6761 , \6768 );
and \U$6581 ( \6770 , \5998 , \6039 );
and \U$6582 ( \6771 , \5967 , \6037 );
nor \U$6583 ( \6772 , \6770 , \6771 );
xnor \U$6584 ( \6773 , \6772 , \6046 );
and \U$6585 ( \6774 , \6018 , \6055 );
and \U$6586 ( \6775 , \5986 , \6053 );
nor \U$6587 ( \6776 , \6774 , \6775 );
xnor \U$6588 ( \6777 , \6776 , \6062 );
xor \U$6589 ( \6778 , \6773 , \6777 );
and \U$6590 ( \6779 , \6041 , \6082 );
and \U$6591 ( \6780 , \6006 , \6066 );
nor \U$6592 ( \6781 , \6779 , \6780 );
xnor \U$6593 ( \6782 , \6781 , \5736 );
xor \U$6594 ( \6783 , \6778 , \6782 );
xor \U$6595 ( \6784 , \6769 , \6783 );
and \U$6596 ( \6785 , \5937 , \5977 );
and \U$6597 ( \6786 , \5906 , \5975 );
nor \U$6598 ( \6787 , \6785 , \6786 );
xnor \U$6599 ( \6788 , \6787 , \5984 );
and \U$6600 ( \6789 , \5957 , \5996 );
and \U$6601 ( \6790 , \5925 , \5994 );
nor \U$6602 ( \6791 , \6789 , \6790 );
xnor \U$6603 ( \6792 , \6791 , \6003 );
xor \U$6604 ( \6793 , \6788 , \6792 );
and \U$6605 ( \6794 , \5979 , \6016 );
and \U$6606 ( \6795 , \5945 , \6014 );
nor \U$6607 ( \6796 , \6794 , \6795 );
xnor \U$6608 ( \6797 , \6796 , \6023 );
xor \U$6609 ( \6798 , \6793 , \6797 );
xor \U$6610 ( \6799 , \6784 , \6798 );
xor \U$6611 ( \6800 , \6757 , \6799 );
xor \U$6612 ( \6801 , \6711 , \6800 );
and \U$6613 ( \6802 , \6560 , \6564 );
and \U$6614 ( \6803 , \6564 , \6569 );
and \U$6615 ( \6804 , \6560 , \6569 );
or \U$6616 ( \6805 , \6802 , \6803 , \6804 );
and \U$6617 ( \6806 , \6548 , \6552 );
and \U$6618 ( \6807 , \6552 , \6554 );
and \U$6619 ( \6808 , \6548 , \6554 );
or \U$6620 ( \6809 , \6806 , \6807 , \6808 );
xor \U$6621 ( \6810 , \6805 , \6809 );
or \U$6622 ( \6811 , \6529 , \6543 );
xor \U$6623 ( \6812 , \6810 , \6811 );
xor \U$6624 ( \6813 , \6801 , \6812 );
xor \U$6625 ( \6814 , \6682 , \6813 );
xor \U$6626 ( \6815 , \6664 , \6814 );
xor \U$6627 ( \6816 , \4668 , \5654 );
buf \U$6628 ( \6817 , \6816 );
buf \U$6629 ( \6818 , \6817 );
xor \U$6630 ( \6819 , \4760 , \5652 );
buf \U$6631 ( \6820 , \6819 );
buf \U$6632 ( \6821 , \6820 );
and \U$6633 ( \6822 , \6818 , \6821 );
not \U$6634 ( \6823 , \6822 );
and \U$6635 ( \6824 , \5747 , \6823 );
not \U$6636 ( \6825 , \6824 );
and \U$6637 ( \6826 , \5770 , \5750 );
and \U$6638 ( \6827 , \5737 , \5748 );
nor \U$6639 ( \6828 , \6826 , \6827 );
xnor \U$6640 ( \6829 , \6828 , \5755 );
and \U$6641 ( \6830 , \6825 , \6829 );
and \U$6642 ( \6831 , \5792 , \5768 );
and \U$6643 ( \6832 , \5758 , \5766 );
nor \U$6644 ( \6833 , \6831 , \6832 );
xnor \U$6645 ( \6834 , \6833 , \5775 );
and \U$6646 ( \6835 , \6829 , \6834 );
and \U$6647 ( \6836 , \6825 , \6834 );
or \U$6648 ( \6837 , \6830 , \6835 , \6836 );
and \U$6649 ( \6838 , \5811 , \5790 );
and \U$6650 ( \6839 , \5780 , \5788 );
nor \U$6651 ( \6840 , \6838 , \6839 );
xnor \U$6652 ( \6841 , \6840 , \5797 );
and \U$6653 ( \6842 , \5831 , \5809 );
and \U$6654 ( \6843 , \5799 , \5807 );
nor \U$6655 ( \6844 , \6842 , \6843 );
xnor \U$6656 ( \6845 , \6844 , \5816 );
and \U$6657 ( \6846 , \6841 , \6845 );
and \U$6658 ( \6847 , \5854 , \5829 );
and \U$6659 ( \6848 , \5819 , \5827 );
nor \U$6660 ( \6849 , \6847 , \6848 );
xnor \U$6661 ( \6850 , \6849 , \5836 );
and \U$6662 ( \6851 , \6845 , \6850 );
and \U$6663 ( \6852 , \6841 , \6850 );
or \U$6664 ( \6853 , \6846 , \6851 , \6852 );
and \U$6665 ( \6854 , \6837 , \6853 );
and \U$6666 ( \6855 , \5873 , \5852 );
and \U$6667 ( \6856 , \5842 , \5850 );
nor \U$6668 ( \6857 , \6855 , \6856 );
xnor \U$6669 ( \6858 , \6857 , \5859 );
and \U$6670 ( \6859 , \5893 , \5871 );
and \U$6671 ( \6860 , \5861 , \5869 );
nor \U$6672 ( \6861 , \6859 , \6860 );
xnor \U$6673 ( \6862 , \6861 , \5878 );
and \U$6674 ( \6863 , \6858 , \6862 );
and \U$6675 ( \6864 , \5918 , \5891 );
and \U$6676 ( \6865 , \5881 , \5889 );
nor \U$6677 ( \6866 , \6864 , \6865 );
xnor \U$6678 ( \6867 , \6866 , \5898 );
and \U$6679 ( \6868 , \6862 , \6867 );
and \U$6680 ( \6869 , \6858 , \6867 );
or \U$6681 ( \6870 , \6863 , \6868 , \6869 );
and \U$6682 ( \6871 , \6853 , \6870 );
and \U$6683 ( \6872 , \6837 , \6870 );
or \U$6684 ( \6873 , \6854 , \6871 , \6872 );
and \U$6685 ( \6874 , \5937 , \5916 );
and \U$6686 ( \6875 , \5906 , \5914 );
nor \U$6687 ( \6876 , \6874 , \6875 );
xnor \U$6688 ( \6877 , \6876 , \5923 );
and \U$6689 ( \6878 , \5957 , \5935 );
and \U$6690 ( \6879 , \5925 , \5933 );
nor \U$6691 ( \6880 , \6878 , \6879 );
xnor \U$6692 ( \6881 , \6880 , \5942 );
and \U$6693 ( \6882 , \6877 , \6881 );
and \U$6694 ( \6883 , \5979 , \5955 );
and \U$6695 ( \6884 , \5945 , \5953 );
nor \U$6696 ( \6885 , \6883 , \6884 );
xnor \U$6697 ( \6886 , \6885 , \5962 );
and \U$6698 ( \6887 , \6881 , \6886 );
and \U$6699 ( \6888 , \6877 , \6886 );
or \U$6700 ( \6889 , \6882 , \6887 , \6888 );
and \U$6701 ( \6890 , \5998 , \5977 );
and \U$6702 ( \6891 , \5967 , \5975 );
nor \U$6703 ( \6892 , \6890 , \6891 );
xnor \U$6704 ( \6893 , \6892 , \5984 );
and \U$6705 ( \6894 , \6018 , \5996 );
and \U$6706 ( \6895 , \5986 , \5994 );
nor \U$6707 ( \6896 , \6894 , \6895 );
xnor \U$6708 ( \6897 , \6896 , \6003 );
and \U$6709 ( \6898 , \6893 , \6897 );
and \U$6710 ( \6899 , \6041 , \6016 );
and \U$6711 ( \6900 , \6006 , \6014 );
nor \U$6712 ( \6901 , \6899 , \6900 );
xnor \U$6713 ( \6902 , \6901 , \6023 );
and \U$6714 ( \6903 , \6897 , \6902 );
and \U$6715 ( \6904 , \6893 , \6902 );
or \U$6716 ( \6905 , \6898 , \6903 , \6904 );
and \U$6717 ( \6906 , \6889 , \6905 );
and \U$6718 ( \6907 , \6057 , \6039 );
and \U$6719 ( \6908 , \6029 , \6037 );
nor \U$6720 ( \6909 , \6907 , \6908 );
xnor \U$6721 ( \6910 , \6909 , \6046 );
and \U$6722 ( \6911 , \6065 , \6055 );
and \U$6723 ( \6912 , \6048 , \6053 );
nor \U$6724 ( \6913 , \6911 , \6912 );
xnor \U$6725 ( \6914 , \6913 , \6062 );
and \U$6726 ( \6915 , \6910 , \6914 );
and \U$6727 ( \6916 , \6905 , \6915 );
and \U$6728 ( \6917 , \6889 , \6915 );
or \U$6729 ( \6918 , \6906 , \6916 , \6917 );
and \U$6730 ( \6919 , \6873 , \6918 );
xor \U$6731 ( \6920 , \6047 , \6063 );
xor \U$6732 ( \6921 , \6920 , \6068 );
xor \U$6733 ( \6922 , \5985 , \6004 );
xor \U$6734 ( \6923 , \6922 , \6024 );
or \U$6735 ( \6924 , \6921 , \6923 );
and \U$6736 ( \6925 , \6918 , \6924 );
and \U$6737 ( \6926 , \6873 , \6924 );
or \U$6738 ( \6927 , \6919 , \6925 , \6926 );
xor \U$6739 ( \6928 , \5924 , \5943 );
xor \U$6740 ( \6929 , \6928 , \5963 );
xor \U$6741 ( \6930 , \5860 , \5879 );
xor \U$6742 ( \6931 , \6930 , \5899 );
and \U$6743 ( \6932 , \6929 , \6931 );
xor \U$6744 ( \6933 , \5798 , \5817 );
xor \U$6745 ( \6934 , \6933 , \5837 );
and \U$6746 ( \6935 , \6931 , \6934 );
and \U$6747 ( \6936 , \6929 , \6934 );
or \U$6748 ( \6937 , \6932 , \6935 , \6936 );
xor \U$6749 ( \6938 , \6136 , \6150 );
xor \U$6750 ( \6939 , \6938 , \6162 );
and \U$6751 ( \6940 , \6937 , \6939 );
xor \U$6752 ( \6941 , \6087 , \6101 );
xor \U$6753 ( \6942 , \6941 , \6116 );
and \U$6754 ( \6943 , \6939 , \6942 );
and \U$6755 ( \6944 , \6937 , \6942 );
or \U$6756 ( \6945 , \6940 , \6943 , \6944 );
and \U$6757 ( \6946 , \6927 , \6945 );
xor \U$6758 ( \6947 , \5966 , \6027 );
xor \U$6759 ( \6948 , \6947 , \6071 );
xor \U$6760 ( \6949 , \5779 , \5840 );
xor \U$6761 ( \6950 , \6949 , \5902 );
and \U$6762 ( \6951 , \6948 , \6950 );
and \U$6763 ( \6952 , \6945 , \6951 );
and \U$6764 ( \6953 , \6927 , \6951 );
or \U$6765 ( \6954 , \6946 , \6952 , \6953 );
xor \U$6766 ( \6955 , \6313 , \6324 );
xor \U$6767 ( \6956 , \6955 , \6339 );
xor \U$6768 ( \6957 , \6165 , \6236 );
xor \U$6769 ( \6958 , \6957 , \6281 );
and \U$6770 ( \6959 , \6956 , \6958 );
xor \U$6771 ( \6960 , \5905 , \6074 );
xor \U$6772 ( \6961 , \6960 , \6119 );
and \U$6773 ( \6962 , \6958 , \6961 );
and \U$6774 ( \6963 , \6956 , \6961 );
or \U$6775 ( \6964 , \6959 , \6962 , \6963 );
and \U$6776 ( \6965 , \6954 , \6964 );
xor \U$6777 ( \6966 , \6374 , \6463 );
xor \U$6778 ( \6967 , \6966 , \6475 );
and \U$6779 ( \6968 , \6964 , \6967 );
and \U$6780 ( \6969 , \6954 , \6967 );
or \U$6781 ( \6970 , \6965 , \6968 , \6969 );
xor \U$6782 ( \6971 , \6668 , \6672 );
xor \U$6783 ( \6972 , \6971 , \6674 );
and \U$6784 ( \6973 , \6970 , \6972 );
xor \U$6785 ( \6974 , \6345 , \6478 );
xor \U$6786 ( \6975 , \6974 , \6646 );
and \U$6787 ( \6976 , \6972 , \6975 );
and \U$6788 ( \6977 , \6970 , \6975 );
or \U$6789 ( \6978 , \6973 , \6976 , \6977 );
nand \U$6790 ( \6979 , \6815 , \6978 );
nor \U$6791 ( \6980 , \6815 , \6978 );
not \U$6792 ( \6981 , \6980 );
nand \U$6793 ( \6982 , \6979 , \6981 );
xor \U$6794 ( \6983 , \5606 , \5609 );
buf \U$6795 ( \6984 , \6983 );
buf \U$6796 ( \6985 , \6984 );
xor \U$6797 ( \6986 , \5608 , \2371 );
buf \U$6798 ( \6987 , \6986 );
buf \U$6799 ( \6988 , \6987 );
xor \U$6800 ( \6989 , \6985 , \6988 );
not \U$6801 ( \6990 , \6988 );
and \U$6802 ( \6991 , \6989 , \6990 );
and \U$6803 ( \6992 , \5799 , \6991 );
and \U$6804 ( \6993 , \5811 , \6988 );
nor \U$6805 ( \6994 , \6992 , \6993 );
xnor \U$6806 ( \6995 , \6994 , \6985 );
and \U$6807 ( \6996 , \5755 , \6995 );
xor \U$6808 ( \6997 , \5597 , \5612 );
buf \U$6809 ( \6998 , \6997 );
buf \U$6810 ( \6999 , \6998 );
xor \U$6811 ( \7000 , \5602 , \5610 );
buf \U$6812 ( \7001 , \7000 );
buf \U$6813 ( \7002 , \7001 );
xor \U$6814 ( \7003 , \6999 , \7002 );
xor \U$6815 ( \7004 , \7002 , \6985 );
not \U$6816 ( \7005 , \7004 );
and \U$6817 ( \7006 , \7003 , \7005 );
and \U$6818 ( \7007 , \5819 , \7006 );
and \U$6819 ( \7008 , \5831 , \7004 );
nor \U$6820 ( \7009 , \7007 , \7008 );
and \U$6821 ( \7010 , \7002 , \6985 );
not \U$6822 ( \7011 , \7010 );
and \U$6823 ( \7012 , \6999 , \7011 );
xnor \U$6824 ( \7013 , \7009 , \7012 );
and \U$6825 ( \7014 , \6995 , \7013 );
and \U$6826 ( \7015 , \5755 , \7013 );
or \U$6827 ( \7016 , \6996 , \7014 , \7015 );
xor \U$6828 ( \7017 , \5577 , \5616 );
buf \U$6829 ( \7018 , \7017 );
buf \U$6830 ( \7019 , \7018 );
xor \U$6831 ( \7020 , \5589 , \5614 );
buf \U$6832 ( \7021 , \7020 );
buf \U$6833 ( \7022 , \7021 );
xor \U$6834 ( \7023 , \7019 , \7022 );
xor \U$6835 ( \7024 , \7022 , \6999 );
not \U$6836 ( \7025 , \7024 );
and \U$6837 ( \7026 , \7023 , \7025 );
and \U$6838 ( \7027 , \5842 , \7026 );
and \U$6839 ( \7028 , \5854 , \7024 );
nor \U$6840 ( \7029 , \7027 , \7028 );
and \U$6841 ( \7030 , \7022 , \6999 );
not \U$6842 ( \7031 , \7030 );
and \U$6843 ( \7032 , \7019 , \7031 );
xnor \U$6844 ( \7033 , \7029 , \7032 );
xor \U$6845 ( \7034 , \5550 , \5620 );
buf \U$6846 ( \7035 , \7034 );
buf \U$6847 ( \7036 , \7035 );
xor \U$6848 ( \7037 , \5569 , \5618 );
buf \U$6849 ( \7038 , \7037 );
buf \U$6850 ( \7039 , \7038 );
xor \U$6851 ( \7040 , \7036 , \7039 );
xor \U$6852 ( \7041 , \7039 , \7019 );
not \U$6853 ( \7042 , \7041 );
and \U$6854 ( \7043 , \7040 , \7042 );
and \U$6855 ( \7044 , \5861 , \7043 );
and \U$6856 ( \7045 , \5873 , \7041 );
nor \U$6857 ( \7046 , \7044 , \7045 );
and \U$6858 ( \7047 , \7039 , \7019 );
not \U$6859 ( \7048 , \7047 );
and \U$6860 ( \7049 , \7036 , \7048 );
xnor \U$6861 ( \7050 , \7046 , \7049 );
and \U$6862 ( \7051 , \7033 , \7050 );
xor \U$6863 ( \7052 , \5516 , \5624 );
buf \U$6864 ( \7053 , \7052 );
buf \U$6865 ( \7054 , \7053 );
xor \U$6866 ( \7055 , \5524 , \5622 );
buf \U$6867 ( \7056 , \7055 );
buf \U$6868 ( \7057 , \7056 );
xor \U$6869 ( \7058 , \7054 , \7057 );
xor \U$6870 ( \7059 , \7057 , \7036 );
not \U$6871 ( \7060 , \7059 );
and \U$6872 ( \7061 , \7058 , \7060 );
and \U$6873 ( \7062 , \5881 , \7061 );
and \U$6874 ( \7063 , \5893 , \7059 );
nor \U$6875 ( \7064 , \7062 , \7063 );
and \U$6876 ( \7065 , \7057 , \7036 );
not \U$6877 ( \7066 , \7065 );
and \U$6878 ( \7067 , \7054 , \7066 );
xnor \U$6879 ( \7068 , \7064 , \7067 );
and \U$6880 ( \7069 , \7050 , \7068 );
and \U$6881 ( \7070 , \7033 , \7068 );
or \U$6882 ( \7071 , \7051 , \7069 , \7070 );
and \U$6883 ( \7072 , \7016 , \7071 );
xor \U$6884 ( \7073 , \5448 , \5628 );
buf \U$6885 ( \7074 , \7073 );
buf \U$6886 ( \7075 , \7074 );
xor \U$6887 ( \7076 , \5482 , \5626 );
buf \U$6888 ( \7077 , \7076 );
buf \U$6889 ( \7078 , \7077 );
xor \U$6890 ( \7079 , \7075 , \7078 );
xor \U$6891 ( \7080 , \7078 , \7054 );
not \U$6892 ( \7081 , \7080 );
and \U$6893 ( \7082 , \7079 , \7081 );
and \U$6894 ( \7083 , \5906 , \7082 );
and \U$6895 ( \7084 , \5918 , \7080 );
nor \U$6896 ( \7085 , \7083 , \7084 );
and \U$6897 ( \7086 , \7078 , \7054 );
not \U$6898 ( \7087 , \7086 );
and \U$6899 ( \7088 , \7075 , \7087 );
xnor \U$6900 ( \7089 , \7085 , \7088 );
xor \U$6901 ( \7090 , \5387 , \5632 );
buf \U$6902 ( \7091 , \7090 );
buf \U$6903 ( \7092 , \7091 );
xor \U$6904 ( \7093 , \5440 , \5630 );
buf \U$6905 ( \7094 , \7093 );
buf \U$6906 ( \7095 , \7094 );
xor \U$6907 ( \7096 , \7092 , \7095 );
xor \U$6908 ( \7097 , \7095 , \7075 );
not \U$6909 ( \7098 , \7097 );
and \U$6910 ( \7099 , \7096 , \7098 );
and \U$6911 ( \7100 , \5925 , \7099 );
and \U$6912 ( \7101 , \5937 , \7097 );
nor \U$6913 ( \7102 , \7100 , \7101 );
and \U$6914 ( \7103 , \7095 , \7075 );
not \U$6915 ( \7104 , \7103 );
and \U$6916 ( \7105 , \7092 , \7104 );
xnor \U$6917 ( \7106 , \7102 , \7105 );
and \U$6918 ( \7107 , \7089 , \7106 );
xor \U$6919 ( \7108 , \5295 , \5636 );
buf \U$6920 ( \7109 , \7108 );
buf \U$6921 ( \7110 , \7109 );
xor \U$6922 ( \7111 , \5348 , \5634 );
buf \U$6923 ( \7112 , \7111 );
buf \U$6924 ( \7113 , \7112 );
xor \U$6925 ( \7114 , \7110 , \7113 );
xor \U$6926 ( \7115 , \7113 , \7092 );
not \U$6927 ( \7116 , \7115 );
and \U$6928 ( \7117 , \7114 , \7116 );
and \U$6929 ( \7118 , \5945 , \7117 );
and \U$6930 ( \7119 , \5957 , \7115 );
nor \U$6931 ( \7120 , \7118 , \7119 );
and \U$6932 ( \7121 , \7113 , \7092 );
not \U$6933 ( \7122 , \7121 );
and \U$6934 ( \7123 , \7110 , \7122 );
xnor \U$6935 ( \7124 , \7120 , \7123 );
and \U$6936 ( \7125 , \7106 , \7124 );
and \U$6937 ( \7126 , \7089 , \7124 );
or \U$6938 ( \7127 , \7107 , \7125 , \7126 );
and \U$6939 ( \7128 , \7071 , \7127 );
and \U$6940 ( \7129 , \7016 , \7127 );
or \U$6941 ( \7130 , \7072 , \7128 , \7129 );
xor \U$6942 ( \7131 , \5169 , \5640 );
buf \U$6943 ( \7132 , \7131 );
buf \U$6944 ( \7133 , \7132 );
xor \U$6945 ( \7134 , \5224 , \5638 );
buf \U$6946 ( \7135 , \7134 );
buf \U$6947 ( \7136 , \7135 );
xor \U$6948 ( \7137 , \7133 , \7136 );
xor \U$6949 ( \7138 , \7136 , \7110 );
not \U$6950 ( \7139 , \7138 );
and \U$6951 ( \7140 , \7137 , \7139 );
and \U$6952 ( \7141 , \5967 , \7140 );
and \U$6953 ( \7142 , \5979 , \7138 );
nor \U$6954 ( \7143 , \7141 , \7142 );
and \U$6955 ( \7144 , \7136 , \7110 );
not \U$6956 ( \7145 , \7144 );
and \U$6957 ( \7146 , \7133 , \7145 );
xnor \U$6958 ( \7147 , \7143 , \7146 );
xor \U$6959 ( \7148 , \5102 , \5644 );
buf \U$6960 ( \7149 , \7148 );
buf \U$6961 ( \7150 , \7149 );
xor \U$6962 ( \7151 , \5110 , \5642 );
buf \U$6963 ( \7152 , \7151 );
buf \U$6964 ( \7153 , \7152 );
xor \U$6965 ( \7154 , \7150 , \7153 );
xor \U$6966 ( \7155 , \7153 , \7133 );
not \U$6967 ( \7156 , \7155 );
and \U$6968 ( \7157 , \7154 , \7156 );
and \U$6969 ( \7158 , \5986 , \7157 );
and \U$6970 ( \7159 , \5998 , \7155 );
nor \U$6971 ( \7160 , \7158 , \7159 );
and \U$6972 ( \7161 , \7153 , \7133 );
not \U$6973 ( \7162 , \7161 );
and \U$6974 ( \7163 , \7150 , \7162 );
xnor \U$6975 ( \7164 , \7160 , \7163 );
and \U$6976 ( \7165 , \7147 , \7164 );
xor \U$6977 ( \7166 , \4943 , \5648 );
buf \U$6978 ( \7167 , \7166 );
buf \U$6979 ( \7168 , \7167 );
xor \U$6980 ( \7169 , \5023 , \5646 );
buf \U$6981 ( \7170 , \7169 );
buf \U$6982 ( \7171 , \7170 );
xor \U$6983 ( \7172 , \7168 , \7171 );
xor \U$6984 ( \7173 , \7171 , \7150 );
not \U$6985 ( \7174 , \7173 );
and \U$6986 ( \7175 , \7172 , \7174 );
and \U$6987 ( \7176 , \6006 , \7175 );
and \U$6988 ( \7177 , \6018 , \7173 );
nor \U$6989 ( \7178 , \7176 , \7177 );
and \U$6990 ( \7179 , \7171 , \7150 );
not \U$6991 ( \7180 , \7179 );
and \U$6992 ( \7181 , \7168 , \7180 );
xnor \U$6993 ( \7182 , \7178 , \7181 );
and \U$6994 ( \7183 , \7164 , \7182 );
and \U$6995 ( \7184 , \7147 , \7182 );
or \U$6996 ( \7185 , \7165 , \7183 , \7184 );
xor \U$6997 ( \7186 , \4848 , \5650 );
buf \U$6998 ( \7187 , \7186 );
buf \U$6999 ( \7188 , \7187 );
xor \U$7000 ( \7189 , \6821 , \7188 );
xor \U$7001 ( \7190 , \7188 , \7168 );
not \U$7002 ( \7191 , \7190 );
and \U$7003 ( \7192 , \7189 , \7191 );
and \U$7004 ( \7193 , \6029 , \7192 );
and \U$7005 ( \7194 , \6041 , \7190 );
nor \U$7006 ( \7195 , \7193 , \7194 );
and \U$7007 ( \7196 , \7188 , \7168 );
not \U$7008 ( \7197 , \7196 );
and \U$7009 ( \7198 , \6821 , \7197 );
xnor \U$7010 ( \7199 , \7195 , \7198 );
xor \U$7011 ( \7200 , \5747 , \6818 );
xor \U$7012 ( \7201 , \6818 , \6821 );
not \U$7013 ( \7202 , \7201 );
and \U$7014 ( \7203 , \7200 , \7202 );
and \U$7015 ( \7204 , \6048 , \7203 );
and \U$7016 ( \7205 , \6057 , \7201 );
nor \U$7017 ( \7206 , \7204 , \7205 );
xnor \U$7018 ( \7207 , \7206 , \6824 );
and \U$7019 ( \7208 , \7199 , \7207 );
nand \U$7020 ( \7209 , \6065 , \5748 );
xnor \U$7021 ( \7210 , \7209 , \5755 );
and \U$7022 ( \7211 , \7207 , \7210 );
and \U$7023 ( \7212 , \7199 , \7210 );
or \U$7024 ( \7213 , \7208 , \7211 , \7212 );
and \U$7025 ( \7214 , \7185 , \7213 );
and \U$7026 ( \7215 , \6057 , \7203 );
and \U$7027 ( \7216 , \6029 , \7201 );
nor \U$7028 ( \7217 , \7215 , \7216 );
xnor \U$7029 ( \7218 , \7217 , \6824 );
and \U$7030 ( \7219 , \7213 , \7218 );
and \U$7031 ( \7220 , \7185 , \7218 );
or \U$7032 ( \7221 , \7214 , \7219 , \7220 );
and \U$7033 ( \7222 , \7130 , \7221 );
and \U$7034 ( \7223 , \6065 , \5750 );
and \U$7035 ( \7224 , \6048 , \5748 );
nor \U$7036 ( \7225 , \7223 , \7224 );
xnor \U$7037 ( \7226 , \7225 , \5755 );
and \U$7038 ( \7227 , \5998 , \7157 );
and \U$7039 ( \7228 , \5967 , \7155 );
nor \U$7040 ( \7229 , \7227 , \7228 );
xnor \U$7041 ( \7230 , \7229 , \7163 );
and \U$7042 ( \7231 , \6018 , \7175 );
and \U$7043 ( \7232 , \5986 , \7173 );
nor \U$7044 ( \7233 , \7231 , \7232 );
xnor \U$7045 ( \7234 , \7233 , \7181 );
xor \U$7046 ( \7235 , \7230 , \7234 );
and \U$7047 ( \7236 , \6041 , \7192 );
and \U$7048 ( \7237 , \6006 , \7190 );
nor \U$7049 ( \7238 , \7236 , \7237 );
xnor \U$7050 ( \7239 , \7238 , \7198 );
xor \U$7051 ( \7240 , \7235 , \7239 );
and \U$7052 ( \7241 , \7226 , \7240 );
and \U$7053 ( \7242 , \5937 , \7099 );
and \U$7054 ( \7243 , \5906 , \7097 );
nor \U$7055 ( \7244 , \7242 , \7243 );
xnor \U$7056 ( \7245 , \7244 , \7105 );
and \U$7057 ( \7246 , \5957 , \7117 );
and \U$7058 ( \7247 , \5925 , \7115 );
nor \U$7059 ( \7248 , \7246 , \7247 );
xnor \U$7060 ( \7249 , \7248 , \7123 );
xor \U$7061 ( \7250 , \7245 , \7249 );
and \U$7062 ( \7251 , \5979 , \7140 );
and \U$7063 ( \7252 , \5945 , \7138 );
nor \U$7064 ( \7253 , \7251 , \7252 );
xnor \U$7065 ( \7254 , \7253 , \7146 );
xor \U$7066 ( \7255 , \7250 , \7254 );
and \U$7067 ( \7256 , \7240 , \7255 );
and \U$7068 ( \7257 , \7226 , \7255 );
or \U$7069 ( \7258 , \7241 , \7256 , \7257 );
and \U$7070 ( \7259 , \7221 , \7258 );
and \U$7071 ( \7260 , \7130 , \7258 );
or \U$7072 ( \7261 , \7222 , \7259 , \7260 );
and \U$7073 ( \7262 , \5780 , \6991 );
and \U$7074 ( \7263 , \5792 , \6988 );
nor \U$7075 ( \7264 , \7262 , \7263 );
xnor \U$7076 ( \7265 , \7264 , \6985 );
xor \U$7077 ( \7266 , \5775 , \7265 );
and \U$7078 ( \7267 , \5799 , \7006 );
and \U$7079 ( \7268 , \5811 , \7004 );
nor \U$7080 ( \7269 , \7267 , \7268 );
xnor \U$7081 ( \7270 , \7269 , \7012 );
xor \U$7082 ( \7271 , \7266 , \7270 );
and \U$7083 ( \7272 , \5945 , \7140 );
and \U$7084 ( \7273 , \5957 , \7138 );
nor \U$7085 ( \7274 , \7272 , \7273 );
xnor \U$7086 ( \7275 , \7274 , \7146 );
and \U$7087 ( \7276 , \5967 , \7157 );
and \U$7088 ( \7277 , \5979 , \7155 );
nor \U$7089 ( \7278 , \7276 , \7277 );
xnor \U$7090 ( \7279 , \7278 , \7163 );
xor \U$7091 ( \7280 , \7275 , \7279 );
and \U$7092 ( \7281 , \5986 , \7175 );
and \U$7093 ( \7282 , \5998 , \7173 );
nor \U$7094 ( \7283 , \7281 , \7282 );
xnor \U$7095 ( \7284 , \7283 , \7181 );
xor \U$7096 ( \7285 , \7280 , \7284 );
and \U$7097 ( \7286 , \5881 , \7082 );
and \U$7098 ( \7287 , \5893 , \7080 );
nor \U$7099 ( \7288 , \7286 , \7287 );
xnor \U$7100 ( \7289 , \7288 , \7088 );
and \U$7101 ( \7290 , \5906 , \7099 );
and \U$7102 ( \7291 , \5918 , \7097 );
nor \U$7103 ( \7292 , \7290 , \7291 );
xnor \U$7104 ( \7293 , \7292 , \7105 );
xor \U$7105 ( \7294 , \7289 , \7293 );
and \U$7106 ( \7295 , \5925 , \7117 );
and \U$7107 ( \7296 , \5937 , \7115 );
nor \U$7108 ( \7297 , \7295 , \7296 );
xnor \U$7109 ( \7298 , \7297 , \7123 );
xor \U$7110 ( \7299 , \7294 , \7298 );
xor \U$7111 ( \7300 , \7285 , \7299 );
and \U$7112 ( \7301 , \5819 , \7026 );
and \U$7113 ( \7302 , \5831 , \7024 );
nor \U$7114 ( \7303 , \7301 , \7302 );
xnor \U$7115 ( \7304 , \7303 , \7032 );
and \U$7116 ( \7305 , \5842 , \7043 );
and \U$7117 ( \7306 , \5854 , \7041 );
nor \U$7118 ( \7307 , \7305 , \7306 );
xnor \U$7119 ( \7308 , \7307 , \7049 );
xor \U$7120 ( \7309 , \7304 , \7308 );
and \U$7121 ( \7310 , \5861 , \7061 );
and \U$7122 ( \7311 , \5873 , \7059 );
nor \U$7123 ( \7312 , \7310 , \7311 );
xnor \U$7124 ( \7313 , \7312 , \7067 );
xor \U$7125 ( \7314 , \7309 , \7313 );
xor \U$7126 ( \7315 , \7300 , \7314 );
and \U$7127 ( \7316 , \7271 , \7315 );
and \U$7128 ( \7317 , \7230 , \7234 );
and \U$7129 ( \7318 , \7234 , \7239 );
and \U$7130 ( \7319 , \7230 , \7239 );
or \U$7131 ( \7320 , \7317 , \7318 , \7319 );
nand \U$7132 ( \7321 , \6065 , \5766 );
xnor \U$7133 ( \7322 , \7321 , \5775 );
xor \U$7134 ( \7323 , \7320 , \7322 );
and \U$7135 ( \7324 , \6006 , \7192 );
and \U$7136 ( \7325 , \6018 , \7190 );
nor \U$7137 ( \7326 , \7324 , \7325 );
xnor \U$7138 ( \7327 , \7326 , \7198 );
and \U$7139 ( \7328 , \6029 , \7203 );
and \U$7140 ( \7329 , \6041 , \7201 );
nor \U$7141 ( \7330 , \7328 , \7329 );
xnor \U$7142 ( \7331 , \7330 , \6824 );
xor \U$7143 ( \7332 , \7327 , \7331 );
and \U$7144 ( \7333 , \6048 , \5750 );
and \U$7145 ( \7334 , \6057 , \5748 );
nor \U$7146 ( \7335 , \7333 , \7334 );
xnor \U$7147 ( \7336 , \7335 , \5755 );
xor \U$7148 ( \7337 , \7332 , \7336 );
xor \U$7149 ( \7338 , \7323 , \7337 );
and \U$7150 ( \7339 , \7315 , \7338 );
and \U$7151 ( \7340 , \7271 , \7338 );
or \U$7152 ( \7341 , \7316 , \7339 , \7340 );
and \U$7153 ( \7342 , \7261 , \7341 );
and \U$7154 ( \7343 , \5775 , \7265 );
and \U$7155 ( \7344 , \7265 , \7270 );
and \U$7156 ( \7345 , \5775 , \7270 );
or \U$7157 ( \7346 , \7343 , \7344 , \7345 );
and \U$7158 ( \7347 , \7304 , \7308 );
and \U$7159 ( \7348 , \7308 , \7313 );
and \U$7160 ( \7349 , \7304 , \7313 );
or \U$7161 ( \7350 , \7347 , \7348 , \7349 );
xor \U$7162 ( \7351 , \7346 , \7350 );
and \U$7163 ( \7352 , \7289 , \7293 );
and \U$7164 ( \7353 , \7293 , \7298 );
and \U$7165 ( \7354 , \7289 , \7298 );
or \U$7166 ( \7355 , \7352 , \7353 , \7354 );
xor \U$7167 ( \7356 , \7351 , \7355 );
and \U$7168 ( \7357 , \7341 , \7356 );
and \U$7169 ( \7358 , \7261 , \7356 );
or \U$7170 ( \7359 , \7342 , \7357 , \7358 );
and \U$7171 ( \7360 , \5792 , \6991 );
and \U$7172 ( \7361 , \5758 , \6988 );
nor \U$7173 ( \7362 , \7360 , \7361 );
xnor \U$7174 ( \7363 , \7362 , \6985 );
and \U$7175 ( \7364 , \5811 , \7006 );
and \U$7176 ( \7365 , \5780 , \7004 );
nor \U$7177 ( \7366 , \7364 , \7365 );
xnor \U$7178 ( \7367 , \7366 , \7012 );
xor \U$7179 ( \7368 , \7363 , \7367 );
and \U$7180 ( \7369 , \5831 , \7026 );
and \U$7181 ( \7370 , \5799 , \7024 );
nor \U$7182 ( \7371 , \7369 , \7370 );
xnor \U$7183 ( \7372 , \7371 , \7032 );
xor \U$7184 ( \7373 , \7368 , \7372 );
and \U$7185 ( \7374 , \5979 , \7157 );
and \U$7186 ( \7375 , \5945 , \7155 );
nor \U$7187 ( \7376 , \7374 , \7375 );
xnor \U$7188 ( \7377 , \7376 , \7163 );
and \U$7189 ( \7378 , \5998 , \7175 );
and \U$7190 ( \7379 , \5967 , \7173 );
nor \U$7191 ( \7380 , \7378 , \7379 );
xnor \U$7192 ( \7381 , \7380 , \7181 );
xor \U$7193 ( \7382 , \7377 , \7381 );
and \U$7194 ( \7383 , \6018 , \7192 );
and \U$7195 ( \7384 , \5986 , \7190 );
nor \U$7196 ( \7385 , \7383 , \7384 );
xnor \U$7197 ( \7386 , \7385 , \7198 );
xor \U$7198 ( \7387 , \7382 , \7386 );
and \U$7199 ( \7388 , \5918 , \7099 );
and \U$7200 ( \7389 , \5881 , \7097 );
nor \U$7201 ( \7390 , \7388 , \7389 );
xnor \U$7202 ( \7391 , \7390 , \7105 );
and \U$7203 ( \7392 , \5937 , \7117 );
and \U$7204 ( \7393 , \5906 , \7115 );
nor \U$7205 ( \7394 , \7392 , \7393 );
xnor \U$7206 ( \7395 , \7394 , \7123 );
xor \U$7207 ( \7396 , \7391 , \7395 );
and \U$7208 ( \7397 , \5957 , \7140 );
and \U$7209 ( \7398 , \5925 , \7138 );
nor \U$7210 ( \7399 , \7397 , \7398 );
xnor \U$7211 ( \7400 , \7399 , \7146 );
xor \U$7212 ( \7401 , \7396 , \7400 );
xor \U$7213 ( \7402 , \7387 , \7401 );
and \U$7214 ( \7403 , \5854 , \7043 );
and \U$7215 ( \7404 , \5819 , \7041 );
nor \U$7216 ( \7405 , \7403 , \7404 );
xnor \U$7217 ( \7406 , \7405 , \7049 );
and \U$7218 ( \7407 , \5873 , \7061 );
and \U$7219 ( \7408 , \5842 , \7059 );
nor \U$7220 ( \7409 , \7407 , \7408 );
xnor \U$7221 ( \7410 , \7409 , \7067 );
xor \U$7222 ( \7411 , \7406 , \7410 );
and \U$7223 ( \7412 , \5893 , \7082 );
and \U$7224 ( \7413 , \5861 , \7080 );
nor \U$7225 ( \7414 , \7412 , \7413 );
xnor \U$7226 ( \7415 , \7414 , \7088 );
xor \U$7227 ( \7416 , \7411 , \7415 );
xor \U$7228 ( \7417 , \7402 , \7416 );
xor \U$7229 ( \7418 , \7373 , \7417 );
and \U$7230 ( \7419 , \7275 , \7279 );
and \U$7231 ( \7420 , \7279 , \7284 );
and \U$7232 ( \7421 , \7275 , \7284 );
or \U$7233 ( \7422 , \7419 , \7420 , \7421 );
and \U$7234 ( \7423 , \7327 , \7331 );
and \U$7235 ( \7424 , \7331 , \7336 );
and \U$7236 ( \7425 , \7327 , \7336 );
or \U$7237 ( \7426 , \7423 , \7424 , \7425 );
xor \U$7238 ( \7427 , \7422 , \7426 );
and \U$7239 ( \7428 , \6041 , \7203 );
and \U$7240 ( \7429 , \6006 , \7201 );
nor \U$7241 ( \7430 , \7428 , \7429 );
xnor \U$7242 ( \7431 , \7430 , \6824 );
and \U$7243 ( \7432 , \6057 , \5750 );
and \U$7244 ( \7433 , \6029 , \5748 );
nor \U$7245 ( \7434 , \7432 , \7433 );
xnor \U$7246 ( \7435 , \7434 , \5755 );
xor \U$7247 ( \7436 , \7431 , \7435 );
and \U$7248 ( \7437 , \6065 , \5768 );
and \U$7249 ( \7438 , \6048 , \5766 );
nor \U$7250 ( \7439 , \7437 , \7438 );
xnor \U$7251 ( \7440 , \7439 , \5775 );
xor \U$7252 ( \7441 , \7436 , \7440 );
xor \U$7253 ( \7442 , \7427 , \7441 );
xor \U$7254 ( \7443 , \7418 , \7442 );
and \U$7255 ( \7444 , \5811 , \6991 );
and \U$7256 ( \7445 , \5780 , \6988 );
nor \U$7257 ( \7446 , \7444 , \7445 );
xnor \U$7258 ( \7447 , \7446 , \6985 );
and \U$7259 ( \7448 , \5831 , \7006 );
and \U$7260 ( \7449 , \5799 , \7004 );
nor \U$7261 ( \7450 , \7448 , \7449 );
xnor \U$7262 ( \7451 , \7450 , \7012 );
and \U$7263 ( \7452 , \7447 , \7451 );
and \U$7264 ( \7453 , \5854 , \7026 );
and \U$7265 ( \7454 , \5819 , \7024 );
nor \U$7266 ( \7455 , \7453 , \7454 );
xnor \U$7267 ( \7456 , \7455 , \7032 );
and \U$7268 ( \7457 , \7451 , \7456 );
and \U$7269 ( \7458 , \7447 , \7456 );
or \U$7270 ( \7459 , \7452 , \7457 , \7458 );
and \U$7271 ( \7460 , \5873 , \7043 );
and \U$7272 ( \7461 , \5842 , \7041 );
nor \U$7273 ( \7462 , \7460 , \7461 );
xnor \U$7274 ( \7463 , \7462 , \7049 );
and \U$7275 ( \7464 , \5893 , \7061 );
and \U$7276 ( \7465 , \5861 , \7059 );
nor \U$7277 ( \7466 , \7464 , \7465 );
xnor \U$7278 ( \7467 , \7466 , \7067 );
and \U$7279 ( \7468 , \7463 , \7467 );
and \U$7280 ( \7469 , \5918 , \7082 );
and \U$7281 ( \7470 , \5881 , \7080 );
nor \U$7282 ( \7471 , \7469 , \7470 );
xnor \U$7283 ( \7472 , \7471 , \7088 );
and \U$7284 ( \7473 , \7467 , \7472 );
and \U$7285 ( \7474 , \7463 , \7472 );
or \U$7286 ( \7475 , \7468 , \7473 , \7474 );
and \U$7287 ( \7476 , \7459 , \7475 );
and \U$7288 ( \7477 , \7245 , \7249 );
and \U$7289 ( \7478 , \7249 , \7254 );
and \U$7290 ( \7479 , \7245 , \7254 );
or \U$7291 ( \7480 , \7477 , \7478 , \7479 );
and \U$7292 ( \7481 , \7475 , \7480 );
and \U$7293 ( \7482 , \7459 , \7480 );
or \U$7294 ( \7483 , \7476 , \7481 , \7482 );
and \U$7295 ( \7484 , \7320 , \7322 );
and \U$7296 ( \7485 , \7322 , \7337 );
and \U$7297 ( \7486 , \7320 , \7337 );
or \U$7298 ( \7487 , \7484 , \7485 , \7486 );
xor \U$7299 ( \7488 , \7483 , \7487 );
and \U$7300 ( \7489 , \7285 , \7299 );
and \U$7301 ( \7490 , \7299 , \7314 );
and \U$7302 ( \7491 , \7285 , \7314 );
or \U$7303 ( \7492 , \7489 , \7490 , \7491 );
xor \U$7304 ( \7493 , \7488 , \7492 );
and \U$7305 ( \7494 , \7443 , \7493 );
and \U$7306 ( \7495 , \7359 , \7494 );
and \U$7307 ( \7496 , \5861 , \7082 );
and \U$7308 ( \7497 , \5873 , \7080 );
nor \U$7309 ( \7498 , \7496 , \7497 );
xnor \U$7310 ( \7499 , \7498 , \7088 );
and \U$7311 ( \7500 , \5881 , \7099 );
and \U$7312 ( \7501 , \5893 , \7097 );
nor \U$7313 ( \7502 , \7500 , \7501 );
xnor \U$7314 ( \7503 , \7502 , \7105 );
xor \U$7315 ( \7504 , \7499 , \7503 );
and \U$7316 ( \7505 , \5906 , \7117 );
and \U$7317 ( \7506 , \5918 , \7115 );
nor \U$7318 ( \7507 , \7505 , \7506 );
xnor \U$7319 ( \7508 , \7507 , \7123 );
xor \U$7320 ( \7509 , \7504 , \7508 );
and \U$7321 ( \7510 , \5799 , \7026 );
and \U$7322 ( \7511 , \5811 , \7024 );
nor \U$7323 ( \7512 , \7510 , \7511 );
xnor \U$7324 ( \7513 , \7512 , \7032 );
and \U$7325 ( \7514 , \5819 , \7043 );
and \U$7326 ( \7515 , \5831 , \7041 );
nor \U$7327 ( \7516 , \7514 , \7515 );
xnor \U$7328 ( \7517 , \7516 , \7049 );
xor \U$7329 ( \7518 , \7513 , \7517 );
and \U$7330 ( \7519 , \5842 , \7061 );
and \U$7331 ( \7520 , \5854 , \7059 );
nor \U$7332 ( \7521 , \7519 , \7520 );
xnor \U$7333 ( \7522 , \7521 , \7067 );
xor \U$7334 ( \7523 , \7518 , \7522 );
xor \U$7335 ( \7524 , \7509 , \7523 );
and \U$7336 ( \7525 , \5758 , \6991 );
and \U$7337 ( \7526 , \5770 , \6988 );
nor \U$7338 ( \7527 , \7525 , \7526 );
xnor \U$7339 ( \7528 , \7527 , \6985 );
xor \U$7340 ( \7529 , \5797 , \7528 );
and \U$7341 ( \7530 , \5780 , \7006 );
and \U$7342 ( \7531 , \5792 , \7004 );
nor \U$7343 ( \7532 , \7530 , \7531 );
xnor \U$7344 ( \7533 , \7532 , \7012 );
xor \U$7345 ( \7534 , \7529 , \7533 );
xor \U$7346 ( \7535 , \7524 , \7534 );
nand \U$7347 ( \7536 , \6065 , \5788 );
xnor \U$7348 ( \7537 , \7536 , \5797 );
and \U$7349 ( \7538 , \5986 , \7192 );
and \U$7350 ( \7539 , \5998 , \7190 );
nor \U$7351 ( \7540 , \7538 , \7539 );
xnor \U$7352 ( \7541 , \7540 , \7198 );
and \U$7353 ( \7542 , \6006 , \7203 );
and \U$7354 ( \7543 , \6018 , \7201 );
nor \U$7355 ( \7544 , \7542 , \7543 );
xnor \U$7356 ( \7545 , \7544 , \6824 );
xor \U$7357 ( \7546 , \7541 , \7545 );
and \U$7358 ( \7547 , \6029 , \5750 );
and \U$7359 ( \7548 , \6041 , \5748 );
nor \U$7360 ( \7549 , \7547 , \7548 );
xnor \U$7361 ( \7550 , \7549 , \5755 );
xor \U$7362 ( \7551 , \7546 , \7550 );
xor \U$7363 ( \7552 , \7537 , \7551 );
and \U$7364 ( \7553 , \5925 , \7140 );
and \U$7365 ( \7554 , \5937 , \7138 );
nor \U$7366 ( \7555 , \7553 , \7554 );
xnor \U$7367 ( \7556 , \7555 , \7146 );
and \U$7368 ( \7557 , \5945 , \7157 );
and \U$7369 ( \7558 , \5957 , \7155 );
nor \U$7370 ( \7559 , \7557 , \7558 );
xnor \U$7371 ( \7560 , \7559 , \7163 );
xor \U$7372 ( \7561 , \7556 , \7560 );
and \U$7373 ( \7562 , \5967 , \7175 );
and \U$7374 ( \7563 , \5979 , \7173 );
nor \U$7375 ( \7564 , \7562 , \7563 );
xnor \U$7376 ( \7565 , \7564 , \7181 );
xor \U$7377 ( \7566 , \7561 , \7565 );
xor \U$7378 ( \7567 , \7552 , \7566 );
xor \U$7379 ( \7568 , \7535 , \7567 );
and \U$7380 ( \7569 , \7377 , \7381 );
and \U$7381 ( \7570 , \7381 , \7386 );
and \U$7382 ( \7571 , \7377 , \7386 );
or \U$7383 ( \7572 , \7569 , \7570 , \7571 );
and \U$7384 ( \7573 , \7431 , \7435 );
and \U$7385 ( \7574 , \7435 , \7440 );
and \U$7386 ( \7575 , \7431 , \7440 );
or \U$7387 ( \7576 , \7573 , \7574 , \7575 );
xor \U$7388 ( \7577 , \7572 , \7576 );
and \U$7389 ( \7578 , \6048 , \5768 );
and \U$7390 ( \7579 , \6057 , \5766 );
nor \U$7391 ( \7580 , \7578 , \7579 );
xnor \U$7392 ( \7581 , \7580 , \5775 );
xor \U$7393 ( \7582 , \7577 , \7581 );
xor \U$7394 ( \7583 , \7568 , \7582 );
and \U$7395 ( \7584 , \7494 , \7583 );
and \U$7396 ( \7585 , \7359 , \7583 );
or \U$7397 ( \7586 , \7495 , \7584 , \7585 );
and \U$7398 ( \7587 , \7346 , \7350 );
and \U$7399 ( \7588 , \7350 , \7355 );
and \U$7400 ( \7589 , \7346 , \7355 );
or \U$7401 ( \7590 , \7587 , \7588 , \7589 );
and \U$7402 ( \7591 , \7422 , \7426 );
and \U$7403 ( \7592 , \7426 , \7441 );
and \U$7404 ( \7593 , \7422 , \7441 );
or \U$7405 ( \7594 , \7591 , \7592 , \7593 );
xor \U$7406 ( \7595 , \7590 , \7594 );
and \U$7407 ( \7596 , \7387 , \7401 );
and \U$7408 ( \7597 , \7401 , \7416 );
and \U$7409 ( \7598 , \7387 , \7416 );
or \U$7410 ( \7599 , \7596 , \7597 , \7598 );
xor \U$7411 ( \7600 , \7595 , \7599 );
and \U$7412 ( \7601 , \7483 , \7487 );
and \U$7413 ( \7602 , \7487 , \7492 );
and \U$7414 ( \7603 , \7483 , \7492 );
or \U$7415 ( \7604 , \7601 , \7602 , \7603 );
and \U$7416 ( \7605 , \7373 , \7417 );
and \U$7417 ( \7606 , \7417 , \7442 );
and \U$7418 ( \7607 , \7373 , \7442 );
or \U$7419 ( \7608 , \7605 , \7606 , \7607 );
xor \U$7420 ( \7609 , \7604 , \7608 );
and \U$7421 ( \7610 , \7363 , \7367 );
and \U$7422 ( \7611 , \7367 , \7372 );
and \U$7423 ( \7612 , \7363 , \7372 );
or \U$7424 ( \7613 , \7610 , \7611 , \7612 );
and \U$7425 ( \7614 , \7406 , \7410 );
and \U$7426 ( \7615 , \7410 , \7415 );
and \U$7427 ( \7616 , \7406 , \7415 );
or \U$7428 ( \7617 , \7614 , \7615 , \7616 );
xor \U$7429 ( \7618 , \7613 , \7617 );
and \U$7430 ( \7619 , \7391 , \7395 );
and \U$7431 ( \7620 , \7395 , \7400 );
and \U$7432 ( \7621 , \7391 , \7400 );
or \U$7433 ( \7622 , \7619 , \7620 , \7621 );
xor \U$7434 ( \7623 , \7618 , \7622 );
xor \U$7435 ( \7624 , \7609 , \7623 );
and \U$7436 ( \7625 , \7600 , \7624 );
xor \U$7437 ( \7626 , \7586 , \7625 );
and \U$7438 ( \7627 , \7604 , \7608 );
and \U$7439 ( \7628 , \7608 , \7623 );
and \U$7440 ( \7629 , \7604 , \7623 );
or \U$7441 ( \7630 , \7627 , \7628 , \7629 );
and \U$7442 ( \7631 , \7509 , \7523 );
and \U$7443 ( \7632 , \7523 , \7534 );
and \U$7444 ( \7633 , \7509 , \7534 );
or \U$7445 ( \7634 , \7631 , \7632 , \7633 );
and \U$7446 ( \7635 , \5831 , \7043 );
and \U$7447 ( \7636 , \5799 , \7041 );
nor \U$7448 ( \7637 , \7635 , \7636 );
xnor \U$7449 ( \7638 , \7637 , \7049 );
and \U$7450 ( \7639 , \5854 , \7061 );
and \U$7451 ( \7640 , \5819 , \7059 );
nor \U$7452 ( \7641 , \7639 , \7640 );
xnor \U$7453 ( \7642 , \7641 , \7067 );
xor \U$7454 ( \7643 , \7638 , \7642 );
and \U$7455 ( \7644 , \5873 , \7082 );
and \U$7456 ( \7645 , \5842 , \7080 );
nor \U$7457 ( \7646 , \7644 , \7645 );
xnor \U$7458 ( \7647 , \7646 , \7088 );
xor \U$7459 ( \7648 , \7643 , \7647 );
xor \U$7460 ( \7649 , \7634 , \7648 );
and \U$7461 ( \7650 , \5770 , \6991 );
and \U$7462 ( \7651 , \5737 , \6988 );
nor \U$7463 ( \7652 , \7650 , \7651 );
xnor \U$7464 ( \7653 , \7652 , \6985 );
and \U$7465 ( \7654 , \5792 , \7006 );
and \U$7466 ( \7655 , \5758 , \7004 );
nor \U$7467 ( \7656 , \7654 , \7655 );
xnor \U$7468 ( \7657 , \7656 , \7012 );
xor \U$7469 ( \7658 , \7653 , \7657 );
and \U$7470 ( \7659 , \5811 , \7026 );
and \U$7471 ( \7660 , \5780 , \7024 );
nor \U$7472 ( \7661 , \7659 , \7660 );
xnor \U$7473 ( \7662 , \7661 , \7032 );
xor \U$7474 ( \7663 , \7658 , \7662 );
xor \U$7475 ( \7664 , \7649 , \7663 );
and \U$7476 ( \7665 , \7613 , \7617 );
and \U$7477 ( \7666 , \7617 , \7622 );
and \U$7478 ( \7667 , \7613 , \7622 );
or \U$7479 ( \7668 , \7665 , \7666 , \7667 );
and \U$7480 ( \7669 , \7572 , \7576 );
and \U$7481 ( \7670 , \7576 , \7581 );
and \U$7482 ( \7671 , \7572 , \7581 );
or \U$7483 ( \7672 , \7669 , \7670 , \7671 );
xor \U$7484 ( \7673 , \7668 , \7672 );
and \U$7485 ( \7674 , \7537 , \7551 );
and \U$7486 ( \7675 , \7551 , \7566 );
and \U$7487 ( \7676 , \7537 , \7566 );
or \U$7488 ( \7677 , \7674 , \7675 , \7676 );
xor \U$7489 ( \7678 , \7673 , \7677 );
xor \U$7490 ( \7679 , \7664 , \7678 );
xor \U$7491 ( \7680 , \7630 , \7679 );
and \U$7492 ( \7681 , \7590 , \7594 );
and \U$7493 ( \7682 , \7594 , \7599 );
and \U$7494 ( \7683 , \7590 , \7599 );
or \U$7495 ( \7684 , \7681 , \7682 , \7683 );
and \U$7496 ( \7685 , \7535 , \7567 );
and \U$7497 ( \7686 , \7567 , \7582 );
and \U$7498 ( \7687 , \7535 , \7582 );
or \U$7499 ( \7688 , \7685 , \7686 , \7687 );
xor \U$7500 ( \7689 , \7684 , \7688 );
and \U$7501 ( \7690 , \6018 , \7203 );
and \U$7502 ( \7691 , \5986 , \7201 );
nor \U$7503 ( \7692 , \7690 , \7691 );
xnor \U$7504 ( \7693 , \7692 , \6824 );
and \U$7505 ( \7694 , \6041 , \5750 );
and \U$7506 ( \7695 , \6006 , \5748 );
nor \U$7507 ( \7696 , \7694 , \7695 );
xnor \U$7508 ( \7697 , \7696 , \5755 );
xor \U$7509 ( \7698 , \7693 , \7697 );
and \U$7510 ( \7699 , \6057 , \5768 );
and \U$7511 ( \7700 , \6029 , \5766 );
nor \U$7512 ( \7701 , \7699 , \7700 );
xnor \U$7513 ( \7702 , \7701 , \5775 );
xor \U$7514 ( \7703 , \7698 , \7702 );
and \U$7515 ( \7704 , \5957 , \7157 );
and \U$7516 ( \7705 , \5925 , \7155 );
nor \U$7517 ( \7706 , \7704 , \7705 );
xnor \U$7518 ( \7707 , \7706 , \7163 );
and \U$7519 ( \7708 , \5979 , \7175 );
and \U$7520 ( \7709 , \5945 , \7173 );
nor \U$7521 ( \7710 , \7708 , \7709 );
xnor \U$7522 ( \7711 , \7710 , \7181 );
xor \U$7523 ( \7712 , \7707 , \7711 );
and \U$7524 ( \7713 , \5998 , \7192 );
and \U$7525 ( \7714 , \5967 , \7190 );
nor \U$7526 ( \7715 , \7713 , \7714 );
xnor \U$7527 ( \7716 , \7715 , \7198 );
xor \U$7528 ( \7717 , \7712 , \7716 );
xor \U$7529 ( \7718 , \7703 , \7717 );
and \U$7530 ( \7719 , \5893 , \7099 );
and \U$7531 ( \7720 , \5861 , \7097 );
nor \U$7532 ( \7721 , \7719 , \7720 );
xnor \U$7533 ( \7722 , \7721 , \7105 );
and \U$7534 ( \7723 , \5918 , \7117 );
and \U$7535 ( \7724 , \5881 , \7115 );
nor \U$7536 ( \7725 , \7723 , \7724 );
xnor \U$7537 ( \7726 , \7725 , \7123 );
xor \U$7538 ( \7727 , \7722 , \7726 );
and \U$7539 ( \7728 , \5937 , \7140 );
and \U$7540 ( \7729 , \5906 , \7138 );
nor \U$7541 ( \7730 , \7728 , \7729 );
xnor \U$7542 ( \7731 , \7730 , \7146 );
xor \U$7543 ( \7732 , \7727 , \7731 );
xor \U$7544 ( \7733 , \7718 , \7732 );
and \U$7545 ( \7734 , \7556 , \7560 );
and \U$7546 ( \7735 , \7560 , \7565 );
and \U$7547 ( \7736 , \7556 , \7565 );
or \U$7548 ( \7737 , \7734 , \7735 , \7736 );
and \U$7549 ( \7738 , \7541 , \7545 );
and \U$7550 ( \7739 , \7545 , \7550 );
and \U$7551 ( \7740 , \7541 , \7550 );
or \U$7552 ( \7741 , \7738 , \7739 , \7740 );
xor \U$7553 ( \7742 , \7737 , \7741 );
and \U$7554 ( \7743 , \6065 , \5790 );
and \U$7555 ( \7744 , \6048 , \5788 );
nor \U$7556 ( \7745 , \7743 , \7744 );
xnor \U$7557 ( \7746 , \7745 , \5797 );
xor \U$7558 ( \7747 , \7742 , \7746 );
xor \U$7559 ( \7748 , \7733 , \7747 );
and \U$7560 ( \7749 , \5797 , \7528 );
and \U$7561 ( \7750 , \7528 , \7533 );
and \U$7562 ( \7751 , \5797 , \7533 );
or \U$7563 ( \7752 , \7749 , \7750 , \7751 );
and \U$7564 ( \7753 , \7513 , \7517 );
and \U$7565 ( \7754 , \7517 , \7522 );
and \U$7566 ( \7755 , \7513 , \7522 );
or \U$7567 ( \7756 , \7753 , \7754 , \7755 );
xor \U$7568 ( \7757 , \7752 , \7756 );
and \U$7569 ( \7758 , \7499 , \7503 );
and \U$7570 ( \7759 , \7503 , \7508 );
and \U$7571 ( \7760 , \7499 , \7508 );
or \U$7572 ( \7761 , \7758 , \7759 , \7760 );
xor \U$7573 ( \7762 , \7757 , \7761 );
xor \U$7574 ( \7763 , \7748 , \7762 );
xor \U$7575 ( \7764 , \7689 , \7763 );
xor \U$7576 ( \7765 , \7680 , \7764 );
xor \U$7577 ( \7766 , \7626 , \7765 );
and \U$7578 ( \7767 , \5831 , \6991 );
and \U$7579 ( \7768 , \5799 , \6988 );
nor \U$7580 ( \7769 , \7767 , \7768 );
xnor \U$7581 ( \7770 , \7769 , \6985 );
and \U$7582 ( \7771 , \5854 , \7006 );
and \U$7583 ( \7772 , \5819 , \7004 );
nor \U$7584 ( \7773 , \7771 , \7772 );
xnor \U$7585 ( \7774 , \7773 , \7012 );
and \U$7586 ( \7775 , \7770 , \7774 );
and \U$7587 ( \7776 , \5873 , \7026 );
and \U$7588 ( \7777 , \5842 , \7024 );
nor \U$7589 ( \7778 , \7776 , \7777 );
xnor \U$7590 ( \7779 , \7778 , \7032 );
and \U$7591 ( \7780 , \7774 , \7779 );
and \U$7592 ( \7781 , \7770 , \7779 );
or \U$7593 ( \7782 , \7775 , \7780 , \7781 );
and \U$7594 ( \7783 , \5893 , \7043 );
and \U$7595 ( \7784 , \5861 , \7041 );
nor \U$7596 ( \7785 , \7783 , \7784 );
xnor \U$7597 ( \7786 , \7785 , \7049 );
and \U$7598 ( \7787 , \5918 , \7061 );
and \U$7599 ( \7788 , \5881 , \7059 );
nor \U$7600 ( \7789 , \7787 , \7788 );
xnor \U$7601 ( \7790 , \7789 , \7067 );
and \U$7602 ( \7791 , \7786 , \7790 );
and \U$7603 ( \7792 , \5937 , \7082 );
and \U$7604 ( \7793 , \5906 , \7080 );
nor \U$7605 ( \7794 , \7792 , \7793 );
xnor \U$7606 ( \7795 , \7794 , \7088 );
and \U$7607 ( \7796 , \7790 , \7795 );
and \U$7608 ( \7797 , \7786 , \7795 );
or \U$7609 ( \7798 , \7791 , \7796 , \7797 );
and \U$7610 ( \7799 , \7782 , \7798 );
and \U$7611 ( \7800 , \5957 , \7099 );
and \U$7612 ( \7801 , \5925 , \7097 );
nor \U$7613 ( \7802 , \7800 , \7801 );
xnor \U$7614 ( \7803 , \7802 , \7105 );
and \U$7615 ( \7804 , \5979 , \7117 );
and \U$7616 ( \7805 , \5945 , \7115 );
nor \U$7617 ( \7806 , \7804 , \7805 );
xnor \U$7618 ( \7807 , \7806 , \7123 );
and \U$7619 ( \7808 , \7803 , \7807 );
and \U$7620 ( \7809 , \5998 , \7140 );
and \U$7621 ( \7810 , \5967 , \7138 );
nor \U$7622 ( \7811 , \7809 , \7810 );
xnor \U$7623 ( \7812 , \7811 , \7146 );
and \U$7624 ( \7813 , \7807 , \7812 );
and \U$7625 ( \7814 , \7803 , \7812 );
or \U$7626 ( \7815 , \7808 , \7813 , \7814 );
and \U$7627 ( \7816 , \7798 , \7815 );
and \U$7628 ( \7817 , \7782 , \7815 );
or \U$7629 ( \7818 , \7799 , \7816 , \7817 );
and \U$7630 ( \7819 , \6018 , \7157 );
and \U$7631 ( \7820 , \5986 , \7155 );
nor \U$7632 ( \7821 , \7819 , \7820 );
xnor \U$7633 ( \7822 , \7821 , \7163 );
and \U$7634 ( \7823 , \6041 , \7175 );
and \U$7635 ( \7824 , \6006 , \7173 );
nor \U$7636 ( \7825 , \7823 , \7824 );
xnor \U$7637 ( \7826 , \7825 , \7181 );
and \U$7638 ( \7827 , \7822 , \7826 );
and \U$7639 ( \7828 , \6057 , \7192 );
and \U$7640 ( \7829 , \6029 , \7190 );
nor \U$7641 ( \7830 , \7828 , \7829 );
xnor \U$7642 ( \7831 , \7830 , \7198 );
and \U$7643 ( \7832 , \7826 , \7831 );
and \U$7644 ( \7833 , \7822 , \7831 );
or \U$7645 ( \7834 , \7827 , \7832 , \7833 );
xor \U$7646 ( \7835 , \7199 , \7207 );
xor \U$7647 ( \7836 , \7835 , \7210 );
and \U$7648 ( \7837 , \7834 , \7836 );
xor \U$7649 ( \7838 , \7147 , \7164 );
xor \U$7650 ( \7839 , \7838 , \7182 );
and \U$7651 ( \7840 , \7836 , \7839 );
and \U$7652 ( \7841 , \7834 , \7839 );
or \U$7653 ( \7842 , \7837 , \7840 , \7841 );
and \U$7654 ( \7843 , \7818 , \7842 );
xor \U$7655 ( \7844 , \7089 , \7106 );
xor \U$7656 ( \7845 , \7844 , \7124 );
xor \U$7657 ( \7846 , \7033 , \7050 );
xor \U$7658 ( \7847 , \7846 , \7068 );
and \U$7659 ( \7848 , \7845 , \7847 );
xor \U$7660 ( \7849 , \5755 , \6995 );
xor \U$7661 ( \7850 , \7849 , \7013 );
and \U$7662 ( \7851 , \7847 , \7850 );
and \U$7663 ( \7852 , \7845 , \7850 );
or \U$7664 ( \7853 , \7848 , \7851 , \7852 );
and \U$7665 ( \7854 , \7842 , \7853 );
and \U$7666 ( \7855 , \7818 , \7853 );
or \U$7667 ( \7856 , \7843 , \7854 , \7855 );
xor \U$7668 ( \7857 , \7463 , \7467 );
xor \U$7669 ( \7858 , \7857 , \7472 );
xor \U$7670 ( \7859 , \7447 , \7451 );
xor \U$7671 ( \7860 , \7859 , \7456 );
and \U$7672 ( \7861 , \7858 , \7860 );
xor \U$7673 ( \7862 , \7226 , \7240 );
xor \U$7674 ( \7863 , \7862 , \7255 );
and \U$7675 ( \7864 , \7860 , \7863 );
and \U$7676 ( \7865 , \7858 , \7863 );
or \U$7677 ( \7866 , \7861 , \7864 , \7865 );
and \U$7678 ( \7867 , \7856 , \7866 );
xor \U$7679 ( \7868 , \7459 , \7475 );
xor \U$7680 ( \7869 , \7868 , \7480 );
and \U$7681 ( \7870 , \7866 , \7869 );
and \U$7682 ( \7871 , \7856 , \7869 );
or \U$7683 ( \7872 , \7867 , \7870 , \7871 );
xor \U$7684 ( \7873 , \7443 , \7493 );
and \U$7685 ( \7874 , \7872 , \7873 );
xor \U$7686 ( \7875 , \7261 , \7341 );
xor \U$7687 ( \7876 , \7875 , \7356 );
and \U$7688 ( \7877 , \7873 , \7876 );
and \U$7689 ( \7878 , \7872 , \7876 );
or \U$7690 ( \7879 , \7874 , \7877 , \7878 );
xor \U$7691 ( \7880 , \7600 , \7624 );
and \U$7692 ( \7881 , \7879 , \7880 );
xor \U$7693 ( \7882 , \7359 , \7494 );
xor \U$7694 ( \7883 , \7882 , \7583 );
and \U$7695 ( \7884 , \7880 , \7883 );
and \U$7696 ( \7885 , \7879 , \7883 );
or \U$7697 ( \7886 , \7881 , \7884 , \7885 );
nor \U$7698 ( \7887 , \7766 , \7886 );
and \U$7699 ( \7888 , \7630 , \7679 );
and \U$7700 ( \7889 , \7679 , \7764 );
and \U$7701 ( \7890 , \7630 , \7764 );
or \U$7702 ( \7891 , \7888 , \7889 , \7890 );
and \U$7703 ( \7892 , \7668 , \7672 );
and \U$7704 ( \7893 , \7672 , \7677 );
and \U$7705 ( \7894 , \7668 , \7677 );
or \U$7706 ( \7895 , \7892 , \7893 , \7894 );
and \U$7707 ( \7896 , \7634 , \7648 );
and \U$7708 ( \7897 , \7648 , \7663 );
and \U$7709 ( \7898 , \7634 , \7663 );
or \U$7710 ( \7899 , \7896 , \7897 , \7898 );
xor \U$7711 ( \7900 , \7895 , \7899 );
and \U$7712 ( \7901 , \7733 , \7747 );
and \U$7713 ( \7902 , \7747 , \7762 );
and \U$7714 ( \7903 , \7733 , \7762 );
or \U$7715 ( \7904 , \7901 , \7902 , \7903 );
xor \U$7716 ( \7905 , \7900 , \7904 );
xor \U$7717 ( \7906 , \7891 , \7905 );
and \U$7718 ( \7907 , \7684 , \7688 );
and \U$7719 ( \7908 , \7688 , \7763 );
and \U$7720 ( \7909 , \7684 , \7763 );
or \U$7721 ( \7910 , \7907 , \7908 , \7909 );
and \U$7722 ( \7911 , \7664 , \7678 );
xor \U$7723 ( \7912 , \7910 , \7911 );
and \U$7724 ( \7913 , \7707 , \7711 );
and \U$7725 ( \7914 , \7711 , \7716 );
and \U$7726 ( \7915 , \7707 , \7716 );
or \U$7727 ( \7916 , \7913 , \7914 , \7915 );
and \U$7728 ( \7917 , \7693 , \7697 );
and \U$7729 ( \7918 , \7697 , \7702 );
and \U$7730 ( \7919 , \7693 , \7702 );
or \U$7731 ( \7920 , \7917 , \7918 , \7919 );
xor \U$7732 ( \7921 , \7916 , \7920 );
and \U$7733 ( \7922 , \6029 , \5768 );
and \U$7734 ( \7923 , \6041 , \5766 );
nor \U$7735 ( \7924 , \7922 , \7923 );
xnor \U$7736 ( \7925 , \7924 , \5775 );
and \U$7737 ( \7926 , \6048 , \5790 );
and \U$7738 ( \7927 , \6057 , \5788 );
nor \U$7739 ( \7928 , \7926 , \7927 );
xnor \U$7740 ( \7929 , \7928 , \5797 );
xor \U$7741 ( \7930 , \7925 , \7929 );
nand \U$7742 ( \7931 , \6065 , \5807 );
xnor \U$7743 ( \7932 , \7931 , \5816 );
xor \U$7744 ( \7933 , \7930 , \7932 );
xor \U$7745 ( \7934 , \7921 , \7933 );
and \U$7746 ( \7935 , \7653 , \7657 );
and \U$7747 ( \7936 , \7657 , \7662 );
and \U$7748 ( \7937 , \7653 , \7662 );
or \U$7749 ( \7938 , \7935 , \7936 , \7937 );
and \U$7750 ( \7939 , \7638 , \7642 );
and \U$7751 ( \7940 , \7642 , \7647 );
and \U$7752 ( \7941 , \7638 , \7647 );
or \U$7753 ( \7942 , \7939 , \7940 , \7941 );
xor \U$7754 ( \7943 , \7938 , \7942 );
and \U$7755 ( \7944 , \7722 , \7726 );
and \U$7756 ( \7945 , \7726 , \7731 );
and \U$7757 ( \7946 , \7722 , \7731 );
or \U$7758 ( \7947 , \7944 , \7945 , \7946 );
xor \U$7759 ( \7948 , \7943 , \7947 );
xor \U$7760 ( \7949 , \7934 , \7948 );
and \U$7761 ( \7950 , \5780 , \7026 );
and \U$7762 ( \7951 , \5792 , \7024 );
nor \U$7763 ( \7952 , \7950 , \7951 );
xnor \U$7764 ( \7953 , \7952 , \7032 );
and \U$7765 ( \7954 , \5799 , \7043 );
and \U$7766 ( \7955 , \5811 , \7041 );
nor \U$7767 ( \7956 , \7954 , \7955 );
xnor \U$7768 ( \7957 , \7956 , \7049 );
xor \U$7769 ( \7958 , \7953 , \7957 );
and \U$7770 ( \7959 , \5819 , \7061 );
and \U$7771 ( \7960 , \5831 , \7059 );
nor \U$7772 ( \7961 , \7959 , \7960 );
xnor \U$7773 ( \7962 , \7961 , \7067 );
xor \U$7774 ( \7963 , \7958 , \7962 );
and \U$7775 ( \7964 , \5737 , \6991 );
not \U$7776 ( \7965 , \7964 );
xnor \U$7777 ( \7966 , \7965 , \6985 );
xor \U$7778 ( \7967 , \5816 , \7966 );
and \U$7779 ( \7968 , \5758 , \7006 );
and \U$7780 ( \7969 , \5770 , \7004 );
nor \U$7781 ( \7970 , \7968 , \7969 );
xnor \U$7782 ( \7971 , \7970 , \7012 );
xor \U$7783 ( \7972 , \7967 , \7971 );
xor \U$7784 ( \7973 , \7963 , \7972 );
and \U$7785 ( \7974 , \5967 , \7192 );
and \U$7786 ( \7975 , \5979 , \7190 );
nor \U$7787 ( \7976 , \7974 , \7975 );
xnor \U$7788 ( \7977 , \7976 , \7198 );
and \U$7789 ( \7978 , \5986 , \7203 );
and \U$7790 ( \7979 , \5998 , \7201 );
nor \U$7791 ( \7980 , \7978 , \7979 );
xnor \U$7792 ( \7981 , \7980 , \6824 );
xor \U$7793 ( \7982 , \7977 , \7981 );
and \U$7794 ( \7983 , \6006 , \5750 );
and \U$7795 ( \7984 , \6018 , \5748 );
nor \U$7796 ( \7985 , \7983 , \7984 );
xnor \U$7797 ( \7986 , \7985 , \5755 );
xor \U$7798 ( \7987 , \7982 , \7986 );
and \U$7799 ( \7988 , \5906 , \7140 );
and \U$7800 ( \7989 , \5918 , \7138 );
nor \U$7801 ( \7990 , \7988 , \7989 );
xnor \U$7802 ( \7991 , \7990 , \7146 );
and \U$7803 ( \7992 , \5925 , \7157 );
and \U$7804 ( \7993 , \5937 , \7155 );
nor \U$7805 ( \7994 , \7992 , \7993 );
xnor \U$7806 ( \7995 , \7994 , \7163 );
xor \U$7807 ( \7996 , \7991 , \7995 );
and \U$7808 ( \7997 , \5945 , \7175 );
and \U$7809 ( \7998 , \5957 , \7173 );
nor \U$7810 ( \7999 , \7997 , \7998 );
xnor \U$7811 ( \8000 , \7999 , \7181 );
xor \U$7812 ( \8001 , \7996 , \8000 );
xor \U$7813 ( \8002 , \7987 , \8001 );
and \U$7814 ( \8003 , \5842 , \7082 );
and \U$7815 ( \8004 , \5854 , \7080 );
nor \U$7816 ( \8005 , \8003 , \8004 );
xnor \U$7817 ( \8006 , \8005 , \7088 );
and \U$7818 ( \8007 , \5861 , \7099 );
and \U$7819 ( \8008 , \5873 , \7097 );
nor \U$7820 ( \8009 , \8007 , \8008 );
xnor \U$7821 ( \8010 , \8009 , \7105 );
xor \U$7822 ( \8011 , \8006 , \8010 );
and \U$7823 ( \8012 , \5881 , \7117 );
and \U$7824 ( \8013 , \5893 , \7115 );
nor \U$7825 ( \8014 , \8012 , \8013 );
xnor \U$7826 ( \8015 , \8014 , \7123 );
xor \U$7827 ( \8016 , \8011 , \8015 );
xor \U$7828 ( \8017 , \8002 , \8016 );
xor \U$7829 ( \8018 , \7973 , \8017 );
xor \U$7830 ( \8019 , \7949 , \8018 );
and \U$7831 ( \8020 , \7752 , \7756 );
and \U$7832 ( \8021 , \7756 , \7761 );
and \U$7833 ( \8022 , \7752 , \7761 );
or \U$7834 ( \8023 , \8020 , \8021 , \8022 );
and \U$7835 ( \8024 , \7737 , \7741 );
and \U$7836 ( \8025 , \7741 , \7746 );
and \U$7837 ( \8026 , \7737 , \7746 );
or \U$7838 ( \8027 , \8024 , \8025 , \8026 );
xor \U$7839 ( \8028 , \8023 , \8027 );
and \U$7840 ( \8029 , \7703 , \7717 );
and \U$7841 ( \8030 , \7717 , \7732 );
and \U$7842 ( \8031 , \7703 , \7732 );
or \U$7843 ( \8032 , \8029 , \8030 , \8031 );
xor \U$7844 ( \8033 , \8028 , \8032 );
xor \U$7845 ( \8034 , \8019 , \8033 );
xor \U$7846 ( \8035 , \7912 , \8034 );
xor \U$7847 ( \8036 , \7906 , \8035 );
and \U$7848 ( \8037 , \7586 , \7625 );
and \U$7849 ( \8038 , \7625 , \7765 );
and \U$7850 ( \8039 , \7586 , \7765 );
or \U$7851 ( \8040 , \8037 , \8038 , \8039 );
nor \U$7852 ( \8041 , \8036 , \8040 );
nor \U$7853 ( \8042 , \7887 , \8041 );
and \U$7854 ( \8043 , \7910 , \7911 );
and \U$7855 ( \8044 , \7911 , \8034 );
and \U$7856 ( \8045 , \7910 , \8034 );
or \U$7857 ( \8046 , \8043 , \8044 , \8045 );
and \U$7858 ( \8047 , \8023 , \8027 );
and \U$7859 ( \8048 , \8027 , \8032 );
and \U$7860 ( \8049 , \8023 , \8032 );
or \U$7861 ( \8050 , \8047 , \8048 , \8049 );
and \U$7862 ( \8051 , \7963 , \7972 );
and \U$7863 ( \8052 , \7972 , \8017 );
and \U$7864 ( \8053 , \7963 , \8017 );
or \U$7865 ( \8054 , \8051 , \8052 , \8053 );
xor \U$7866 ( \8055 , \8050 , \8054 );
and \U$7867 ( \8056 , \7934 , \7948 );
xor \U$7868 ( \8057 , \8055 , \8056 );
xor \U$7869 ( \8058 , \8046 , \8057 );
and \U$7870 ( \8059 , \7895 , \7899 );
and \U$7871 ( \8060 , \7899 , \7904 );
and \U$7872 ( \8061 , \7895 , \7904 );
or \U$7873 ( \8062 , \8059 , \8060 , \8061 );
and \U$7874 ( \8063 , \7949 , \8018 );
and \U$7875 ( \8064 , \8018 , \8033 );
and \U$7876 ( \8065 , \7949 , \8033 );
or \U$7877 ( \8066 , \8063 , \8064 , \8065 );
xor \U$7878 ( \8067 , \8062 , \8066 );
and \U$7879 ( \8068 , \5816 , \7966 );
and \U$7880 ( \8069 , \7966 , \7971 );
and \U$7881 ( \8070 , \5816 , \7971 );
or \U$7882 ( \8071 , \8068 , \8069 , \8070 );
and \U$7883 ( \8072 , \7953 , \7957 );
and \U$7884 ( \8073 , \7957 , \7962 );
and \U$7885 ( \8074 , \7953 , \7962 );
or \U$7886 ( \8075 , \8072 , \8073 , \8074 );
xor \U$7887 ( \8076 , \8071 , \8075 );
and \U$7888 ( \8077 , \8006 , \8010 );
and \U$7889 ( \8078 , \8010 , \8015 );
and \U$7890 ( \8079 , \8006 , \8015 );
or \U$7891 ( \8080 , \8077 , \8078 , \8079 );
xor \U$7892 ( \8081 , \8076 , \8080 );
and \U$7893 ( \8082 , \5873 , \7099 );
and \U$7894 ( \8083 , \5842 , \7097 );
nor \U$7895 ( \8084 , \8082 , \8083 );
xnor \U$7896 ( \8085 , \8084 , \7105 );
and \U$7897 ( \8086 , \5893 , \7117 );
and \U$7898 ( \8087 , \5861 , \7115 );
nor \U$7899 ( \8088 , \8086 , \8087 );
xnor \U$7900 ( \8089 , \8088 , \7123 );
xor \U$7901 ( \8090 , \8085 , \8089 );
and \U$7902 ( \8091 , \5918 , \7140 );
and \U$7903 ( \8092 , \5881 , \7138 );
nor \U$7904 ( \8093 , \8091 , \8092 );
xnor \U$7905 ( \8094 , \8093 , \7146 );
xor \U$7906 ( \8095 , \8090 , \8094 );
and \U$7907 ( \8096 , \5811 , \7043 );
and \U$7908 ( \8097 , \5780 , \7041 );
nor \U$7909 ( \8098 , \8096 , \8097 );
xnor \U$7910 ( \8099 , \8098 , \7049 );
and \U$7911 ( \8100 , \5831 , \7061 );
and \U$7912 ( \8101 , \5799 , \7059 );
nor \U$7913 ( \8102 , \8100 , \8101 );
xnor \U$7914 ( \8103 , \8102 , \7067 );
xor \U$7915 ( \8104 , \8099 , \8103 );
and \U$7916 ( \8105 , \5854 , \7082 );
and \U$7917 ( \8106 , \5819 , \7080 );
nor \U$7918 ( \8107 , \8105 , \8106 );
xnor \U$7919 ( \8108 , \8107 , \7088 );
xor \U$7920 ( \8109 , \8104 , \8108 );
xor \U$7921 ( \8110 , \8095 , \8109 );
not \U$7922 ( \8111 , \6985 );
and \U$7923 ( \8112 , \5770 , \7006 );
and \U$7924 ( \8113 , \5737 , \7004 );
nor \U$7925 ( \8114 , \8112 , \8113 );
xnor \U$7926 ( \8115 , \8114 , \7012 );
xor \U$7927 ( \8116 , \8111 , \8115 );
and \U$7928 ( \8117 , \5792 , \7026 );
and \U$7929 ( \8118 , \5758 , \7024 );
nor \U$7930 ( \8119 , \8117 , \8118 );
xnor \U$7931 ( \8120 , \8119 , \7032 );
xor \U$7932 ( \8121 , \8116 , \8120 );
xor \U$7933 ( \8122 , \8110 , \8121 );
and \U$7934 ( \8123 , \6057 , \5790 );
and \U$7935 ( \8124 , \6029 , \5788 );
nor \U$7936 ( \8125 , \8123 , \8124 );
xnor \U$7937 ( \8126 , \8125 , \5797 );
and \U$7938 ( \8127 , \6065 , \5809 );
and \U$7939 ( \8128 , \6048 , \5807 );
nor \U$7940 ( \8129 , \8127 , \8128 );
xnor \U$7941 ( \8130 , \8129 , \5816 );
xnor \U$7942 ( \8131 , \8126 , \8130 );
and \U$7943 ( \8132 , \5998 , \7203 );
and \U$7944 ( \8133 , \5967 , \7201 );
nor \U$7945 ( \8134 , \8132 , \8133 );
xnor \U$7946 ( \8135 , \8134 , \6824 );
and \U$7947 ( \8136 , \6018 , \5750 );
and \U$7948 ( \8137 , \5986 , \5748 );
nor \U$7949 ( \8138 , \8136 , \8137 );
xnor \U$7950 ( \8139 , \8138 , \5755 );
xor \U$7951 ( \8140 , \8135 , \8139 );
and \U$7952 ( \8141 , \6041 , \5768 );
and \U$7953 ( \8142 , \6006 , \5766 );
nor \U$7954 ( \8143 , \8141 , \8142 );
xnor \U$7955 ( \8144 , \8143 , \5775 );
xor \U$7956 ( \8145 , \8140 , \8144 );
xor \U$7957 ( \8146 , \8131 , \8145 );
and \U$7958 ( \8147 , \5937 , \7157 );
and \U$7959 ( \8148 , \5906 , \7155 );
nor \U$7960 ( \8149 , \8147 , \8148 );
xnor \U$7961 ( \8150 , \8149 , \7163 );
and \U$7962 ( \8151 , \5957 , \7175 );
and \U$7963 ( \8152 , \5925 , \7173 );
nor \U$7964 ( \8153 , \8151 , \8152 );
xnor \U$7965 ( \8154 , \8153 , \7181 );
xor \U$7966 ( \8155 , \8150 , \8154 );
and \U$7967 ( \8156 , \5979 , \7192 );
and \U$7968 ( \8157 , \5945 , \7190 );
nor \U$7969 ( \8158 , \8156 , \8157 );
xnor \U$7970 ( \8159 , \8158 , \7198 );
xor \U$7971 ( \8160 , \8155 , \8159 );
xor \U$7972 ( \8161 , \8146 , \8160 );
xor \U$7973 ( \8162 , \8122 , \8161 );
and \U$7974 ( \8163 , \7991 , \7995 );
and \U$7975 ( \8164 , \7995 , \8000 );
and \U$7976 ( \8165 , \7991 , \8000 );
or \U$7977 ( \8166 , \8163 , \8164 , \8165 );
and \U$7978 ( \8167 , \7977 , \7981 );
and \U$7979 ( \8168 , \7981 , \7986 );
and \U$7980 ( \8169 , \7977 , \7986 );
or \U$7981 ( \8170 , \8167 , \8168 , \8169 );
xor \U$7982 ( \8171 , \8166 , \8170 );
and \U$7983 ( \8172 , \7925 , \7929 );
and \U$7984 ( \8173 , \7929 , \7932 );
and \U$7985 ( \8174 , \7925 , \7932 );
or \U$7986 ( \8175 , \8172 , \8173 , \8174 );
xor \U$7987 ( \8176 , \8171 , \8175 );
xor \U$7988 ( \8177 , \8162 , \8176 );
xor \U$7989 ( \8178 , \8081 , \8177 );
and \U$7990 ( \8179 , \7938 , \7942 );
and \U$7991 ( \8180 , \7942 , \7947 );
and \U$7992 ( \8181 , \7938 , \7947 );
or \U$7993 ( \8182 , \8179 , \8180 , \8181 );
and \U$7994 ( \8183 , \7916 , \7920 );
and \U$7995 ( \8184 , \7920 , \7933 );
and \U$7996 ( \8185 , \7916 , \7933 );
or \U$7997 ( \8186 , \8183 , \8184 , \8185 );
xor \U$7998 ( \8187 , \8182 , \8186 );
and \U$7999 ( \8188 , \7987 , \8001 );
and \U$8000 ( \8189 , \8001 , \8016 );
and \U$8001 ( \8190 , \7987 , \8016 );
or \U$8002 ( \8191 , \8188 , \8189 , \8190 );
xor \U$8003 ( \8192 , \8187 , \8191 );
xor \U$8004 ( \8193 , \8178 , \8192 );
xor \U$8005 ( \8194 , \8067 , \8193 );
xor \U$8006 ( \8195 , \8058 , \8194 );
and \U$8007 ( \8196 , \7891 , \7905 );
and \U$8008 ( \8197 , \7905 , \8035 );
and \U$8009 ( \8198 , \7891 , \8035 );
or \U$8010 ( \8199 , \8196 , \8197 , \8198 );
nor \U$8011 ( \8200 , \8195 , \8199 );
and \U$8012 ( \8201 , \8062 , \8066 );
and \U$8013 ( \8202 , \8066 , \8193 );
and \U$8014 ( \8203 , \8062 , \8193 );
or \U$8015 ( \8204 , \8201 , \8202 , \8203 );
and \U$8016 ( \8205 , \8071 , \8075 );
and \U$8017 ( \8206 , \8075 , \8080 );
and \U$8018 ( \8207 , \8071 , \8080 );
or \U$8019 ( \8208 , \8205 , \8206 , \8207 );
and \U$8020 ( \8209 , \8166 , \8170 );
and \U$8021 ( \8210 , \8170 , \8175 );
and \U$8022 ( \8211 , \8166 , \8175 );
or \U$8023 ( \8212 , \8209 , \8210 , \8211 );
xor \U$8024 ( \8213 , \8208 , \8212 );
and \U$8025 ( \8214 , \8131 , \8145 );
and \U$8026 ( \8215 , \8145 , \8160 );
and \U$8027 ( \8216 , \8131 , \8160 );
or \U$8028 ( \8217 , \8214 , \8215 , \8216 );
xor \U$8029 ( \8218 , \8213 , \8217 );
and \U$8030 ( \8219 , \8182 , \8186 );
and \U$8031 ( \8220 , \8186 , \8191 );
and \U$8032 ( \8221 , \8182 , \8191 );
or \U$8033 ( \8222 , \8219 , \8220 , \8221 );
and \U$8034 ( \8223 , \8122 , \8161 );
and \U$8035 ( \8224 , \8161 , \8176 );
and \U$8036 ( \8225 , \8122 , \8176 );
or \U$8037 ( \8226 , \8223 , \8224 , \8225 );
xor \U$8038 ( \8227 , \8222 , \8226 );
and \U$8039 ( \8228 , \6029 , \5790 );
and \U$8040 ( \8229 , \6041 , \5788 );
nor \U$8041 ( \8230 , \8228 , \8229 );
xnor \U$8042 ( \8231 , \8230 , \5797 );
and \U$8043 ( \8232 , \6048 , \5809 );
and \U$8044 ( \8233 , \6057 , \5807 );
nor \U$8045 ( \8234 , \8232 , \8233 );
xnor \U$8046 ( \8235 , \8234 , \5816 );
xor \U$8047 ( \8236 , \8231 , \8235 );
nand \U$8048 ( \8237 , \6065 , \5827 );
xnor \U$8049 ( \8238 , \8237 , \5836 );
xor \U$8050 ( \8239 , \8236 , \8238 );
and \U$8051 ( \8240 , \5967 , \7203 );
and \U$8052 ( \8241 , \5979 , \7201 );
nor \U$8053 ( \8242 , \8240 , \8241 );
xnor \U$8054 ( \8243 , \8242 , \6824 );
and \U$8055 ( \8244 , \5986 , \5750 );
and \U$8056 ( \8245 , \5998 , \5748 );
nor \U$8057 ( \8246 , \8244 , \8245 );
xnor \U$8058 ( \8247 , \8246 , \5755 );
xor \U$8059 ( \8248 , \8243 , \8247 );
and \U$8060 ( \8249 , \6006 , \5768 );
and \U$8061 ( \8250 , \6018 , \5766 );
nor \U$8062 ( \8251 , \8249 , \8250 );
xnor \U$8063 ( \8252 , \8251 , \5775 );
xor \U$8064 ( \8253 , \8248 , \8252 );
xnor \U$8065 ( \8254 , \8239 , \8253 );
and \U$8066 ( \8255 , \8150 , \8154 );
and \U$8067 ( \8256 , \8154 , \8159 );
and \U$8068 ( \8257 , \8150 , \8159 );
or \U$8069 ( \8258 , \8255 , \8256 , \8257 );
and \U$8070 ( \8259 , \8135 , \8139 );
and \U$8071 ( \8260 , \8139 , \8144 );
and \U$8072 ( \8261 , \8135 , \8144 );
or \U$8073 ( \8262 , \8259 , \8260 , \8261 );
xor \U$8074 ( \8263 , \8258 , \8262 );
or \U$8075 ( \8264 , \8126 , \8130 );
xor \U$8076 ( \8265 , \8263 , \8264 );
xor \U$8077 ( \8266 , \8254 , \8265 );
and \U$8078 ( \8267 , \8111 , \8115 );
and \U$8079 ( \8268 , \8115 , \8120 );
and \U$8080 ( \8269 , \8111 , \8120 );
or \U$8081 ( \8270 , \8267 , \8268 , \8269 );
and \U$8082 ( \8271 , \8099 , \8103 );
and \U$8083 ( \8272 , \8103 , \8108 );
and \U$8084 ( \8273 , \8099 , \8108 );
or \U$8085 ( \8274 , \8271 , \8272 , \8273 );
xor \U$8086 ( \8275 , \8270 , \8274 );
and \U$8087 ( \8276 , \8085 , \8089 );
and \U$8088 ( \8277 , \8089 , \8094 );
and \U$8089 ( \8278 , \8085 , \8094 );
or \U$8090 ( \8279 , \8276 , \8277 , \8278 );
xor \U$8091 ( \8280 , \8275 , \8279 );
xor \U$8092 ( \8281 , \8266 , \8280 );
xor \U$8093 ( \8282 , \8227 , \8281 );
xor \U$8094 ( \8283 , \8218 , \8282 );
xor \U$8095 ( \8284 , \8204 , \8283 );
and \U$8096 ( \8285 , \8050 , \8054 );
and \U$8097 ( \8286 , \8054 , \8056 );
and \U$8098 ( \8287 , \8050 , \8056 );
or \U$8099 ( \8288 , \8285 , \8286 , \8287 );
and \U$8100 ( \8289 , \8081 , \8177 );
and \U$8101 ( \8290 , \8177 , \8192 );
and \U$8102 ( \8291 , \8081 , \8192 );
or \U$8103 ( \8292 , \8289 , \8290 , \8291 );
xor \U$8104 ( \8293 , \8288 , \8292 );
and \U$8105 ( \8294 , \8095 , \8109 );
and \U$8106 ( \8295 , \8109 , \8121 );
and \U$8107 ( \8296 , \8095 , \8121 );
or \U$8108 ( \8297 , \8294 , \8295 , \8296 );
and \U$8109 ( \8298 , \5737 , \7006 );
not \U$8110 ( \8299 , \8298 );
xnor \U$8111 ( \8300 , \8299 , \7012 );
xor \U$8112 ( \8301 , \5836 , \8300 );
and \U$8113 ( \8302 , \5758 , \7026 );
and \U$8114 ( \8303 , \5770 , \7024 );
nor \U$8115 ( \8304 , \8302 , \8303 );
xnor \U$8116 ( \8305 , \8304 , \7032 );
xor \U$8117 ( \8306 , \8301 , \8305 );
xor \U$8118 ( \8307 , \8297 , \8306 );
and \U$8119 ( \8308 , \5906 , \7157 );
and \U$8120 ( \8309 , \5918 , \7155 );
nor \U$8121 ( \8310 , \8308 , \8309 );
xnor \U$8122 ( \8311 , \8310 , \7163 );
and \U$8123 ( \8312 , \5925 , \7175 );
and \U$8124 ( \8313 , \5937 , \7173 );
nor \U$8125 ( \8314 , \8312 , \8313 );
xnor \U$8126 ( \8315 , \8314 , \7181 );
xor \U$8127 ( \8316 , \8311 , \8315 );
and \U$8128 ( \8317 , \5945 , \7192 );
and \U$8129 ( \8318 , \5957 , \7190 );
nor \U$8130 ( \8319 , \8317 , \8318 );
xnor \U$8131 ( \8320 , \8319 , \7198 );
xor \U$8132 ( \8321 , \8316 , \8320 );
and \U$8133 ( \8322 , \5842 , \7099 );
and \U$8134 ( \8323 , \5854 , \7097 );
nor \U$8135 ( \8324 , \8322 , \8323 );
xnor \U$8136 ( \8325 , \8324 , \7105 );
and \U$8137 ( \8326 , \5861 , \7117 );
and \U$8138 ( \8327 , \5873 , \7115 );
nor \U$8139 ( \8328 , \8326 , \8327 );
xnor \U$8140 ( \8329 , \8328 , \7123 );
xor \U$8141 ( \8330 , \8325 , \8329 );
and \U$8142 ( \8331 , \5881 , \7140 );
and \U$8143 ( \8332 , \5893 , \7138 );
nor \U$8144 ( \8333 , \8331 , \8332 );
xnor \U$8145 ( \8334 , \8333 , \7146 );
xor \U$8146 ( \8335 , \8330 , \8334 );
xor \U$8147 ( \8336 , \8321 , \8335 );
and \U$8148 ( \8337 , \5780 , \7043 );
and \U$8149 ( \8338 , \5792 , \7041 );
nor \U$8150 ( \8339 , \8337 , \8338 );
xnor \U$8151 ( \8340 , \8339 , \7049 );
and \U$8152 ( \8341 , \5799 , \7061 );
and \U$8153 ( \8342 , \5811 , \7059 );
nor \U$8154 ( \8343 , \8341 , \8342 );
xnor \U$8155 ( \8344 , \8343 , \7067 );
xor \U$8156 ( \8345 , \8340 , \8344 );
and \U$8157 ( \8346 , \5819 , \7082 );
and \U$8158 ( \8347 , \5831 , \7080 );
nor \U$8159 ( \8348 , \8346 , \8347 );
xnor \U$8160 ( \8349 , \8348 , \7088 );
xor \U$8161 ( \8350 , \8345 , \8349 );
xor \U$8162 ( \8351 , \8336 , \8350 );
xor \U$8163 ( \8352 , \8307 , \8351 );
xor \U$8164 ( \8353 , \8293 , \8352 );
xor \U$8165 ( \8354 , \8284 , \8353 );
and \U$8166 ( \8355 , \8046 , \8057 );
and \U$8167 ( \8356 , \8057 , \8194 );
and \U$8168 ( \8357 , \8046 , \8194 );
or \U$8169 ( \8358 , \8355 , \8356 , \8357 );
nor \U$8170 ( \8359 , \8354 , \8358 );
nor \U$8171 ( \8360 , \8200 , \8359 );
nand \U$8172 ( \8361 , \8042 , \8360 );
and \U$8173 ( \8362 , \8288 , \8292 );
and \U$8174 ( \8363 , \8292 , \8352 );
and \U$8175 ( \8364 , \8288 , \8352 );
or \U$8176 ( \8365 , \8362 , \8363 , \8364 );
and \U$8177 ( \8366 , \8218 , \8282 );
xor \U$8178 ( \8367 , \8365 , \8366 );
and \U$8179 ( \8368 , \8222 , \8226 );
and \U$8180 ( \8369 , \8226 , \8281 );
and \U$8181 ( \8370 , \8222 , \8281 );
or \U$8182 ( \8371 , \8368 , \8369 , \8370 );
and \U$8183 ( \8372 , \8311 , \8315 );
and \U$8184 ( \8373 , \8315 , \8320 );
and \U$8185 ( \8374 , \8311 , \8320 );
or \U$8186 ( \8375 , \8372 , \8373 , \8374 );
and \U$8187 ( \8376 , \8243 , \8247 );
and \U$8188 ( \8377 , \8247 , \8252 );
and \U$8189 ( \8378 , \8243 , \8252 );
or \U$8190 ( \8379 , \8376 , \8377 , \8378 );
xor \U$8191 ( \8380 , \8375 , \8379 );
and \U$8192 ( \8381 , \8231 , \8235 );
and \U$8193 ( \8382 , \8235 , \8238 );
and \U$8194 ( \8383 , \8231 , \8238 );
or \U$8195 ( \8384 , \8381 , \8382 , \8383 );
xor \U$8196 ( \8385 , \8380 , \8384 );
and \U$8197 ( \8386 , \5836 , \8300 );
and \U$8198 ( \8387 , \8300 , \8305 );
and \U$8199 ( \8388 , \5836 , \8305 );
or \U$8200 ( \8389 , \8386 , \8387 , \8388 );
and \U$8201 ( \8390 , \8340 , \8344 );
and \U$8202 ( \8391 , \8344 , \8349 );
and \U$8203 ( \8392 , \8340 , \8349 );
or \U$8204 ( \8393 , \8390 , \8391 , \8392 );
xor \U$8205 ( \8394 , \8389 , \8393 );
and \U$8206 ( \8395 , \8325 , \8329 );
and \U$8207 ( \8396 , \8329 , \8334 );
and \U$8208 ( \8397 , \8325 , \8334 );
or \U$8209 ( \8398 , \8395 , \8396 , \8397 );
xor \U$8210 ( \8399 , \8394 , \8398 );
xor \U$8211 ( \8400 , \8385 , \8399 );
and \U$8212 ( \8401 , \8321 , \8335 );
and \U$8213 ( \8402 , \8335 , \8350 );
and \U$8214 ( \8403 , \8321 , \8350 );
or \U$8215 ( \8404 , \8401 , \8402 , \8403 );
and \U$8216 ( \8405 , \5873 , \7117 );
and \U$8217 ( \8406 , \5842 , \7115 );
nor \U$8218 ( \8407 , \8405 , \8406 );
xnor \U$8219 ( \8408 , \8407 , \7123 );
and \U$8220 ( \8409 , \5893 , \7140 );
and \U$8221 ( \8410 , \5861 , \7138 );
nor \U$8222 ( \8411 , \8409 , \8410 );
xnor \U$8223 ( \8412 , \8411 , \7146 );
xor \U$8224 ( \8413 , \8408 , \8412 );
and \U$8225 ( \8414 , \5918 , \7157 );
and \U$8226 ( \8415 , \5881 , \7155 );
nor \U$8227 ( \8416 , \8414 , \8415 );
xnor \U$8228 ( \8417 , \8416 , \7163 );
xor \U$8229 ( \8418 , \8413 , \8417 );
and \U$8230 ( \8419 , \5811 , \7061 );
and \U$8231 ( \8420 , \5780 , \7059 );
nor \U$8232 ( \8421 , \8419 , \8420 );
xnor \U$8233 ( \8422 , \8421 , \7067 );
and \U$8234 ( \8423 , \5831 , \7082 );
and \U$8235 ( \8424 , \5799 , \7080 );
nor \U$8236 ( \8425 , \8423 , \8424 );
xnor \U$8237 ( \8426 , \8425 , \7088 );
xor \U$8238 ( \8427 , \8422 , \8426 );
and \U$8239 ( \8428 , \5854 , \7099 );
and \U$8240 ( \8429 , \5819 , \7097 );
nor \U$8241 ( \8430 , \8428 , \8429 );
xnor \U$8242 ( \8431 , \8430 , \7105 );
xor \U$8243 ( \8432 , \8427 , \8431 );
xor \U$8244 ( \8433 , \8418 , \8432 );
not \U$8245 ( \8434 , \7012 );
and \U$8246 ( \8435 , \5770 , \7026 );
and \U$8247 ( \8436 , \5737 , \7024 );
nor \U$8248 ( \8437 , \8435 , \8436 );
xnor \U$8249 ( \8438 , \8437 , \7032 );
xor \U$8250 ( \8439 , \8434 , \8438 );
and \U$8251 ( \8440 , \5792 , \7043 );
and \U$8252 ( \8441 , \5758 , \7041 );
nor \U$8253 ( \8442 , \8440 , \8441 );
xnor \U$8254 ( \8443 , \8442 , \7049 );
xor \U$8255 ( \8444 , \8439 , \8443 );
xor \U$8256 ( \8445 , \8433 , \8444 );
xor \U$8257 ( \8446 , \8404 , \8445 );
and \U$8258 ( \8447 , \6057 , \5809 );
and \U$8259 ( \8448 , \6029 , \5807 );
nor \U$8260 ( \8449 , \8447 , \8448 );
xnor \U$8261 ( \8450 , \8449 , \5816 );
and \U$8262 ( \8451 , \6065 , \5829 );
and \U$8263 ( \8452 , \6048 , \5827 );
nor \U$8264 ( \8453 , \8451 , \8452 );
xnor \U$8265 ( \8454 , \8453 , \5836 );
xor \U$8266 ( \8455 , \8450 , \8454 );
and \U$8267 ( \8456 , \5998 , \5750 );
and \U$8268 ( \8457 , \5967 , \5748 );
nor \U$8269 ( \8458 , \8456 , \8457 );
xnor \U$8270 ( \8459 , \8458 , \5755 );
and \U$8271 ( \8460 , \6018 , \5768 );
and \U$8272 ( \8461 , \5986 , \5766 );
nor \U$8273 ( \8462 , \8460 , \8461 );
xnor \U$8274 ( \8463 , \8462 , \5775 );
xor \U$8275 ( \8464 , \8459 , \8463 );
and \U$8276 ( \8465 , \6041 , \5790 );
and \U$8277 ( \8466 , \6006 , \5788 );
nor \U$8278 ( \8467 , \8465 , \8466 );
xnor \U$8279 ( \8468 , \8467 , \5797 );
xor \U$8280 ( \8469 , \8464 , \8468 );
xor \U$8281 ( \8470 , \8455 , \8469 );
and \U$8282 ( \8471 , \5937 , \7175 );
and \U$8283 ( \8472 , \5906 , \7173 );
nor \U$8284 ( \8473 , \8471 , \8472 );
xnor \U$8285 ( \8474 , \8473 , \7181 );
and \U$8286 ( \8475 , \5957 , \7192 );
and \U$8287 ( \8476 , \5925 , \7190 );
nor \U$8288 ( \8477 , \8475 , \8476 );
xnor \U$8289 ( \8478 , \8477 , \7198 );
xor \U$8290 ( \8479 , \8474 , \8478 );
and \U$8291 ( \8480 , \5979 , \7203 );
and \U$8292 ( \8481 , \5945 , \7201 );
nor \U$8293 ( \8482 , \8480 , \8481 );
xnor \U$8294 ( \8483 , \8482 , \6824 );
xor \U$8295 ( \8484 , \8479 , \8483 );
xor \U$8296 ( \8485 , \8470 , \8484 );
xor \U$8297 ( \8486 , \8446 , \8485 );
xor \U$8298 ( \8487 , \8400 , \8486 );
and \U$8299 ( \8488 , \8270 , \8274 );
and \U$8300 ( \8489 , \8274 , \8279 );
and \U$8301 ( \8490 , \8270 , \8279 );
or \U$8302 ( \8491 , \8488 , \8489 , \8490 );
and \U$8303 ( \8492 , \8258 , \8262 );
and \U$8304 ( \8493 , \8262 , \8264 );
and \U$8305 ( \8494 , \8258 , \8264 );
or \U$8306 ( \8495 , \8492 , \8493 , \8494 );
xor \U$8307 ( \8496 , \8491 , \8495 );
or \U$8308 ( \8497 , \8239 , \8253 );
xor \U$8309 ( \8498 , \8496 , \8497 );
xor \U$8310 ( \8499 , \8487 , \8498 );
xor \U$8311 ( \8500 , \8371 , \8499 );
and \U$8312 ( \8501 , \8208 , \8212 );
and \U$8313 ( \8502 , \8212 , \8217 );
and \U$8314 ( \8503 , \8208 , \8217 );
or \U$8315 ( \8504 , \8501 , \8502 , \8503 );
and \U$8316 ( \8505 , \8297 , \8306 );
and \U$8317 ( \8506 , \8306 , \8351 );
and \U$8318 ( \8507 , \8297 , \8351 );
or \U$8319 ( \8508 , \8505 , \8506 , \8507 );
xor \U$8320 ( \8509 , \8504 , \8508 );
and \U$8321 ( \8510 , \8254 , \8265 );
and \U$8322 ( \8511 , \8265 , \8280 );
and \U$8323 ( \8512 , \8254 , \8280 );
or \U$8324 ( \8513 , \8510 , \8511 , \8512 );
xor \U$8325 ( \8514 , \8509 , \8513 );
xor \U$8326 ( \8515 , \8500 , \8514 );
xor \U$8327 ( \8516 , \8367 , \8515 );
and \U$8328 ( \8517 , \8204 , \8283 );
and \U$8329 ( \8518 , \8283 , \8353 );
and \U$8330 ( \8519 , \8204 , \8353 );
or \U$8331 ( \8520 , \8517 , \8518 , \8519 );
nor \U$8332 ( \8521 , \8516 , \8520 );
and \U$8333 ( \8522 , \8371 , \8499 );
and \U$8334 ( \8523 , \8499 , \8514 );
and \U$8335 ( \8524 , \8371 , \8514 );
or \U$8336 ( \8525 , \8522 , \8523 , \8524 );
and \U$8337 ( \8526 , \8491 , \8495 );
and \U$8338 ( \8527 , \8495 , \8497 );
and \U$8339 ( \8528 , \8491 , \8497 );
or \U$8340 ( \8529 , \8526 , \8527 , \8528 );
and \U$8341 ( \8530 , \8404 , \8445 );
and \U$8342 ( \8531 , \8445 , \8485 );
and \U$8343 ( \8532 , \8404 , \8485 );
or \U$8344 ( \8533 , \8530 , \8531 , \8532 );
xor \U$8345 ( \8534 , \8529 , \8533 );
and \U$8346 ( \8535 , \8385 , \8399 );
xor \U$8347 ( \8536 , \8534 , \8535 );
xor \U$8348 ( \8537 , \8525 , \8536 );
and \U$8349 ( \8538 , \8504 , \8508 );
and \U$8350 ( \8539 , \8508 , \8513 );
and \U$8351 ( \8540 , \8504 , \8513 );
or \U$8352 ( \8541 , \8538 , \8539 , \8540 );
and \U$8353 ( \8542 , \8400 , \8486 );
and \U$8354 ( \8543 , \8486 , \8498 );
and \U$8355 ( \8544 , \8400 , \8498 );
or \U$8356 ( \8545 , \8542 , \8543 , \8544 );
xor \U$8357 ( \8546 , \8541 , \8545 );
and \U$8358 ( \8547 , \6029 , \5809 );
and \U$8359 ( \8548 , \6041 , \5807 );
nor \U$8360 ( \8549 , \8547 , \8548 );
xnor \U$8361 ( \8550 , \8549 , \5816 );
and \U$8362 ( \8551 , \6048 , \5829 );
and \U$8363 ( \8552 , \6057 , \5827 );
nor \U$8364 ( \8553 , \8551 , \8552 );
xnor \U$8365 ( \8554 , \8553 , \5836 );
xor \U$8366 ( \8555 , \8550 , \8554 );
nand \U$8367 ( \8556 , \6065 , \5850 );
xnor \U$8368 ( \8557 , \8556 , \5859 );
xor \U$8369 ( \8558 , \8555 , \8557 );
and \U$8370 ( \8559 , \5967 , \5750 );
and \U$8371 ( \8560 , \5979 , \5748 );
nor \U$8372 ( \8561 , \8559 , \8560 );
xnor \U$8373 ( \8562 , \8561 , \5755 );
and \U$8374 ( \8563 , \5986 , \5768 );
and \U$8375 ( \8564 , \5998 , \5766 );
nor \U$8376 ( \8565 , \8563 , \8564 );
xnor \U$8377 ( \8566 , \8565 , \5775 );
xor \U$8378 ( \8567 , \8562 , \8566 );
and \U$8379 ( \8568 , \6006 , \5790 );
and \U$8380 ( \8569 , \6018 , \5788 );
nor \U$8381 ( \8570 , \8568 , \8569 );
xnor \U$8382 ( \8571 , \8570 , \5797 );
xor \U$8383 ( \8572 , \8567 , \8571 );
xnor \U$8384 ( \8573 , \8558 , \8572 );
and \U$8385 ( \8574 , \8474 , \8478 );
and \U$8386 ( \8575 , \8478 , \8483 );
and \U$8387 ( \8576 , \8474 , \8483 );
or \U$8388 ( \8577 , \8574 , \8575 , \8576 );
and \U$8389 ( \8578 , \8459 , \8463 );
and \U$8390 ( \8579 , \8463 , \8468 );
and \U$8391 ( \8580 , \8459 , \8468 );
or \U$8392 ( \8581 , \8578 , \8579 , \8580 );
xor \U$8393 ( \8582 , \8577 , \8581 );
and \U$8394 ( \8583 , \8450 , \8454 );
xor \U$8395 ( \8584 , \8582 , \8583 );
xor \U$8396 ( \8585 , \8573 , \8584 );
and \U$8397 ( \8586 , \8434 , \8438 );
and \U$8398 ( \8587 , \8438 , \8443 );
and \U$8399 ( \8588 , \8434 , \8443 );
or \U$8400 ( \8589 , \8586 , \8587 , \8588 );
and \U$8401 ( \8590 , \8422 , \8426 );
and \U$8402 ( \8591 , \8426 , \8431 );
and \U$8403 ( \8592 , \8422 , \8431 );
or \U$8404 ( \8593 , \8590 , \8591 , \8592 );
xor \U$8405 ( \8594 , \8589 , \8593 );
and \U$8406 ( \8595 , \8408 , \8412 );
and \U$8407 ( \8596 , \8412 , \8417 );
and \U$8408 ( \8597 , \8408 , \8417 );
or \U$8409 ( \8598 , \8595 , \8596 , \8597 );
xor \U$8410 ( \8599 , \8594 , \8598 );
xor \U$8411 ( \8600 , \8585 , \8599 );
and \U$8412 ( \8601 , \8418 , \8432 );
and \U$8413 ( \8602 , \8432 , \8444 );
and \U$8414 ( \8603 , \8418 , \8444 );
or \U$8415 ( \8604 , \8601 , \8602 , \8603 );
and \U$8416 ( \8605 , \5737 , \7026 );
not \U$8417 ( \8606 , \8605 );
xnor \U$8418 ( \8607 , \8606 , \7032 );
xor \U$8419 ( \8608 , \5859 , \8607 );
and \U$8420 ( \8609 , \5758 , \7043 );
and \U$8421 ( \8610 , \5770 , \7041 );
nor \U$8422 ( \8611 , \8609 , \8610 );
xnor \U$8423 ( \8612 , \8611 , \7049 );
xor \U$8424 ( \8613 , \8608 , \8612 );
xor \U$8425 ( \8614 , \8604 , \8613 );
and \U$8426 ( \8615 , \5906 , \7175 );
and \U$8427 ( \8616 , \5918 , \7173 );
nor \U$8428 ( \8617 , \8615 , \8616 );
xnor \U$8429 ( \8618 , \8617 , \7181 );
and \U$8430 ( \8619 , \5925 , \7192 );
and \U$8431 ( \8620 , \5937 , \7190 );
nor \U$8432 ( \8621 , \8619 , \8620 );
xnor \U$8433 ( \8622 , \8621 , \7198 );
xor \U$8434 ( \8623 , \8618 , \8622 );
and \U$8435 ( \8624 , \5945 , \7203 );
and \U$8436 ( \8625 , \5957 , \7201 );
nor \U$8437 ( \8626 , \8624 , \8625 );
xnor \U$8438 ( \8627 , \8626 , \6824 );
xor \U$8439 ( \8628 , \8623 , \8627 );
and \U$8440 ( \8629 , \5842 , \7117 );
and \U$8441 ( \8630 , \5854 , \7115 );
nor \U$8442 ( \8631 , \8629 , \8630 );
xnor \U$8443 ( \8632 , \8631 , \7123 );
and \U$8444 ( \8633 , \5861 , \7140 );
and \U$8445 ( \8634 , \5873 , \7138 );
nor \U$8446 ( \8635 , \8633 , \8634 );
xnor \U$8447 ( \8636 , \8635 , \7146 );
xor \U$8448 ( \8637 , \8632 , \8636 );
and \U$8449 ( \8638 , \5881 , \7157 );
and \U$8450 ( \8639 , \5893 , \7155 );
nor \U$8451 ( \8640 , \8638 , \8639 );
xnor \U$8452 ( \8641 , \8640 , \7163 );
xor \U$8453 ( \8642 , \8637 , \8641 );
xor \U$8454 ( \8643 , \8628 , \8642 );
and \U$8455 ( \8644 , \5780 , \7061 );
and \U$8456 ( \8645 , \5792 , \7059 );
nor \U$8457 ( \8646 , \8644 , \8645 );
xnor \U$8458 ( \8647 , \8646 , \7067 );
and \U$8459 ( \8648 , \5799 , \7082 );
and \U$8460 ( \8649 , \5811 , \7080 );
nor \U$8461 ( \8650 , \8648 , \8649 );
xnor \U$8462 ( \8651 , \8650 , \7088 );
xor \U$8463 ( \8652 , \8647 , \8651 );
and \U$8464 ( \8653 , \5819 , \7099 );
and \U$8465 ( \8654 , \5831 , \7097 );
nor \U$8466 ( \8655 , \8653 , \8654 );
xnor \U$8467 ( \8656 , \8655 , \7105 );
xor \U$8468 ( \8657 , \8652 , \8656 );
xor \U$8469 ( \8658 , \8643 , \8657 );
xor \U$8470 ( \8659 , \8614 , \8658 );
xor \U$8471 ( \8660 , \8600 , \8659 );
and \U$8472 ( \8661 , \8389 , \8393 );
and \U$8473 ( \8662 , \8393 , \8398 );
and \U$8474 ( \8663 , \8389 , \8398 );
or \U$8475 ( \8664 , \8661 , \8662 , \8663 );
and \U$8476 ( \8665 , \8375 , \8379 );
and \U$8477 ( \8666 , \8379 , \8384 );
and \U$8478 ( \8667 , \8375 , \8384 );
or \U$8479 ( \8668 , \8665 , \8666 , \8667 );
xor \U$8480 ( \8669 , \8664 , \8668 );
and \U$8481 ( \8670 , \8455 , \8469 );
and \U$8482 ( \8671 , \8469 , \8484 );
and \U$8483 ( \8672 , \8455 , \8484 );
or \U$8484 ( \8673 , \8670 , \8671 , \8672 );
xor \U$8485 ( \8674 , \8669 , \8673 );
xor \U$8486 ( \8675 , \8660 , \8674 );
xor \U$8487 ( \8676 , \8546 , \8675 );
xor \U$8488 ( \8677 , \8537 , \8676 );
and \U$8489 ( \8678 , \8365 , \8366 );
and \U$8490 ( \8679 , \8366 , \8515 );
and \U$8491 ( \8680 , \8365 , \8515 );
or \U$8492 ( \8681 , \8678 , \8679 , \8680 );
nor \U$8493 ( \8682 , \8677 , \8681 );
nor \U$8494 ( \8683 , \8521 , \8682 );
and \U$8495 ( \8684 , \8541 , \8545 );
and \U$8496 ( \8685 , \8545 , \8675 );
and \U$8497 ( \8686 , \8541 , \8675 );
or \U$8498 ( \8687 , \8684 , \8685 , \8686 );
and \U$8499 ( \8688 , \8664 , \8668 );
and \U$8500 ( \8689 , \8668 , \8673 );
and \U$8501 ( \8690 , \8664 , \8673 );
or \U$8502 ( \8691 , \8688 , \8689 , \8690 );
and \U$8503 ( \8692 , \8604 , \8613 );
and \U$8504 ( \8693 , \8613 , \8658 );
and \U$8505 ( \8694 , \8604 , \8658 );
or \U$8506 ( \8695 , \8692 , \8693 , \8694 );
xor \U$8507 ( \8696 , \8691 , \8695 );
and \U$8508 ( \8697 , \8573 , \8584 );
and \U$8509 ( \8698 , \8584 , \8599 );
and \U$8510 ( \8699 , \8573 , \8599 );
or \U$8511 ( \8700 , \8697 , \8698 , \8699 );
xor \U$8512 ( \8701 , \8696 , \8700 );
xor \U$8513 ( \8702 , \8687 , \8701 );
and \U$8514 ( \8703 , \8529 , \8533 );
and \U$8515 ( \8704 , \8533 , \8535 );
and \U$8516 ( \8705 , \8529 , \8535 );
or \U$8517 ( \8706 , \8703 , \8704 , \8705 );
and \U$8518 ( \8707 , \8600 , \8659 );
and \U$8519 ( \8708 , \8659 , \8674 );
and \U$8520 ( \8709 , \8600 , \8674 );
or \U$8521 ( \8710 , \8707 , \8708 , \8709 );
xor \U$8522 ( \8711 , \8706 , \8710 );
and \U$8523 ( \8712 , \8618 , \8622 );
and \U$8524 ( \8713 , \8622 , \8627 );
and \U$8525 ( \8714 , \8618 , \8627 );
or \U$8526 ( \8715 , \8712 , \8713 , \8714 );
and \U$8527 ( \8716 , \8562 , \8566 );
and \U$8528 ( \8717 , \8566 , \8571 );
and \U$8529 ( \8718 , \8562 , \8571 );
or \U$8530 ( \8719 , \8716 , \8717 , \8718 );
xor \U$8531 ( \8720 , \8715 , \8719 );
and \U$8532 ( \8721 , \8550 , \8554 );
and \U$8533 ( \8722 , \8554 , \8557 );
and \U$8534 ( \8723 , \8550 , \8557 );
or \U$8535 ( \8724 , \8721 , \8722 , \8723 );
xor \U$8536 ( \8725 , \8720 , \8724 );
and \U$8537 ( \8726 , \5859 , \8607 );
and \U$8538 ( \8727 , \8607 , \8612 );
and \U$8539 ( \8728 , \5859 , \8612 );
or \U$8540 ( \8729 , \8726 , \8727 , \8728 );
and \U$8541 ( \8730 , \8647 , \8651 );
and \U$8542 ( \8731 , \8651 , \8656 );
and \U$8543 ( \8732 , \8647 , \8656 );
or \U$8544 ( \8733 , \8730 , \8731 , \8732 );
xor \U$8545 ( \8734 , \8729 , \8733 );
and \U$8546 ( \8735 , \8632 , \8636 );
and \U$8547 ( \8736 , \8636 , \8641 );
and \U$8548 ( \8737 , \8632 , \8641 );
or \U$8549 ( \8738 , \8735 , \8736 , \8737 );
xor \U$8550 ( \8739 , \8734 , \8738 );
xor \U$8551 ( \8740 , \8725 , \8739 );
and \U$8552 ( \8741 , \8628 , \8642 );
and \U$8553 ( \8742 , \8642 , \8657 );
and \U$8554 ( \8743 , \8628 , \8657 );
or \U$8555 ( \8744 , \8741 , \8742 , \8743 );
and \U$8556 ( \8745 , \5873 , \7140 );
and \U$8557 ( \8746 , \5842 , \7138 );
nor \U$8558 ( \8747 , \8745 , \8746 );
xnor \U$8559 ( \8748 , \8747 , \7146 );
and \U$8560 ( \8749 , \5893 , \7157 );
and \U$8561 ( \8750 , \5861 , \7155 );
nor \U$8562 ( \8751 , \8749 , \8750 );
xnor \U$8563 ( \8752 , \8751 , \7163 );
xor \U$8564 ( \8753 , \8748 , \8752 );
and \U$8565 ( \8754 , \5918 , \7175 );
and \U$8566 ( \8755 , \5881 , \7173 );
nor \U$8567 ( \8756 , \8754 , \8755 );
xnor \U$8568 ( \8757 , \8756 , \7181 );
xor \U$8569 ( \8758 , \8753 , \8757 );
and \U$8570 ( \8759 , \5811 , \7082 );
and \U$8571 ( \8760 , \5780 , \7080 );
nor \U$8572 ( \8761 , \8759 , \8760 );
xnor \U$8573 ( \8762 , \8761 , \7088 );
and \U$8574 ( \8763 , \5831 , \7099 );
and \U$8575 ( \8764 , \5799 , \7097 );
nor \U$8576 ( \8765 , \8763 , \8764 );
xnor \U$8577 ( \8766 , \8765 , \7105 );
xor \U$8578 ( \8767 , \8762 , \8766 );
and \U$8579 ( \8768 , \5854 , \7117 );
and \U$8580 ( \8769 , \5819 , \7115 );
nor \U$8581 ( \8770 , \8768 , \8769 );
xnor \U$8582 ( \8771 , \8770 , \7123 );
xor \U$8583 ( \8772 , \8767 , \8771 );
xor \U$8584 ( \8773 , \8758 , \8772 );
not \U$8585 ( \8774 , \7032 );
and \U$8586 ( \8775 , \5770 , \7043 );
and \U$8587 ( \8776 , \5737 , \7041 );
nor \U$8588 ( \8777 , \8775 , \8776 );
xnor \U$8589 ( \8778 , \8777 , \7049 );
xor \U$8590 ( \8779 , \8774 , \8778 );
and \U$8591 ( \8780 , \5792 , \7061 );
and \U$8592 ( \8781 , \5758 , \7059 );
nor \U$8593 ( \8782 , \8780 , \8781 );
xnor \U$8594 ( \8783 , \8782 , \7067 );
xor \U$8595 ( \8784 , \8779 , \8783 );
xor \U$8596 ( \8785 , \8773 , \8784 );
xor \U$8597 ( \8786 , \8744 , \8785 );
and \U$8598 ( \8787 , \6057 , \5829 );
and \U$8599 ( \8788 , \6029 , \5827 );
nor \U$8600 ( \8789 , \8787 , \8788 );
xnor \U$8601 ( \8790 , \8789 , \5836 );
and \U$8602 ( \8791 , \6065 , \5852 );
and \U$8603 ( \8792 , \6048 , \5850 );
nor \U$8604 ( \8793 , \8791 , \8792 );
xnor \U$8605 ( \8794 , \8793 , \5859 );
xor \U$8606 ( \8795 , \8790 , \8794 );
and \U$8607 ( \8796 , \5998 , \5768 );
and \U$8608 ( \8797 , \5967 , \5766 );
nor \U$8609 ( \8798 , \8796 , \8797 );
xnor \U$8610 ( \8799 , \8798 , \5775 );
and \U$8611 ( \8800 , \6018 , \5790 );
and \U$8612 ( \8801 , \5986 , \5788 );
nor \U$8613 ( \8802 , \8800 , \8801 );
xnor \U$8614 ( \8803 , \8802 , \5797 );
xor \U$8615 ( \8804 , \8799 , \8803 );
and \U$8616 ( \8805 , \6041 , \5809 );
and \U$8617 ( \8806 , \6006 , \5807 );
nor \U$8618 ( \8807 , \8805 , \8806 );
xnor \U$8619 ( \8808 , \8807 , \5816 );
xor \U$8620 ( \8809 , \8804 , \8808 );
xor \U$8621 ( \8810 , \8795 , \8809 );
and \U$8622 ( \8811 , \5937 , \7192 );
and \U$8623 ( \8812 , \5906 , \7190 );
nor \U$8624 ( \8813 , \8811 , \8812 );
xnor \U$8625 ( \8814 , \8813 , \7198 );
and \U$8626 ( \8815 , \5957 , \7203 );
and \U$8627 ( \8816 , \5925 , \7201 );
nor \U$8628 ( \8817 , \8815 , \8816 );
xnor \U$8629 ( \8818 , \8817 , \6824 );
xor \U$8630 ( \8819 , \8814 , \8818 );
and \U$8631 ( \8820 , \5979 , \5750 );
and \U$8632 ( \8821 , \5945 , \5748 );
nor \U$8633 ( \8822 , \8820 , \8821 );
xnor \U$8634 ( \8823 , \8822 , \5755 );
xor \U$8635 ( \8824 , \8819 , \8823 );
xor \U$8636 ( \8825 , \8810 , \8824 );
xor \U$8637 ( \8826 , \8786 , \8825 );
xor \U$8638 ( \8827 , \8740 , \8826 );
and \U$8639 ( \8828 , \8589 , \8593 );
and \U$8640 ( \8829 , \8593 , \8598 );
and \U$8641 ( \8830 , \8589 , \8598 );
or \U$8642 ( \8831 , \8828 , \8829 , \8830 );
and \U$8643 ( \8832 , \8577 , \8581 );
and \U$8644 ( \8833 , \8581 , \8583 );
and \U$8645 ( \8834 , \8577 , \8583 );
or \U$8646 ( \8835 , \8832 , \8833 , \8834 );
xor \U$8647 ( \8836 , \8831 , \8835 );
or \U$8648 ( \8837 , \8558 , \8572 );
xor \U$8649 ( \8838 , \8836 , \8837 );
xor \U$8650 ( \8839 , \8827 , \8838 );
xor \U$8651 ( \8840 , \8711 , \8839 );
xor \U$8652 ( \8841 , \8702 , \8840 );
and \U$8653 ( \8842 , \8525 , \8536 );
and \U$8654 ( \8843 , \8536 , \8676 );
and \U$8655 ( \8844 , \8525 , \8676 );
or \U$8656 ( \8845 , \8842 , \8843 , \8844 );
nor \U$8657 ( \8846 , \8841 , \8845 );
and \U$8658 ( \8847 , \8706 , \8710 );
and \U$8659 ( \8848 , \8710 , \8839 );
and \U$8660 ( \8849 , \8706 , \8839 );
or \U$8661 ( \8850 , \8847 , \8848 , \8849 );
and \U$8662 ( \8851 , \8831 , \8835 );
and \U$8663 ( \8852 , \8835 , \8837 );
and \U$8664 ( \8853 , \8831 , \8837 );
or \U$8665 ( \8854 , \8851 , \8852 , \8853 );
and \U$8666 ( \8855 , \8744 , \8785 );
and \U$8667 ( \8856 , \8785 , \8825 );
and \U$8668 ( \8857 , \8744 , \8825 );
or \U$8669 ( \8858 , \8855 , \8856 , \8857 );
xor \U$8670 ( \8859 , \8854 , \8858 );
and \U$8671 ( \8860 , \8725 , \8739 );
xor \U$8672 ( \8861 , \8859 , \8860 );
xor \U$8673 ( \8862 , \8850 , \8861 );
and \U$8674 ( \8863 , \8691 , \8695 );
and \U$8675 ( \8864 , \8695 , \8700 );
and \U$8676 ( \8865 , \8691 , \8700 );
or \U$8677 ( \8866 , \8863 , \8864 , \8865 );
and \U$8678 ( \8867 , \8740 , \8826 );
and \U$8679 ( \8868 , \8826 , \8838 );
and \U$8680 ( \8869 , \8740 , \8838 );
or \U$8681 ( \8870 , \8867 , \8868 , \8869 );
xor \U$8682 ( \8871 , \8866 , \8870 );
and \U$8683 ( \8872 , \6029 , \5829 );
and \U$8684 ( \8873 , \6041 , \5827 );
nor \U$8685 ( \8874 , \8872 , \8873 );
xnor \U$8686 ( \8875 , \8874 , \5836 );
and \U$8687 ( \8876 , \6048 , \5852 );
and \U$8688 ( \8877 , \6057 , \5850 );
nor \U$8689 ( \8878 , \8876 , \8877 );
xnor \U$8690 ( \8879 , \8878 , \5859 );
xor \U$8691 ( \8880 , \8875 , \8879 );
nand \U$8692 ( \8881 , \6065 , \5869 );
xnor \U$8693 ( \8882 , \8881 , \5878 );
xor \U$8694 ( \8883 , \8880 , \8882 );
and \U$8695 ( \8884 , \5967 , \5768 );
and \U$8696 ( \8885 , \5979 , \5766 );
nor \U$8697 ( \8886 , \8884 , \8885 );
xnor \U$8698 ( \8887 , \8886 , \5775 );
and \U$8699 ( \8888 , \5986 , \5790 );
and \U$8700 ( \8889 , \5998 , \5788 );
nor \U$8701 ( \8890 , \8888 , \8889 );
xnor \U$8702 ( \8891 , \8890 , \5797 );
xor \U$8703 ( \8892 , \8887 , \8891 );
and \U$8704 ( \8893 , \6006 , \5809 );
and \U$8705 ( \8894 , \6018 , \5807 );
nor \U$8706 ( \8895 , \8893 , \8894 );
xnor \U$8707 ( \8896 , \8895 , \5816 );
xor \U$8708 ( \8897 , \8892 , \8896 );
xnor \U$8709 ( \8898 , \8883 , \8897 );
and \U$8710 ( \8899 , \8814 , \8818 );
and \U$8711 ( \8900 , \8818 , \8823 );
and \U$8712 ( \8901 , \8814 , \8823 );
or \U$8713 ( \8902 , \8899 , \8900 , \8901 );
and \U$8714 ( \8903 , \8799 , \8803 );
and \U$8715 ( \8904 , \8803 , \8808 );
and \U$8716 ( \8905 , \8799 , \8808 );
or \U$8717 ( \8906 , \8903 , \8904 , \8905 );
xor \U$8718 ( \8907 , \8902 , \8906 );
and \U$8719 ( \8908 , \8790 , \8794 );
xor \U$8720 ( \8909 , \8907 , \8908 );
xor \U$8721 ( \8910 , \8898 , \8909 );
and \U$8722 ( \8911 , \8774 , \8778 );
and \U$8723 ( \8912 , \8778 , \8783 );
and \U$8724 ( \8913 , \8774 , \8783 );
or \U$8725 ( \8914 , \8911 , \8912 , \8913 );
and \U$8726 ( \8915 , \8762 , \8766 );
and \U$8727 ( \8916 , \8766 , \8771 );
and \U$8728 ( \8917 , \8762 , \8771 );
or \U$8729 ( \8918 , \8915 , \8916 , \8917 );
xor \U$8730 ( \8919 , \8914 , \8918 );
and \U$8731 ( \8920 , \8748 , \8752 );
and \U$8732 ( \8921 , \8752 , \8757 );
and \U$8733 ( \8922 , \8748 , \8757 );
or \U$8734 ( \8923 , \8920 , \8921 , \8922 );
xor \U$8735 ( \8924 , \8919 , \8923 );
xor \U$8736 ( \8925 , \8910 , \8924 );
and \U$8737 ( \8926 , \8758 , \8772 );
and \U$8738 ( \8927 , \8772 , \8784 );
and \U$8739 ( \8928 , \8758 , \8784 );
or \U$8740 ( \8929 , \8926 , \8927 , \8928 );
and \U$8741 ( \8930 , \5737 , \7043 );
not \U$8742 ( \8931 , \8930 );
xnor \U$8743 ( \8932 , \8931 , \7049 );
xor \U$8744 ( \8933 , \5878 , \8932 );
and \U$8745 ( \8934 , \5758 , \7061 );
and \U$8746 ( \8935 , \5770 , \7059 );
nor \U$8747 ( \8936 , \8934 , \8935 );
xnor \U$8748 ( \8937 , \8936 , \7067 );
xor \U$8749 ( \8938 , \8933 , \8937 );
xor \U$8750 ( \8939 , \8929 , \8938 );
and \U$8751 ( \8940 , \5906 , \7192 );
and \U$8752 ( \8941 , \5918 , \7190 );
nor \U$8753 ( \8942 , \8940 , \8941 );
xnor \U$8754 ( \8943 , \8942 , \7198 );
and \U$8755 ( \8944 , \5925 , \7203 );
and \U$8756 ( \8945 , \5937 , \7201 );
nor \U$8757 ( \8946 , \8944 , \8945 );
xnor \U$8758 ( \8947 , \8946 , \6824 );
xor \U$8759 ( \8948 , \8943 , \8947 );
and \U$8760 ( \8949 , \5945 , \5750 );
and \U$8761 ( \8950 , \5957 , \5748 );
nor \U$8762 ( \8951 , \8949 , \8950 );
xnor \U$8763 ( \8952 , \8951 , \5755 );
xor \U$8764 ( \8953 , \8948 , \8952 );
and \U$8765 ( \8954 , \5842 , \7140 );
and \U$8766 ( \8955 , \5854 , \7138 );
nor \U$8767 ( \8956 , \8954 , \8955 );
xnor \U$8768 ( \8957 , \8956 , \7146 );
and \U$8769 ( \8958 , \5861 , \7157 );
and \U$8770 ( \8959 , \5873 , \7155 );
nor \U$8771 ( \8960 , \8958 , \8959 );
xnor \U$8772 ( \8961 , \8960 , \7163 );
xor \U$8773 ( \8962 , \8957 , \8961 );
and \U$8774 ( \8963 , \5881 , \7175 );
and \U$8775 ( \8964 , \5893 , \7173 );
nor \U$8776 ( \8965 , \8963 , \8964 );
xnor \U$8777 ( \8966 , \8965 , \7181 );
xor \U$8778 ( \8967 , \8962 , \8966 );
xor \U$8779 ( \8968 , \8953 , \8967 );
and \U$8780 ( \8969 , \5780 , \7082 );
and \U$8781 ( \8970 , \5792 , \7080 );
nor \U$8782 ( \8971 , \8969 , \8970 );
xnor \U$8783 ( \8972 , \8971 , \7088 );
and \U$8784 ( \8973 , \5799 , \7099 );
and \U$8785 ( \8974 , \5811 , \7097 );
nor \U$8786 ( \8975 , \8973 , \8974 );
xnor \U$8787 ( \8976 , \8975 , \7105 );
xor \U$8788 ( \8977 , \8972 , \8976 );
and \U$8789 ( \8978 , \5819 , \7117 );
and \U$8790 ( \8979 , \5831 , \7115 );
nor \U$8791 ( \8980 , \8978 , \8979 );
xnor \U$8792 ( \8981 , \8980 , \7123 );
xor \U$8793 ( \8982 , \8977 , \8981 );
xor \U$8794 ( \8983 , \8968 , \8982 );
xor \U$8795 ( \8984 , \8939 , \8983 );
xor \U$8796 ( \8985 , \8925 , \8984 );
and \U$8797 ( \8986 , \8729 , \8733 );
and \U$8798 ( \8987 , \8733 , \8738 );
and \U$8799 ( \8988 , \8729 , \8738 );
or \U$8800 ( \8989 , \8986 , \8987 , \8988 );
and \U$8801 ( \8990 , \8715 , \8719 );
and \U$8802 ( \8991 , \8719 , \8724 );
and \U$8803 ( \8992 , \8715 , \8724 );
or \U$8804 ( \8993 , \8990 , \8991 , \8992 );
xor \U$8805 ( \8994 , \8989 , \8993 );
and \U$8806 ( \8995 , \8795 , \8809 );
and \U$8807 ( \8996 , \8809 , \8824 );
and \U$8808 ( \8997 , \8795 , \8824 );
or \U$8809 ( \8998 , \8995 , \8996 , \8997 );
xor \U$8810 ( \8999 , \8994 , \8998 );
xor \U$8811 ( \9000 , \8985 , \8999 );
xor \U$8812 ( \9001 , \8871 , \9000 );
xor \U$8813 ( \9002 , \8862 , \9001 );
and \U$8814 ( \9003 , \8687 , \8701 );
and \U$8815 ( \9004 , \8701 , \8840 );
and \U$8816 ( \9005 , \8687 , \8840 );
or \U$8817 ( \9006 , \9003 , \9004 , \9005 );
nor \U$8818 ( \9007 , \9002 , \9006 );
nor \U$8819 ( \9008 , \8846 , \9007 );
nand \U$8820 ( \9009 , \8683 , \9008 );
nor \U$8821 ( \9010 , \8361 , \9009 );
and \U$8822 ( \9011 , \8866 , \8870 );
and \U$8823 ( \9012 , \8870 , \9000 );
and \U$8824 ( \9013 , \8866 , \9000 );
or \U$8825 ( \9014 , \9011 , \9012 , \9013 );
and \U$8826 ( \9015 , \8989 , \8993 );
and \U$8827 ( \9016 , \8993 , \8998 );
and \U$8828 ( \9017 , \8989 , \8998 );
or \U$8829 ( \9018 , \9015 , \9016 , \9017 );
and \U$8830 ( \9019 , \8929 , \8938 );
and \U$8831 ( \9020 , \8938 , \8983 );
and \U$8832 ( \9021 , \8929 , \8983 );
or \U$8833 ( \9022 , \9019 , \9020 , \9021 );
xor \U$8834 ( \9023 , \9018 , \9022 );
and \U$8835 ( \9024 , \8898 , \8909 );
and \U$8836 ( \9025 , \8909 , \8924 );
and \U$8837 ( \9026 , \8898 , \8924 );
or \U$8838 ( \9027 , \9024 , \9025 , \9026 );
xor \U$8839 ( \9028 , \9023 , \9027 );
xor \U$8840 ( \9029 , \9014 , \9028 );
and \U$8841 ( \9030 , \8854 , \8858 );
and \U$8842 ( \9031 , \8858 , \8860 );
and \U$8843 ( \9032 , \8854 , \8860 );
or \U$8844 ( \9033 , \9030 , \9031 , \9032 );
and \U$8845 ( \9034 , \8925 , \8984 );
and \U$8846 ( \9035 , \8984 , \8999 );
and \U$8847 ( \9036 , \8925 , \8999 );
or \U$8848 ( \9037 , \9034 , \9035 , \9036 );
xor \U$8849 ( \9038 , \9033 , \9037 );
and \U$8850 ( \9039 , \8943 , \8947 );
and \U$8851 ( \9040 , \8947 , \8952 );
and \U$8852 ( \9041 , \8943 , \8952 );
or \U$8853 ( \9042 , \9039 , \9040 , \9041 );
and \U$8854 ( \9043 , \8887 , \8891 );
and \U$8855 ( \9044 , \8891 , \8896 );
and \U$8856 ( \9045 , \8887 , \8896 );
or \U$8857 ( \9046 , \9043 , \9044 , \9045 );
xor \U$8858 ( \9047 , \9042 , \9046 );
and \U$8859 ( \9048 , \8875 , \8879 );
and \U$8860 ( \9049 , \8879 , \8882 );
and \U$8861 ( \9050 , \8875 , \8882 );
or \U$8862 ( \9051 , \9048 , \9049 , \9050 );
xor \U$8863 ( \9052 , \9047 , \9051 );
and \U$8864 ( \9053 , \5878 , \8932 );
and \U$8865 ( \9054 , \8932 , \8937 );
and \U$8866 ( \9055 , \5878 , \8937 );
or \U$8867 ( \9056 , \9053 , \9054 , \9055 );
and \U$8868 ( \9057 , \8972 , \8976 );
and \U$8869 ( \9058 , \8976 , \8981 );
and \U$8870 ( \9059 , \8972 , \8981 );
or \U$8871 ( \9060 , \9057 , \9058 , \9059 );
xor \U$8872 ( \9061 , \9056 , \9060 );
and \U$8873 ( \9062 , \8957 , \8961 );
and \U$8874 ( \9063 , \8961 , \8966 );
and \U$8875 ( \9064 , \8957 , \8966 );
or \U$8876 ( \9065 , \9062 , \9063 , \9064 );
xor \U$8877 ( \9066 , \9061 , \9065 );
xor \U$8878 ( \9067 , \9052 , \9066 );
and \U$8879 ( \9068 , \8953 , \8967 );
and \U$8880 ( \9069 , \8967 , \8982 );
and \U$8881 ( \9070 , \8953 , \8982 );
or \U$8882 ( \9071 , \9068 , \9069 , \9070 );
and \U$8883 ( \9072 , \5873 , \7157 );
and \U$8884 ( \9073 , \5842 , \7155 );
nor \U$8885 ( \9074 , \9072 , \9073 );
xnor \U$8886 ( \9075 , \9074 , \7163 );
and \U$8887 ( \9076 , \5893 , \7175 );
and \U$8888 ( \9077 , \5861 , \7173 );
nor \U$8889 ( \9078 , \9076 , \9077 );
xnor \U$8890 ( \9079 , \9078 , \7181 );
xor \U$8891 ( \9080 , \9075 , \9079 );
and \U$8892 ( \9081 , \5918 , \7192 );
and \U$8893 ( \9082 , \5881 , \7190 );
nor \U$8894 ( \9083 , \9081 , \9082 );
xnor \U$8895 ( \9084 , \9083 , \7198 );
xor \U$8896 ( \9085 , \9080 , \9084 );
and \U$8897 ( \9086 , \5811 , \7099 );
and \U$8898 ( \9087 , \5780 , \7097 );
nor \U$8899 ( \9088 , \9086 , \9087 );
xnor \U$8900 ( \9089 , \9088 , \7105 );
and \U$8901 ( \9090 , \5831 , \7117 );
and \U$8902 ( \9091 , \5799 , \7115 );
nor \U$8903 ( \9092 , \9090 , \9091 );
xnor \U$8904 ( \9093 , \9092 , \7123 );
xor \U$8905 ( \9094 , \9089 , \9093 );
and \U$8906 ( \9095 , \5854 , \7140 );
and \U$8907 ( \9096 , \5819 , \7138 );
nor \U$8908 ( \9097 , \9095 , \9096 );
xnor \U$8909 ( \9098 , \9097 , \7146 );
xor \U$8910 ( \9099 , \9094 , \9098 );
xor \U$8911 ( \9100 , \9085 , \9099 );
not \U$8912 ( \9101 , \7049 );
and \U$8913 ( \9102 , \5770 , \7061 );
and \U$8914 ( \9103 , \5737 , \7059 );
nor \U$8915 ( \9104 , \9102 , \9103 );
xnor \U$8916 ( \9105 , \9104 , \7067 );
xor \U$8917 ( \9106 , \9101 , \9105 );
and \U$8918 ( \9107 , \5792 , \7082 );
and \U$8919 ( \9108 , \5758 , \7080 );
nor \U$8920 ( \9109 , \9107 , \9108 );
xnor \U$8921 ( \9110 , \9109 , \7088 );
xor \U$8922 ( \9111 , \9106 , \9110 );
xor \U$8923 ( \9112 , \9100 , \9111 );
xor \U$8924 ( \9113 , \9071 , \9112 );
and \U$8925 ( \9114 , \6057 , \5852 );
and \U$8926 ( \9115 , \6029 , \5850 );
nor \U$8927 ( \9116 , \9114 , \9115 );
xnor \U$8928 ( \9117 , \9116 , \5859 );
and \U$8929 ( \9118 , \6065 , \5871 );
and \U$8930 ( \9119 , \6048 , \5869 );
nor \U$8931 ( \9120 , \9118 , \9119 );
xnor \U$8932 ( \9121 , \9120 , \5878 );
xor \U$8933 ( \9122 , \9117 , \9121 );
and \U$8934 ( \9123 , \5998 , \5790 );
and \U$8935 ( \9124 , \5967 , \5788 );
nor \U$8936 ( \9125 , \9123 , \9124 );
xnor \U$8937 ( \9126 , \9125 , \5797 );
and \U$8938 ( \9127 , \6018 , \5809 );
and \U$8939 ( \9128 , \5986 , \5807 );
nor \U$8940 ( \9129 , \9127 , \9128 );
xnor \U$8941 ( \9130 , \9129 , \5816 );
xor \U$8942 ( \9131 , \9126 , \9130 );
and \U$8943 ( \9132 , \6041 , \5829 );
and \U$8944 ( \9133 , \6006 , \5827 );
nor \U$8945 ( \9134 , \9132 , \9133 );
xnor \U$8946 ( \9135 , \9134 , \5836 );
xor \U$8947 ( \9136 , \9131 , \9135 );
xor \U$8948 ( \9137 , \9122 , \9136 );
and \U$8949 ( \9138 , \5937 , \7203 );
and \U$8950 ( \9139 , \5906 , \7201 );
nor \U$8951 ( \9140 , \9138 , \9139 );
xnor \U$8952 ( \9141 , \9140 , \6824 );
and \U$8953 ( \9142 , \5957 , \5750 );
and \U$8954 ( \9143 , \5925 , \5748 );
nor \U$8955 ( \9144 , \9142 , \9143 );
xnor \U$8956 ( \9145 , \9144 , \5755 );
xor \U$8957 ( \9146 , \9141 , \9145 );
and \U$8958 ( \9147 , \5979 , \5768 );
and \U$8959 ( \9148 , \5945 , \5766 );
nor \U$8960 ( \9149 , \9147 , \9148 );
xnor \U$8961 ( \9150 , \9149 , \5775 );
xor \U$8962 ( \9151 , \9146 , \9150 );
xor \U$8963 ( \9152 , \9137 , \9151 );
xor \U$8964 ( \9153 , \9113 , \9152 );
xor \U$8965 ( \9154 , \9067 , \9153 );
and \U$8966 ( \9155 , \8914 , \8918 );
and \U$8967 ( \9156 , \8918 , \8923 );
and \U$8968 ( \9157 , \8914 , \8923 );
or \U$8969 ( \9158 , \9155 , \9156 , \9157 );
and \U$8970 ( \9159 , \8902 , \8906 );
and \U$8971 ( \9160 , \8906 , \8908 );
and \U$8972 ( \9161 , \8902 , \8908 );
or \U$8973 ( \9162 , \9159 , \9160 , \9161 );
xor \U$8974 ( \9163 , \9158 , \9162 );
or \U$8975 ( \9164 , \8883 , \8897 );
xor \U$8976 ( \9165 , \9163 , \9164 );
xor \U$8977 ( \9166 , \9154 , \9165 );
xor \U$8978 ( \9167 , \9038 , \9166 );
xor \U$8979 ( \9168 , \9029 , \9167 );
and \U$8980 ( \9169 , \8850 , \8861 );
and \U$8981 ( \9170 , \8861 , \9001 );
and \U$8982 ( \9171 , \8850 , \9001 );
or \U$8983 ( \9172 , \9169 , \9170 , \9171 );
nor \U$8984 ( \9173 , \9168 , \9172 );
and \U$8985 ( \9174 , \9033 , \9037 );
and \U$8986 ( \9175 , \9037 , \9166 );
and \U$8987 ( \9176 , \9033 , \9166 );
or \U$8988 ( \9177 , \9174 , \9175 , \9176 );
and \U$8989 ( \9178 , \9158 , \9162 );
and \U$8990 ( \9179 , \9162 , \9164 );
and \U$8991 ( \9180 , \9158 , \9164 );
or \U$8992 ( \9181 , \9178 , \9179 , \9180 );
and \U$8993 ( \9182 , \9071 , \9112 );
and \U$8994 ( \9183 , \9112 , \9152 );
and \U$8995 ( \9184 , \9071 , \9152 );
or \U$8996 ( \9185 , \9182 , \9183 , \9184 );
xor \U$8997 ( \9186 , \9181 , \9185 );
and \U$8998 ( \9187 , \9052 , \9066 );
xor \U$8999 ( \9188 , \9186 , \9187 );
xor \U$9000 ( \9189 , \9177 , \9188 );
and \U$9001 ( \9190 , \9018 , \9022 );
and \U$9002 ( \9191 , \9022 , \9027 );
and \U$9003 ( \9192 , \9018 , \9027 );
or \U$9004 ( \9193 , \9190 , \9191 , \9192 );
and \U$9005 ( \9194 , \9067 , \9153 );
and \U$9006 ( \9195 , \9153 , \9165 );
and \U$9007 ( \9196 , \9067 , \9165 );
or \U$9008 ( \9197 , \9194 , \9195 , \9196 );
xor \U$9009 ( \9198 , \9193 , \9197 );
and \U$9010 ( \9199 , \6029 , \5852 );
and \U$9011 ( \9200 , \6041 , \5850 );
nor \U$9012 ( \9201 , \9199 , \9200 );
xnor \U$9013 ( \9202 , \9201 , \5859 );
and \U$9014 ( \9203 , \6048 , \5871 );
and \U$9015 ( \9204 , \6057 , \5869 );
nor \U$9016 ( \9205 , \9203 , \9204 );
xnor \U$9017 ( \9206 , \9205 , \5878 );
xor \U$9018 ( \9207 , \9202 , \9206 );
nand \U$9019 ( \9208 , \6065 , \5889 );
xnor \U$9020 ( \9209 , \9208 , \5898 );
xor \U$9021 ( \9210 , \9207 , \9209 );
and \U$9022 ( \9211 , \5967 , \5790 );
and \U$9023 ( \9212 , \5979 , \5788 );
nor \U$9024 ( \9213 , \9211 , \9212 );
xnor \U$9025 ( \9214 , \9213 , \5797 );
and \U$9026 ( \9215 , \5986 , \5809 );
and \U$9027 ( \9216 , \5998 , \5807 );
nor \U$9028 ( \9217 , \9215 , \9216 );
xnor \U$9029 ( \9218 , \9217 , \5816 );
xor \U$9030 ( \9219 , \9214 , \9218 );
and \U$9031 ( \9220 , \6006 , \5829 );
and \U$9032 ( \9221 , \6018 , \5827 );
nor \U$9033 ( \9222 , \9220 , \9221 );
xnor \U$9034 ( \9223 , \9222 , \5836 );
xor \U$9035 ( \9224 , \9219 , \9223 );
xnor \U$9036 ( \9225 , \9210 , \9224 );
and \U$9037 ( \9226 , \9141 , \9145 );
and \U$9038 ( \9227 , \9145 , \9150 );
and \U$9039 ( \9228 , \9141 , \9150 );
or \U$9040 ( \9229 , \9226 , \9227 , \9228 );
and \U$9041 ( \9230 , \9126 , \9130 );
and \U$9042 ( \9231 , \9130 , \9135 );
and \U$9043 ( \9232 , \9126 , \9135 );
or \U$9044 ( \9233 , \9230 , \9231 , \9232 );
xor \U$9045 ( \9234 , \9229 , \9233 );
and \U$9046 ( \9235 , \9117 , \9121 );
xor \U$9047 ( \9236 , \9234 , \9235 );
xor \U$9048 ( \9237 , \9225 , \9236 );
and \U$9049 ( \9238 , \9101 , \9105 );
and \U$9050 ( \9239 , \9105 , \9110 );
and \U$9051 ( \9240 , \9101 , \9110 );
or \U$9052 ( \9241 , \9238 , \9239 , \9240 );
and \U$9053 ( \9242 , \9089 , \9093 );
and \U$9054 ( \9243 , \9093 , \9098 );
and \U$9055 ( \9244 , \9089 , \9098 );
or \U$9056 ( \9245 , \9242 , \9243 , \9244 );
xor \U$9057 ( \9246 , \9241 , \9245 );
and \U$9058 ( \9247 , \9075 , \9079 );
and \U$9059 ( \9248 , \9079 , \9084 );
and \U$9060 ( \9249 , \9075 , \9084 );
or \U$9061 ( \9250 , \9247 , \9248 , \9249 );
xor \U$9062 ( \9251 , \9246 , \9250 );
xor \U$9063 ( \9252 , \9237 , \9251 );
and \U$9064 ( \9253 , \9085 , \9099 );
and \U$9065 ( \9254 , \9099 , \9111 );
and \U$9066 ( \9255 , \9085 , \9111 );
or \U$9067 ( \9256 , \9253 , \9254 , \9255 );
and \U$9068 ( \9257 , \5737 , \7061 );
not \U$9069 ( \9258 , \9257 );
xnor \U$9070 ( \9259 , \9258 , \7067 );
xor \U$9071 ( \9260 , \5898 , \9259 );
and \U$9072 ( \9261 , \5758 , \7082 );
and \U$9073 ( \9262 , \5770 , \7080 );
nor \U$9074 ( \9263 , \9261 , \9262 );
xnor \U$9075 ( \9264 , \9263 , \7088 );
xor \U$9076 ( \9265 , \9260 , \9264 );
xor \U$9077 ( \9266 , \9256 , \9265 );
and \U$9078 ( \9267 , \5906 , \7203 );
and \U$9079 ( \9268 , \5918 , \7201 );
nor \U$9080 ( \9269 , \9267 , \9268 );
xnor \U$9081 ( \9270 , \9269 , \6824 );
and \U$9082 ( \9271 , \5925 , \5750 );
and \U$9083 ( \9272 , \5937 , \5748 );
nor \U$9084 ( \9273 , \9271 , \9272 );
xnor \U$9085 ( \9274 , \9273 , \5755 );
xor \U$9086 ( \9275 , \9270 , \9274 );
and \U$9087 ( \9276 , \5945 , \5768 );
and \U$9088 ( \9277 , \5957 , \5766 );
nor \U$9089 ( \9278 , \9276 , \9277 );
xnor \U$9090 ( \9279 , \9278 , \5775 );
xor \U$9091 ( \9280 , \9275 , \9279 );
and \U$9092 ( \9281 , \5842 , \7157 );
and \U$9093 ( \9282 , \5854 , \7155 );
nor \U$9094 ( \9283 , \9281 , \9282 );
xnor \U$9095 ( \9284 , \9283 , \7163 );
and \U$9096 ( \9285 , \5861 , \7175 );
and \U$9097 ( \9286 , \5873 , \7173 );
nor \U$9098 ( \9287 , \9285 , \9286 );
xnor \U$9099 ( \9288 , \9287 , \7181 );
xor \U$9100 ( \9289 , \9284 , \9288 );
and \U$9101 ( \9290 , \5881 , \7192 );
and \U$9102 ( \9291 , \5893 , \7190 );
nor \U$9103 ( \9292 , \9290 , \9291 );
xnor \U$9104 ( \9293 , \9292 , \7198 );
xor \U$9105 ( \9294 , \9289 , \9293 );
xor \U$9106 ( \9295 , \9280 , \9294 );
and \U$9107 ( \9296 , \5780 , \7099 );
and \U$9108 ( \9297 , \5792 , \7097 );
nor \U$9109 ( \9298 , \9296 , \9297 );
xnor \U$9110 ( \9299 , \9298 , \7105 );
and \U$9111 ( \9300 , \5799 , \7117 );
and \U$9112 ( \9301 , \5811 , \7115 );
nor \U$9113 ( \9302 , \9300 , \9301 );
xnor \U$9114 ( \9303 , \9302 , \7123 );
xor \U$9115 ( \9304 , \9299 , \9303 );
and \U$9116 ( \9305 , \5819 , \7140 );
and \U$9117 ( \9306 , \5831 , \7138 );
nor \U$9118 ( \9307 , \9305 , \9306 );
xnor \U$9119 ( \9308 , \9307 , \7146 );
xor \U$9120 ( \9309 , \9304 , \9308 );
xor \U$9121 ( \9310 , \9295 , \9309 );
xor \U$9122 ( \9311 , \9266 , \9310 );
xor \U$9123 ( \9312 , \9252 , \9311 );
and \U$9124 ( \9313 , \9056 , \9060 );
and \U$9125 ( \9314 , \9060 , \9065 );
and \U$9126 ( \9315 , \9056 , \9065 );
or \U$9127 ( \9316 , \9313 , \9314 , \9315 );
and \U$9128 ( \9317 , \9042 , \9046 );
and \U$9129 ( \9318 , \9046 , \9051 );
and \U$9130 ( \9319 , \9042 , \9051 );
or \U$9131 ( \9320 , \9317 , \9318 , \9319 );
xor \U$9132 ( \9321 , \9316 , \9320 );
and \U$9133 ( \9322 , \9122 , \9136 );
and \U$9134 ( \9323 , \9136 , \9151 );
and \U$9135 ( \9324 , \9122 , \9151 );
or \U$9136 ( \9325 , \9322 , \9323 , \9324 );
xor \U$9137 ( \9326 , \9321 , \9325 );
xor \U$9138 ( \9327 , \9312 , \9326 );
xor \U$9139 ( \9328 , \9198 , \9327 );
xor \U$9140 ( \9329 , \9189 , \9328 );
and \U$9141 ( \9330 , \9014 , \9028 );
and \U$9142 ( \9331 , \9028 , \9167 );
and \U$9143 ( \9332 , \9014 , \9167 );
or \U$9144 ( \9333 , \9330 , \9331 , \9332 );
nor \U$9145 ( \9334 , \9329 , \9333 );
nor \U$9146 ( \9335 , \9173 , \9334 );
and \U$9147 ( \9336 , \9193 , \9197 );
and \U$9148 ( \9337 , \9197 , \9327 );
and \U$9149 ( \9338 , \9193 , \9327 );
or \U$9150 ( \9339 , \9336 , \9337 , \9338 );
and \U$9151 ( \9340 , \9316 , \9320 );
and \U$9152 ( \9341 , \9320 , \9325 );
and \U$9153 ( \9342 , \9316 , \9325 );
or \U$9154 ( \9343 , \9340 , \9341 , \9342 );
and \U$9155 ( \9344 , \9256 , \9265 );
and \U$9156 ( \9345 , \9265 , \9310 );
and \U$9157 ( \9346 , \9256 , \9310 );
or \U$9158 ( \9347 , \9344 , \9345 , \9346 );
xor \U$9159 ( \9348 , \9343 , \9347 );
and \U$9160 ( \9349 , \9225 , \9236 );
and \U$9161 ( \9350 , \9236 , \9251 );
and \U$9162 ( \9351 , \9225 , \9251 );
or \U$9163 ( \9352 , \9349 , \9350 , \9351 );
xor \U$9164 ( \9353 , \9348 , \9352 );
xor \U$9165 ( \9354 , \9339 , \9353 );
and \U$9166 ( \9355 , \9181 , \9185 );
and \U$9167 ( \9356 , \9185 , \9187 );
and \U$9168 ( \9357 , \9181 , \9187 );
or \U$9169 ( \9358 , \9355 , \9356 , \9357 );
and \U$9170 ( \9359 , \9252 , \9311 );
and \U$9171 ( \9360 , \9311 , \9326 );
and \U$9172 ( \9361 , \9252 , \9326 );
or \U$9173 ( \9362 , \9359 , \9360 , \9361 );
xor \U$9174 ( \9363 , \9358 , \9362 );
and \U$9175 ( \9364 , \9270 , \9274 );
and \U$9176 ( \9365 , \9274 , \9279 );
and \U$9177 ( \9366 , \9270 , \9279 );
or \U$9178 ( \9367 , \9364 , \9365 , \9366 );
and \U$9179 ( \9368 , \9214 , \9218 );
and \U$9180 ( \9369 , \9218 , \9223 );
and \U$9181 ( \9370 , \9214 , \9223 );
or \U$9182 ( \9371 , \9368 , \9369 , \9370 );
xor \U$9183 ( \9372 , \9367 , \9371 );
and \U$9184 ( \9373 , \9202 , \9206 );
and \U$9185 ( \9374 , \9206 , \9209 );
and \U$9186 ( \9375 , \9202 , \9209 );
or \U$9187 ( \9376 , \9373 , \9374 , \9375 );
xor \U$9188 ( \9377 , \9372 , \9376 );
and \U$9189 ( \9378 , \5898 , \9259 );
and \U$9190 ( \9379 , \9259 , \9264 );
and \U$9191 ( \9380 , \5898 , \9264 );
or \U$9192 ( \9381 , \9378 , \9379 , \9380 );
and \U$9193 ( \9382 , \9299 , \9303 );
and \U$9194 ( \9383 , \9303 , \9308 );
and \U$9195 ( \9384 , \9299 , \9308 );
or \U$9196 ( \9385 , \9382 , \9383 , \9384 );
xor \U$9197 ( \9386 , \9381 , \9385 );
and \U$9198 ( \9387 , \9284 , \9288 );
and \U$9199 ( \9388 , \9288 , \9293 );
and \U$9200 ( \9389 , \9284 , \9293 );
or \U$9201 ( \9390 , \9387 , \9388 , \9389 );
xor \U$9202 ( \9391 , \9386 , \9390 );
xor \U$9203 ( \9392 , \9377 , \9391 );
and \U$9204 ( \9393 , \9280 , \9294 );
and \U$9205 ( \9394 , \9294 , \9309 );
and \U$9206 ( \9395 , \9280 , \9309 );
or \U$9207 ( \9396 , \9393 , \9394 , \9395 );
and \U$9208 ( \9397 , \5873 , \7175 );
and \U$9209 ( \9398 , \5842 , \7173 );
nor \U$9210 ( \9399 , \9397 , \9398 );
xnor \U$9211 ( \9400 , \9399 , \7181 );
and \U$9212 ( \9401 , \5893 , \7192 );
and \U$9213 ( \9402 , \5861 , \7190 );
nor \U$9214 ( \9403 , \9401 , \9402 );
xnor \U$9215 ( \9404 , \9403 , \7198 );
xor \U$9216 ( \9405 , \9400 , \9404 );
and \U$9217 ( \9406 , \5918 , \7203 );
and \U$9218 ( \9407 , \5881 , \7201 );
nor \U$9219 ( \9408 , \9406 , \9407 );
xnor \U$9220 ( \9409 , \9408 , \6824 );
xor \U$9221 ( \9410 , \9405 , \9409 );
and \U$9222 ( \9411 , \5811 , \7117 );
and \U$9223 ( \9412 , \5780 , \7115 );
nor \U$9224 ( \9413 , \9411 , \9412 );
xnor \U$9225 ( \9414 , \9413 , \7123 );
and \U$9226 ( \9415 , \5831 , \7140 );
and \U$9227 ( \9416 , \5799 , \7138 );
nor \U$9228 ( \9417 , \9415 , \9416 );
xnor \U$9229 ( \9418 , \9417 , \7146 );
xor \U$9230 ( \9419 , \9414 , \9418 );
and \U$9231 ( \9420 , \5854 , \7157 );
and \U$9232 ( \9421 , \5819 , \7155 );
nor \U$9233 ( \9422 , \9420 , \9421 );
xnor \U$9234 ( \9423 , \9422 , \7163 );
xor \U$9235 ( \9424 , \9419 , \9423 );
xor \U$9236 ( \9425 , \9410 , \9424 );
not \U$9237 ( \9426 , \7067 );
and \U$9238 ( \9427 , \5770 , \7082 );
and \U$9239 ( \9428 , \5737 , \7080 );
nor \U$9240 ( \9429 , \9427 , \9428 );
xnor \U$9241 ( \9430 , \9429 , \7088 );
xor \U$9242 ( \9431 , \9426 , \9430 );
and \U$9243 ( \9432 , \5792 , \7099 );
and \U$9244 ( \9433 , \5758 , \7097 );
nor \U$9245 ( \9434 , \9432 , \9433 );
xnor \U$9246 ( \9435 , \9434 , \7105 );
xor \U$9247 ( \9436 , \9431 , \9435 );
xor \U$9248 ( \9437 , \9425 , \9436 );
xor \U$9249 ( \9438 , \9396 , \9437 );
and \U$9250 ( \9439 , \6057 , \5871 );
and \U$9251 ( \9440 , \6029 , \5869 );
nor \U$9252 ( \9441 , \9439 , \9440 );
xnor \U$9253 ( \9442 , \9441 , \5878 );
and \U$9254 ( \9443 , \6065 , \5891 );
and \U$9255 ( \9444 , \6048 , \5889 );
nor \U$9256 ( \9445 , \9443 , \9444 );
xnor \U$9257 ( \9446 , \9445 , \5898 );
xor \U$9258 ( \9447 , \9442 , \9446 );
and \U$9259 ( \9448 , \5998 , \5809 );
and \U$9260 ( \9449 , \5967 , \5807 );
nor \U$9261 ( \9450 , \9448 , \9449 );
xnor \U$9262 ( \9451 , \9450 , \5816 );
and \U$9263 ( \9452 , \6018 , \5829 );
and \U$9264 ( \9453 , \5986 , \5827 );
nor \U$9265 ( \9454 , \9452 , \9453 );
xnor \U$9266 ( \9455 , \9454 , \5836 );
xor \U$9267 ( \9456 , \9451 , \9455 );
and \U$9268 ( \9457 , \6041 , \5852 );
and \U$9269 ( \9458 , \6006 , \5850 );
nor \U$9270 ( \9459 , \9457 , \9458 );
xnor \U$9271 ( \9460 , \9459 , \5859 );
xor \U$9272 ( \9461 , \9456 , \9460 );
xor \U$9273 ( \9462 , \9447 , \9461 );
and \U$9274 ( \9463 , \5937 , \5750 );
and \U$9275 ( \9464 , \5906 , \5748 );
nor \U$9276 ( \9465 , \9463 , \9464 );
xnor \U$9277 ( \9466 , \9465 , \5755 );
and \U$9278 ( \9467 , \5957 , \5768 );
and \U$9279 ( \9468 , \5925 , \5766 );
nor \U$9280 ( \9469 , \9467 , \9468 );
xnor \U$9281 ( \9470 , \9469 , \5775 );
xor \U$9282 ( \9471 , \9466 , \9470 );
and \U$9283 ( \9472 , \5979 , \5790 );
and \U$9284 ( \9473 , \5945 , \5788 );
nor \U$9285 ( \9474 , \9472 , \9473 );
xnor \U$9286 ( \9475 , \9474 , \5797 );
xor \U$9287 ( \9476 , \9471 , \9475 );
xor \U$9288 ( \9477 , \9462 , \9476 );
xor \U$9289 ( \9478 , \9438 , \9477 );
xor \U$9290 ( \9479 , \9392 , \9478 );
and \U$9291 ( \9480 , \9241 , \9245 );
and \U$9292 ( \9481 , \9245 , \9250 );
and \U$9293 ( \9482 , \9241 , \9250 );
or \U$9294 ( \9483 , \9480 , \9481 , \9482 );
and \U$9295 ( \9484 , \9229 , \9233 );
and \U$9296 ( \9485 , \9233 , \9235 );
and \U$9297 ( \9486 , \9229 , \9235 );
or \U$9298 ( \9487 , \9484 , \9485 , \9486 );
xor \U$9299 ( \9488 , \9483 , \9487 );
or \U$9300 ( \9489 , \9210 , \9224 );
xor \U$9301 ( \9490 , \9488 , \9489 );
xor \U$9302 ( \9491 , \9479 , \9490 );
xor \U$9303 ( \9492 , \9363 , \9491 );
xor \U$9304 ( \9493 , \9354 , \9492 );
and \U$9305 ( \9494 , \9177 , \9188 );
and \U$9306 ( \9495 , \9188 , \9328 );
and \U$9307 ( \9496 , \9177 , \9328 );
or \U$9308 ( \9497 , \9494 , \9495 , \9496 );
nor \U$9309 ( \9498 , \9493 , \9497 );
and \U$9310 ( \9499 , \9358 , \9362 );
and \U$9311 ( \9500 , \9362 , \9491 );
and \U$9312 ( \9501 , \9358 , \9491 );
or \U$9313 ( \9502 , \9499 , \9500 , \9501 );
and \U$9314 ( \9503 , \9483 , \9487 );
and \U$9315 ( \9504 , \9487 , \9489 );
and \U$9316 ( \9505 , \9483 , \9489 );
or \U$9317 ( \9506 , \9503 , \9504 , \9505 );
and \U$9318 ( \9507 , \9396 , \9437 );
and \U$9319 ( \9508 , \9437 , \9477 );
and \U$9320 ( \9509 , \9396 , \9477 );
or \U$9321 ( \9510 , \9507 , \9508 , \9509 );
xor \U$9322 ( \9511 , \9506 , \9510 );
and \U$9323 ( \9512 , \9377 , \9391 );
xor \U$9324 ( \9513 , \9511 , \9512 );
xor \U$9325 ( \9514 , \9502 , \9513 );
and \U$9326 ( \9515 , \9343 , \9347 );
and \U$9327 ( \9516 , \9347 , \9352 );
and \U$9328 ( \9517 , \9343 , \9352 );
or \U$9329 ( \9518 , \9515 , \9516 , \9517 );
and \U$9330 ( \9519 , \9392 , \9478 );
and \U$9331 ( \9520 , \9478 , \9490 );
and \U$9332 ( \9521 , \9392 , \9490 );
or \U$9333 ( \9522 , \9519 , \9520 , \9521 );
xor \U$9334 ( \9523 , \9518 , \9522 );
and \U$9335 ( \9524 , \6029 , \5871 );
and \U$9336 ( \9525 , \6041 , \5869 );
nor \U$9337 ( \9526 , \9524 , \9525 );
xnor \U$9338 ( \9527 , \9526 , \5878 );
and \U$9339 ( \9528 , \6048 , \5891 );
and \U$9340 ( \9529 , \6057 , \5889 );
nor \U$9341 ( \9530 , \9528 , \9529 );
xnor \U$9342 ( \9531 , \9530 , \5898 );
xor \U$9343 ( \9532 , \9527 , \9531 );
nand \U$9344 ( \9533 , \6065 , \5914 );
xnor \U$9345 ( \9534 , \9533 , \5923 );
xor \U$9346 ( \9535 , \9532 , \9534 );
and \U$9347 ( \9536 , \5967 , \5809 );
and \U$9348 ( \9537 , \5979 , \5807 );
nor \U$9349 ( \9538 , \9536 , \9537 );
xnor \U$9350 ( \9539 , \9538 , \5816 );
and \U$9351 ( \9540 , \5986 , \5829 );
and \U$9352 ( \9541 , \5998 , \5827 );
nor \U$9353 ( \9542 , \9540 , \9541 );
xnor \U$9354 ( \9543 , \9542 , \5836 );
xor \U$9355 ( \9544 , \9539 , \9543 );
and \U$9356 ( \9545 , \6006 , \5852 );
and \U$9357 ( \9546 , \6018 , \5850 );
nor \U$9358 ( \9547 , \9545 , \9546 );
xnor \U$9359 ( \9548 , \9547 , \5859 );
xor \U$9360 ( \9549 , \9544 , \9548 );
xnor \U$9361 ( \9550 , \9535 , \9549 );
and \U$9362 ( \9551 , \9466 , \9470 );
and \U$9363 ( \9552 , \9470 , \9475 );
and \U$9364 ( \9553 , \9466 , \9475 );
or \U$9365 ( \9554 , \9551 , \9552 , \9553 );
and \U$9366 ( \9555 , \9451 , \9455 );
and \U$9367 ( \9556 , \9455 , \9460 );
and \U$9368 ( \9557 , \9451 , \9460 );
or \U$9369 ( \9558 , \9555 , \9556 , \9557 );
xor \U$9370 ( \9559 , \9554 , \9558 );
and \U$9371 ( \9560 , \9442 , \9446 );
xor \U$9372 ( \9561 , \9559 , \9560 );
xor \U$9373 ( \9562 , \9550 , \9561 );
and \U$9374 ( \9563 , \9426 , \9430 );
and \U$9375 ( \9564 , \9430 , \9435 );
and \U$9376 ( \9565 , \9426 , \9435 );
or \U$9377 ( \9566 , \9563 , \9564 , \9565 );
and \U$9378 ( \9567 , \9414 , \9418 );
and \U$9379 ( \9568 , \9418 , \9423 );
and \U$9380 ( \9569 , \9414 , \9423 );
or \U$9381 ( \9570 , \9567 , \9568 , \9569 );
xor \U$9382 ( \9571 , \9566 , \9570 );
and \U$9383 ( \9572 , \9400 , \9404 );
and \U$9384 ( \9573 , \9404 , \9409 );
and \U$9385 ( \9574 , \9400 , \9409 );
or \U$9386 ( \9575 , \9572 , \9573 , \9574 );
xor \U$9387 ( \9576 , \9571 , \9575 );
xor \U$9388 ( \9577 , \9562 , \9576 );
and \U$9389 ( \9578 , \9410 , \9424 );
and \U$9390 ( \9579 , \9424 , \9436 );
and \U$9391 ( \9580 , \9410 , \9436 );
or \U$9392 ( \9581 , \9578 , \9579 , \9580 );
and \U$9393 ( \9582 , \5737 , \7082 );
not \U$9394 ( \9583 , \9582 );
xnor \U$9395 ( \9584 , \9583 , \7088 );
xor \U$9396 ( \9585 , \5923 , \9584 );
and \U$9397 ( \9586 , \5758 , \7099 );
and \U$9398 ( \9587 , \5770 , \7097 );
nor \U$9399 ( \9588 , \9586 , \9587 );
xnor \U$9400 ( \9589 , \9588 , \7105 );
xor \U$9401 ( \9590 , \9585 , \9589 );
xor \U$9402 ( \9591 , \9581 , \9590 );
and \U$9403 ( \9592 , \5906 , \5750 );
and \U$9404 ( \9593 , \5918 , \5748 );
nor \U$9405 ( \9594 , \9592 , \9593 );
xnor \U$9406 ( \9595 , \9594 , \5755 );
and \U$9407 ( \9596 , \5925 , \5768 );
and \U$9408 ( \9597 , \5937 , \5766 );
nor \U$9409 ( \9598 , \9596 , \9597 );
xnor \U$9410 ( \9599 , \9598 , \5775 );
xor \U$9411 ( \9600 , \9595 , \9599 );
and \U$9412 ( \9601 , \5945 , \5790 );
and \U$9413 ( \9602 , \5957 , \5788 );
nor \U$9414 ( \9603 , \9601 , \9602 );
xnor \U$9415 ( \9604 , \9603 , \5797 );
xor \U$9416 ( \9605 , \9600 , \9604 );
and \U$9417 ( \9606 , \5842 , \7175 );
and \U$9418 ( \9607 , \5854 , \7173 );
nor \U$9419 ( \9608 , \9606 , \9607 );
xnor \U$9420 ( \9609 , \9608 , \7181 );
and \U$9421 ( \9610 , \5861 , \7192 );
and \U$9422 ( \9611 , \5873 , \7190 );
nor \U$9423 ( \9612 , \9610 , \9611 );
xnor \U$9424 ( \9613 , \9612 , \7198 );
xor \U$9425 ( \9614 , \9609 , \9613 );
and \U$9426 ( \9615 , \5881 , \7203 );
and \U$9427 ( \9616 , \5893 , \7201 );
nor \U$9428 ( \9617 , \9615 , \9616 );
xnor \U$9429 ( \9618 , \9617 , \6824 );
xor \U$9430 ( \9619 , \9614 , \9618 );
xor \U$9431 ( \9620 , \9605 , \9619 );
and \U$9432 ( \9621 , \5780 , \7117 );
and \U$9433 ( \9622 , \5792 , \7115 );
nor \U$9434 ( \9623 , \9621 , \9622 );
xnor \U$9435 ( \9624 , \9623 , \7123 );
and \U$9436 ( \9625 , \5799 , \7140 );
and \U$9437 ( \9626 , \5811 , \7138 );
nor \U$9438 ( \9627 , \9625 , \9626 );
xnor \U$9439 ( \9628 , \9627 , \7146 );
xor \U$9440 ( \9629 , \9624 , \9628 );
and \U$9441 ( \9630 , \5819 , \7157 );
and \U$9442 ( \9631 , \5831 , \7155 );
nor \U$9443 ( \9632 , \9630 , \9631 );
xnor \U$9444 ( \9633 , \9632 , \7163 );
xor \U$9445 ( \9634 , \9629 , \9633 );
xor \U$9446 ( \9635 , \9620 , \9634 );
xor \U$9447 ( \9636 , \9591 , \9635 );
xor \U$9448 ( \9637 , \9577 , \9636 );
and \U$9449 ( \9638 , \9381 , \9385 );
and \U$9450 ( \9639 , \9385 , \9390 );
and \U$9451 ( \9640 , \9381 , \9390 );
or \U$9452 ( \9641 , \9638 , \9639 , \9640 );
and \U$9453 ( \9642 , \9367 , \9371 );
and \U$9454 ( \9643 , \9371 , \9376 );
and \U$9455 ( \9644 , \9367 , \9376 );
or \U$9456 ( \9645 , \9642 , \9643 , \9644 );
xor \U$9457 ( \9646 , \9641 , \9645 );
and \U$9458 ( \9647 , \9447 , \9461 );
and \U$9459 ( \9648 , \9461 , \9476 );
and \U$9460 ( \9649 , \9447 , \9476 );
or \U$9461 ( \9650 , \9647 , \9648 , \9649 );
xor \U$9462 ( \9651 , \9646 , \9650 );
xor \U$9463 ( \9652 , \9637 , \9651 );
xor \U$9464 ( \9653 , \9523 , \9652 );
xor \U$9465 ( \9654 , \9514 , \9653 );
and \U$9466 ( \9655 , \9339 , \9353 );
and \U$9467 ( \9656 , \9353 , \9492 );
and \U$9468 ( \9657 , \9339 , \9492 );
or \U$9469 ( \9658 , \9655 , \9656 , \9657 );
nor \U$9470 ( \9659 , \9654 , \9658 );
nor \U$9471 ( \9660 , \9498 , \9659 );
nand \U$9472 ( \9661 , \9335 , \9660 );
and \U$9473 ( \9662 , \9518 , \9522 );
and \U$9474 ( \9663 , \9522 , \9652 );
and \U$9475 ( \9664 , \9518 , \9652 );
or \U$9476 ( \9665 , \9662 , \9663 , \9664 );
and \U$9477 ( \9666 , \9641 , \9645 );
and \U$9478 ( \9667 , \9645 , \9650 );
and \U$9479 ( \9668 , \9641 , \9650 );
or \U$9480 ( \9669 , \9666 , \9667 , \9668 );
and \U$9481 ( \9670 , \9581 , \9590 );
and \U$9482 ( \9671 , \9590 , \9635 );
and \U$9483 ( \9672 , \9581 , \9635 );
or \U$9484 ( \9673 , \9670 , \9671 , \9672 );
xor \U$9485 ( \9674 , \9669 , \9673 );
and \U$9486 ( \9675 , \9550 , \9561 );
and \U$9487 ( \9676 , \9561 , \9576 );
and \U$9488 ( \9677 , \9550 , \9576 );
or \U$9489 ( \9678 , \9675 , \9676 , \9677 );
xor \U$9490 ( \9679 , \9674 , \9678 );
xor \U$9491 ( \9680 , \9665 , \9679 );
and \U$9492 ( \9681 , \9506 , \9510 );
and \U$9493 ( \9682 , \9510 , \9512 );
and \U$9494 ( \9683 , \9506 , \9512 );
or \U$9495 ( \9684 , \9681 , \9682 , \9683 );
and \U$9496 ( \9685 , \9577 , \9636 );
and \U$9497 ( \9686 , \9636 , \9651 );
and \U$9498 ( \9687 , \9577 , \9651 );
or \U$9499 ( \9688 , \9685 , \9686 , \9687 );
xor \U$9500 ( \9689 , \9684 , \9688 );
and \U$9501 ( \9690 , \9595 , \9599 );
and \U$9502 ( \9691 , \9599 , \9604 );
and \U$9503 ( \9692 , \9595 , \9604 );
or \U$9504 ( \9693 , \9690 , \9691 , \9692 );
and \U$9505 ( \9694 , \9539 , \9543 );
and \U$9506 ( \9695 , \9543 , \9548 );
and \U$9507 ( \9696 , \9539 , \9548 );
or \U$9508 ( \9697 , \9694 , \9695 , \9696 );
xor \U$9509 ( \9698 , \9693 , \9697 );
and \U$9510 ( \9699 , \9527 , \9531 );
and \U$9511 ( \9700 , \9531 , \9534 );
and \U$9512 ( \9701 , \9527 , \9534 );
or \U$9513 ( \9702 , \9699 , \9700 , \9701 );
xor \U$9514 ( \9703 , \9698 , \9702 );
and \U$9515 ( \9704 , \5923 , \9584 );
and \U$9516 ( \9705 , \9584 , \9589 );
and \U$9517 ( \9706 , \5923 , \9589 );
or \U$9518 ( \9707 , \9704 , \9705 , \9706 );
and \U$9519 ( \9708 , \9624 , \9628 );
and \U$9520 ( \9709 , \9628 , \9633 );
and \U$9521 ( \9710 , \9624 , \9633 );
or \U$9522 ( \9711 , \9708 , \9709 , \9710 );
xor \U$9523 ( \9712 , \9707 , \9711 );
and \U$9524 ( \9713 , \9609 , \9613 );
and \U$9525 ( \9714 , \9613 , \9618 );
and \U$9526 ( \9715 , \9609 , \9618 );
or \U$9527 ( \9716 , \9713 , \9714 , \9715 );
xor \U$9528 ( \9717 , \9712 , \9716 );
xor \U$9529 ( \9718 , \9703 , \9717 );
and \U$9530 ( \9719 , \9605 , \9619 );
and \U$9531 ( \9720 , \9619 , \9634 );
and \U$9532 ( \9721 , \9605 , \9634 );
or \U$9533 ( \9722 , \9719 , \9720 , \9721 );
and \U$9534 ( \9723 , \5873 , \7192 );
and \U$9535 ( \9724 , \5842 , \7190 );
nor \U$9536 ( \9725 , \9723 , \9724 );
xnor \U$9537 ( \9726 , \9725 , \7198 );
and \U$9538 ( \9727 , \5893 , \7203 );
and \U$9539 ( \9728 , \5861 , \7201 );
nor \U$9540 ( \9729 , \9727 , \9728 );
xnor \U$9541 ( \9730 , \9729 , \6824 );
xor \U$9542 ( \9731 , \9726 , \9730 );
and \U$9543 ( \9732 , \5918 , \5750 );
and \U$9544 ( \9733 , \5881 , \5748 );
nor \U$9545 ( \9734 , \9732 , \9733 );
xnor \U$9546 ( \9735 , \9734 , \5755 );
xor \U$9547 ( \9736 , \9731 , \9735 );
and \U$9548 ( \9737 , \5811 , \7140 );
and \U$9549 ( \9738 , \5780 , \7138 );
nor \U$9550 ( \9739 , \9737 , \9738 );
xnor \U$9551 ( \9740 , \9739 , \7146 );
and \U$9552 ( \9741 , \5831 , \7157 );
and \U$9553 ( \9742 , \5799 , \7155 );
nor \U$9554 ( \9743 , \9741 , \9742 );
xnor \U$9555 ( \9744 , \9743 , \7163 );
xor \U$9556 ( \9745 , \9740 , \9744 );
and \U$9557 ( \9746 , \5854 , \7175 );
and \U$9558 ( \9747 , \5819 , \7173 );
nor \U$9559 ( \9748 , \9746 , \9747 );
xnor \U$9560 ( \9749 , \9748 , \7181 );
xor \U$9561 ( \9750 , \9745 , \9749 );
xor \U$9562 ( \9751 , \9736 , \9750 );
not \U$9563 ( \9752 , \7088 );
and \U$9564 ( \9753 , \5770 , \7099 );
and \U$9565 ( \9754 , \5737 , \7097 );
nor \U$9566 ( \9755 , \9753 , \9754 );
xnor \U$9567 ( \9756 , \9755 , \7105 );
xor \U$9568 ( \9757 , \9752 , \9756 );
and \U$9569 ( \9758 , \5792 , \7117 );
and \U$9570 ( \9759 , \5758 , \7115 );
nor \U$9571 ( \9760 , \9758 , \9759 );
xnor \U$9572 ( \9761 , \9760 , \7123 );
xor \U$9573 ( \9762 , \9757 , \9761 );
xor \U$9574 ( \9763 , \9751 , \9762 );
xor \U$9575 ( \9764 , \9722 , \9763 );
and \U$9576 ( \9765 , \6057 , \5891 );
and \U$9577 ( \9766 , \6029 , \5889 );
nor \U$9578 ( \9767 , \9765 , \9766 );
xnor \U$9579 ( \9768 , \9767 , \5898 );
and \U$9580 ( \9769 , \6065 , \5916 );
and \U$9581 ( \9770 , \6048 , \5914 );
nor \U$9582 ( \9771 , \9769 , \9770 );
xnor \U$9583 ( \9772 , \9771 , \5923 );
xor \U$9584 ( \9773 , \9768 , \9772 );
and \U$9585 ( \9774 , \5998 , \5829 );
and \U$9586 ( \9775 , \5967 , \5827 );
nor \U$9587 ( \9776 , \9774 , \9775 );
xnor \U$9588 ( \9777 , \9776 , \5836 );
and \U$9589 ( \9778 , \6018 , \5852 );
and \U$9590 ( \9779 , \5986 , \5850 );
nor \U$9591 ( \9780 , \9778 , \9779 );
xnor \U$9592 ( \9781 , \9780 , \5859 );
xor \U$9593 ( \9782 , \9777 , \9781 );
and \U$9594 ( \9783 , \6041 , \5871 );
and \U$9595 ( \9784 , \6006 , \5869 );
nor \U$9596 ( \9785 , \9783 , \9784 );
xnor \U$9597 ( \9786 , \9785 , \5878 );
xor \U$9598 ( \9787 , \9782 , \9786 );
xor \U$9599 ( \9788 , \9773 , \9787 );
and \U$9600 ( \9789 , \5937 , \5768 );
and \U$9601 ( \9790 , \5906 , \5766 );
nor \U$9602 ( \9791 , \9789 , \9790 );
xnor \U$9603 ( \9792 , \9791 , \5775 );
and \U$9604 ( \9793 , \5957 , \5790 );
and \U$9605 ( \9794 , \5925 , \5788 );
nor \U$9606 ( \9795 , \9793 , \9794 );
xnor \U$9607 ( \9796 , \9795 , \5797 );
xor \U$9608 ( \9797 , \9792 , \9796 );
and \U$9609 ( \9798 , \5979 , \5809 );
and \U$9610 ( \9799 , \5945 , \5807 );
nor \U$9611 ( \9800 , \9798 , \9799 );
xnor \U$9612 ( \9801 , \9800 , \5816 );
xor \U$9613 ( \9802 , \9797 , \9801 );
xor \U$9614 ( \9803 , \9788 , \9802 );
xor \U$9615 ( \9804 , \9764 , \9803 );
xor \U$9616 ( \9805 , \9718 , \9804 );
and \U$9617 ( \9806 , \9566 , \9570 );
and \U$9618 ( \9807 , \9570 , \9575 );
and \U$9619 ( \9808 , \9566 , \9575 );
or \U$9620 ( \9809 , \9806 , \9807 , \9808 );
and \U$9621 ( \9810 , \9554 , \9558 );
and \U$9622 ( \9811 , \9558 , \9560 );
and \U$9623 ( \9812 , \9554 , \9560 );
or \U$9624 ( \9813 , \9810 , \9811 , \9812 );
xor \U$9625 ( \9814 , \9809 , \9813 );
or \U$9626 ( \9815 , \9535 , \9549 );
xor \U$9627 ( \9816 , \9814 , \9815 );
xor \U$9628 ( \9817 , \9805 , \9816 );
xor \U$9629 ( \9818 , \9689 , \9817 );
xor \U$9630 ( \9819 , \9680 , \9818 );
and \U$9631 ( \9820 , \9502 , \9513 );
and \U$9632 ( \9821 , \9513 , \9653 );
and \U$9633 ( \9822 , \9502 , \9653 );
or \U$9634 ( \9823 , \9820 , \9821 , \9822 );
nor \U$9635 ( \9824 , \9819 , \9823 );
and \U$9636 ( \9825 , \9684 , \9688 );
and \U$9637 ( \9826 , \9688 , \9817 );
and \U$9638 ( \9827 , \9684 , \9817 );
or \U$9639 ( \9828 , \9825 , \9826 , \9827 );
and \U$9640 ( \9829 , \9809 , \9813 );
and \U$9641 ( \9830 , \9813 , \9815 );
and \U$9642 ( \9831 , \9809 , \9815 );
or \U$9643 ( \9832 , \9829 , \9830 , \9831 );
and \U$9644 ( \9833 , \9722 , \9763 );
and \U$9645 ( \9834 , \9763 , \9803 );
and \U$9646 ( \9835 , \9722 , \9803 );
or \U$9647 ( \9836 , \9833 , \9834 , \9835 );
xor \U$9648 ( \9837 , \9832 , \9836 );
and \U$9649 ( \9838 , \9703 , \9717 );
xor \U$9650 ( \9839 , \9837 , \9838 );
xor \U$9651 ( \9840 , \9828 , \9839 );
and \U$9652 ( \9841 , \9669 , \9673 );
and \U$9653 ( \9842 , \9673 , \9678 );
and \U$9654 ( \9843 , \9669 , \9678 );
or \U$9655 ( \9844 , \9841 , \9842 , \9843 );
and \U$9656 ( \9845 , \9718 , \9804 );
and \U$9657 ( \9846 , \9804 , \9816 );
and \U$9658 ( \9847 , \9718 , \9816 );
or \U$9659 ( \9848 , \9845 , \9846 , \9847 );
xor \U$9660 ( \9849 , \9844 , \9848 );
and \U$9661 ( \9850 , \6029 , \5891 );
and \U$9662 ( \9851 , \6041 , \5889 );
nor \U$9663 ( \9852 , \9850 , \9851 );
xnor \U$9664 ( \9853 , \9852 , \5898 );
and \U$9665 ( \9854 , \6048 , \5916 );
and \U$9666 ( \9855 , \6057 , \5914 );
nor \U$9667 ( \9856 , \9854 , \9855 );
xnor \U$9668 ( \9857 , \9856 , \5923 );
xor \U$9669 ( \9858 , \9853 , \9857 );
nand \U$9670 ( \9859 , \6065 , \5933 );
xnor \U$9671 ( \9860 , \9859 , \5942 );
xor \U$9672 ( \9861 , \9858 , \9860 );
and \U$9673 ( \9862 , \5967 , \5829 );
and \U$9674 ( \9863 , \5979 , \5827 );
nor \U$9675 ( \9864 , \9862 , \9863 );
xnor \U$9676 ( \9865 , \9864 , \5836 );
and \U$9677 ( \9866 , \5986 , \5852 );
and \U$9678 ( \9867 , \5998 , \5850 );
nor \U$9679 ( \9868 , \9866 , \9867 );
xnor \U$9680 ( \9869 , \9868 , \5859 );
xor \U$9681 ( \9870 , \9865 , \9869 );
and \U$9682 ( \9871 , \6006 , \5871 );
and \U$9683 ( \9872 , \6018 , \5869 );
nor \U$9684 ( \9873 , \9871 , \9872 );
xnor \U$9685 ( \9874 , \9873 , \5878 );
xor \U$9686 ( \9875 , \9870 , \9874 );
xnor \U$9687 ( \9876 , \9861 , \9875 );
and \U$9688 ( \9877 , \9792 , \9796 );
and \U$9689 ( \9878 , \9796 , \9801 );
and \U$9690 ( \9879 , \9792 , \9801 );
or \U$9691 ( \9880 , \9877 , \9878 , \9879 );
and \U$9692 ( \9881 , \9777 , \9781 );
and \U$9693 ( \9882 , \9781 , \9786 );
and \U$9694 ( \9883 , \9777 , \9786 );
or \U$9695 ( \9884 , \9881 , \9882 , \9883 );
xor \U$9696 ( \9885 , \9880 , \9884 );
and \U$9697 ( \9886 , \9768 , \9772 );
xor \U$9698 ( \9887 , \9885 , \9886 );
xor \U$9699 ( \9888 , \9876 , \9887 );
and \U$9700 ( \9889 , \9752 , \9756 );
and \U$9701 ( \9890 , \9756 , \9761 );
and \U$9702 ( \9891 , \9752 , \9761 );
or \U$9703 ( \9892 , \9889 , \9890 , \9891 );
and \U$9704 ( \9893 , \9740 , \9744 );
and \U$9705 ( \9894 , \9744 , \9749 );
and \U$9706 ( \9895 , \9740 , \9749 );
or \U$9707 ( \9896 , \9893 , \9894 , \9895 );
xor \U$9708 ( \9897 , \9892 , \9896 );
and \U$9709 ( \9898 , \9726 , \9730 );
and \U$9710 ( \9899 , \9730 , \9735 );
and \U$9711 ( \9900 , \9726 , \9735 );
or \U$9712 ( \9901 , \9898 , \9899 , \9900 );
xor \U$9713 ( \9902 , \9897 , \9901 );
xor \U$9714 ( \9903 , \9888 , \9902 );
and \U$9715 ( \9904 , \9736 , \9750 );
and \U$9716 ( \9905 , \9750 , \9762 );
and \U$9717 ( \9906 , \9736 , \9762 );
or \U$9718 ( \9907 , \9904 , \9905 , \9906 );
and \U$9719 ( \9908 , \5737 , \7099 );
not \U$9720 ( \9909 , \9908 );
xnor \U$9721 ( \9910 , \9909 , \7105 );
xor \U$9722 ( \9911 , \5942 , \9910 );
and \U$9723 ( \9912 , \5758 , \7117 );
and \U$9724 ( \9913 , \5770 , \7115 );
nor \U$9725 ( \9914 , \9912 , \9913 );
xnor \U$9726 ( \9915 , \9914 , \7123 );
xor \U$9727 ( \9916 , \9911 , \9915 );
xor \U$9728 ( \9917 , \9907 , \9916 );
and \U$9729 ( \9918 , \5906 , \5768 );
and \U$9730 ( \9919 , \5918 , \5766 );
nor \U$9731 ( \9920 , \9918 , \9919 );
xnor \U$9732 ( \9921 , \9920 , \5775 );
and \U$9733 ( \9922 , \5925 , \5790 );
and \U$9734 ( \9923 , \5937 , \5788 );
nor \U$9735 ( \9924 , \9922 , \9923 );
xnor \U$9736 ( \9925 , \9924 , \5797 );
xor \U$9737 ( \9926 , \9921 , \9925 );
and \U$9738 ( \9927 , \5945 , \5809 );
and \U$9739 ( \9928 , \5957 , \5807 );
nor \U$9740 ( \9929 , \9927 , \9928 );
xnor \U$9741 ( \9930 , \9929 , \5816 );
xor \U$9742 ( \9931 , \9926 , \9930 );
and \U$9743 ( \9932 , \5842 , \7192 );
and \U$9744 ( \9933 , \5854 , \7190 );
nor \U$9745 ( \9934 , \9932 , \9933 );
xnor \U$9746 ( \9935 , \9934 , \7198 );
and \U$9747 ( \9936 , \5861 , \7203 );
and \U$9748 ( \9937 , \5873 , \7201 );
nor \U$9749 ( \9938 , \9936 , \9937 );
xnor \U$9750 ( \9939 , \9938 , \6824 );
xor \U$9751 ( \9940 , \9935 , \9939 );
and \U$9752 ( \9941 , \5881 , \5750 );
and \U$9753 ( \9942 , \5893 , \5748 );
nor \U$9754 ( \9943 , \9941 , \9942 );
xnor \U$9755 ( \9944 , \9943 , \5755 );
xor \U$9756 ( \9945 , \9940 , \9944 );
xor \U$9757 ( \9946 , \9931 , \9945 );
and \U$9758 ( \9947 , \5780 , \7140 );
and \U$9759 ( \9948 , \5792 , \7138 );
nor \U$9760 ( \9949 , \9947 , \9948 );
xnor \U$9761 ( \9950 , \9949 , \7146 );
and \U$9762 ( \9951 , \5799 , \7157 );
and \U$9763 ( \9952 , \5811 , \7155 );
nor \U$9764 ( \9953 , \9951 , \9952 );
xnor \U$9765 ( \9954 , \9953 , \7163 );
xor \U$9766 ( \9955 , \9950 , \9954 );
and \U$9767 ( \9956 , \5819 , \7175 );
and \U$9768 ( \9957 , \5831 , \7173 );
nor \U$9769 ( \9958 , \9956 , \9957 );
xnor \U$9770 ( \9959 , \9958 , \7181 );
xor \U$9771 ( \9960 , \9955 , \9959 );
xor \U$9772 ( \9961 , \9946 , \9960 );
xor \U$9773 ( \9962 , \9917 , \9961 );
xor \U$9774 ( \9963 , \9903 , \9962 );
and \U$9775 ( \9964 , \9707 , \9711 );
and \U$9776 ( \9965 , \9711 , \9716 );
and \U$9777 ( \9966 , \9707 , \9716 );
or \U$9778 ( \9967 , \9964 , \9965 , \9966 );
and \U$9779 ( \9968 , \9693 , \9697 );
and \U$9780 ( \9969 , \9697 , \9702 );
and \U$9781 ( \9970 , \9693 , \9702 );
or \U$9782 ( \9971 , \9968 , \9969 , \9970 );
xor \U$9783 ( \9972 , \9967 , \9971 );
and \U$9784 ( \9973 , \9773 , \9787 );
and \U$9785 ( \9974 , \9787 , \9802 );
and \U$9786 ( \9975 , \9773 , \9802 );
or \U$9787 ( \9976 , \9973 , \9974 , \9975 );
xor \U$9788 ( \9977 , \9972 , \9976 );
xor \U$9789 ( \9978 , \9963 , \9977 );
xor \U$9790 ( \9979 , \9849 , \9978 );
xor \U$9791 ( \9980 , \9840 , \9979 );
and \U$9792 ( \9981 , \9665 , \9679 );
and \U$9793 ( \9982 , \9679 , \9818 );
and \U$9794 ( \9983 , \9665 , \9818 );
or \U$9795 ( \9984 , \9981 , \9982 , \9983 );
nor \U$9796 ( \9985 , \9980 , \9984 );
nor \U$9797 ( \9986 , \9824 , \9985 );
and \U$9798 ( \9987 , \9844 , \9848 );
and \U$9799 ( \9988 , \9848 , \9978 );
and \U$9800 ( \9989 , \9844 , \9978 );
or \U$9801 ( \9990 , \9987 , \9988 , \9989 );
and \U$9802 ( \9991 , \9967 , \9971 );
and \U$9803 ( \9992 , \9971 , \9976 );
and \U$9804 ( \9993 , \9967 , \9976 );
or \U$9805 ( \9994 , \9991 , \9992 , \9993 );
and \U$9806 ( \9995 , \9907 , \9916 );
and \U$9807 ( \9996 , \9916 , \9961 );
and \U$9808 ( \9997 , \9907 , \9961 );
or \U$9809 ( \9998 , \9995 , \9996 , \9997 );
xor \U$9810 ( \9999 , \9994 , \9998 );
and \U$9811 ( \10000 , \9876 , \9887 );
and \U$9812 ( \10001 , \9887 , \9902 );
and \U$9813 ( \10002 , \9876 , \9902 );
or \U$9814 ( \10003 , \10000 , \10001 , \10002 );
xor \U$9815 ( \10004 , \9999 , \10003 );
xor \U$9816 ( \10005 , \9990 , \10004 );
and \U$9817 ( \10006 , \9832 , \9836 );
and \U$9818 ( \10007 , \9836 , \9838 );
and \U$9819 ( \10008 , \9832 , \9838 );
or \U$9820 ( \10009 , \10006 , \10007 , \10008 );
and \U$9821 ( \10010 , \9903 , \9962 );
and \U$9822 ( \10011 , \9962 , \9977 );
and \U$9823 ( \10012 , \9903 , \9977 );
or \U$9824 ( \10013 , \10010 , \10011 , \10012 );
xor \U$9825 ( \10014 , \10009 , \10013 );
and \U$9826 ( \10015 , \9921 , \9925 );
and \U$9827 ( \10016 , \9925 , \9930 );
and \U$9828 ( \10017 , \9921 , \9930 );
or \U$9829 ( \10018 , \10015 , \10016 , \10017 );
and \U$9830 ( \10019 , \9865 , \9869 );
and \U$9831 ( \10020 , \9869 , \9874 );
and \U$9832 ( \10021 , \9865 , \9874 );
or \U$9833 ( \10022 , \10019 , \10020 , \10021 );
xor \U$9834 ( \10023 , \10018 , \10022 );
and \U$9835 ( \10024 , \9853 , \9857 );
and \U$9836 ( \10025 , \9857 , \9860 );
and \U$9837 ( \10026 , \9853 , \9860 );
or \U$9838 ( \10027 , \10024 , \10025 , \10026 );
xor \U$9839 ( \10028 , \10023 , \10027 );
and \U$9840 ( \10029 , \5942 , \9910 );
and \U$9841 ( \10030 , \9910 , \9915 );
and \U$9842 ( \10031 , \5942 , \9915 );
or \U$9843 ( \10032 , \10029 , \10030 , \10031 );
and \U$9844 ( \10033 , \9950 , \9954 );
and \U$9845 ( \10034 , \9954 , \9959 );
and \U$9846 ( \10035 , \9950 , \9959 );
or \U$9847 ( \10036 , \10033 , \10034 , \10035 );
xor \U$9848 ( \10037 , \10032 , \10036 );
and \U$9849 ( \10038 , \9935 , \9939 );
and \U$9850 ( \10039 , \9939 , \9944 );
and \U$9851 ( \10040 , \9935 , \9944 );
or \U$9852 ( \10041 , \10038 , \10039 , \10040 );
xor \U$9853 ( \10042 , \10037 , \10041 );
xor \U$9854 ( \10043 , \10028 , \10042 );
and \U$9855 ( \10044 , \9931 , \9945 );
and \U$9856 ( \10045 , \9945 , \9960 );
and \U$9857 ( \10046 , \9931 , \9960 );
or \U$9858 ( \10047 , \10044 , \10045 , \10046 );
and \U$9859 ( \10048 , \5873 , \7203 );
and \U$9860 ( \10049 , \5842 , \7201 );
nor \U$9861 ( \10050 , \10048 , \10049 );
xnor \U$9862 ( \10051 , \10050 , \6824 );
and \U$9863 ( \10052 , \5893 , \5750 );
and \U$9864 ( \10053 , \5861 , \5748 );
nor \U$9865 ( \10054 , \10052 , \10053 );
xnor \U$9866 ( \10055 , \10054 , \5755 );
xor \U$9867 ( \10056 , \10051 , \10055 );
and \U$9868 ( \10057 , \5918 , \5768 );
and \U$9869 ( \10058 , \5881 , \5766 );
nor \U$9870 ( \10059 , \10057 , \10058 );
xnor \U$9871 ( \10060 , \10059 , \5775 );
xor \U$9872 ( \10061 , \10056 , \10060 );
and \U$9873 ( \10062 , \5811 , \7157 );
and \U$9874 ( \10063 , \5780 , \7155 );
nor \U$9875 ( \10064 , \10062 , \10063 );
xnor \U$9876 ( \10065 , \10064 , \7163 );
and \U$9877 ( \10066 , \5831 , \7175 );
and \U$9878 ( \10067 , \5799 , \7173 );
nor \U$9879 ( \10068 , \10066 , \10067 );
xnor \U$9880 ( \10069 , \10068 , \7181 );
xor \U$9881 ( \10070 , \10065 , \10069 );
and \U$9882 ( \10071 , \5854 , \7192 );
and \U$9883 ( \10072 , \5819 , \7190 );
nor \U$9884 ( \10073 , \10071 , \10072 );
xnor \U$9885 ( \10074 , \10073 , \7198 );
xor \U$9886 ( \10075 , \10070 , \10074 );
xor \U$9887 ( \10076 , \10061 , \10075 );
not \U$9888 ( \10077 , \7105 );
and \U$9889 ( \10078 , \5770 , \7117 );
and \U$9890 ( \10079 , \5737 , \7115 );
nor \U$9891 ( \10080 , \10078 , \10079 );
xnor \U$9892 ( \10081 , \10080 , \7123 );
xor \U$9893 ( \10082 , \10077 , \10081 );
and \U$9894 ( \10083 , \5792 , \7140 );
and \U$9895 ( \10084 , \5758 , \7138 );
nor \U$9896 ( \10085 , \10083 , \10084 );
xnor \U$9897 ( \10086 , \10085 , \7146 );
xor \U$9898 ( \10087 , \10082 , \10086 );
xor \U$9899 ( \10088 , \10076 , \10087 );
xor \U$9900 ( \10089 , \10047 , \10088 );
and \U$9901 ( \10090 , \6057 , \5916 );
and \U$9902 ( \10091 , \6029 , \5914 );
nor \U$9903 ( \10092 , \10090 , \10091 );
xnor \U$9904 ( \10093 , \10092 , \5923 );
and \U$9905 ( \10094 , \6065 , \5935 );
and \U$9906 ( \10095 , \6048 , \5933 );
nor \U$9907 ( \10096 , \10094 , \10095 );
xnor \U$9908 ( \10097 , \10096 , \5942 );
xor \U$9909 ( \10098 , \10093 , \10097 );
and \U$9910 ( \10099 , \5998 , \5852 );
and \U$9911 ( \10100 , \5967 , \5850 );
nor \U$9912 ( \10101 , \10099 , \10100 );
xnor \U$9913 ( \10102 , \10101 , \5859 );
and \U$9914 ( \10103 , \6018 , \5871 );
and \U$9915 ( \10104 , \5986 , \5869 );
nor \U$9916 ( \10105 , \10103 , \10104 );
xnor \U$9917 ( \10106 , \10105 , \5878 );
xor \U$9918 ( \10107 , \10102 , \10106 );
and \U$9919 ( \10108 , \6041 , \5891 );
and \U$9920 ( \10109 , \6006 , \5889 );
nor \U$9921 ( \10110 , \10108 , \10109 );
xnor \U$9922 ( \10111 , \10110 , \5898 );
xor \U$9923 ( \10112 , \10107 , \10111 );
xor \U$9924 ( \10113 , \10098 , \10112 );
and \U$9925 ( \10114 , \5937 , \5790 );
and \U$9926 ( \10115 , \5906 , \5788 );
nor \U$9927 ( \10116 , \10114 , \10115 );
xnor \U$9928 ( \10117 , \10116 , \5797 );
and \U$9929 ( \10118 , \5957 , \5809 );
and \U$9930 ( \10119 , \5925 , \5807 );
nor \U$9931 ( \10120 , \10118 , \10119 );
xnor \U$9932 ( \10121 , \10120 , \5816 );
xor \U$9933 ( \10122 , \10117 , \10121 );
and \U$9934 ( \10123 , \5979 , \5829 );
and \U$9935 ( \10124 , \5945 , \5827 );
nor \U$9936 ( \10125 , \10123 , \10124 );
xnor \U$9937 ( \10126 , \10125 , \5836 );
xor \U$9938 ( \10127 , \10122 , \10126 );
xor \U$9939 ( \10128 , \10113 , \10127 );
xor \U$9940 ( \10129 , \10089 , \10128 );
xor \U$9941 ( \10130 , \10043 , \10129 );
and \U$9942 ( \10131 , \9892 , \9896 );
and \U$9943 ( \10132 , \9896 , \9901 );
and \U$9944 ( \10133 , \9892 , \9901 );
or \U$9945 ( \10134 , \10131 , \10132 , \10133 );
and \U$9946 ( \10135 , \9880 , \9884 );
and \U$9947 ( \10136 , \9884 , \9886 );
and \U$9948 ( \10137 , \9880 , \9886 );
or \U$9949 ( \10138 , \10135 , \10136 , \10137 );
xor \U$9950 ( \10139 , \10134 , \10138 );
or \U$9951 ( \10140 , \9861 , \9875 );
xor \U$9952 ( \10141 , \10139 , \10140 );
xor \U$9953 ( \10142 , \10130 , \10141 );
xor \U$9954 ( \10143 , \10014 , \10142 );
xor \U$9955 ( \10144 , \10005 , \10143 );
and \U$9956 ( \10145 , \9828 , \9839 );
and \U$9957 ( \10146 , \9839 , \9979 );
and \U$9958 ( \10147 , \9828 , \9979 );
or \U$9959 ( \10148 , \10145 , \10146 , \10147 );
nor \U$9960 ( \10149 , \10144 , \10148 );
and \U$9961 ( \10150 , \10009 , \10013 );
and \U$9962 ( \10151 , \10013 , \10142 );
and \U$9963 ( \10152 , \10009 , \10142 );
or \U$9964 ( \10153 , \10150 , \10151 , \10152 );
and \U$9965 ( \10154 , \10134 , \10138 );
and \U$9966 ( \10155 , \10138 , \10140 );
and \U$9967 ( \10156 , \10134 , \10140 );
or \U$9968 ( \10157 , \10154 , \10155 , \10156 );
and \U$9969 ( \10158 , \10047 , \10088 );
and \U$9970 ( \10159 , \10088 , \10128 );
and \U$9971 ( \10160 , \10047 , \10128 );
or \U$9972 ( \10161 , \10158 , \10159 , \10160 );
xor \U$9973 ( \10162 , \10157 , \10161 );
and \U$9974 ( \10163 , \10028 , \10042 );
xor \U$9975 ( \10164 , \10162 , \10163 );
xor \U$9976 ( \10165 , \10153 , \10164 );
and \U$9977 ( \10166 , \9994 , \9998 );
and \U$9978 ( \10167 , \9998 , \10003 );
and \U$9979 ( \10168 , \9994 , \10003 );
or \U$9980 ( \10169 , \10166 , \10167 , \10168 );
and \U$9981 ( \10170 , \10043 , \10129 );
and \U$9982 ( \10171 , \10129 , \10141 );
and \U$9983 ( \10172 , \10043 , \10141 );
or \U$9984 ( \10173 , \10170 , \10171 , \10172 );
xor \U$9985 ( \10174 , \10169 , \10173 );
and \U$9986 ( \10175 , \6029 , \5916 );
and \U$9987 ( \10176 , \6041 , \5914 );
nor \U$9988 ( \10177 , \10175 , \10176 );
xnor \U$9989 ( \10178 , \10177 , \5923 );
and \U$9990 ( \10179 , \6048 , \5935 );
and \U$9991 ( \10180 , \6057 , \5933 );
nor \U$9992 ( \10181 , \10179 , \10180 );
xnor \U$9993 ( \10182 , \10181 , \5942 );
xor \U$9994 ( \10183 , \10178 , \10182 );
nand \U$9995 ( \10184 , \6065 , \5953 );
xnor \U$9996 ( \10185 , \10184 , \5962 );
xor \U$9997 ( \10186 , \10183 , \10185 );
and \U$9998 ( \10187 , \5967 , \5852 );
and \U$9999 ( \10188 , \5979 , \5850 );
nor \U$10000 ( \10189 , \10187 , \10188 );
xnor \U$10001 ( \10190 , \10189 , \5859 );
and \U$10002 ( \10191 , \5986 , \5871 );
and \U$10003 ( \10192 , \5998 , \5869 );
nor \U$10004 ( \10193 , \10191 , \10192 );
xnor \U$10005 ( \10194 , \10193 , \5878 );
xor \U$10006 ( \10195 , \10190 , \10194 );
and \U$10007 ( \10196 , \6006 , \5891 );
and \U$10008 ( \10197 , \6018 , \5889 );
nor \U$10009 ( \10198 , \10196 , \10197 );
xnor \U$10010 ( \10199 , \10198 , \5898 );
xor \U$10011 ( \10200 , \10195 , \10199 );
xnor \U$10012 ( \10201 , \10186 , \10200 );
and \U$10013 ( \10202 , \10117 , \10121 );
and \U$10014 ( \10203 , \10121 , \10126 );
and \U$10015 ( \10204 , \10117 , \10126 );
or \U$10016 ( \10205 , \10202 , \10203 , \10204 );
and \U$10017 ( \10206 , \10102 , \10106 );
and \U$10018 ( \10207 , \10106 , \10111 );
and \U$10019 ( \10208 , \10102 , \10111 );
or \U$10020 ( \10209 , \10206 , \10207 , \10208 );
xor \U$10021 ( \10210 , \10205 , \10209 );
and \U$10022 ( \10211 , \10093 , \10097 );
xor \U$10023 ( \10212 , \10210 , \10211 );
xor \U$10024 ( \10213 , \10201 , \10212 );
and \U$10025 ( \10214 , \10077 , \10081 );
and \U$10026 ( \10215 , \10081 , \10086 );
and \U$10027 ( \10216 , \10077 , \10086 );
or \U$10028 ( \10217 , \10214 , \10215 , \10216 );
and \U$10029 ( \10218 , \10065 , \10069 );
and \U$10030 ( \10219 , \10069 , \10074 );
and \U$10031 ( \10220 , \10065 , \10074 );
or \U$10032 ( \10221 , \10218 , \10219 , \10220 );
xor \U$10033 ( \10222 , \10217 , \10221 );
and \U$10034 ( \10223 , \10051 , \10055 );
and \U$10035 ( \10224 , \10055 , \10060 );
and \U$10036 ( \10225 , \10051 , \10060 );
or \U$10037 ( \10226 , \10223 , \10224 , \10225 );
xor \U$10038 ( \10227 , \10222 , \10226 );
xor \U$10039 ( \10228 , \10213 , \10227 );
and \U$10040 ( \10229 , \10061 , \10075 );
and \U$10041 ( \10230 , \10075 , \10087 );
and \U$10042 ( \10231 , \10061 , \10087 );
or \U$10043 ( \10232 , \10229 , \10230 , \10231 );
and \U$10044 ( \10233 , \5737 , \7117 );
not \U$10045 ( \10234 , \10233 );
xnor \U$10046 ( \10235 , \10234 , \7123 );
xor \U$10047 ( \10236 , \5962 , \10235 );
and \U$10048 ( \10237 , \5758 , \7140 );
and \U$10049 ( \10238 , \5770 , \7138 );
nor \U$10050 ( \10239 , \10237 , \10238 );
xnor \U$10051 ( \10240 , \10239 , \7146 );
xor \U$10052 ( \10241 , \10236 , \10240 );
xor \U$10053 ( \10242 , \10232 , \10241 );
and \U$10054 ( \10243 , \5906 , \5790 );
and \U$10055 ( \10244 , \5918 , \5788 );
nor \U$10056 ( \10245 , \10243 , \10244 );
xnor \U$10057 ( \10246 , \10245 , \5797 );
and \U$10058 ( \10247 , \5925 , \5809 );
and \U$10059 ( \10248 , \5937 , \5807 );
nor \U$10060 ( \10249 , \10247 , \10248 );
xnor \U$10061 ( \10250 , \10249 , \5816 );
xor \U$10062 ( \10251 , \10246 , \10250 );
and \U$10063 ( \10252 , \5945 , \5829 );
and \U$10064 ( \10253 , \5957 , \5827 );
nor \U$10065 ( \10254 , \10252 , \10253 );
xnor \U$10066 ( \10255 , \10254 , \5836 );
xor \U$10067 ( \10256 , \10251 , \10255 );
and \U$10068 ( \10257 , \5842 , \7203 );
and \U$10069 ( \10258 , \5854 , \7201 );
nor \U$10070 ( \10259 , \10257 , \10258 );
xnor \U$10071 ( \10260 , \10259 , \6824 );
and \U$10072 ( \10261 , \5861 , \5750 );
and \U$10073 ( \10262 , \5873 , \5748 );
nor \U$10074 ( \10263 , \10261 , \10262 );
xnor \U$10075 ( \10264 , \10263 , \5755 );
xor \U$10076 ( \10265 , \10260 , \10264 );
and \U$10077 ( \10266 , \5881 , \5768 );
and \U$10078 ( \10267 , \5893 , \5766 );
nor \U$10079 ( \10268 , \10266 , \10267 );
xnor \U$10080 ( \10269 , \10268 , \5775 );
xor \U$10081 ( \10270 , \10265 , \10269 );
xor \U$10082 ( \10271 , \10256 , \10270 );
and \U$10083 ( \10272 , \5780 , \7157 );
and \U$10084 ( \10273 , \5792 , \7155 );
nor \U$10085 ( \10274 , \10272 , \10273 );
xnor \U$10086 ( \10275 , \10274 , \7163 );
and \U$10087 ( \10276 , \5799 , \7175 );
and \U$10088 ( \10277 , \5811 , \7173 );
nor \U$10089 ( \10278 , \10276 , \10277 );
xnor \U$10090 ( \10279 , \10278 , \7181 );
xor \U$10091 ( \10280 , \10275 , \10279 );
and \U$10092 ( \10281 , \5819 , \7192 );
and \U$10093 ( \10282 , \5831 , \7190 );
nor \U$10094 ( \10283 , \10281 , \10282 );
xnor \U$10095 ( \10284 , \10283 , \7198 );
xor \U$10096 ( \10285 , \10280 , \10284 );
xor \U$10097 ( \10286 , \10271 , \10285 );
xor \U$10098 ( \10287 , \10242 , \10286 );
xor \U$10099 ( \10288 , \10228 , \10287 );
and \U$10100 ( \10289 , \10032 , \10036 );
and \U$10101 ( \10290 , \10036 , \10041 );
and \U$10102 ( \10291 , \10032 , \10041 );
or \U$10103 ( \10292 , \10289 , \10290 , \10291 );
and \U$10104 ( \10293 , \10018 , \10022 );
and \U$10105 ( \10294 , \10022 , \10027 );
and \U$10106 ( \10295 , \10018 , \10027 );
or \U$10107 ( \10296 , \10293 , \10294 , \10295 );
xor \U$10108 ( \10297 , \10292 , \10296 );
and \U$10109 ( \10298 , \10098 , \10112 );
and \U$10110 ( \10299 , \10112 , \10127 );
and \U$10111 ( \10300 , \10098 , \10127 );
or \U$10112 ( \10301 , \10298 , \10299 , \10300 );
xor \U$10113 ( \10302 , \10297 , \10301 );
xor \U$10114 ( \10303 , \10288 , \10302 );
xor \U$10115 ( \10304 , \10174 , \10303 );
xor \U$10116 ( \10305 , \10165 , \10304 );
and \U$10117 ( \10306 , \9990 , \10004 );
and \U$10118 ( \10307 , \10004 , \10143 );
and \U$10119 ( \10308 , \9990 , \10143 );
or \U$10120 ( \10309 , \10306 , \10307 , \10308 );
nor \U$10121 ( \10310 , \10305 , \10309 );
nor \U$10122 ( \10311 , \10149 , \10310 );
nand \U$10123 ( \10312 , \9986 , \10311 );
nor \U$10124 ( \10313 , \9661 , \10312 );
nand \U$10125 ( \10314 , \9010 , \10313 );
and \U$10126 ( \10315 , \10169 , \10173 );
and \U$10127 ( \10316 , \10173 , \10303 );
and \U$10128 ( \10317 , \10169 , \10303 );
or \U$10129 ( \10318 , \10315 , \10316 , \10317 );
and \U$10130 ( \10319 , \10292 , \10296 );
and \U$10131 ( \10320 , \10296 , \10301 );
and \U$10132 ( \10321 , \10292 , \10301 );
or \U$10133 ( \10322 , \10319 , \10320 , \10321 );
and \U$10134 ( \10323 , \10232 , \10241 );
and \U$10135 ( \10324 , \10241 , \10286 );
and \U$10136 ( \10325 , \10232 , \10286 );
or \U$10137 ( \10326 , \10323 , \10324 , \10325 );
xor \U$10138 ( \10327 , \10322 , \10326 );
and \U$10139 ( \10328 , \10201 , \10212 );
and \U$10140 ( \10329 , \10212 , \10227 );
and \U$10141 ( \10330 , \10201 , \10227 );
or \U$10142 ( \10331 , \10328 , \10329 , \10330 );
xor \U$10143 ( \10332 , \10327 , \10331 );
xor \U$10144 ( \10333 , \10318 , \10332 );
and \U$10145 ( \10334 , \10157 , \10161 );
and \U$10146 ( \10335 , \10161 , \10163 );
and \U$10147 ( \10336 , \10157 , \10163 );
or \U$10148 ( \10337 , \10334 , \10335 , \10336 );
and \U$10149 ( \10338 , \10228 , \10287 );
and \U$10150 ( \10339 , \10287 , \10302 );
and \U$10151 ( \10340 , \10228 , \10302 );
or \U$10152 ( \10341 , \10338 , \10339 , \10340 );
xor \U$10153 ( \10342 , \10337 , \10341 );
and \U$10154 ( \10343 , \10246 , \10250 );
and \U$10155 ( \10344 , \10250 , \10255 );
and \U$10156 ( \10345 , \10246 , \10255 );
or \U$10157 ( \10346 , \10343 , \10344 , \10345 );
and \U$10158 ( \10347 , \10190 , \10194 );
and \U$10159 ( \10348 , \10194 , \10199 );
and \U$10160 ( \10349 , \10190 , \10199 );
or \U$10161 ( \10350 , \10347 , \10348 , \10349 );
xor \U$10162 ( \10351 , \10346 , \10350 );
and \U$10163 ( \10352 , \10178 , \10182 );
and \U$10164 ( \10353 , \10182 , \10185 );
and \U$10165 ( \10354 , \10178 , \10185 );
or \U$10166 ( \10355 , \10352 , \10353 , \10354 );
xor \U$10167 ( \10356 , \10351 , \10355 );
and \U$10168 ( \10357 , \5962 , \10235 );
and \U$10169 ( \10358 , \10235 , \10240 );
and \U$10170 ( \10359 , \5962 , \10240 );
or \U$10171 ( \10360 , \10357 , \10358 , \10359 );
and \U$10172 ( \10361 , \10275 , \10279 );
and \U$10173 ( \10362 , \10279 , \10284 );
and \U$10174 ( \10363 , \10275 , \10284 );
or \U$10175 ( \10364 , \10361 , \10362 , \10363 );
xor \U$10176 ( \10365 , \10360 , \10364 );
and \U$10177 ( \10366 , \10260 , \10264 );
and \U$10178 ( \10367 , \10264 , \10269 );
and \U$10179 ( \10368 , \10260 , \10269 );
or \U$10180 ( \10369 , \10366 , \10367 , \10368 );
xor \U$10181 ( \10370 , \10365 , \10369 );
xor \U$10182 ( \10371 , \10356 , \10370 );
and \U$10183 ( \10372 , \10256 , \10270 );
and \U$10184 ( \10373 , \10270 , \10285 );
and \U$10185 ( \10374 , \10256 , \10285 );
or \U$10186 ( \10375 , \10372 , \10373 , \10374 );
and \U$10187 ( \10376 , \5873 , \5750 );
and \U$10188 ( \10377 , \5842 , \5748 );
nor \U$10189 ( \10378 , \10376 , \10377 );
xnor \U$10190 ( \10379 , \10378 , \5755 );
and \U$10191 ( \10380 , \5893 , \5768 );
and \U$10192 ( \10381 , \5861 , \5766 );
nor \U$10193 ( \10382 , \10380 , \10381 );
xnor \U$10194 ( \10383 , \10382 , \5775 );
xor \U$10195 ( \10384 , \10379 , \10383 );
and \U$10196 ( \10385 , \5918 , \5790 );
and \U$10197 ( \10386 , \5881 , \5788 );
nor \U$10198 ( \10387 , \10385 , \10386 );
xnor \U$10199 ( \10388 , \10387 , \5797 );
xor \U$10200 ( \10389 , \10384 , \10388 );
and \U$10201 ( \10390 , \5811 , \7175 );
and \U$10202 ( \10391 , \5780 , \7173 );
nor \U$10203 ( \10392 , \10390 , \10391 );
xnor \U$10204 ( \10393 , \10392 , \7181 );
and \U$10205 ( \10394 , \5831 , \7192 );
and \U$10206 ( \10395 , \5799 , \7190 );
nor \U$10207 ( \10396 , \10394 , \10395 );
xnor \U$10208 ( \10397 , \10396 , \7198 );
xor \U$10209 ( \10398 , \10393 , \10397 );
and \U$10210 ( \10399 , \5854 , \7203 );
and \U$10211 ( \10400 , \5819 , \7201 );
nor \U$10212 ( \10401 , \10399 , \10400 );
xnor \U$10213 ( \10402 , \10401 , \6824 );
xor \U$10214 ( \10403 , \10398 , \10402 );
xor \U$10215 ( \10404 , \10389 , \10403 );
not \U$10216 ( \10405 , \7123 );
and \U$10217 ( \10406 , \5770 , \7140 );
and \U$10218 ( \10407 , \5737 , \7138 );
nor \U$10219 ( \10408 , \10406 , \10407 );
xnor \U$10220 ( \10409 , \10408 , \7146 );
xor \U$10221 ( \10410 , \10405 , \10409 );
and \U$10222 ( \10411 , \5792 , \7157 );
and \U$10223 ( \10412 , \5758 , \7155 );
nor \U$10224 ( \10413 , \10411 , \10412 );
xnor \U$10225 ( \10414 , \10413 , \7163 );
xor \U$10226 ( \10415 , \10410 , \10414 );
xor \U$10227 ( \10416 , \10404 , \10415 );
xor \U$10228 ( \10417 , \10375 , \10416 );
and \U$10229 ( \10418 , \6057 , \5935 );
and \U$10230 ( \10419 , \6029 , \5933 );
nor \U$10231 ( \10420 , \10418 , \10419 );
xnor \U$10232 ( \10421 , \10420 , \5942 );
and \U$10233 ( \10422 , \6065 , \5955 );
and \U$10234 ( \10423 , \6048 , \5953 );
nor \U$10235 ( \10424 , \10422 , \10423 );
xnor \U$10236 ( \10425 , \10424 , \5962 );
xor \U$10237 ( \10426 , \10421 , \10425 );
and \U$10238 ( \10427 , \5998 , \5871 );
and \U$10239 ( \10428 , \5967 , \5869 );
nor \U$10240 ( \10429 , \10427 , \10428 );
xnor \U$10241 ( \10430 , \10429 , \5878 );
and \U$10242 ( \10431 , \6018 , \5891 );
and \U$10243 ( \10432 , \5986 , \5889 );
nor \U$10244 ( \10433 , \10431 , \10432 );
xnor \U$10245 ( \10434 , \10433 , \5898 );
xor \U$10246 ( \10435 , \10430 , \10434 );
and \U$10247 ( \10436 , \6041 , \5916 );
and \U$10248 ( \10437 , \6006 , \5914 );
nor \U$10249 ( \10438 , \10436 , \10437 );
xnor \U$10250 ( \10439 , \10438 , \5923 );
xor \U$10251 ( \10440 , \10435 , \10439 );
xor \U$10252 ( \10441 , \10426 , \10440 );
and \U$10253 ( \10442 , \5937 , \5809 );
and \U$10254 ( \10443 , \5906 , \5807 );
nor \U$10255 ( \10444 , \10442 , \10443 );
xnor \U$10256 ( \10445 , \10444 , \5816 );
and \U$10257 ( \10446 , \5957 , \5829 );
and \U$10258 ( \10447 , \5925 , \5827 );
nor \U$10259 ( \10448 , \10446 , \10447 );
xnor \U$10260 ( \10449 , \10448 , \5836 );
xor \U$10261 ( \10450 , \10445 , \10449 );
and \U$10262 ( \10451 , \5979 , \5852 );
and \U$10263 ( \10452 , \5945 , \5850 );
nor \U$10264 ( \10453 , \10451 , \10452 );
xnor \U$10265 ( \10454 , \10453 , \5859 );
xor \U$10266 ( \10455 , \10450 , \10454 );
xor \U$10267 ( \10456 , \10441 , \10455 );
xor \U$10268 ( \10457 , \10417 , \10456 );
xor \U$10269 ( \10458 , \10371 , \10457 );
and \U$10270 ( \10459 , \10217 , \10221 );
and \U$10271 ( \10460 , \10221 , \10226 );
and \U$10272 ( \10461 , \10217 , \10226 );
or \U$10273 ( \10462 , \10459 , \10460 , \10461 );
and \U$10274 ( \10463 , \10205 , \10209 );
and \U$10275 ( \10464 , \10209 , \10211 );
and \U$10276 ( \10465 , \10205 , \10211 );
or \U$10277 ( \10466 , \10463 , \10464 , \10465 );
xor \U$10278 ( \10467 , \10462 , \10466 );
or \U$10279 ( \10468 , \10186 , \10200 );
xor \U$10280 ( \10469 , \10467 , \10468 );
xor \U$10281 ( \10470 , \10458 , \10469 );
xor \U$10282 ( \10471 , \10342 , \10470 );
xor \U$10283 ( \10472 , \10333 , \10471 );
and \U$10284 ( \10473 , \10153 , \10164 );
and \U$10285 ( \10474 , \10164 , \10304 );
and \U$10286 ( \10475 , \10153 , \10304 );
or \U$10287 ( \10476 , \10473 , \10474 , \10475 );
nor \U$10288 ( \10477 , \10472 , \10476 );
and \U$10289 ( \10478 , \10337 , \10341 );
and \U$10290 ( \10479 , \10341 , \10470 );
and \U$10291 ( \10480 , \10337 , \10470 );
or \U$10292 ( \10481 , \10478 , \10479 , \10480 );
and \U$10293 ( \10482 , \10462 , \10466 );
and \U$10294 ( \10483 , \10466 , \10468 );
and \U$10295 ( \10484 , \10462 , \10468 );
or \U$10296 ( \10485 , \10482 , \10483 , \10484 );
and \U$10297 ( \10486 , \10375 , \10416 );
and \U$10298 ( \10487 , \10416 , \10456 );
and \U$10299 ( \10488 , \10375 , \10456 );
or \U$10300 ( \10489 , \10486 , \10487 , \10488 );
xor \U$10301 ( \10490 , \10485 , \10489 );
and \U$10302 ( \10491 , \10356 , \10370 );
xor \U$10303 ( \10492 , \10490 , \10491 );
xor \U$10304 ( \10493 , \10481 , \10492 );
and \U$10305 ( \10494 , \10322 , \10326 );
and \U$10306 ( \10495 , \10326 , \10331 );
and \U$10307 ( \10496 , \10322 , \10331 );
or \U$10308 ( \10497 , \10494 , \10495 , \10496 );
and \U$10309 ( \10498 , \10371 , \10457 );
and \U$10310 ( \10499 , \10457 , \10469 );
and \U$10311 ( \10500 , \10371 , \10469 );
or \U$10312 ( \10501 , \10498 , \10499 , \10500 );
xor \U$10313 ( \10502 , \10497 , \10501 );
and \U$10314 ( \10503 , \6029 , \5935 );
and \U$10315 ( \10504 , \6041 , \5933 );
nor \U$10316 ( \10505 , \10503 , \10504 );
xnor \U$10317 ( \10506 , \10505 , \5942 );
and \U$10318 ( \10507 , \6048 , \5955 );
and \U$10319 ( \10508 , \6057 , \5953 );
nor \U$10320 ( \10509 , \10507 , \10508 );
xnor \U$10321 ( \10510 , \10509 , \5962 );
xor \U$10322 ( \10511 , \10506 , \10510 );
nand \U$10323 ( \10512 , \6065 , \5975 );
xnor \U$10324 ( \10513 , \10512 , \5984 );
xor \U$10325 ( \10514 , \10511 , \10513 );
and \U$10326 ( \10515 , \5967 , \5871 );
and \U$10327 ( \10516 , \5979 , \5869 );
nor \U$10328 ( \10517 , \10515 , \10516 );
xnor \U$10329 ( \10518 , \10517 , \5878 );
and \U$10330 ( \10519 , \5986 , \5891 );
and \U$10331 ( \10520 , \5998 , \5889 );
nor \U$10332 ( \10521 , \10519 , \10520 );
xnor \U$10333 ( \10522 , \10521 , \5898 );
xor \U$10334 ( \10523 , \10518 , \10522 );
and \U$10335 ( \10524 , \6006 , \5916 );
and \U$10336 ( \10525 , \6018 , \5914 );
nor \U$10337 ( \10526 , \10524 , \10525 );
xnor \U$10338 ( \10527 , \10526 , \5923 );
xor \U$10339 ( \10528 , \10523 , \10527 );
xnor \U$10340 ( \10529 , \10514 , \10528 );
and \U$10341 ( \10530 , \10445 , \10449 );
and \U$10342 ( \10531 , \10449 , \10454 );
and \U$10343 ( \10532 , \10445 , \10454 );
or \U$10344 ( \10533 , \10530 , \10531 , \10532 );
and \U$10345 ( \10534 , \10430 , \10434 );
and \U$10346 ( \10535 , \10434 , \10439 );
and \U$10347 ( \10536 , \10430 , \10439 );
or \U$10348 ( \10537 , \10534 , \10535 , \10536 );
xor \U$10349 ( \10538 , \10533 , \10537 );
and \U$10350 ( \10539 , \10421 , \10425 );
xor \U$10351 ( \10540 , \10538 , \10539 );
xor \U$10352 ( \10541 , \10529 , \10540 );
and \U$10353 ( \10542 , \10405 , \10409 );
and \U$10354 ( \10543 , \10409 , \10414 );
and \U$10355 ( \10544 , \10405 , \10414 );
or \U$10356 ( \10545 , \10542 , \10543 , \10544 );
and \U$10357 ( \10546 , \10393 , \10397 );
and \U$10358 ( \10547 , \10397 , \10402 );
and \U$10359 ( \10548 , \10393 , \10402 );
or \U$10360 ( \10549 , \10546 , \10547 , \10548 );
xor \U$10361 ( \10550 , \10545 , \10549 );
and \U$10362 ( \10551 , \10379 , \10383 );
and \U$10363 ( \10552 , \10383 , \10388 );
and \U$10364 ( \10553 , \10379 , \10388 );
or \U$10365 ( \10554 , \10551 , \10552 , \10553 );
xor \U$10366 ( \10555 , \10550 , \10554 );
xor \U$10367 ( \10556 , \10541 , \10555 );
and \U$10368 ( \10557 , \10389 , \10403 );
and \U$10369 ( \10558 , \10403 , \10415 );
and \U$10370 ( \10559 , \10389 , \10415 );
or \U$10371 ( \10560 , \10557 , \10558 , \10559 );
and \U$10372 ( \10561 , \5737 , \7140 );
not \U$10373 ( \10562 , \10561 );
xnor \U$10374 ( \10563 , \10562 , \7146 );
xor \U$10375 ( \10564 , \5984 , \10563 );
and \U$10376 ( \10565 , \5758 , \7157 );
and \U$10377 ( \10566 , \5770 , \7155 );
nor \U$10378 ( \10567 , \10565 , \10566 );
xnor \U$10379 ( \10568 , \10567 , \7163 );
xor \U$10380 ( \10569 , \10564 , \10568 );
xor \U$10381 ( \10570 , \10560 , \10569 );
and \U$10382 ( \10571 , \5906 , \5809 );
and \U$10383 ( \10572 , \5918 , \5807 );
nor \U$10384 ( \10573 , \10571 , \10572 );
xnor \U$10385 ( \10574 , \10573 , \5816 );
and \U$10386 ( \10575 , \5925 , \5829 );
and \U$10387 ( \10576 , \5937 , \5827 );
nor \U$10388 ( \10577 , \10575 , \10576 );
xnor \U$10389 ( \10578 , \10577 , \5836 );
xor \U$10390 ( \10579 , \10574 , \10578 );
and \U$10391 ( \10580 , \5945 , \5852 );
and \U$10392 ( \10581 , \5957 , \5850 );
nor \U$10393 ( \10582 , \10580 , \10581 );
xnor \U$10394 ( \10583 , \10582 , \5859 );
xor \U$10395 ( \10584 , \10579 , \10583 );
and \U$10396 ( \10585 , \5842 , \5750 );
and \U$10397 ( \10586 , \5854 , \5748 );
nor \U$10398 ( \10587 , \10585 , \10586 );
xnor \U$10399 ( \10588 , \10587 , \5755 );
and \U$10400 ( \10589 , \5861 , \5768 );
and \U$10401 ( \10590 , \5873 , \5766 );
nor \U$10402 ( \10591 , \10589 , \10590 );
xnor \U$10403 ( \10592 , \10591 , \5775 );
xor \U$10404 ( \10593 , \10588 , \10592 );
and \U$10405 ( \10594 , \5881 , \5790 );
and \U$10406 ( \10595 , \5893 , \5788 );
nor \U$10407 ( \10596 , \10594 , \10595 );
xnor \U$10408 ( \10597 , \10596 , \5797 );
xor \U$10409 ( \10598 , \10593 , \10597 );
xor \U$10410 ( \10599 , \10584 , \10598 );
and \U$10411 ( \10600 , \5780 , \7175 );
and \U$10412 ( \10601 , \5792 , \7173 );
nor \U$10413 ( \10602 , \10600 , \10601 );
xnor \U$10414 ( \10603 , \10602 , \7181 );
and \U$10415 ( \10604 , \5799 , \7192 );
and \U$10416 ( \10605 , \5811 , \7190 );
nor \U$10417 ( \10606 , \10604 , \10605 );
xnor \U$10418 ( \10607 , \10606 , \7198 );
xor \U$10419 ( \10608 , \10603 , \10607 );
and \U$10420 ( \10609 , \5819 , \7203 );
and \U$10421 ( \10610 , \5831 , \7201 );
nor \U$10422 ( \10611 , \10609 , \10610 );
xnor \U$10423 ( \10612 , \10611 , \6824 );
xor \U$10424 ( \10613 , \10608 , \10612 );
xor \U$10425 ( \10614 , \10599 , \10613 );
xor \U$10426 ( \10615 , \10570 , \10614 );
xor \U$10427 ( \10616 , \10556 , \10615 );
and \U$10428 ( \10617 , \10360 , \10364 );
and \U$10429 ( \10618 , \10364 , \10369 );
and \U$10430 ( \10619 , \10360 , \10369 );
or \U$10431 ( \10620 , \10617 , \10618 , \10619 );
and \U$10432 ( \10621 , \10346 , \10350 );
and \U$10433 ( \10622 , \10350 , \10355 );
and \U$10434 ( \10623 , \10346 , \10355 );
or \U$10435 ( \10624 , \10621 , \10622 , \10623 );
xor \U$10436 ( \10625 , \10620 , \10624 );
and \U$10437 ( \10626 , \10426 , \10440 );
and \U$10438 ( \10627 , \10440 , \10455 );
and \U$10439 ( \10628 , \10426 , \10455 );
or \U$10440 ( \10629 , \10626 , \10627 , \10628 );
xor \U$10441 ( \10630 , \10625 , \10629 );
xor \U$10442 ( \10631 , \10616 , \10630 );
xor \U$10443 ( \10632 , \10502 , \10631 );
xor \U$10444 ( \10633 , \10493 , \10632 );
and \U$10445 ( \10634 , \10318 , \10332 );
and \U$10446 ( \10635 , \10332 , \10471 );
and \U$10447 ( \10636 , \10318 , \10471 );
or \U$10448 ( \10637 , \10634 , \10635 , \10636 );
nor \U$10449 ( \10638 , \10633 , \10637 );
nor \U$10450 ( \10639 , \10477 , \10638 );
and \U$10451 ( \10640 , \10497 , \10501 );
and \U$10452 ( \10641 , \10501 , \10631 );
and \U$10453 ( \10642 , \10497 , \10631 );
or \U$10454 ( \10643 , \10640 , \10641 , \10642 );
and \U$10455 ( \10644 , \10620 , \10624 );
and \U$10456 ( \10645 , \10624 , \10629 );
and \U$10457 ( \10646 , \10620 , \10629 );
or \U$10458 ( \10647 , \10644 , \10645 , \10646 );
and \U$10459 ( \10648 , \10560 , \10569 );
and \U$10460 ( \10649 , \10569 , \10614 );
and \U$10461 ( \10650 , \10560 , \10614 );
or \U$10462 ( \10651 , \10648 , \10649 , \10650 );
xor \U$10463 ( \10652 , \10647 , \10651 );
and \U$10464 ( \10653 , \10529 , \10540 );
and \U$10465 ( \10654 , \10540 , \10555 );
and \U$10466 ( \10655 , \10529 , \10555 );
or \U$10467 ( \10656 , \10653 , \10654 , \10655 );
xor \U$10468 ( \10657 , \10652 , \10656 );
xor \U$10469 ( \10658 , \10643 , \10657 );
and \U$10470 ( \10659 , \10485 , \10489 );
and \U$10471 ( \10660 , \10489 , \10491 );
and \U$10472 ( \10661 , \10485 , \10491 );
or \U$10473 ( \10662 , \10659 , \10660 , \10661 );
and \U$10474 ( \10663 , \10556 , \10615 );
and \U$10475 ( \10664 , \10615 , \10630 );
and \U$10476 ( \10665 , \10556 , \10630 );
or \U$10477 ( \10666 , \10663 , \10664 , \10665 );
xor \U$10478 ( \10667 , \10662 , \10666 );
and \U$10479 ( \10668 , \10574 , \10578 );
and \U$10480 ( \10669 , \10578 , \10583 );
and \U$10481 ( \10670 , \10574 , \10583 );
or \U$10482 ( \10671 , \10668 , \10669 , \10670 );
and \U$10483 ( \10672 , \10518 , \10522 );
and \U$10484 ( \10673 , \10522 , \10527 );
and \U$10485 ( \10674 , \10518 , \10527 );
or \U$10486 ( \10675 , \10672 , \10673 , \10674 );
xor \U$10487 ( \10676 , \10671 , \10675 );
and \U$10488 ( \10677 , \10506 , \10510 );
and \U$10489 ( \10678 , \10510 , \10513 );
and \U$10490 ( \10679 , \10506 , \10513 );
or \U$10491 ( \10680 , \10677 , \10678 , \10679 );
xor \U$10492 ( \10681 , \10676 , \10680 );
and \U$10493 ( \10682 , \5984 , \10563 );
and \U$10494 ( \10683 , \10563 , \10568 );
and \U$10495 ( \10684 , \5984 , \10568 );
or \U$10496 ( \10685 , \10682 , \10683 , \10684 );
and \U$10497 ( \10686 , \10603 , \10607 );
and \U$10498 ( \10687 , \10607 , \10612 );
and \U$10499 ( \10688 , \10603 , \10612 );
or \U$10500 ( \10689 , \10686 , \10687 , \10688 );
xor \U$10501 ( \10690 , \10685 , \10689 );
and \U$10502 ( \10691 , \10588 , \10592 );
and \U$10503 ( \10692 , \10592 , \10597 );
and \U$10504 ( \10693 , \10588 , \10597 );
or \U$10505 ( \10694 , \10691 , \10692 , \10693 );
xor \U$10506 ( \10695 , \10690 , \10694 );
xor \U$10507 ( \10696 , \10681 , \10695 );
and \U$10508 ( \10697 , \10584 , \10598 );
and \U$10509 ( \10698 , \10598 , \10613 );
and \U$10510 ( \10699 , \10584 , \10613 );
or \U$10511 ( \10700 , \10697 , \10698 , \10699 );
and \U$10512 ( \10701 , \5873 , \5768 );
and \U$10513 ( \10702 , \5842 , \5766 );
nor \U$10514 ( \10703 , \10701 , \10702 );
xnor \U$10515 ( \10704 , \10703 , \5775 );
and \U$10516 ( \10705 , \5893 , \5790 );
and \U$10517 ( \10706 , \5861 , \5788 );
nor \U$10518 ( \10707 , \10705 , \10706 );
xnor \U$10519 ( \10708 , \10707 , \5797 );
xor \U$10520 ( \10709 , \10704 , \10708 );
and \U$10521 ( \10710 , \5918 , \5809 );
and \U$10522 ( \10711 , \5881 , \5807 );
nor \U$10523 ( \10712 , \10710 , \10711 );
xnor \U$10524 ( \10713 , \10712 , \5816 );
xor \U$10525 ( \10714 , \10709 , \10713 );
and \U$10526 ( \10715 , \5811 , \7192 );
and \U$10527 ( \10716 , \5780 , \7190 );
nor \U$10528 ( \10717 , \10715 , \10716 );
xnor \U$10529 ( \10718 , \10717 , \7198 );
and \U$10530 ( \10719 , \5831 , \7203 );
and \U$10531 ( \10720 , \5799 , \7201 );
nor \U$10532 ( \10721 , \10719 , \10720 );
xnor \U$10533 ( \10722 , \10721 , \6824 );
xor \U$10534 ( \10723 , \10718 , \10722 );
and \U$10535 ( \10724 , \5854 , \5750 );
and \U$10536 ( \10725 , \5819 , \5748 );
nor \U$10537 ( \10726 , \10724 , \10725 );
xnor \U$10538 ( \10727 , \10726 , \5755 );
xor \U$10539 ( \10728 , \10723 , \10727 );
xor \U$10540 ( \10729 , \10714 , \10728 );
not \U$10541 ( \10730 , \7146 );
and \U$10542 ( \10731 , \5770 , \7157 );
and \U$10543 ( \10732 , \5737 , \7155 );
nor \U$10544 ( \10733 , \10731 , \10732 );
xnor \U$10545 ( \10734 , \10733 , \7163 );
xor \U$10546 ( \10735 , \10730 , \10734 );
and \U$10547 ( \10736 , \5792 , \7175 );
and \U$10548 ( \10737 , \5758 , \7173 );
nor \U$10549 ( \10738 , \10736 , \10737 );
xnor \U$10550 ( \10739 , \10738 , \7181 );
xor \U$10551 ( \10740 , \10735 , \10739 );
xor \U$10552 ( \10741 , \10729 , \10740 );
xor \U$10553 ( \10742 , \10700 , \10741 );
and \U$10554 ( \10743 , \6057 , \5955 );
and \U$10555 ( \10744 , \6029 , \5953 );
nor \U$10556 ( \10745 , \10743 , \10744 );
xnor \U$10557 ( \10746 , \10745 , \5962 );
and \U$10558 ( \10747 , \6065 , \5977 );
and \U$10559 ( \10748 , \6048 , \5975 );
nor \U$10560 ( \10749 , \10747 , \10748 );
xnor \U$10561 ( \10750 , \10749 , \5984 );
xor \U$10562 ( \10751 , \10746 , \10750 );
and \U$10563 ( \10752 , \5998 , \5891 );
and \U$10564 ( \10753 , \5967 , \5889 );
nor \U$10565 ( \10754 , \10752 , \10753 );
xnor \U$10566 ( \10755 , \10754 , \5898 );
and \U$10567 ( \10756 , \6018 , \5916 );
and \U$10568 ( \10757 , \5986 , \5914 );
nor \U$10569 ( \10758 , \10756 , \10757 );
xnor \U$10570 ( \10759 , \10758 , \5923 );
xor \U$10571 ( \10760 , \10755 , \10759 );
and \U$10572 ( \10761 , \6041 , \5935 );
and \U$10573 ( \10762 , \6006 , \5933 );
nor \U$10574 ( \10763 , \10761 , \10762 );
xnor \U$10575 ( \10764 , \10763 , \5942 );
xor \U$10576 ( \10765 , \10760 , \10764 );
xor \U$10577 ( \10766 , \10751 , \10765 );
and \U$10578 ( \10767 , \5937 , \5829 );
and \U$10579 ( \10768 , \5906 , \5827 );
nor \U$10580 ( \10769 , \10767 , \10768 );
xnor \U$10581 ( \10770 , \10769 , \5836 );
and \U$10582 ( \10771 , \5957 , \5852 );
and \U$10583 ( \10772 , \5925 , \5850 );
nor \U$10584 ( \10773 , \10771 , \10772 );
xnor \U$10585 ( \10774 , \10773 , \5859 );
xor \U$10586 ( \10775 , \10770 , \10774 );
and \U$10587 ( \10776 , \5979 , \5871 );
and \U$10588 ( \10777 , \5945 , \5869 );
nor \U$10589 ( \10778 , \10776 , \10777 );
xnor \U$10590 ( \10779 , \10778 , \5878 );
xor \U$10591 ( \10780 , \10775 , \10779 );
xor \U$10592 ( \10781 , \10766 , \10780 );
xor \U$10593 ( \10782 , \10742 , \10781 );
xor \U$10594 ( \10783 , \10696 , \10782 );
and \U$10595 ( \10784 , \10545 , \10549 );
and \U$10596 ( \10785 , \10549 , \10554 );
and \U$10597 ( \10786 , \10545 , \10554 );
or \U$10598 ( \10787 , \10784 , \10785 , \10786 );
and \U$10599 ( \10788 , \10533 , \10537 );
and \U$10600 ( \10789 , \10537 , \10539 );
and \U$10601 ( \10790 , \10533 , \10539 );
or \U$10602 ( \10791 , \10788 , \10789 , \10790 );
xor \U$10603 ( \10792 , \10787 , \10791 );
or \U$10604 ( \10793 , \10514 , \10528 );
xor \U$10605 ( \10794 , \10792 , \10793 );
xor \U$10606 ( \10795 , \10783 , \10794 );
xor \U$10607 ( \10796 , \10667 , \10795 );
xor \U$10608 ( \10797 , \10658 , \10796 );
and \U$10609 ( \10798 , \10481 , \10492 );
and \U$10610 ( \10799 , \10492 , \10632 );
and \U$10611 ( \10800 , \10481 , \10632 );
or \U$10612 ( \10801 , \10798 , \10799 , \10800 );
nor \U$10613 ( \10802 , \10797 , \10801 );
and \U$10614 ( \10803 , \10662 , \10666 );
and \U$10615 ( \10804 , \10666 , \10795 );
and \U$10616 ( \10805 , \10662 , \10795 );
or \U$10617 ( \10806 , \10803 , \10804 , \10805 );
and \U$10618 ( \10807 , \10787 , \10791 );
and \U$10619 ( \10808 , \10791 , \10793 );
and \U$10620 ( \10809 , \10787 , \10793 );
or \U$10621 ( \10810 , \10807 , \10808 , \10809 );
and \U$10622 ( \10811 , \10700 , \10741 );
and \U$10623 ( \10812 , \10741 , \10781 );
and \U$10624 ( \10813 , \10700 , \10781 );
or \U$10625 ( \10814 , \10811 , \10812 , \10813 );
xor \U$10626 ( \10815 , \10810 , \10814 );
and \U$10627 ( \10816 , \10681 , \10695 );
xor \U$10628 ( \10817 , \10815 , \10816 );
xor \U$10629 ( \10818 , \10806 , \10817 );
and \U$10630 ( \10819 , \10647 , \10651 );
and \U$10631 ( \10820 , \10651 , \10656 );
and \U$10632 ( \10821 , \10647 , \10656 );
or \U$10633 ( \10822 , \10819 , \10820 , \10821 );
and \U$10634 ( \10823 , \10696 , \10782 );
and \U$10635 ( \10824 , \10782 , \10794 );
and \U$10636 ( \10825 , \10696 , \10794 );
or \U$10637 ( \10826 , \10823 , \10824 , \10825 );
xor \U$10638 ( \10827 , \10822 , \10826 );
and \U$10639 ( \10828 , \6029 , \5955 );
and \U$10640 ( \10829 , \6041 , \5953 );
nor \U$10641 ( \10830 , \10828 , \10829 );
xnor \U$10642 ( \10831 , \10830 , \5962 );
and \U$10643 ( \10832 , \6048 , \5977 );
and \U$10644 ( \10833 , \6057 , \5975 );
nor \U$10645 ( \10834 , \10832 , \10833 );
xnor \U$10646 ( \10835 , \10834 , \5984 );
xor \U$10647 ( \10836 , \10831 , \10835 );
nand \U$10648 ( \10837 , \6065 , \5994 );
xnor \U$10649 ( \10838 , \10837 , \6003 );
xor \U$10650 ( \10839 , \10836 , \10838 );
and \U$10651 ( \10840 , \5967 , \5891 );
and \U$10652 ( \10841 , \5979 , \5889 );
nor \U$10653 ( \10842 , \10840 , \10841 );
xnor \U$10654 ( \10843 , \10842 , \5898 );
and \U$10655 ( \10844 , \5986 , \5916 );
and \U$10656 ( \10845 , \5998 , \5914 );
nor \U$10657 ( \10846 , \10844 , \10845 );
xnor \U$10658 ( \10847 , \10846 , \5923 );
xor \U$10659 ( \10848 , \10843 , \10847 );
and \U$10660 ( \10849 , \6006 , \5935 );
and \U$10661 ( \10850 , \6018 , \5933 );
nor \U$10662 ( \10851 , \10849 , \10850 );
xnor \U$10663 ( \10852 , \10851 , \5942 );
xor \U$10664 ( \10853 , \10848 , \10852 );
xnor \U$10665 ( \10854 , \10839 , \10853 );
and \U$10666 ( \10855 , \10770 , \10774 );
and \U$10667 ( \10856 , \10774 , \10779 );
and \U$10668 ( \10857 , \10770 , \10779 );
or \U$10669 ( \10858 , \10855 , \10856 , \10857 );
and \U$10670 ( \10859 , \10755 , \10759 );
and \U$10671 ( \10860 , \10759 , \10764 );
and \U$10672 ( \10861 , \10755 , \10764 );
or \U$10673 ( \10862 , \10859 , \10860 , \10861 );
xor \U$10674 ( \10863 , \10858 , \10862 );
and \U$10675 ( \10864 , \10746 , \10750 );
xor \U$10676 ( \10865 , \10863 , \10864 );
xor \U$10677 ( \10866 , \10854 , \10865 );
and \U$10678 ( \10867 , \10730 , \10734 );
and \U$10679 ( \10868 , \10734 , \10739 );
and \U$10680 ( \10869 , \10730 , \10739 );
or \U$10681 ( \10870 , \10867 , \10868 , \10869 );
and \U$10682 ( \10871 , \10718 , \10722 );
and \U$10683 ( \10872 , \10722 , \10727 );
and \U$10684 ( \10873 , \10718 , \10727 );
or \U$10685 ( \10874 , \10871 , \10872 , \10873 );
xor \U$10686 ( \10875 , \10870 , \10874 );
and \U$10687 ( \10876 , \10704 , \10708 );
and \U$10688 ( \10877 , \10708 , \10713 );
and \U$10689 ( \10878 , \10704 , \10713 );
or \U$10690 ( \10879 , \10876 , \10877 , \10878 );
xor \U$10691 ( \10880 , \10875 , \10879 );
xor \U$10692 ( \10881 , \10866 , \10880 );
and \U$10693 ( \10882 , \10714 , \10728 );
and \U$10694 ( \10883 , \10728 , \10740 );
and \U$10695 ( \10884 , \10714 , \10740 );
or \U$10696 ( \10885 , \10882 , \10883 , \10884 );
and \U$10697 ( \10886 , \5737 , \7157 );
not \U$10698 ( \10887 , \10886 );
xnor \U$10699 ( \10888 , \10887 , \7163 );
xor \U$10700 ( \10889 , \6003 , \10888 );
and \U$10701 ( \10890 , \5758 , \7175 );
and \U$10702 ( \10891 , \5770 , \7173 );
nor \U$10703 ( \10892 , \10890 , \10891 );
xnor \U$10704 ( \10893 , \10892 , \7181 );
xor \U$10705 ( \10894 , \10889 , \10893 );
xor \U$10706 ( \10895 , \10885 , \10894 );
and \U$10707 ( \10896 , \5906 , \5829 );
and \U$10708 ( \10897 , \5918 , \5827 );
nor \U$10709 ( \10898 , \10896 , \10897 );
xnor \U$10710 ( \10899 , \10898 , \5836 );
and \U$10711 ( \10900 , \5925 , \5852 );
and \U$10712 ( \10901 , \5937 , \5850 );
nor \U$10713 ( \10902 , \10900 , \10901 );
xnor \U$10714 ( \10903 , \10902 , \5859 );
xor \U$10715 ( \10904 , \10899 , \10903 );
and \U$10716 ( \10905 , \5945 , \5871 );
and \U$10717 ( \10906 , \5957 , \5869 );
nor \U$10718 ( \10907 , \10905 , \10906 );
xnor \U$10719 ( \10908 , \10907 , \5878 );
xor \U$10720 ( \10909 , \10904 , \10908 );
and \U$10721 ( \10910 , \5842 , \5768 );
and \U$10722 ( \10911 , \5854 , \5766 );
nor \U$10723 ( \10912 , \10910 , \10911 );
xnor \U$10724 ( \10913 , \10912 , \5775 );
and \U$10725 ( \10914 , \5861 , \5790 );
and \U$10726 ( \10915 , \5873 , \5788 );
nor \U$10727 ( \10916 , \10914 , \10915 );
xnor \U$10728 ( \10917 , \10916 , \5797 );
xor \U$10729 ( \10918 , \10913 , \10917 );
and \U$10730 ( \10919 , \5881 , \5809 );
and \U$10731 ( \10920 , \5893 , \5807 );
nor \U$10732 ( \10921 , \10919 , \10920 );
xnor \U$10733 ( \10922 , \10921 , \5816 );
xor \U$10734 ( \10923 , \10918 , \10922 );
xor \U$10735 ( \10924 , \10909 , \10923 );
and \U$10736 ( \10925 , \5780 , \7192 );
and \U$10737 ( \10926 , \5792 , \7190 );
nor \U$10738 ( \10927 , \10925 , \10926 );
xnor \U$10739 ( \10928 , \10927 , \7198 );
and \U$10740 ( \10929 , \5799 , \7203 );
and \U$10741 ( \10930 , \5811 , \7201 );
nor \U$10742 ( \10931 , \10929 , \10930 );
xnor \U$10743 ( \10932 , \10931 , \6824 );
xor \U$10744 ( \10933 , \10928 , \10932 );
and \U$10745 ( \10934 , \5819 , \5750 );
and \U$10746 ( \10935 , \5831 , \5748 );
nor \U$10747 ( \10936 , \10934 , \10935 );
xnor \U$10748 ( \10937 , \10936 , \5755 );
xor \U$10749 ( \10938 , \10933 , \10937 );
xor \U$10750 ( \10939 , \10924 , \10938 );
xor \U$10751 ( \10940 , \10895 , \10939 );
xor \U$10752 ( \10941 , \10881 , \10940 );
and \U$10753 ( \10942 , \10685 , \10689 );
and \U$10754 ( \10943 , \10689 , \10694 );
and \U$10755 ( \10944 , \10685 , \10694 );
or \U$10756 ( \10945 , \10942 , \10943 , \10944 );
and \U$10757 ( \10946 , \10671 , \10675 );
and \U$10758 ( \10947 , \10675 , \10680 );
and \U$10759 ( \10948 , \10671 , \10680 );
or \U$10760 ( \10949 , \10946 , \10947 , \10948 );
xor \U$10761 ( \10950 , \10945 , \10949 );
and \U$10762 ( \10951 , \10751 , \10765 );
and \U$10763 ( \10952 , \10765 , \10780 );
and \U$10764 ( \10953 , \10751 , \10780 );
or \U$10765 ( \10954 , \10951 , \10952 , \10953 );
xor \U$10766 ( \10955 , \10950 , \10954 );
xor \U$10767 ( \10956 , \10941 , \10955 );
xor \U$10768 ( \10957 , \10827 , \10956 );
xor \U$10769 ( \10958 , \10818 , \10957 );
and \U$10770 ( \10959 , \10643 , \10657 );
and \U$10771 ( \10960 , \10657 , \10796 );
and \U$10772 ( \10961 , \10643 , \10796 );
or \U$10773 ( \10962 , \10959 , \10960 , \10961 );
nor \U$10774 ( \10963 , \10958 , \10962 );
nor \U$10775 ( \10964 , \10802 , \10963 );
nand \U$10776 ( \10965 , \10639 , \10964 );
and \U$10777 ( \10966 , \10822 , \10826 );
and \U$10778 ( \10967 , \10826 , \10956 );
and \U$10779 ( \10968 , \10822 , \10956 );
or \U$10780 ( \10969 , \10966 , \10967 , \10968 );
and \U$10781 ( \10970 , \10945 , \10949 );
and \U$10782 ( \10971 , \10949 , \10954 );
and \U$10783 ( \10972 , \10945 , \10954 );
or \U$10784 ( \10973 , \10970 , \10971 , \10972 );
and \U$10785 ( \10974 , \10885 , \10894 );
and \U$10786 ( \10975 , \10894 , \10939 );
and \U$10787 ( \10976 , \10885 , \10939 );
or \U$10788 ( \10977 , \10974 , \10975 , \10976 );
xor \U$10789 ( \10978 , \10973 , \10977 );
and \U$10790 ( \10979 , \10854 , \10865 );
and \U$10791 ( \10980 , \10865 , \10880 );
and \U$10792 ( \10981 , \10854 , \10880 );
or \U$10793 ( \10982 , \10979 , \10980 , \10981 );
xor \U$10794 ( \10983 , \10978 , \10982 );
xor \U$10795 ( \10984 , \10969 , \10983 );
and \U$10796 ( \10985 , \10810 , \10814 );
and \U$10797 ( \10986 , \10814 , \10816 );
and \U$10798 ( \10987 , \10810 , \10816 );
or \U$10799 ( \10988 , \10985 , \10986 , \10987 );
and \U$10800 ( \10989 , \10881 , \10940 );
and \U$10801 ( \10990 , \10940 , \10955 );
and \U$10802 ( \10991 , \10881 , \10955 );
or \U$10803 ( \10992 , \10989 , \10990 , \10991 );
xor \U$10804 ( \10993 , \10988 , \10992 );
and \U$10805 ( \10994 , \10899 , \10903 );
and \U$10806 ( \10995 , \10903 , \10908 );
and \U$10807 ( \10996 , \10899 , \10908 );
or \U$10808 ( \10997 , \10994 , \10995 , \10996 );
and \U$10809 ( \10998 , \10843 , \10847 );
and \U$10810 ( \10999 , \10847 , \10852 );
and \U$10811 ( \11000 , \10843 , \10852 );
or \U$10812 ( \11001 , \10998 , \10999 , \11000 );
xor \U$10813 ( \11002 , \10997 , \11001 );
and \U$10814 ( \11003 , \10831 , \10835 );
and \U$10815 ( \11004 , \10835 , \10838 );
and \U$10816 ( \11005 , \10831 , \10838 );
or \U$10817 ( \11006 , \11003 , \11004 , \11005 );
xor \U$10818 ( \11007 , \11002 , \11006 );
and \U$10819 ( \11008 , \6003 , \10888 );
and \U$10820 ( \11009 , \10888 , \10893 );
and \U$10821 ( \11010 , \6003 , \10893 );
or \U$10822 ( \11011 , \11008 , \11009 , \11010 );
and \U$10823 ( \11012 , \10928 , \10932 );
and \U$10824 ( \11013 , \10932 , \10937 );
and \U$10825 ( \11014 , \10928 , \10937 );
or \U$10826 ( \11015 , \11012 , \11013 , \11014 );
xor \U$10827 ( \11016 , \11011 , \11015 );
and \U$10828 ( \11017 , \10913 , \10917 );
and \U$10829 ( \11018 , \10917 , \10922 );
and \U$10830 ( \11019 , \10913 , \10922 );
or \U$10831 ( \11020 , \11017 , \11018 , \11019 );
xor \U$10832 ( \11021 , \11016 , \11020 );
xor \U$10833 ( \11022 , \11007 , \11021 );
and \U$10834 ( \11023 , \10909 , \10923 );
and \U$10835 ( \11024 , \10923 , \10938 );
and \U$10836 ( \11025 , \10909 , \10938 );
or \U$10837 ( \11026 , \11023 , \11024 , \11025 );
and \U$10838 ( \11027 , \5873 , \5790 );
and \U$10839 ( \11028 , \5842 , \5788 );
nor \U$10840 ( \11029 , \11027 , \11028 );
xnor \U$10841 ( \11030 , \11029 , \5797 );
and \U$10842 ( \11031 , \5893 , \5809 );
and \U$10843 ( \11032 , \5861 , \5807 );
nor \U$10844 ( \11033 , \11031 , \11032 );
xnor \U$10845 ( \11034 , \11033 , \5816 );
xor \U$10846 ( \11035 , \11030 , \11034 );
and \U$10847 ( \11036 , \5918 , \5829 );
and \U$10848 ( \11037 , \5881 , \5827 );
nor \U$10849 ( \11038 , \11036 , \11037 );
xnor \U$10850 ( \11039 , \11038 , \5836 );
xor \U$10851 ( \11040 , \11035 , \11039 );
and \U$10852 ( \11041 , \5811 , \7203 );
and \U$10853 ( \11042 , \5780 , \7201 );
nor \U$10854 ( \11043 , \11041 , \11042 );
xnor \U$10855 ( \11044 , \11043 , \6824 );
and \U$10856 ( \11045 , \5831 , \5750 );
and \U$10857 ( \11046 , \5799 , \5748 );
nor \U$10858 ( \11047 , \11045 , \11046 );
xnor \U$10859 ( \11048 , \11047 , \5755 );
xor \U$10860 ( \11049 , \11044 , \11048 );
and \U$10861 ( \11050 , \5854 , \5768 );
and \U$10862 ( \11051 , \5819 , \5766 );
nor \U$10863 ( \11052 , \11050 , \11051 );
xnor \U$10864 ( \11053 , \11052 , \5775 );
xor \U$10865 ( \11054 , \11049 , \11053 );
xor \U$10866 ( \11055 , \11040 , \11054 );
not \U$10867 ( \11056 , \7163 );
and \U$10868 ( \11057 , \5770 , \7175 );
and \U$10869 ( \11058 , \5737 , \7173 );
nor \U$10870 ( \11059 , \11057 , \11058 );
xnor \U$10871 ( \11060 , \11059 , \7181 );
xor \U$10872 ( \11061 , \11056 , \11060 );
and \U$10873 ( \11062 , \5792 , \7192 );
and \U$10874 ( \11063 , \5758 , \7190 );
nor \U$10875 ( \11064 , \11062 , \11063 );
xnor \U$10876 ( \11065 , \11064 , \7198 );
xor \U$10877 ( \11066 , \11061 , \11065 );
xor \U$10878 ( \11067 , \11055 , \11066 );
xor \U$10879 ( \11068 , \11026 , \11067 );
and \U$10880 ( \11069 , \6057 , \5977 );
and \U$10881 ( \11070 , \6029 , \5975 );
nor \U$10882 ( \11071 , \11069 , \11070 );
xnor \U$10883 ( \11072 , \11071 , \5984 );
and \U$10884 ( \11073 , \6065 , \5996 );
and \U$10885 ( \11074 , \6048 , \5994 );
nor \U$10886 ( \11075 , \11073 , \11074 );
xnor \U$10887 ( \11076 , \11075 , \6003 );
xor \U$10888 ( \11077 , \11072 , \11076 );
and \U$10889 ( \11078 , \5998 , \5916 );
and \U$10890 ( \11079 , \5967 , \5914 );
nor \U$10891 ( \11080 , \11078 , \11079 );
xnor \U$10892 ( \11081 , \11080 , \5923 );
and \U$10893 ( \11082 , \6018 , \5935 );
and \U$10894 ( \11083 , \5986 , \5933 );
nor \U$10895 ( \11084 , \11082 , \11083 );
xnor \U$10896 ( \11085 , \11084 , \5942 );
xor \U$10897 ( \11086 , \11081 , \11085 );
and \U$10898 ( \11087 , \6041 , \5955 );
and \U$10899 ( \11088 , \6006 , \5953 );
nor \U$10900 ( \11089 , \11087 , \11088 );
xnor \U$10901 ( \11090 , \11089 , \5962 );
xor \U$10902 ( \11091 , \11086 , \11090 );
xor \U$10903 ( \11092 , \11077 , \11091 );
and \U$10904 ( \11093 , \5937 , \5852 );
and \U$10905 ( \11094 , \5906 , \5850 );
nor \U$10906 ( \11095 , \11093 , \11094 );
xnor \U$10907 ( \11096 , \11095 , \5859 );
and \U$10908 ( \11097 , \5957 , \5871 );
and \U$10909 ( \11098 , \5925 , \5869 );
nor \U$10910 ( \11099 , \11097 , \11098 );
xnor \U$10911 ( \11100 , \11099 , \5878 );
xor \U$10912 ( \11101 , \11096 , \11100 );
and \U$10913 ( \11102 , \5979 , \5891 );
and \U$10914 ( \11103 , \5945 , \5889 );
nor \U$10915 ( \11104 , \11102 , \11103 );
xnor \U$10916 ( \11105 , \11104 , \5898 );
xor \U$10917 ( \11106 , \11101 , \11105 );
xor \U$10918 ( \11107 , \11092 , \11106 );
xor \U$10919 ( \11108 , \11068 , \11107 );
xor \U$10920 ( \11109 , \11022 , \11108 );
and \U$10921 ( \11110 , \10870 , \10874 );
and \U$10922 ( \11111 , \10874 , \10879 );
and \U$10923 ( \11112 , \10870 , \10879 );
or \U$10924 ( \11113 , \11110 , \11111 , \11112 );
and \U$10925 ( \11114 , \10858 , \10862 );
and \U$10926 ( \11115 , \10862 , \10864 );
and \U$10927 ( \11116 , \10858 , \10864 );
or \U$10928 ( \11117 , \11114 , \11115 , \11116 );
xor \U$10929 ( \11118 , \11113 , \11117 );
or \U$10930 ( \11119 , \10839 , \10853 );
xor \U$10931 ( \11120 , \11118 , \11119 );
xor \U$10932 ( \11121 , \11109 , \11120 );
xor \U$10933 ( \11122 , \10993 , \11121 );
xor \U$10934 ( \11123 , \10984 , \11122 );
and \U$10935 ( \11124 , \10806 , \10817 );
and \U$10936 ( \11125 , \10817 , \10957 );
and \U$10937 ( \11126 , \10806 , \10957 );
or \U$10938 ( \11127 , \11124 , \11125 , \11126 );
nor \U$10939 ( \11128 , \11123 , \11127 );
and \U$10940 ( \11129 , \10988 , \10992 );
and \U$10941 ( \11130 , \10992 , \11121 );
and \U$10942 ( \11131 , \10988 , \11121 );
or \U$10943 ( \11132 , \11129 , \11130 , \11131 );
and \U$10944 ( \11133 , \11113 , \11117 );
and \U$10945 ( \11134 , \11117 , \11119 );
and \U$10946 ( \11135 , \11113 , \11119 );
or \U$10947 ( \11136 , \11133 , \11134 , \11135 );
and \U$10948 ( \11137 , \11026 , \11067 );
and \U$10949 ( \11138 , \11067 , \11107 );
and \U$10950 ( \11139 , \11026 , \11107 );
or \U$10951 ( \11140 , \11137 , \11138 , \11139 );
xor \U$10952 ( \11141 , \11136 , \11140 );
and \U$10953 ( \11142 , \11007 , \11021 );
xor \U$10954 ( \11143 , \11141 , \11142 );
xor \U$10955 ( \11144 , \11132 , \11143 );
and \U$10956 ( \11145 , \10973 , \10977 );
and \U$10957 ( \11146 , \10977 , \10982 );
and \U$10958 ( \11147 , \10973 , \10982 );
or \U$10959 ( \11148 , \11145 , \11146 , \11147 );
and \U$10960 ( \11149 , \11022 , \11108 );
and \U$10961 ( \11150 , \11108 , \11120 );
and \U$10962 ( \11151 , \11022 , \11120 );
or \U$10963 ( \11152 , \11149 , \11150 , \11151 );
xor \U$10964 ( \11153 , \11148 , \11152 );
and \U$10965 ( \11154 , \6029 , \5977 );
and \U$10966 ( \11155 , \6041 , \5975 );
nor \U$10967 ( \11156 , \11154 , \11155 );
xnor \U$10968 ( \11157 , \11156 , \5984 );
and \U$10969 ( \11158 , \6048 , \5996 );
and \U$10970 ( \11159 , \6057 , \5994 );
nor \U$10971 ( \11160 , \11158 , \11159 );
xnor \U$10972 ( \11161 , \11160 , \6003 );
xor \U$10973 ( \11162 , \11157 , \11161 );
nand \U$10974 ( \11163 , \6065 , \6014 );
xnor \U$10975 ( \11164 , \11163 , \6023 );
xor \U$10976 ( \11165 , \11162 , \11164 );
and \U$10977 ( \11166 , \5967 , \5916 );
and \U$10978 ( \11167 , \5979 , \5914 );
nor \U$10979 ( \11168 , \11166 , \11167 );
xnor \U$10980 ( \11169 , \11168 , \5923 );
and \U$10981 ( \11170 , \5986 , \5935 );
and \U$10982 ( \11171 , \5998 , \5933 );
nor \U$10983 ( \11172 , \11170 , \11171 );
xnor \U$10984 ( \11173 , \11172 , \5942 );
xor \U$10985 ( \11174 , \11169 , \11173 );
and \U$10986 ( \11175 , \6006 , \5955 );
and \U$10987 ( \11176 , \6018 , \5953 );
nor \U$10988 ( \11177 , \11175 , \11176 );
xnor \U$10989 ( \11178 , \11177 , \5962 );
xor \U$10990 ( \11179 , \11174 , \11178 );
xnor \U$10991 ( \11180 , \11165 , \11179 );
and \U$10992 ( \11181 , \11096 , \11100 );
and \U$10993 ( \11182 , \11100 , \11105 );
and \U$10994 ( \11183 , \11096 , \11105 );
or \U$10995 ( \11184 , \11181 , \11182 , \11183 );
and \U$10996 ( \11185 , \11081 , \11085 );
and \U$10997 ( \11186 , \11085 , \11090 );
and \U$10998 ( \11187 , \11081 , \11090 );
or \U$10999 ( \11188 , \11185 , \11186 , \11187 );
xor \U$11000 ( \11189 , \11184 , \11188 );
and \U$11001 ( \11190 , \11072 , \11076 );
xor \U$11002 ( \11191 , \11189 , \11190 );
xor \U$11003 ( \11192 , \11180 , \11191 );
and \U$11004 ( \11193 , \11056 , \11060 );
and \U$11005 ( \11194 , \11060 , \11065 );
and \U$11006 ( \11195 , \11056 , \11065 );
or \U$11007 ( \11196 , \11193 , \11194 , \11195 );
and \U$11008 ( \11197 , \11044 , \11048 );
and \U$11009 ( \11198 , \11048 , \11053 );
and \U$11010 ( \11199 , \11044 , \11053 );
or \U$11011 ( \11200 , \11197 , \11198 , \11199 );
xor \U$11012 ( \11201 , \11196 , \11200 );
and \U$11013 ( \11202 , \11030 , \11034 );
and \U$11014 ( \11203 , \11034 , \11039 );
and \U$11015 ( \11204 , \11030 , \11039 );
or \U$11016 ( \11205 , \11202 , \11203 , \11204 );
xor \U$11017 ( \11206 , \11201 , \11205 );
xor \U$11018 ( \11207 , \11192 , \11206 );
and \U$11019 ( \11208 , \11040 , \11054 );
and \U$11020 ( \11209 , \11054 , \11066 );
and \U$11021 ( \11210 , \11040 , \11066 );
or \U$11022 ( \11211 , \11208 , \11209 , \11210 );
and \U$11023 ( \11212 , \5737 , \7175 );
not \U$11024 ( \11213 , \11212 );
xnor \U$11025 ( \11214 , \11213 , \7181 );
xor \U$11026 ( \11215 , \6023 , \11214 );
and \U$11027 ( \11216 , \5758 , \7192 );
and \U$11028 ( \11217 , \5770 , \7190 );
nor \U$11029 ( \11218 , \11216 , \11217 );
xnor \U$11030 ( \11219 , \11218 , \7198 );
xor \U$11031 ( \11220 , \11215 , \11219 );
xor \U$11032 ( \11221 , \11211 , \11220 );
and \U$11033 ( \11222 , \5906 , \5852 );
and \U$11034 ( \11223 , \5918 , \5850 );
nor \U$11035 ( \11224 , \11222 , \11223 );
xnor \U$11036 ( \11225 , \11224 , \5859 );
and \U$11037 ( \11226 , \5925 , \5871 );
and \U$11038 ( \11227 , \5937 , \5869 );
nor \U$11039 ( \11228 , \11226 , \11227 );
xnor \U$11040 ( \11229 , \11228 , \5878 );
xor \U$11041 ( \11230 , \11225 , \11229 );
and \U$11042 ( \11231 , \5945 , \5891 );
and \U$11043 ( \11232 , \5957 , \5889 );
nor \U$11044 ( \11233 , \11231 , \11232 );
xnor \U$11045 ( \11234 , \11233 , \5898 );
xor \U$11046 ( \11235 , \11230 , \11234 );
and \U$11047 ( \11236 , \5842 , \5790 );
and \U$11048 ( \11237 , \5854 , \5788 );
nor \U$11049 ( \11238 , \11236 , \11237 );
xnor \U$11050 ( \11239 , \11238 , \5797 );
and \U$11051 ( \11240 , \5861 , \5809 );
and \U$11052 ( \11241 , \5873 , \5807 );
nor \U$11053 ( \11242 , \11240 , \11241 );
xnor \U$11054 ( \11243 , \11242 , \5816 );
xor \U$11055 ( \11244 , \11239 , \11243 );
and \U$11056 ( \11245 , \5881 , \5829 );
and \U$11057 ( \11246 , \5893 , \5827 );
nor \U$11058 ( \11247 , \11245 , \11246 );
xnor \U$11059 ( \11248 , \11247 , \5836 );
xor \U$11060 ( \11249 , \11244 , \11248 );
xor \U$11061 ( \11250 , \11235 , \11249 );
and \U$11062 ( \11251 , \5780 , \7203 );
and \U$11063 ( \11252 , \5792 , \7201 );
nor \U$11064 ( \11253 , \11251 , \11252 );
xnor \U$11065 ( \11254 , \11253 , \6824 );
and \U$11066 ( \11255 , \5799 , \5750 );
and \U$11067 ( \11256 , \5811 , \5748 );
nor \U$11068 ( \11257 , \11255 , \11256 );
xnor \U$11069 ( \11258 , \11257 , \5755 );
xor \U$11070 ( \11259 , \11254 , \11258 );
and \U$11071 ( \11260 , \5819 , \5768 );
and \U$11072 ( \11261 , \5831 , \5766 );
nor \U$11073 ( \11262 , \11260 , \11261 );
xnor \U$11074 ( \11263 , \11262 , \5775 );
xor \U$11075 ( \11264 , \11259 , \11263 );
xor \U$11076 ( \11265 , \11250 , \11264 );
xor \U$11077 ( \11266 , \11221 , \11265 );
xor \U$11078 ( \11267 , \11207 , \11266 );
and \U$11079 ( \11268 , \11011 , \11015 );
and \U$11080 ( \11269 , \11015 , \11020 );
and \U$11081 ( \11270 , \11011 , \11020 );
or \U$11082 ( \11271 , \11268 , \11269 , \11270 );
and \U$11083 ( \11272 , \10997 , \11001 );
and \U$11084 ( \11273 , \11001 , \11006 );
and \U$11085 ( \11274 , \10997 , \11006 );
or \U$11086 ( \11275 , \11272 , \11273 , \11274 );
xor \U$11087 ( \11276 , \11271 , \11275 );
and \U$11088 ( \11277 , \11077 , \11091 );
and \U$11089 ( \11278 , \11091 , \11106 );
and \U$11090 ( \11279 , \11077 , \11106 );
or \U$11091 ( \11280 , \11277 , \11278 , \11279 );
xor \U$11092 ( \11281 , \11276 , \11280 );
xor \U$11093 ( \11282 , \11267 , \11281 );
xor \U$11094 ( \11283 , \11153 , \11282 );
xor \U$11095 ( \11284 , \11144 , \11283 );
and \U$11096 ( \11285 , \10969 , \10983 );
and \U$11097 ( \11286 , \10983 , \11122 );
and \U$11098 ( \11287 , \10969 , \11122 );
or \U$11099 ( \11288 , \11285 , \11286 , \11287 );
nor \U$11100 ( \11289 , \11284 , \11288 );
nor \U$11101 ( \11290 , \11128 , \11289 );
and \U$11102 ( \11291 , \11148 , \11152 );
and \U$11103 ( \11292 , \11152 , \11282 );
and \U$11104 ( \11293 , \11148 , \11282 );
or \U$11105 ( \11294 , \11291 , \11292 , \11293 );
and \U$11106 ( \11295 , \11271 , \11275 );
and \U$11107 ( \11296 , \11275 , \11280 );
and \U$11108 ( \11297 , \11271 , \11280 );
or \U$11109 ( \11298 , \11295 , \11296 , \11297 );
and \U$11110 ( \11299 , \11211 , \11220 );
and \U$11111 ( \11300 , \11220 , \11265 );
and \U$11112 ( \11301 , \11211 , \11265 );
or \U$11113 ( \11302 , \11299 , \11300 , \11301 );
xor \U$11114 ( \11303 , \11298 , \11302 );
and \U$11115 ( \11304 , \11180 , \11191 );
and \U$11116 ( \11305 , \11191 , \11206 );
and \U$11117 ( \11306 , \11180 , \11206 );
or \U$11118 ( \11307 , \11304 , \11305 , \11306 );
xor \U$11119 ( \11308 , \11303 , \11307 );
xor \U$11120 ( \11309 , \11294 , \11308 );
and \U$11121 ( \11310 , \11136 , \11140 );
and \U$11122 ( \11311 , \11140 , \11142 );
and \U$11123 ( \11312 , \11136 , \11142 );
or \U$11124 ( \11313 , \11310 , \11311 , \11312 );
and \U$11125 ( \11314 , \11207 , \11266 );
and \U$11126 ( \11315 , \11266 , \11281 );
and \U$11127 ( \11316 , \11207 , \11281 );
or \U$11128 ( \11317 , \11314 , \11315 , \11316 );
xor \U$11129 ( \11318 , \11313 , \11317 );
and \U$11130 ( \11319 , \11225 , \11229 );
and \U$11131 ( \11320 , \11229 , \11234 );
and \U$11132 ( \11321 , \11225 , \11234 );
or \U$11133 ( \11322 , \11319 , \11320 , \11321 );
and \U$11134 ( \11323 , \11169 , \11173 );
and \U$11135 ( \11324 , \11173 , \11178 );
and \U$11136 ( \11325 , \11169 , \11178 );
or \U$11137 ( \11326 , \11323 , \11324 , \11325 );
xor \U$11138 ( \11327 , \11322 , \11326 );
and \U$11139 ( \11328 , \11157 , \11161 );
and \U$11140 ( \11329 , \11161 , \11164 );
and \U$11141 ( \11330 , \11157 , \11164 );
or \U$11142 ( \11331 , \11328 , \11329 , \11330 );
xor \U$11143 ( \11332 , \11327 , \11331 );
and \U$11144 ( \11333 , \6023 , \11214 );
and \U$11145 ( \11334 , \11214 , \11219 );
and \U$11146 ( \11335 , \6023 , \11219 );
or \U$11147 ( \11336 , \11333 , \11334 , \11335 );
and \U$11148 ( \11337 , \11254 , \11258 );
and \U$11149 ( \11338 , \11258 , \11263 );
and \U$11150 ( \11339 , \11254 , \11263 );
or \U$11151 ( \11340 , \11337 , \11338 , \11339 );
xor \U$11152 ( \11341 , \11336 , \11340 );
and \U$11153 ( \11342 , \11239 , \11243 );
and \U$11154 ( \11343 , \11243 , \11248 );
and \U$11155 ( \11344 , \11239 , \11248 );
or \U$11156 ( \11345 , \11342 , \11343 , \11344 );
xor \U$11157 ( \11346 , \11341 , \11345 );
xor \U$11158 ( \11347 , \11332 , \11346 );
and \U$11159 ( \11348 , \11235 , \11249 );
and \U$11160 ( \11349 , \11249 , \11264 );
and \U$11161 ( \11350 , \11235 , \11264 );
or \U$11162 ( \11351 , \11348 , \11349 , \11350 );
and \U$11163 ( \11352 , \5873 , \5809 );
and \U$11164 ( \11353 , \5842 , \5807 );
nor \U$11165 ( \11354 , \11352 , \11353 );
xnor \U$11166 ( \11355 , \11354 , \5816 );
and \U$11167 ( \11356 , \5893 , \5829 );
and \U$11168 ( \11357 , \5861 , \5827 );
nor \U$11169 ( \11358 , \11356 , \11357 );
xnor \U$11170 ( \11359 , \11358 , \5836 );
xor \U$11171 ( \11360 , \11355 , \11359 );
and \U$11172 ( \11361 , \5918 , \5852 );
and \U$11173 ( \11362 , \5881 , \5850 );
nor \U$11174 ( \11363 , \11361 , \11362 );
xnor \U$11175 ( \11364 , \11363 , \5859 );
xor \U$11176 ( \11365 , \11360 , \11364 );
and \U$11177 ( \11366 , \5811 , \5750 );
and \U$11178 ( \11367 , \5780 , \5748 );
nor \U$11179 ( \11368 , \11366 , \11367 );
xnor \U$11180 ( \11369 , \11368 , \5755 );
and \U$11181 ( \11370 , \5831 , \5768 );
and \U$11182 ( \11371 , \5799 , \5766 );
nor \U$11183 ( \11372 , \11370 , \11371 );
xnor \U$11184 ( \11373 , \11372 , \5775 );
xor \U$11185 ( \11374 , \11369 , \11373 );
and \U$11186 ( \11375 , \5854 , \5790 );
and \U$11187 ( \11376 , \5819 , \5788 );
nor \U$11188 ( \11377 , \11375 , \11376 );
xnor \U$11189 ( \11378 , \11377 , \5797 );
xor \U$11190 ( \11379 , \11374 , \11378 );
xor \U$11191 ( \11380 , \11365 , \11379 );
not \U$11192 ( \11381 , \7181 );
and \U$11193 ( \11382 , \5770 , \7192 );
and \U$11194 ( \11383 , \5737 , \7190 );
nor \U$11195 ( \11384 , \11382 , \11383 );
xnor \U$11196 ( \11385 , \11384 , \7198 );
xor \U$11197 ( \11386 , \11381 , \11385 );
and \U$11198 ( \11387 , \5792 , \7203 );
and \U$11199 ( \11388 , \5758 , \7201 );
nor \U$11200 ( \11389 , \11387 , \11388 );
xnor \U$11201 ( \11390 , \11389 , \6824 );
xor \U$11202 ( \11391 , \11386 , \11390 );
xor \U$11203 ( \11392 , \11380 , \11391 );
xor \U$11204 ( \11393 , \11351 , \11392 );
and \U$11205 ( \11394 , \6057 , \5996 );
and \U$11206 ( \11395 , \6029 , \5994 );
nor \U$11207 ( \11396 , \11394 , \11395 );
xnor \U$11208 ( \11397 , \11396 , \6003 );
and \U$11209 ( \11398 , \6065 , \6016 );
and \U$11210 ( \11399 , \6048 , \6014 );
nor \U$11211 ( \11400 , \11398 , \11399 );
xnor \U$11212 ( \11401 , \11400 , \6023 );
xor \U$11213 ( \11402 , \11397 , \11401 );
and \U$11214 ( \11403 , \5998 , \5935 );
and \U$11215 ( \11404 , \5967 , \5933 );
nor \U$11216 ( \11405 , \11403 , \11404 );
xnor \U$11217 ( \11406 , \11405 , \5942 );
and \U$11218 ( \11407 , \6018 , \5955 );
and \U$11219 ( \11408 , \5986 , \5953 );
nor \U$11220 ( \11409 , \11407 , \11408 );
xnor \U$11221 ( \11410 , \11409 , \5962 );
xor \U$11222 ( \11411 , \11406 , \11410 );
and \U$11223 ( \11412 , \6041 , \5977 );
and \U$11224 ( \11413 , \6006 , \5975 );
nor \U$11225 ( \11414 , \11412 , \11413 );
xnor \U$11226 ( \11415 , \11414 , \5984 );
xor \U$11227 ( \11416 , \11411 , \11415 );
xor \U$11228 ( \11417 , \11402 , \11416 );
and \U$11229 ( \11418 , \5937 , \5871 );
and \U$11230 ( \11419 , \5906 , \5869 );
nor \U$11231 ( \11420 , \11418 , \11419 );
xnor \U$11232 ( \11421 , \11420 , \5878 );
and \U$11233 ( \11422 , \5957 , \5891 );
and \U$11234 ( \11423 , \5925 , \5889 );
nor \U$11235 ( \11424 , \11422 , \11423 );
xnor \U$11236 ( \11425 , \11424 , \5898 );
xor \U$11237 ( \11426 , \11421 , \11425 );
and \U$11238 ( \11427 , \5979 , \5916 );
and \U$11239 ( \11428 , \5945 , \5914 );
nor \U$11240 ( \11429 , \11427 , \11428 );
xnor \U$11241 ( \11430 , \11429 , \5923 );
xor \U$11242 ( \11431 , \11426 , \11430 );
xor \U$11243 ( \11432 , \11417 , \11431 );
xor \U$11244 ( \11433 , \11393 , \11432 );
xor \U$11245 ( \11434 , \11347 , \11433 );
and \U$11246 ( \11435 , \11196 , \11200 );
and \U$11247 ( \11436 , \11200 , \11205 );
and \U$11248 ( \11437 , \11196 , \11205 );
or \U$11249 ( \11438 , \11435 , \11436 , \11437 );
and \U$11250 ( \11439 , \11184 , \11188 );
and \U$11251 ( \11440 , \11188 , \11190 );
and \U$11252 ( \11441 , \11184 , \11190 );
or \U$11253 ( \11442 , \11439 , \11440 , \11441 );
xor \U$11254 ( \11443 , \11438 , \11442 );
or \U$11255 ( \11444 , \11165 , \11179 );
xor \U$11256 ( \11445 , \11443 , \11444 );
xor \U$11257 ( \11446 , \11434 , \11445 );
xor \U$11258 ( \11447 , \11318 , \11446 );
xor \U$11259 ( \11448 , \11309 , \11447 );
and \U$11260 ( \11449 , \11132 , \11143 );
and \U$11261 ( \11450 , \11143 , \11283 );
and \U$11262 ( \11451 , \11132 , \11283 );
or \U$11263 ( \11452 , \11449 , \11450 , \11451 );
nor \U$11264 ( \11453 , \11448 , \11452 );
and \U$11265 ( \11454 , \11313 , \11317 );
and \U$11266 ( \11455 , \11317 , \11446 );
and \U$11267 ( \11456 , \11313 , \11446 );
or \U$11268 ( \11457 , \11454 , \11455 , \11456 );
and \U$11269 ( \11458 , \11438 , \11442 );
and \U$11270 ( \11459 , \11442 , \11444 );
and \U$11271 ( \11460 , \11438 , \11444 );
or \U$11272 ( \11461 , \11458 , \11459 , \11460 );
and \U$11273 ( \11462 , \11351 , \11392 );
and \U$11274 ( \11463 , \11392 , \11432 );
and \U$11275 ( \11464 , \11351 , \11432 );
or \U$11276 ( \11465 , \11462 , \11463 , \11464 );
xor \U$11277 ( \11466 , \11461 , \11465 );
and \U$11278 ( \11467 , \11332 , \11346 );
xor \U$11279 ( \11468 , \11466 , \11467 );
xor \U$11280 ( \11469 , \11457 , \11468 );
and \U$11281 ( \11470 , \11298 , \11302 );
and \U$11282 ( \11471 , \11302 , \11307 );
and \U$11283 ( \11472 , \11298 , \11307 );
or \U$11284 ( \11473 , \11470 , \11471 , \11472 );
and \U$11285 ( \11474 , \11347 , \11433 );
and \U$11286 ( \11475 , \11433 , \11445 );
and \U$11287 ( \11476 , \11347 , \11445 );
or \U$11288 ( \11477 , \11474 , \11475 , \11476 );
xor \U$11289 ( \11478 , \11473 , \11477 );
and \U$11290 ( \11479 , \6029 , \5996 );
and \U$11291 ( \11480 , \6041 , \5994 );
nor \U$11292 ( \11481 , \11479 , \11480 );
xnor \U$11293 ( \11482 , \11481 , \6003 );
and \U$11294 ( \11483 , \6048 , \6016 );
and \U$11295 ( \11484 , \6057 , \6014 );
nor \U$11296 ( \11485 , \11483 , \11484 );
xnor \U$11297 ( \11486 , \11485 , \6023 );
xor \U$11298 ( \11487 , \11482 , \11486 );
nand \U$11299 ( \11488 , \6065 , \6037 );
xnor \U$11300 ( \11489 , \11488 , \6046 );
xor \U$11301 ( \11490 , \11487 , \11489 );
and \U$11302 ( \11491 , \5967 , \5935 );
and \U$11303 ( \11492 , \5979 , \5933 );
nor \U$11304 ( \11493 , \11491 , \11492 );
xnor \U$11305 ( \11494 , \11493 , \5942 );
and \U$11306 ( \11495 , \5986 , \5955 );
and \U$11307 ( \11496 , \5998 , \5953 );
nor \U$11308 ( \11497 , \11495 , \11496 );
xnor \U$11309 ( \11498 , \11497 , \5962 );
xor \U$11310 ( \11499 , \11494 , \11498 );
and \U$11311 ( \11500 , \6006 , \5977 );
and \U$11312 ( \11501 , \6018 , \5975 );
nor \U$11313 ( \11502 , \11500 , \11501 );
xnor \U$11314 ( \11503 , \11502 , \5984 );
xor \U$11315 ( \11504 , \11499 , \11503 );
xnor \U$11316 ( \11505 , \11490 , \11504 );
and \U$11317 ( \11506 , \11421 , \11425 );
and \U$11318 ( \11507 , \11425 , \11430 );
and \U$11319 ( \11508 , \11421 , \11430 );
or \U$11320 ( \11509 , \11506 , \11507 , \11508 );
and \U$11321 ( \11510 , \11406 , \11410 );
and \U$11322 ( \11511 , \11410 , \11415 );
and \U$11323 ( \11512 , \11406 , \11415 );
or \U$11324 ( \11513 , \11510 , \11511 , \11512 );
xor \U$11325 ( \11514 , \11509 , \11513 );
and \U$11326 ( \11515 , \11397 , \11401 );
xor \U$11327 ( \11516 , \11514 , \11515 );
xor \U$11328 ( \11517 , \11505 , \11516 );
and \U$11329 ( \11518 , \11381 , \11385 );
and \U$11330 ( \11519 , \11385 , \11390 );
and \U$11331 ( \11520 , \11381 , \11390 );
or \U$11332 ( \11521 , \11518 , \11519 , \11520 );
and \U$11333 ( \11522 , \11369 , \11373 );
and \U$11334 ( \11523 , \11373 , \11378 );
and \U$11335 ( \11524 , \11369 , \11378 );
or \U$11336 ( \11525 , \11522 , \11523 , \11524 );
xor \U$11337 ( \11526 , \11521 , \11525 );
and \U$11338 ( \11527 , \11355 , \11359 );
and \U$11339 ( \11528 , \11359 , \11364 );
and \U$11340 ( \11529 , \11355 , \11364 );
or \U$11341 ( \11530 , \11527 , \11528 , \11529 );
xor \U$11342 ( \11531 , \11526 , \11530 );
xor \U$11343 ( \11532 , \11517 , \11531 );
and \U$11344 ( \11533 , \11365 , \11379 );
and \U$11345 ( \11534 , \11379 , \11391 );
and \U$11346 ( \11535 , \11365 , \11391 );
or \U$11347 ( \11536 , \11533 , \11534 , \11535 );
and \U$11348 ( \11537 , \5737 , \7192 );
not \U$11349 ( \11538 , \11537 );
xnor \U$11350 ( \11539 , \11538 , \7198 );
xor \U$11351 ( \11540 , \6046 , \11539 );
and \U$11352 ( \11541 , \5758 , \7203 );
and \U$11353 ( \11542 , \5770 , \7201 );
nor \U$11354 ( \11543 , \11541 , \11542 );
xnor \U$11355 ( \11544 , \11543 , \6824 );
xor \U$11356 ( \11545 , \11540 , \11544 );
xor \U$11357 ( \11546 , \11536 , \11545 );
and \U$11358 ( \11547 , \5906 , \5871 );
and \U$11359 ( \11548 , \5918 , \5869 );
nor \U$11360 ( \11549 , \11547 , \11548 );
xnor \U$11361 ( \11550 , \11549 , \5878 );
and \U$11362 ( \11551 , \5925 , \5891 );
and \U$11363 ( \11552 , \5937 , \5889 );
nor \U$11364 ( \11553 , \11551 , \11552 );
xnor \U$11365 ( \11554 , \11553 , \5898 );
xor \U$11366 ( \11555 , \11550 , \11554 );
and \U$11367 ( \11556 , \5945 , \5916 );
and \U$11368 ( \11557 , \5957 , \5914 );
nor \U$11369 ( \11558 , \11556 , \11557 );
xnor \U$11370 ( \11559 , \11558 , \5923 );
xor \U$11371 ( \11560 , \11555 , \11559 );
and \U$11372 ( \11561 , \5842 , \5809 );
and \U$11373 ( \11562 , \5854 , \5807 );
nor \U$11374 ( \11563 , \11561 , \11562 );
xnor \U$11375 ( \11564 , \11563 , \5816 );
and \U$11376 ( \11565 , \5861 , \5829 );
and \U$11377 ( \11566 , \5873 , \5827 );
nor \U$11378 ( \11567 , \11565 , \11566 );
xnor \U$11379 ( \11568 , \11567 , \5836 );
xor \U$11380 ( \11569 , \11564 , \11568 );
and \U$11381 ( \11570 , \5881 , \5852 );
and \U$11382 ( \11571 , \5893 , \5850 );
nor \U$11383 ( \11572 , \11570 , \11571 );
xnor \U$11384 ( \11573 , \11572 , \5859 );
xor \U$11385 ( \11574 , \11569 , \11573 );
xor \U$11386 ( \11575 , \11560 , \11574 );
and \U$11387 ( \11576 , \5780 , \5750 );
and \U$11388 ( \11577 , \5792 , \5748 );
nor \U$11389 ( \11578 , \11576 , \11577 );
xnor \U$11390 ( \11579 , \11578 , \5755 );
and \U$11391 ( \11580 , \5799 , \5768 );
and \U$11392 ( \11581 , \5811 , \5766 );
nor \U$11393 ( \11582 , \11580 , \11581 );
xnor \U$11394 ( \11583 , \11582 , \5775 );
xor \U$11395 ( \11584 , \11579 , \11583 );
and \U$11396 ( \11585 , \5819 , \5790 );
and \U$11397 ( \11586 , \5831 , \5788 );
nor \U$11398 ( \11587 , \11585 , \11586 );
xnor \U$11399 ( \11588 , \11587 , \5797 );
xor \U$11400 ( \11589 , \11584 , \11588 );
xor \U$11401 ( \11590 , \11575 , \11589 );
xor \U$11402 ( \11591 , \11546 , \11590 );
xor \U$11403 ( \11592 , \11532 , \11591 );
and \U$11404 ( \11593 , \11336 , \11340 );
and \U$11405 ( \11594 , \11340 , \11345 );
and \U$11406 ( \11595 , \11336 , \11345 );
or \U$11407 ( \11596 , \11593 , \11594 , \11595 );
and \U$11408 ( \11597 , \11322 , \11326 );
and \U$11409 ( \11598 , \11326 , \11331 );
and \U$11410 ( \11599 , \11322 , \11331 );
or \U$11411 ( \11600 , \11597 , \11598 , \11599 );
xor \U$11412 ( \11601 , \11596 , \11600 );
and \U$11413 ( \11602 , \11402 , \11416 );
and \U$11414 ( \11603 , \11416 , \11431 );
and \U$11415 ( \11604 , \11402 , \11431 );
or \U$11416 ( \11605 , \11602 , \11603 , \11604 );
xor \U$11417 ( \11606 , \11601 , \11605 );
xor \U$11418 ( \11607 , \11592 , \11606 );
xor \U$11419 ( \11608 , \11478 , \11607 );
xor \U$11420 ( \11609 , \11469 , \11608 );
and \U$11421 ( \11610 , \11294 , \11308 );
and \U$11422 ( \11611 , \11308 , \11447 );
and \U$11423 ( \11612 , \11294 , \11447 );
or \U$11424 ( \11613 , \11610 , \11611 , \11612 );
nor \U$11425 ( \11614 , \11609 , \11613 );
nor \U$11426 ( \11615 , \11453 , \11614 );
nand \U$11427 ( \11616 , \11290 , \11615 );
nor \U$11428 ( \11617 , \10965 , \11616 );
and \U$11429 ( \11618 , \11473 , \11477 );
and \U$11430 ( \11619 , \11477 , \11607 );
and \U$11431 ( \11620 , \11473 , \11607 );
or \U$11432 ( \11621 , \11618 , \11619 , \11620 );
and \U$11433 ( \11622 , \11596 , \11600 );
and \U$11434 ( \11623 , \11600 , \11605 );
and \U$11435 ( \11624 , \11596 , \11605 );
or \U$11436 ( \11625 , \11622 , \11623 , \11624 );
and \U$11437 ( \11626 , \11536 , \11545 );
and \U$11438 ( \11627 , \11545 , \11590 );
and \U$11439 ( \11628 , \11536 , \11590 );
or \U$11440 ( \11629 , \11626 , \11627 , \11628 );
xor \U$11441 ( \11630 , \11625 , \11629 );
and \U$11442 ( \11631 , \11505 , \11516 );
and \U$11443 ( \11632 , \11516 , \11531 );
and \U$11444 ( \11633 , \11505 , \11531 );
or \U$11445 ( \11634 , \11631 , \11632 , \11633 );
xor \U$11446 ( \11635 , \11630 , \11634 );
xor \U$11447 ( \11636 , \11621 , \11635 );
and \U$11448 ( \11637 , \11461 , \11465 );
and \U$11449 ( \11638 , \11465 , \11467 );
and \U$11450 ( \11639 , \11461 , \11467 );
or \U$11451 ( \11640 , \11637 , \11638 , \11639 );
and \U$11452 ( \11641 , \11532 , \11591 );
and \U$11453 ( \11642 , \11591 , \11606 );
and \U$11454 ( \11643 , \11532 , \11606 );
or \U$11455 ( \11644 , \11641 , \11642 , \11643 );
xor \U$11456 ( \11645 , \11640 , \11644 );
and \U$11457 ( \11646 , \11550 , \11554 );
and \U$11458 ( \11647 , \11554 , \11559 );
and \U$11459 ( \11648 , \11550 , \11559 );
or \U$11460 ( \11649 , \11646 , \11647 , \11648 );
and \U$11461 ( \11650 , \11494 , \11498 );
and \U$11462 ( \11651 , \11498 , \11503 );
and \U$11463 ( \11652 , \11494 , \11503 );
or \U$11464 ( \11653 , \11650 , \11651 , \11652 );
xor \U$11465 ( \11654 , \11649 , \11653 );
and \U$11466 ( \11655 , \11482 , \11486 );
and \U$11467 ( \11656 , \11486 , \11489 );
and \U$11468 ( \11657 , \11482 , \11489 );
or \U$11469 ( \11658 , \11655 , \11656 , \11657 );
xor \U$11470 ( \11659 , \11654 , \11658 );
and \U$11471 ( \11660 , \6046 , \11539 );
and \U$11472 ( \11661 , \11539 , \11544 );
and \U$11473 ( \11662 , \6046 , \11544 );
or \U$11474 ( \11663 , \11660 , \11661 , \11662 );
and \U$11475 ( \11664 , \11579 , \11583 );
and \U$11476 ( \11665 , \11583 , \11588 );
and \U$11477 ( \11666 , \11579 , \11588 );
or \U$11478 ( \11667 , \11664 , \11665 , \11666 );
xor \U$11479 ( \11668 , \11663 , \11667 );
and \U$11480 ( \11669 , \11564 , \11568 );
and \U$11481 ( \11670 , \11568 , \11573 );
and \U$11482 ( \11671 , \11564 , \11573 );
or \U$11483 ( \11672 , \11669 , \11670 , \11671 );
xor \U$11484 ( \11673 , \11668 , \11672 );
xor \U$11485 ( \11674 , \11659 , \11673 );
and \U$11486 ( \11675 , \11560 , \11574 );
and \U$11487 ( \11676 , \11574 , \11589 );
and \U$11488 ( \11677 , \11560 , \11589 );
or \U$11489 ( \11678 , \11675 , \11676 , \11677 );
and \U$11490 ( \11679 , \5873 , \5829 );
and \U$11491 ( \11680 , \5842 , \5827 );
nor \U$11492 ( \11681 , \11679 , \11680 );
xnor \U$11493 ( \11682 , \11681 , \5836 );
and \U$11494 ( \11683 , \5893 , \5852 );
and \U$11495 ( \11684 , \5861 , \5850 );
nor \U$11496 ( \11685 , \11683 , \11684 );
xnor \U$11497 ( \11686 , \11685 , \5859 );
xor \U$11498 ( \11687 , \11682 , \11686 );
and \U$11499 ( \11688 , \5918 , \5871 );
and \U$11500 ( \11689 , \5881 , \5869 );
nor \U$11501 ( \11690 , \11688 , \11689 );
xnor \U$11502 ( \11691 , \11690 , \5878 );
xor \U$11503 ( \11692 , \11687 , \11691 );
and \U$11504 ( \11693 , \5811 , \5768 );
and \U$11505 ( \11694 , \5780 , \5766 );
nor \U$11506 ( \11695 , \11693 , \11694 );
xnor \U$11507 ( \11696 , \11695 , \5775 );
and \U$11508 ( \11697 , \5831 , \5790 );
and \U$11509 ( \11698 , \5799 , \5788 );
nor \U$11510 ( \11699 , \11697 , \11698 );
xnor \U$11511 ( \11700 , \11699 , \5797 );
xor \U$11512 ( \11701 , \11696 , \11700 );
and \U$11513 ( \11702 , \5854 , \5809 );
and \U$11514 ( \11703 , \5819 , \5807 );
nor \U$11515 ( \11704 , \11702 , \11703 );
xnor \U$11516 ( \11705 , \11704 , \5816 );
xor \U$11517 ( \11706 , \11701 , \11705 );
xor \U$11518 ( \11707 , \11692 , \11706 );
not \U$11519 ( \11708 , \7198 );
and \U$11520 ( \11709 , \5770 , \7203 );
and \U$11521 ( \11710 , \5737 , \7201 );
nor \U$11522 ( \11711 , \11709 , \11710 );
xnor \U$11523 ( \11712 , \11711 , \6824 );
xor \U$11524 ( \11713 , \11708 , \11712 );
and \U$11525 ( \11714 , \5792 , \5750 );
and \U$11526 ( \11715 , \5758 , \5748 );
nor \U$11527 ( \11716 , \11714 , \11715 );
xnor \U$11528 ( \11717 , \11716 , \5755 );
xor \U$11529 ( \11718 , \11713 , \11717 );
xor \U$11530 ( \11719 , \11707 , \11718 );
xor \U$11531 ( \11720 , \11678 , \11719 );
and \U$11532 ( \11721 , \6057 , \6016 );
and \U$11533 ( \11722 , \6029 , \6014 );
nor \U$11534 ( \11723 , \11721 , \11722 );
xnor \U$11535 ( \11724 , \11723 , \6023 );
and \U$11536 ( \11725 , \6065 , \6039 );
and \U$11537 ( \11726 , \6048 , \6037 );
nor \U$11538 ( \11727 , \11725 , \11726 );
xnor \U$11539 ( \11728 , \11727 , \6046 );
xor \U$11540 ( \11729 , \11724 , \11728 );
and \U$11541 ( \11730 , \5998 , \5955 );
and \U$11542 ( \11731 , \5967 , \5953 );
nor \U$11543 ( \11732 , \11730 , \11731 );
xnor \U$11544 ( \11733 , \11732 , \5962 );
and \U$11545 ( \11734 , \6018 , \5977 );
and \U$11546 ( \11735 , \5986 , \5975 );
nor \U$11547 ( \11736 , \11734 , \11735 );
xnor \U$11548 ( \11737 , \11736 , \5984 );
xor \U$11549 ( \11738 , \11733 , \11737 );
and \U$11550 ( \11739 , \6041 , \5996 );
and \U$11551 ( \11740 , \6006 , \5994 );
nor \U$11552 ( \11741 , \11739 , \11740 );
xnor \U$11553 ( \11742 , \11741 , \6003 );
xor \U$11554 ( \11743 , \11738 , \11742 );
xor \U$11555 ( \11744 , \11729 , \11743 );
and \U$11556 ( \11745 , \5937 , \5891 );
and \U$11557 ( \11746 , \5906 , \5889 );
nor \U$11558 ( \11747 , \11745 , \11746 );
xnor \U$11559 ( \11748 , \11747 , \5898 );
and \U$11560 ( \11749 , \5957 , \5916 );
and \U$11561 ( \11750 , \5925 , \5914 );
nor \U$11562 ( \11751 , \11749 , \11750 );
xnor \U$11563 ( \11752 , \11751 , \5923 );
xor \U$11564 ( \11753 , \11748 , \11752 );
and \U$11565 ( \11754 , \5979 , \5935 );
and \U$11566 ( \11755 , \5945 , \5933 );
nor \U$11567 ( \11756 , \11754 , \11755 );
xnor \U$11568 ( \11757 , \11756 , \5942 );
xor \U$11569 ( \11758 , \11753 , \11757 );
xor \U$11570 ( \11759 , \11744 , \11758 );
xor \U$11571 ( \11760 , \11720 , \11759 );
xor \U$11572 ( \11761 , \11674 , \11760 );
and \U$11573 ( \11762 , \11521 , \11525 );
and \U$11574 ( \11763 , \11525 , \11530 );
and \U$11575 ( \11764 , \11521 , \11530 );
or \U$11576 ( \11765 , \11762 , \11763 , \11764 );
and \U$11577 ( \11766 , \11509 , \11513 );
and \U$11578 ( \11767 , \11513 , \11515 );
and \U$11579 ( \11768 , \11509 , \11515 );
or \U$11580 ( \11769 , \11766 , \11767 , \11768 );
xor \U$11581 ( \11770 , \11765 , \11769 );
or \U$11582 ( \11771 , \11490 , \11504 );
xor \U$11583 ( \11772 , \11770 , \11771 );
xor \U$11584 ( \11773 , \11761 , \11772 );
xor \U$11585 ( \11774 , \11645 , \11773 );
xor \U$11586 ( \11775 , \11636 , \11774 );
and \U$11587 ( \11776 , \11457 , \11468 );
and \U$11588 ( \11777 , \11468 , \11608 );
and \U$11589 ( \11778 , \11457 , \11608 );
or \U$11590 ( \11779 , \11776 , \11777 , \11778 );
nor \U$11591 ( \11780 , \11775 , \11779 );
and \U$11592 ( \11781 , \11640 , \11644 );
and \U$11593 ( \11782 , \11644 , \11773 );
and \U$11594 ( \11783 , \11640 , \11773 );
or \U$11595 ( \11784 , \11781 , \11782 , \11783 );
and \U$11596 ( \11785 , \11765 , \11769 );
and \U$11597 ( \11786 , \11769 , \11771 );
and \U$11598 ( \11787 , \11765 , \11771 );
or \U$11599 ( \11788 , \11785 , \11786 , \11787 );
and \U$11600 ( \11789 , \11678 , \11719 );
and \U$11601 ( \11790 , \11719 , \11759 );
and \U$11602 ( \11791 , \11678 , \11759 );
or \U$11603 ( \11792 , \11789 , \11790 , \11791 );
xor \U$11604 ( \11793 , \11788 , \11792 );
and \U$11605 ( \11794 , \11659 , \11673 );
xor \U$11606 ( \11795 , \11793 , \11794 );
xor \U$11607 ( \11796 , \11784 , \11795 );
and \U$11608 ( \11797 , \11625 , \11629 );
and \U$11609 ( \11798 , \11629 , \11634 );
and \U$11610 ( \11799 , \11625 , \11634 );
or \U$11611 ( \11800 , \11797 , \11798 , \11799 );
and \U$11612 ( \11801 , \11674 , \11760 );
and \U$11613 ( \11802 , \11760 , \11772 );
and \U$11614 ( \11803 , \11674 , \11772 );
or \U$11615 ( \11804 , \11801 , \11802 , \11803 );
xor \U$11616 ( \11805 , \11800 , \11804 );
and \U$11617 ( \11806 , \6029 , \6016 );
and \U$11618 ( \11807 , \6041 , \6014 );
nor \U$11619 ( \11808 , \11806 , \11807 );
xnor \U$11620 ( \11809 , \11808 , \6023 );
and \U$11621 ( \11810 , \6048 , \6039 );
and \U$11622 ( \11811 , \6057 , \6037 );
nor \U$11623 ( \11812 , \11810 , \11811 );
xnor \U$11624 ( \11813 , \11812 , \6046 );
xor \U$11625 ( \11814 , \11809 , \11813 );
nand \U$11626 ( \11815 , \6065 , \6053 );
xnor \U$11627 ( \11816 , \11815 , \6062 );
xor \U$11628 ( \11817 , \11814 , \11816 );
and \U$11629 ( \11818 , \5967 , \5955 );
and \U$11630 ( \11819 , \5979 , \5953 );
nor \U$11631 ( \11820 , \11818 , \11819 );
xnor \U$11632 ( \11821 , \11820 , \5962 );
and \U$11633 ( \11822 , \5986 , \5977 );
and \U$11634 ( \11823 , \5998 , \5975 );
nor \U$11635 ( \11824 , \11822 , \11823 );
xnor \U$11636 ( \11825 , \11824 , \5984 );
xor \U$11637 ( \11826 , \11821 , \11825 );
and \U$11638 ( \11827 , \6006 , \5996 );
and \U$11639 ( \11828 , \6018 , \5994 );
nor \U$11640 ( \11829 , \11827 , \11828 );
xnor \U$11641 ( \11830 , \11829 , \6003 );
xor \U$11642 ( \11831 , \11826 , \11830 );
xnor \U$11643 ( \11832 , \11817 , \11831 );
and \U$11644 ( \11833 , \11748 , \11752 );
and \U$11645 ( \11834 , \11752 , \11757 );
and \U$11646 ( \11835 , \11748 , \11757 );
or \U$11647 ( \11836 , \11833 , \11834 , \11835 );
and \U$11648 ( \11837 , \11733 , \11737 );
and \U$11649 ( \11838 , \11737 , \11742 );
and \U$11650 ( \11839 , \11733 , \11742 );
or \U$11651 ( \11840 , \11837 , \11838 , \11839 );
xor \U$11652 ( \11841 , \11836 , \11840 );
and \U$11653 ( \11842 , \11724 , \11728 );
xor \U$11654 ( \11843 , \11841 , \11842 );
xor \U$11655 ( \11844 , \11832 , \11843 );
and \U$11656 ( \11845 , \11708 , \11712 );
and \U$11657 ( \11846 , \11712 , \11717 );
and \U$11658 ( \11847 , \11708 , \11717 );
or \U$11659 ( \11848 , \11845 , \11846 , \11847 );
and \U$11660 ( \11849 , \11696 , \11700 );
and \U$11661 ( \11850 , \11700 , \11705 );
and \U$11662 ( \11851 , \11696 , \11705 );
or \U$11663 ( \11852 , \11849 , \11850 , \11851 );
xor \U$11664 ( \11853 , \11848 , \11852 );
and \U$11665 ( \11854 , \11682 , \11686 );
and \U$11666 ( \11855 , \11686 , \11691 );
and \U$11667 ( \11856 , \11682 , \11691 );
or \U$11668 ( \11857 , \11854 , \11855 , \11856 );
xor \U$11669 ( \11858 , \11853 , \11857 );
xor \U$11670 ( \11859 , \11844 , \11858 );
and \U$11671 ( \11860 , \11692 , \11706 );
and \U$11672 ( \11861 , \11706 , \11718 );
and \U$11673 ( \11862 , \11692 , \11718 );
or \U$11674 ( \11863 , \11860 , \11861 , \11862 );
and \U$11675 ( \11864 , \5737 , \7203 );
not \U$11676 ( \11865 , \11864 );
xnor \U$11677 ( \11866 , \11865 , \6824 );
xor \U$11678 ( \11867 , \6062 , \11866 );
and \U$11679 ( \11868 , \5758 , \5750 );
and \U$11680 ( \11869 , \5770 , \5748 );
nor \U$11681 ( \11870 , \11868 , \11869 );
xnor \U$11682 ( \11871 , \11870 , \5755 );
xor \U$11683 ( \11872 , \11867 , \11871 );
xor \U$11684 ( \11873 , \11863 , \11872 );
and \U$11685 ( \11874 , \5906 , \5891 );
and \U$11686 ( \11875 , \5918 , \5889 );
nor \U$11687 ( \11876 , \11874 , \11875 );
xnor \U$11688 ( \11877 , \11876 , \5898 );
and \U$11689 ( \11878 , \5925 , \5916 );
and \U$11690 ( \11879 , \5937 , \5914 );
nor \U$11691 ( \11880 , \11878 , \11879 );
xnor \U$11692 ( \11881 , \11880 , \5923 );
xor \U$11693 ( \11882 , \11877 , \11881 );
and \U$11694 ( \11883 , \5945 , \5935 );
and \U$11695 ( \11884 , \5957 , \5933 );
nor \U$11696 ( \11885 , \11883 , \11884 );
xnor \U$11697 ( \11886 , \11885 , \5942 );
xor \U$11698 ( \11887 , \11882 , \11886 );
and \U$11699 ( \11888 , \5842 , \5829 );
and \U$11700 ( \11889 , \5854 , \5827 );
nor \U$11701 ( \11890 , \11888 , \11889 );
xnor \U$11702 ( \11891 , \11890 , \5836 );
and \U$11703 ( \11892 , \5861 , \5852 );
and \U$11704 ( \11893 , \5873 , \5850 );
nor \U$11705 ( \11894 , \11892 , \11893 );
xnor \U$11706 ( \11895 , \11894 , \5859 );
xor \U$11707 ( \11896 , \11891 , \11895 );
and \U$11708 ( \11897 , \5881 , \5871 );
and \U$11709 ( \11898 , \5893 , \5869 );
nor \U$11710 ( \11899 , \11897 , \11898 );
xnor \U$11711 ( \11900 , \11899 , \5878 );
xor \U$11712 ( \11901 , \11896 , \11900 );
xor \U$11713 ( \11902 , \11887 , \11901 );
and \U$11714 ( \11903 , \5780 , \5768 );
and \U$11715 ( \11904 , \5792 , \5766 );
nor \U$11716 ( \11905 , \11903 , \11904 );
xnor \U$11717 ( \11906 , \11905 , \5775 );
and \U$11718 ( \11907 , \5799 , \5790 );
and \U$11719 ( \11908 , \5811 , \5788 );
nor \U$11720 ( \11909 , \11907 , \11908 );
xnor \U$11721 ( \11910 , \11909 , \5797 );
xor \U$11722 ( \11911 , \11906 , \11910 );
and \U$11723 ( \11912 , \5819 , \5809 );
and \U$11724 ( \11913 , \5831 , \5807 );
nor \U$11725 ( \11914 , \11912 , \11913 );
xnor \U$11726 ( \11915 , \11914 , \5816 );
xor \U$11727 ( \11916 , \11911 , \11915 );
xor \U$11728 ( \11917 , \11902 , \11916 );
xor \U$11729 ( \11918 , \11873 , \11917 );
xor \U$11730 ( \11919 , \11859 , \11918 );
and \U$11731 ( \11920 , \11663 , \11667 );
and \U$11732 ( \11921 , \11667 , \11672 );
and \U$11733 ( \11922 , \11663 , \11672 );
or \U$11734 ( \11923 , \11920 , \11921 , \11922 );
and \U$11735 ( \11924 , \11649 , \11653 );
and \U$11736 ( \11925 , \11653 , \11658 );
and \U$11737 ( \11926 , \11649 , \11658 );
or \U$11738 ( \11927 , \11924 , \11925 , \11926 );
xor \U$11739 ( \11928 , \11923 , \11927 );
and \U$11740 ( \11929 , \11729 , \11743 );
and \U$11741 ( \11930 , \11743 , \11758 );
and \U$11742 ( \11931 , \11729 , \11758 );
or \U$11743 ( \11932 , \11929 , \11930 , \11931 );
xor \U$11744 ( \11933 , \11928 , \11932 );
xor \U$11745 ( \11934 , \11919 , \11933 );
xor \U$11746 ( \11935 , \11805 , \11934 );
xor \U$11747 ( \11936 , \11796 , \11935 );
and \U$11748 ( \11937 , \11621 , \11635 );
and \U$11749 ( \11938 , \11635 , \11774 );
and \U$11750 ( \11939 , \11621 , \11774 );
or \U$11751 ( \11940 , \11937 , \11938 , \11939 );
nor \U$11752 ( \11941 , \11936 , \11940 );
nor \U$11753 ( \11942 , \11780 , \11941 );
and \U$11754 ( \11943 , \11800 , \11804 );
and \U$11755 ( \11944 , \11804 , \11934 );
and \U$11756 ( \11945 , \11800 , \11934 );
or \U$11757 ( \11946 , \11943 , \11944 , \11945 );
and \U$11758 ( \11947 , \11923 , \11927 );
and \U$11759 ( \11948 , \11927 , \11932 );
and \U$11760 ( \11949 , \11923 , \11932 );
or \U$11761 ( \11950 , \11947 , \11948 , \11949 );
and \U$11762 ( \11951 , \11863 , \11872 );
and \U$11763 ( \11952 , \11872 , \11917 );
and \U$11764 ( \11953 , \11863 , \11917 );
or \U$11765 ( \11954 , \11951 , \11952 , \11953 );
xor \U$11766 ( \11955 , \11950 , \11954 );
and \U$11767 ( \11956 , \11832 , \11843 );
and \U$11768 ( \11957 , \11843 , \11858 );
and \U$11769 ( \11958 , \11832 , \11858 );
or \U$11770 ( \11959 , \11956 , \11957 , \11958 );
xor \U$11771 ( \11960 , \11955 , \11959 );
xor \U$11772 ( \11961 , \11946 , \11960 );
and \U$11773 ( \11962 , \11788 , \11792 );
and \U$11774 ( \11963 , \11792 , \11794 );
and \U$11775 ( \11964 , \11788 , \11794 );
or \U$11776 ( \11965 , \11962 , \11963 , \11964 );
and \U$11777 ( \11966 , \11859 , \11918 );
and \U$11778 ( \11967 , \11918 , \11933 );
and \U$11779 ( \11968 , \11859 , \11933 );
or \U$11780 ( \11969 , \11966 , \11967 , \11968 );
xor \U$11781 ( \11970 , \11965 , \11969 );
and \U$11782 ( \11971 , \11877 , \11881 );
and \U$11783 ( \11972 , \11881 , \11886 );
and \U$11784 ( \11973 , \11877 , \11886 );
or \U$11785 ( \11974 , \11971 , \11972 , \11973 );
and \U$11786 ( \11975 , \11821 , \11825 );
and \U$11787 ( \11976 , \11825 , \11830 );
and \U$11788 ( \11977 , \11821 , \11830 );
or \U$11789 ( \11978 , \11975 , \11976 , \11977 );
xor \U$11790 ( \11979 , \11974 , \11978 );
and \U$11791 ( \11980 , \11809 , \11813 );
and \U$11792 ( \11981 , \11813 , \11816 );
and \U$11793 ( \11982 , \11809 , \11816 );
or \U$11794 ( \11983 , \11980 , \11981 , \11982 );
xor \U$11795 ( \11984 , \11979 , \11983 );
and \U$11796 ( \11985 , \6062 , \11866 );
and \U$11797 ( \11986 , \11866 , \11871 );
and \U$11798 ( \11987 , \6062 , \11871 );
or \U$11799 ( \11988 , \11985 , \11986 , \11987 );
and \U$11800 ( \11989 , \11906 , \11910 );
and \U$11801 ( \11990 , \11910 , \11915 );
and \U$11802 ( \11991 , \11906 , \11915 );
or \U$11803 ( \11992 , \11989 , \11990 , \11991 );
xor \U$11804 ( \11993 , \11988 , \11992 );
and \U$11805 ( \11994 , \11891 , \11895 );
and \U$11806 ( \11995 , \11895 , \11900 );
and \U$11807 ( \11996 , \11891 , \11900 );
or \U$11808 ( \11997 , \11994 , \11995 , \11996 );
xor \U$11809 ( \11998 , \11993 , \11997 );
xor \U$11810 ( \11999 , \11984 , \11998 );
and \U$11811 ( \12000 , \11887 , \11901 );
and \U$11812 ( \12001 , \11901 , \11916 );
and \U$11813 ( \12002 , \11887 , \11916 );
or \U$11814 ( \12003 , \12000 , \12001 , \12002 );
xor \U$11815 ( \12004 , \6858 , \6862 );
xor \U$11816 ( \12005 , \12004 , \6867 );
xor \U$11817 ( \12006 , \6841 , \6845 );
xor \U$11818 ( \12007 , \12006 , \6850 );
xor \U$11819 ( \12008 , \12005 , \12007 );
xor \U$11820 ( \12009 , \6825 , \6829 );
xor \U$11821 ( \12010 , \12009 , \6834 );
xor \U$11822 ( \12011 , \12008 , \12010 );
xor \U$11823 ( \12012 , \12003 , \12011 );
xor \U$11824 ( \12013 , \6910 , \6914 );
xor \U$11825 ( \12014 , \6893 , \6897 );
xor \U$11826 ( \12015 , \12014 , \6902 );
xor \U$11827 ( \12016 , \12013 , \12015 );
xor \U$11828 ( \12017 , \6877 , \6881 );
xor \U$11829 ( \12018 , \12017 , \6886 );
xor \U$11830 ( \12019 , \12016 , \12018 );
xor \U$11831 ( \12020 , \12012 , \12019 );
xor \U$11832 ( \12021 , \11999 , \12020 );
and \U$11833 ( \12022 , \11848 , \11852 );
and \U$11834 ( \12023 , \11852 , \11857 );
and \U$11835 ( \12024 , \11848 , \11857 );
or \U$11836 ( \12025 , \12022 , \12023 , \12024 );
and \U$11837 ( \12026 , \11836 , \11840 );
and \U$11838 ( \12027 , \11840 , \11842 );
and \U$11839 ( \12028 , \11836 , \11842 );
or \U$11840 ( \12029 , \12026 , \12027 , \12028 );
xor \U$11841 ( \12030 , \12025 , \12029 );
or \U$11842 ( \12031 , \11817 , \11831 );
xor \U$11843 ( \12032 , \12030 , \12031 );
xor \U$11844 ( \12033 , \12021 , \12032 );
xor \U$11845 ( \12034 , \11970 , \12033 );
xor \U$11846 ( \12035 , \11961 , \12034 );
and \U$11847 ( \12036 , \11784 , \11795 );
and \U$11848 ( \12037 , \11795 , \11935 );
and \U$11849 ( \12038 , \11784 , \11935 );
or \U$11850 ( \12039 , \12036 , \12037 , \12038 );
nor \U$11851 ( \12040 , \12035 , \12039 );
and \U$11852 ( \12041 , \11965 , \11969 );
and \U$11853 ( \12042 , \11969 , \12033 );
and \U$11854 ( \12043 , \11965 , \12033 );
or \U$11855 ( \12044 , \12041 , \12042 , \12043 );
and \U$11856 ( \12045 , \12025 , \12029 );
and \U$11857 ( \12046 , \12029 , \12031 );
and \U$11858 ( \12047 , \12025 , \12031 );
or \U$11859 ( \12048 , \12045 , \12046 , \12047 );
and \U$11860 ( \12049 , \12003 , \12011 );
and \U$11861 ( \12050 , \12011 , \12019 );
and \U$11862 ( \12051 , \12003 , \12019 );
or \U$11863 ( \12052 , \12049 , \12050 , \12051 );
xor \U$11864 ( \12053 , \12048 , \12052 );
and \U$11865 ( \12054 , \11984 , \11998 );
xor \U$11866 ( \12055 , \12053 , \12054 );
xor \U$11867 ( \12056 , \12044 , \12055 );
and \U$11868 ( \12057 , \11950 , \11954 );
and \U$11869 ( \12058 , \11954 , \11959 );
and \U$11870 ( \12059 , \11950 , \11959 );
or \U$11871 ( \12060 , \12057 , \12058 , \12059 );
and \U$11872 ( \12061 , \11999 , \12020 );
and \U$11873 ( \12062 , \12020 , \12032 );
and \U$11874 ( \12063 , \11999 , \12032 );
or \U$11875 ( \12064 , \12061 , \12062 , \12063 );
xor \U$11876 ( \12065 , \12060 , \12064 );
xnor \U$11877 ( \12066 , \6921 , \6923 );
xor \U$11878 ( \12067 , \6889 , \6905 );
xor \U$11879 ( \12068 , \12067 , \6915 );
xor \U$11880 ( \12069 , \12066 , \12068 );
xor \U$11881 ( \12070 , \6837 , \6853 );
xor \U$11882 ( \12071 , \12070 , \6870 );
xor \U$11883 ( \12072 , \12069 , \12071 );
and \U$11884 ( \12073 , \12005 , \12007 );
and \U$11885 ( \12074 , \12007 , \12010 );
and \U$11886 ( \12075 , \12005 , \12010 );
or \U$11887 ( \12076 , \12073 , \12074 , \12075 );
xor \U$11888 ( \12077 , \5736 , \5756 );
xor \U$11889 ( \12078 , \12077 , \5776 );
xor \U$11890 ( \12079 , \12076 , \12078 );
xor \U$11891 ( \12080 , \6929 , \6931 );
xor \U$11892 ( \12081 , \12080 , \6934 );
xor \U$11893 ( \12082 , \12079 , \12081 );
xor \U$11894 ( \12083 , \12072 , \12082 );
and \U$11895 ( \12084 , \11988 , \11992 );
and \U$11896 ( \12085 , \11992 , \11997 );
and \U$11897 ( \12086 , \11988 , \11997 );
or \U$11898 ( \12087 , \12084 , \12085 , \12086 );
and \U$11899 ( \12088 , \11974 , \11978 );
and \U$11900 ( \12089 , \11978 , \11983 );
and \U$11901 ( \12090 , \11974 , \11983 );
or \U$11902 ( \12091 , \12088 , \12089 , \12090 );
xor \U$11903 ( \12092 , \12087 , \12091 );
and \U$11904 ( \12093 , \12013 , \12015 );
and \U$11905 ( \12094 , \12015 , \12018 );
and \U$11906 ( \12095 , \12013 , \12018 );
or \U$11907 ( \12096 , \12093 , \12094 , \12095 );
xor \U$11908 ( \12097 , \12092 , \12096 );
xor \U$11909 ( \12098 , \12083 , \12097 );
xor \U$11910 ( \12099 , \12065 , \12098 );
xor \U$11911 ( \12100 , \12056 , \12099 );
and \U$11912 ( \12101 , \11946 , \11960 );
and \U$11913 ( \12102 , \11960 , \12034 );
and \U$11914 ( \12103 , \11946 , \12034 );
or \U$11915 ( \12104 , \12101 , \12102 , \12103 );
nor \U$11916 ( \12105 , \12100 , \12104 );
nor \U$11917 ( \12106 , \12040 , \12105 );
nand \U$11918 ( \12107 , \11942 , \12106 );
and \U$11919 ( \12108 , \12060 , \12064 );
and \U$11920 ( \12109 , \12064 , \12098 );
and \U$11921 ( \12110 , \12060 , \12098 );
or \U$11922 ( \12111 , \12108 , \12109 , \12110 );
and \U$11923 ( \12112 , \12087 , \12091 );
and \U$11924 ( \12113 , \12091 , \12096 );
and \U$11925 ( \12114 , \12087 , \12096 );
or \U$11926 ( \12115 , \12112 , \12113 , \12114 );
and \U$11927 ( \12116 , \12076 , \12078 );
and \U$11928 ( \12117 , \12078 , \12081 );
and \U$11929 ( \12118 , \12076 , \12081 );
or \U$11930 ( \12119 , \12116 , \12117 , \12118 );
xor \U$11931 ( \12120 , \12115 , \12119 );
and \U$11932 ( \12121 , \12066 , \12068 );
and \U$11933 ( \12122 , \12068 , \12071 );
and \U$11934 ( \12123 , \12066 , \12071 );
or \U$11935 ( \12124 , \12121 , \12122 , \12123 );
xor \U$11936 ( \12125 , \12120 , \12124 );
xor \U$11937 ( \12126 , \12111 , \12125 );
and \U$11938 ( \12127 , \12048 , \12052 );
and \U$11939 ( \12128 , \12052 , \12054 );
and \U$11940 ( \12129 , \12048 , \12054 );
or \U$11941 ( \12130 , \12127 , \12128 , \12129 );
and \U$11942 ( \12131 , \12072 , \12082 );
and \U$11943 ( \12132 , \12082 , \12097 );
and \U$11944 ( \12133 , \12072 , \12097 );
or \U$11945 ( \12134 , \12131 , \12132 , \12133 );
xor \U$11946 ( \12135 , \12130 , \12134 );
xor \U$11947 ( \12136 , \6948 , \6950 );
xor \U$11948 ( \12137 , \6937 , \6939 );
xor \U$11949 ( \12138 , \12137 , \6942 );
xor \U$11950 ( \12139 , \12136 , \12138 );
xor \U$11951 ( \12140 , \6873 , \6918 );
xor \U$11952 ( \12141 , \12140 , \6924 );
xor \U$11953 ( \12142 , \12139 , \12141 );
xor \U$11954 ( \12143 , \12135 , \12142 );
xor \U$11955 ( \12144 , \12126 , \12143 );
and \U$11956 ( \12145 , \12044 , \12055 );
and \U$11957 ( \12146 , \12055 , \12099 );
and \U$11958 ( \12147 , \12044 , \12099 );
or \U$11959 ( \12148 , \12145 , \12146 , \12147 );
nor \U$11960 ( \12149 , \12144 , \12148 );
and \U$11961 ( \12150 , \12130 , \12134 );
and \U$11962 ( \12151 , \12134 , \12142 );
and \U$11963 ( \12152 , \12130 , \12142 );
or \U$11964 ( \12153 , \12150 , \12151 , \12152 );
xor \U$11965 ( \12154 , \6927 , \6945 );
xor \U$11966 ( \12155 , \12154 , \6951 );
xor \U$11967 ( \12156 , \12153 , \12155 );
and \U$11968 ( \12157 , \12115 , \12119 );
and \U$11969 ( \12158 , \12119 , \12124 );
and \U$11970 ( \12159 , \12115 , \12124 );
or \U$11971 ( \12160 , \12157 , \12158 , \12159 );
and \U$11972 ( \12161 , \12136 , \12138 );
and \U$11973 ( \12162 , \12138 , \12141 );
and \U$11974 ( \12163 , \12136 , \12141 );
or \U$11975 ( \12164 , \12161 , \12162 , \12163 );
xor \U$11976 ( \12165 , \12160 , \12164 );
xor \U$11977 ( \12166 , \6956 , \6958 );
xor \U$11978 ( \12167 , \12166 , \6961 );
xor \U$11979 ( \12168 , \12165 , \12167 );
xor \U$11980 ( \12169 , \12156 , \12168 );
and \U$11981 ( \12170 , \12111 , \12125 );
and \U$11982 ( \12171 , \12125 , \12143 );
and \U$11983 ( \12172 , \12111 , \12143 );
or \U$11984 ( \12173 , \12170 , \12171 , \12172 );
nor \U$11985 ( \12174 , \12169 , \12173 );
nor \U$11986 ( \12175 , \12149 , \12174 );
and \U$11987 ( \12176 , \12160 , \12164 );
and \U$11988 ( \12177 , \12164 , \12167 );
and \U$11989 ( \12178 , \12160 , \12167 );
or \U$11990 ( \12179 , \12176 , \12177 , \12178 );
xor \U$11991 ( \12180 , \6122 , \6284 );
xor \U$11992 ( \12181 , \12180 , \6342 );
xor \U$11993 ( \12182 , \12179 , \12181 );
xor \U$11994 ( \12183 , \6954 , \6964 );
xor \U$11995 ( \12184 , \12183 , \6967 );
xor \U$11996 ( \12185 , \12182 , \12184 );
and \U$11997 ( \12186 , \12153 , \12155 );
and \U$11998 ( \12187 , \12155 , \12168 );
and \U$11999 ( \12188 , \12153 , \12168 );
or \U$12000 ( \12189 , \12186 , \12187 , \12188 );
nor \U$12001 ( \12190 , \12185 , \12189 );
xor \U$12002 ( \12191 , \6970 , \6972 );
xor \U$12003 ( \12192 , \12191 , \6975 );
and \U$12004 ( \12193 , \12179 , \12181 );
and \U$12005 ( \12194 , \12181 , \12184 );
and \U$12006 ( \12195 , \12179 , \12184 );
or \U$12007 ( \12196 , \12193 , \12194 , \12195 );
nor \U$12008 ( \12197 , \12192 , \12196 );
nor \U$12009 ( \12198 , \12190 , \12197 );
nand \U$12010 ( \12199 , \12175 , \12198 );
nor \U$12011 ( \12200 , \12107 , \12199 );
nand \U$12012 ( \12201 , \11617 , \12200 );
nor \U$12013 ( \12202 , \10314 , \12201 );
and \U$12014 ( \12203 , \5945 , \6991 );
and \U$12015 ( \12204 , \5957 , \6988 );
nor \U$12016 ( \12205 , \12203 , \12204 );
xnor \U$12017 ( \12206 , \12205 , \6985 );
and \U$12018 ( \12207 , \7105 , \12206 );
and \U$12019 ( \12208 , \5967 , \7006 );
and \U$12020 ( \12209 , \5979 , \7004 );
nor \U$12021 ( \12210 , \12208 , \12209 );
xnor \U$12022 ( \12211 , \12210 , \7012 );
and \U$12023 ( \12212 , \12206 , \12211 );
and \U$12024 ( \12213 , \7105 , \12211 );
or \U$12025 ( \12214 , \12207 , \12212 , \12213 );
and \U$12026 ( \12215 , \5986 , \7026 );
and \U$12027 ( \12216 , \5998 , \7024 );
nor \U$12028 ( \12217 , \12215 , \12216 );
xnor \U$12029 ( \12218 , \12217 , \7032 );
and \U$12030 ( \12219 , \6006 , \7043 );
and \U$12031 ( \12220 , \6018 , \7041 );
nor \U$12032 ( \12221 , \12219 , \12220 );
xnor \U$12033 ( \12222 , \12221 , \7049 );
and \U$12034 ( \12223 , \12218 , \12222 );
and \U$12035 ( \12224 , \6029 , \7061 );
and \U$12036 ( \12225 , \6041 , \7059 );
nor \U$12037 ( \12226 , \12224 , \12225 );
xnor \U$12038 ( \12227 , \12226 , \7067 );
and \U$12039 ( \12228 , \12222 , \12227 );
and \U$12040 ( \12229 , \12218 , \12227 );
or \U$12041 ( \12230 , \12223 , \12228 , \12229 );
and \U$12042 ( \12231 , \12214 , \12230 );
and \U$12043 ( \12232 , \6065 , \7099 );
and \U$12044 ( \12233 , \6048 , \7097 );
nor \U$12045 ( \12234 , \12232 , \12233 );
xnor \U$12046 ( \12235 , \12234 , \7105 );
and \U$12047 ( \12236 , \12230 , \12235 );
and \U$12048 ( \12237 , \12214 , \12235 );
or \U$12049 ( \12238 , \12231 , \12236 , \12237 );
and \U$12050 ( \12239 , \5967 , \7026 );
and \U$12051 ( \12240 , \5979 , \7024 );
nor \U$12052 ( \12241 , \12239 , \12240 );
xnor \U$12053 ( \12242 , \12241 , \7032 );
and \U$12054 ( \12243 , \5986 , \7043 );
and \U$12055 ( \12244 , \5998 , \7041 );
nor \U$12056 ( \12245 , \12243 , \12244 );
xnor \U$12057 ( \12246 , \12245 , \7049 );
xor \U$12058 ( \12247 , \12242 , \12246 );
and \U$12059 ( \12248 , \6006 , \7061 );
and \U$12060 ( \12249 , \6018 , \7059 );
nor \U$12061 ( \12250 , \12248 , \12249 );
xnor \U$12062 ( \12251 , \12250 , \7067 );
xor \U$12063 ( \12252 , \12247 , \12251 );
and \U$12064 ( \12253 , \5925 , \6991 );
and \U$12065 ( \12254 , \5937 , \6988 );
nor \U$12066 ( \12255 , \12253 , \12254 );
xnor \U$12067 ( \12256 , \12255 , \6985 );
xor \U$12068 ( \12257 , \7123 , \12256 );
and \U$12069 ( \12258 , \5945 , \7006 );
and \U$12070 ( \12259 , \5957 , \7004 );
nor \U$12071 ( \12260 , \12258 , \12259 );
xnor \U$12072 ( \12261 , \12260 , \7012 );
xor \U$12073 ( \12262 , \12257 , \12261 );
xor \U$12074 ( \12263 , \12252 , \12262 );
and \U$12075 ( \12264 , \12238 , \12263 );
and \U$12076 ( \12265 , \5957 , \6991 );
and \U$12077 ( \12266 , \5925 , \6988 );
nor \U$12078 ( \12267 , \12265 , \12266 );
xnor \U$12079 ( \12268 , \12267 , \6985 );
and \U$12080 ( \12269 , \5979 , \7006 );
and \U$12081 ( \12270 , \5945 , \7004 );
nor \U$12082 ( \12271 , \12269 , \12270 );
xnor \U$12083 ( \12272 , \12271 , \7012 );
and \U$12084 ( \12273 , \12268 , \12272 );
and \U$12085 ( \12274 , \5998 , \7026 );
and \U$12086 ( \12275 , \5967 , \7024 );
nor \U$12087 ( \12276 , \12274 , \12275 );
xnor \U$12088 ( \12277 , \12276 , \7032 );
and \U$12089 ( \12278 , \12272 , \12277 );
and \U$12090 ( \12279 , \12268 , \12277 );
or \U$12091 ( \12280 , \12273 , \12278 , \12279 );
and \U$12092 ( \12281 , \6018 , \7043 );
and \U$12093 ( \12282 , \5986 , \7041 );
nor \U$12094 ( \12283 , \12281 , \12282 );
xnor \U$12095 ( \12284 , \12283 , \7049 );
and \U$12096 ( \12285 , \6041 , \7061 );
and \U$12097 ( \12286 , \6006 , \7059 );
nor \U$12098 ( \12287 , \12285 , \12286 );
xnor \U$12099 ( \12288 , \12287 , \7067 );
and \U$12100 ( \12289 , \12284 , \12288 );
and \U$12101 ( \12290 , \6057 , \7082 );
and \U$12102 ( \12291 , \6029 , \7080 );
nor \U$12103 ( \12292 , \12290 , \12291 );
xnor \U$12104 ( \12293 , \12292 , \7088 );
and \U$12105 ( \12294 , \12288 , \12293 );
and \U$12106 ( \12295 , \12284 , \12293 );
or \U$12107 ( \12296 , \12289 , \12294 , \12295 );
xor \U$12108 ( \12297 , \12280 , \12296 );
and \U$12109 ( \12298 , \6029 , \7082 );
and \U$12110 ( \12299 , \6041 , \7080 );
nor \U$12111 ( \12300 , \12298 , \12299 );
xnor \U$12112 ( \12301 , \12300 , \7088 );
and \U$12113 ( \12302 , \6048 , \7099 );
and \U$12114 ( \12303 , \6057 , \7097 );
nor \U$12115 ( \12304 , \12302 , \12303 );
xnor \U$12116 ( \12305 , \12304 , \7105 );
xor \U$12117 ( \12306 , \12301 , \12305 );
nand \U$12118 ( \12307 , \6065 , \7115 );
xnor \U$12119 ( \12308 , \12307 , \7123 );
xor \U$12120 ( \12309 , \12306 , \12308 );
xor \U$12121 ( \12310 , \12297 , \12309 );
and \U$12122 ( \12311 , \12263 , \12310 );
and \U$12123 ( \12312 , \12238 , \12310 );
or \U$12124 ( \12313 , \12264 , \12311 , \12312 );
and \U$12125 ( \12314 , \7123 , \12256 );
and \U$12126 ( \12315 , \12256 , \12261 );
and \U$12127 ( \12316 , \7123 , \12261 );
or \U$12128 ( \12317 , \12314 , \12315 , \12316 );
and \U$12129 ( \12318 , \12242 , \12246 );
and \U$12130 ( \12319 , \12246 , \12251 );
and \U$12131 ( \12320 , \12242 , \12251 );
or \U$12132 ( \12321 , \12318 , \12319 , \12320 );
xor \U$12133 ( \12322 , \12317 , \12321 );
and \U$12134 ( \12323 , \12301 , \12305 );
and \U$12135 ( \12324 , \12305 , \12308 );
and \U$12136 ( \12325 , \12301 , \12308 );
or \U$12137 ( \12326 , \12323 , \12324 , \12325 );
xor \U$12138 ( \12327 , \12322 , \12326 );
xor \U$12139 ( \12328 , \12313 , \12327 );
and \U$12140 ( \12329 , \12280 , \12296 );
and \U$12141 ( \12330 , \12296 , \12309 );
and \U$12142 ( \12331 , \12280 , \12309 );
or \U$12143 ( \12332 , \12329 , \12330 , \12331 );
and \U$12144 ( \12333 , \12252 , \12262 );
xor \U$12145 ( \12334 , \12332 , \12333 );
and \U$12146 ( \12335 , \6057 , \7099 );
and \U$12147 ( \12336 , \6029 , \7097 );
nor \U$12148 ( \12337 , \12335 , \12336 );
xnor \U$12149 ( \12338 , \12337 , \7105 );
and \U$12150 ( \12339 , \6065 , \7117 );
and \U$12151 ( \12340 , \6048 , \7115 );
nor \U$12152 ( \12341 , \12339 , \12340 );
xnor \U$12153 ( \12342 , \12341 , \7123 );
xor \U$12154 ( \12343 , \12338 , \12342 );
and \U$12155 ( \12344 , \5998 , \7043 );
and \U$12156 ( \12345 , \5967 , \7041 );
nor \U$12157 ( \12346 , \12344 , \12345 );
xnor \U$12158 ( \12347 , \12346 , \7049 );
and \U$12159 ( \12348 , \6018 , \7061 );
and \U$12160 ( \12349 , \5986 , \7059 );
nor \U$12161 ( \12350 , \12348 , \12349 );
xnor \U$12162 ( \12351 , \12350 , \7067 );
xor \U$12163 ( \12352 , \12347 , \12351 );
and \U$12164 ( \12353 , \6041 , \7082 );
and \U$12165 ( \12354 , \6006 , \7080 );
nor \U$12166 ( \12355 , \12353 , \12354 );
xnor \U$12167 ( \12356 , \12355 , \7088 );
xor \U$12168 ( \12357 , \12352 , \12356 );
xor \U$12169 ( \12358 , \12343 , \12357 );
and \U$12170 ( \12359 , \5937 , \6991 );
and \U$12171 ( \12360 , \5906 , \6988 );
nor \U$12172 ( \12361 , \12359 , \12360 );
xnor \U$12173 ( \12362 , \12361 , \6985 );
and \U$12174 ( \12363 , \5957 , \7006 );
and \U$12175 ( \12364 , \5925 , \7004 );
nor \U$12176 ( \12365 , \12363 , \12364 );
xnor \U$12177 ( \12366 , \12365 , \7012 );
xor \U$12178 ( \12367 , \12362 , \12366 );
and \U$12179 ( \12368 , \5979 , \7026 );
and \U$12180 ( \12369 , \5945 , \7024 );
nor \U$12181 ( \12370 , \12368 , \12369 );
xnor \U$12182 ( \12371 , \12370 , \7032 );
xor \U$12183 ( \12372 , \12367 , \12371 );
xor \U$12184 ( \12373 , \12358 , \12372 );
xor \U$12185 ( \12374 , \12334 , \12373 );
xor \U$12186 ( \12375 , \12328 , \12374 );
and \U$12187 ( \12376 , \5979 , \6991 );
and \U$12188 ( \12377 , \5945 , \6988 );
nor \U$12189 ( \12378 , \12376 , \12377 );
xnor \U$12190 ( \12379 , \12378 , \6985 );
and \U$12191 ( \12380 , \5998 , \7006 );
and \U$12192 ( \12381 , \5967 , \7004 );
nor \U$12193 ( \12382 , \12380 , \12381 );
xnor \U$12194 ( \12383 , \12382 , \7012 );
and \U$12195 ( \12384 , \12379 , \12383 );
and \U$12196 ( \12385 , \6018 , \7026 );
and \U$12197 ( \12386 , \5986 , \7024 );
nor \U$12198 ( \12387 , \12385 , \12386 );
xnor \U$12199 ( \12388 , \12387 , \7032 );
and \U$12200 ( \12389 , \12383 , \12388 );
and \U$12201 ( \12390 , \12379 , \12388 );
or \U$12202 ( \12391 , \12384 , \12389 , \12390 );
and \U$12203 ( \12392 , \6041 , \7043 );
and \U$12204 ( \12393 , \6006 , \7041 );
nor \U$12205 ( \12394 , \12392 , \12393 );
xnor \U$12206 ( \12395 , \12394 , \7049 );
and \U$12207 ( \12396 , \6057 , \7061 );
and \U$12208 ( \12397 , \6029 , \7059 );
nor \U$12209 ( \12398 , \12396 , \12397 );
xnor \U$12210 ( \12399 , \12398 , \7067 );
and \U$12211 ( \12400 , \12395 , \12399 );
and \U$12212 ( \12401 , \6065 , \7082 );
and \U$12213 ( \12402 , \6048 , \7080 );
nor \U$12214 ( \12403 , \12401 , \12402 );
xnor \U$12215 ( \12404 , \12403 , \7088 );
and \U$12216 ( \12405 , \12399 , \12404 );
and \U$12217 ( \12406 , \12395 , \12404 );
or \U$12218 ( \12407 , \12400 , \12405 , \12406 );
and \U$12219 ( \12408 , \12391 , \12407 );
and \U$12220 ( \12409 , \6048 , \7082 );
and \U$12221 ( \12410 , \6057 , \7080 );
nor \U$12222 ( \12411 , \12409 , \12410 );
xnor \U$12223 ( \12412 , \12411 , \7088 );
and \U$12224 ( \12413 , \12407 , \12412 );
and \U$12225 ( \12414 , \12391 , \12412 );
or \U$12226 ( \12415 , \12408 , \12413 , \12414 );
nand \U$12227 ( \12416 , \6065 , \7097 );
xnor \U$12228 ( \12417 , \12416 , \7105 );
xor \U$12229 ( \12418 , \12218 , \12222 );
xor \U$12230 ( \12419 , \12418 , \12227 );
and \U$12231 ( \12420 , \12417 , \12419 );
xor \U$12232 ( \12421 , \7105 , \12206 );
xor \U$12233 ( \12422 , \12421 , \12211 );
and \U$12234 ( \12423 , \12419 , \12422 );
and \U$12235 ( \12424 , \12417 , \12422 );
or \U$12236 ( \12425 , \12420 , \12423 , \12424 );
and \U$12237 ( \12426 , \12415 , \12425 );
xor \U$12238 ( \12427 , \12284 , \12288 );
xor \U$12239 ( \12428 , \12427 , \12293 );
and \U$12240 ( \12429 , \12425 , \12428 );
and \U$12241 ( \12430 , \12415 , \12428 );
or \U$12242 ( \12431 , \12426 , \12429 , \12430 );
xor \U$12243 ( \12432 , \12268 , \12272 );
xor \U$12244 ( \12433 , \12432 , \12277 );
xor \U$12245 ( \12434 , \12214 , \12230 );
xor \U$12246 ( \12435 , \12434 , \12235 );
and \U$12247 ( \12436 , \12433 , \12435 );
and \U$12248 ( \12437 , \12431 , \12436 );
xor \U$12249 ( \12438 , \12238 , \12263 );
xor \U$12250 ( \12439 , \12438 , \12310 );
and \U$12251 ( \12440 , \12436 , \12439 );
and \U$12252 ( \12441 , \12431 , \12439 );
or \U$12253 ( \12442 , \12437 , \12440 , \12441 );
nor \U$12254 ( \12443 , \12375 , \12442 );
and \U$12255 ( \12444 , \12332 , \12333 );
and \U$12256 ( \12445 , \12333 , \12373 );
and \U$12257 ( \12446 , \12332 , \12373 );
or \U$12258 ( \12447 , \12444 , \12445 , \12446 );
nand \U$12259 ( \12448 , \6065 , \7138 );
xnor \U$12260 ( \12449 , \12448 , \7146 );
and \U$12261 ( \12450 , \6006 , \7082 );
and \U$12262 ( \12451 , \6018 , \7080 );
nor \U$12263 ( \12452 , \12450 , \12451 );
xnor \U$12264 ( \12453 , \12452 , \7088 );
and \U$12265 ( \12454 , \6029 , \7099 );
and \U$12266 ( \12455 , \6041 , \7097 );
nor \U$12267 ( \12456 , \12454 , \12455 );
xnor \U$12268 ( \12457 , \12456 , \7105 );
xor \U$12269 ( \12458 , \12453 , \12457 );
and \U$12270 ( \12459 , \6048 , \7117 );
and \U$12271 ( \12460 , \6057 , \7115 );
nor \U$12272 ( \12461 , \12459 , \12460 );
xnor \U$12273 ( \12462 , \12461 , \7123 );
xor \U$12274 ( \12463 , \12458 , \12462 );
xor \U$12275 ( \12464 , \12449 , \12463 );
and \U$12276 ( \12465 , \5945 , \7026 );
and \U$12277 ( \12466 , \5957 , \7024 );
nor \U$12278 ( \12467 , \12465 , \12466 );
xnor \U$12279 ( \12468 , \12467 , \7032 );
and \U$12280 ( \12469 , \5967 , \7043 );
and \U$12281 ( \12470 , \5979 , \7041 );
nor \U$12282 ( \12471 , \12469 , \12470 );
xnor \U$12283 ( \12472 , \12471 , \7049 );
xor \U$12284 ( \12473 , \12468 , \12472 );
and \U$12285 ( \12474 , \5986 , \7061 );
and \U$12286 ( \12475 , \5998 , \7059 );
nor \U$12287 ( \12476 , \12474 , \12475 );
xnor \U$12288 ( \12477 , \12476 , \7067 );
xor \U$12289 ( \12478 , \12473 , \12477 );
xor \U$12290 ( \12479 , \12464 , \12478 );
and \U$12291 ( \12480 , \12362 , \12366 );
and \U$12292 ( \12481 , \12366 , \12371 );
and \U$12293 ( \12482 , \12362 , \12371 );
or \U$12294 ( \12483 , \12480 , \12481 , \12482 );
and \U$12295 ( \12484 , \12347 , \12351 );
and \U$12296 ( \12485 , \12351 , \12356 );
and \U$12297 ( \12486 , \12347 , \12356 );
or \U$12298 ( \12487 , \12484 , \12485 , \12486 );
xor \U$12299 ( \12488 , \12483 , \12487 );
and \U$12300 ( \12489 , \12338 , \12342 );
xor \U$12301 ( \12490 , \12488 , \12489 );
xor \U$12302 ( \12491 , \12479 , \12490 );
xor \U$12303 ( \12492 , \12447 , \12491 );
and \U$12304 ( \12493 , \12317 , \12321 );
and \U$12305 ( \12494 , \12321 , \12326 );
and \U$12306 ( \12495 , \12317 , \12326 );
or \U$12307 ( \12496 , \12493 , \12494 , \12495 );
and \U$12308 ( \12497 , \12343 , \12357 );
and \U$12309 ( \12498 , \12357 , \12372 );
and \U$12310 ( \12499 , \12343 , \12372 );
or \U$12311 ( \12500 , \12497 , \12498 , \12499 );
xor \U$12312 ( \12501 , \12496 , \12500 );
and \U$12313 ( \12502 , \5906 , \6991 );
and \U$12314 ( \12503 , \5918 , \6988 );
nor \U$12315 ( \12504 , \12502 , \12503 );
xnor \U$12316 ( \12505 , \12504 , \6985 );
xor \U$12317 ( \12506 , \7146 , \12505 );
and \U$12318 ( \12507 , \5925 , \7006 );
and \U$12319 ( \12508 , \5937 , \7004 );
nor \U$12320 ( \12509 , \12507 , \12508 );
xnor \U$12321 ( \12510 , \12509 , \7012 );
xor \U$12322 ( \12511 , \12506 , \12510 );
xor \U$12323 ( \12512 , \12501 , \12511 );
xor \U$12324 ( \12513 , \12492 , \12512 );
and \U$12325 ( \12514 , \12313 , \12327 );
and \U$12326 ( \12515 , \12327 , \12374 );
and \U$12327 ( \12516 , \12313 , \12374 );
or \U$12328 ( \12517 , \12514 , \12515 , \12516 );
nor \U$12329 ( \12518 , \12513 , \12517 );
nor \U$12330 ( \12519 , \12443 , \12518 );
and \U$12331 ( \12520 , \12483 , \12487 );
and \U$12332 ( \12521 , \12487 , \12489 );
and \U$12333 ( \12522 , \12483 , \12489 );
or \U$12334 ( \12523 , \12520 , \12521 , \12522 );
and \U$12335 ( \12524 , \12449 , \12463 );
and \U$12336 ( \12525 , \12463 , \12478 );
and \U$12337 ( \12526 , \12449 , \12478 );
or \U$12338 ( \12527 , \12524 , \12525 , \12526 );
xor \U$12339 ( \12528 , \12523 , \12527 );
and \U$12340 ( \12529 , \6041 , \7099 );
and \U$12341 ( \12530 , \6006 , \7097 );
nor \U$12342 ( \12531 , \12529 , \12530 );
xnor \U$12343 ( \12532 , \12531 , \7105 );
and \U$12344 ( \12533 , \6057 , \7117 );
and \U$12345 ( \12534 , \6029 , \7115 );
nor \U$12346 ( \12535 , \12533 , \12534 );
xnor \U$12347 ( \12536 , \12535 , \7123 );
xor \U$12348 ( \12537 , \12532 , \12536 );
and \U$12349 ( \12538 , \6065 , \7140 );
and \U$12350 ( \12539 , \6048 , \7138 );
nor \U$12351 ( \12540 , \12538 , \12539 );
xnor \U$12352 ( \12541 , \12540 , \7146 );
xor \U$12353 ( \12542 , \12537 , \12541 );
and \U$12354 ( \12543 , \5979 , \7043 );
and \U$12355 ( \12544 , \5945 , \7041 );
nor \U$12356 ( \12545 , \12543 , \12544 );
xnor \U$12357 ( \12546 , \12545 , \7049 );
and \U$12358 ( \12547 , \5998 , \7061 );
and \U$12359 ( \12548 , \5967 , \7059 );
nor \U$12360 ( \12549 , \12547 , \12548 );
xnor \U$12361 ( \12550 , \12549 , \7067 );
xor \U$12362 ( \12551 , \12546 , \12550 );
and \U$12363 ( \12552 , \6018 , \7082 );
and \U$12364 ( \12553 , \5986 , \7080 );
nor \U$12365 ( \12554 , \12552 , \12553 );
xnor \U$12366 ( \12555 , \12554 , \7088 );
xor \U$12367 ( \12556 , \12551 , \12555 );
xor \U$12368 ( \12557 , \12542 , \12556 );
and \U$12369 ( \12558 , \5918 , \6991 );
and \U$12370 ( \12559 , \5881 , \6988 );
nor \U$12371 ( \12560 , \12558 , \12559 );
xnor \U$12372 ( \12561 , \12560 , \6985 );
and \U$12373 ( \12562 , \5937 , \7006 );
and \U$12374 ( \12563 , \5906 , \7004 );
nor \U$12375 ( \12564 , \12562 , \12563 );
xnor \U$12376 ( \12565 , \12564 , \7012 );
xor \U$12377 ( \12566 , \12561 , \12565 );
and \U$12378 ( \12567 , \5957 , \7026 );
and \U$12379 ( \12568 , \5925 , \7024 );
nor \U$12380 ( \12569 , \12567 , \12568 );
xnor \U$12381 ( \12570 , \12569 , \7032 );
xor \U$12382 ( \12571 , \12566 , \12570 );
xor \U$12383 ( \12572 , \12557 , \12571 );
xor \U$12384 ( \12573 , \12528 , \12572 );
and \U$12385 ( \12574 , \12496 , \12500 );
and \U$12386 ( \12575 , \12500 , \12511 );
and \U$12387 ( \12576 , \12496 , \12511 );
or \U$12388 ( \12577 , \12574 , \12575 , \12576 );
and \U$12389 ( \12578 , \12479 , \12490 );
xor \U$12390 ( \12579 , \12577 , \12578 );
and \U$12391 ( \12580 , \7146 , \12505 );
and \U$12392 ( \12581 , \12505 , \12510 );
and \U$12393 ( \12582 , \7146 , \12510 );
or \U$12394 ( \12583 , \12580 , \12581 , \12582 );
and \U$12395 ( \12584 , \12468 , \12472 );
and \U$12396 ( \12585 , \12472 , \12477 );
and \U$12397 ( \12586 , \12468 , \12477 );
or \U$12398 ( \12587 , \12584 , \12585 , \12586 );
xor \U$12399 ( \12588 , \12583 , \12587 );
and \U$12400 ( \12589 , \12453 , \12457 );
and \U$12401 ( \12590 , \12457 , \12462 );
and \U$12402 ( \12591 , \12453 , \12462 );
or \U$12403 ( \12592 , \12589 , \12590 , \12591 );
xor \U$12404 ( \12593 , \12588 , \12592 );
xor \U$12405 ( \12594 , \12579 , \12593 );
xor \U$12406 ( \12595 , \12573 , \12594 );
and \U$12407 ( \12596 , \12447 , \12491 );
and \U$12408 ( \12597 , \12491 , \12512 );
and \U$12409 ( \12598 , \12447 , \12512 );
or \U$12410 ( \12599 , \12596 , \12597 , \12598 );
nor \U$12411 ( \12600 , \12595 , \12599 );
and \U$12412 ( \12601 , \12577 , \12578 );
and \U$12413 ( \12602 , \12578 , \12593 );
and \U$12414 ( \12603 , \12577 , \12593 );
or \U$12415 ( \12604 , \12601 , \12602 , \12603 );
and \U$12416 ( \12605 , \12523 , \12527 );
and \U$12417 ( \12606 , \12527 , \12572 );
and \U$12418 ( \12607 , \12523 , \12572 );
or \U$12419 ( \12608 , \12605 , \12606 , \12607 );
and \U$12420 ( \12609 , \5881 , \6991 );
and \U$12421 ( \12610 , \5893 , \6988 );
nor \U$12422 ( \12611 , \12609 , \12610 );
xnor \U$12423 ( \12612 , \12611 , \6985 );
xor \U$12424 ( \12613 , \7163 , \12612 );
and \U$12425 ( \12614 , \5906 , \7006 );
and \U$12426 ( \12615 , \5918 , \7004 );
nor \U$12427 ( \12616 , \12614 , \12615 );
xnor \U$12428 ( \12617 , \12616 , \7012 );
xor \U$12429 ( \12618 , \12613 , \12617 );
and \U$12430 ( \12619 , \6048 , \7140 );
and \U$12431 ( \12620 , \6057 , \7138 );
nor \U$12432 ( \12621 , \12619 , \12620 );
xnor \U$12433 ( \12622 , \12621 , \7146 );
nand \U$12434 ( \12623 , \6065 , \7155 );
xnor \U$12435 ( \12624 , \12623 , \7163 );
xor \U$12436 ( \12625 , \12622 , \12624 );
and \U$12437 ( \12626 , \5986 , \7082 );
and \U$12438 ( \12627 , \5998 , \7080 );
nor \U$12439 ( \12628 , \12626 , \12627 );
xnor \U$12440 ( \12629 , \12628 , \7088 );
and \U$12441 ( \12630 , \6006 , \7099 );
and \U$12442 ( \12631 , \6018 , \7097 );
nor \U$12443 ( \12632 , \12630 , \12631 );
xnor \U$12444 ( \12633 , \12632 , \7105 );
xor \U$12445 ( \12634 , \12629 , \12633 );
and \U$12446 ( \12635 , \6029 , \7117 );
and \U$12447 ( \12636 , \6041 , \7115 );
nor \U$12448 ( \12637 , \12635 , \12636 );
xnor \U$12449 ( \12638 , \12637 , \7123 );
xor \U$12450 ( \12639 , \12634 , \12638 );
xor \U$12451 ( \12640 , \12625 , \12639 );
xor \U$12452 ( \12641 , \12618 , \12640 );
and \U$12453 ( \12642 , \12561 , \12565 );
and \U$12454 ( \12643 , \12565 , \12570 );
and \U$12455 ( \12644 , \12561 , \12570 );
or \U$12456 ( \12645 , \12642 , \12643 , \12644 );
and \U$12457 ( \12646 , \12546 , \12550 );
and \U$12458 ( \12647 , \12550 , \12555 );
and \U$12459 ( \12648 , \12546 , \12555 );
or \U$12460 ( \12649 , \12646 , \12647 , \12648 );
xor \U$12461 ( \12650 , \12645 , \12649 );
and \U$12462 ( \12651 , \12532 , \12536 );
and \U$12463 ( \12652 , \12536 , \12541 );
and \U$12464 ( \12653 , \12532 , \12541 );
or \U$12465 ( \12654 , \12651 , \12652 , \12653 );
xor \U$12466 ( \12655 , \12650 , \12654 );
xor \U$12467 ( \12656 , \12641 , \12655 );
xor \U$12468 ( \12657 , \12608 , \12656 );
and \U$12469 ( \12658 , \12583 , \12587 );
and \U$12470 ( \12659 , \12587 , \12592 );
and \U$12471 ( \12660 , \12583 , \12592 );
or \U$12472 ( \12661 , \12658 , \12659 , \12660 );
and \U$12473 ( \12662 , \12542 , \12556 );
and \U$12474 ( \12663 , \12556 , \12571 );
and \U$12475 ( \12664 , \12542 , \12571 );
or \U$12476 ( \12665 , \12662 , \12663 , \12664 );
xor \U$12477 ( \12666 , \12661 , \12665 );
and \U$12478 ( \12667 , \5925 , \7026 );
and \U$12479 ( \12668 , \5937 , \7024 );
nor \U$12480 ( \12669 , \12667 , \12668 );
xnor \U$12481 ( \12670 , \12669 , \7032 );
and \U$12482 ( \12671 , \5945 , \7043 );
and \U$12483 ( \12672 , \5957 , \7041 );
nor \U$12484 ( \12673 , \12671 , \12672 );
xnor \U$12485 ( \12674 , \12673 , \7049 );
xor \U$12486 ( \12675 , \12670 , \12674 );
and \U$12487 ( \12676 , \5967 , \7061 );
and \U$12488 ( \12677 , \5979 , \7059 );
nor \U$12489 ( \12678 , \12676 , \12677 );
xnor \U$12490 ( \12679 , \12678 , \7067 );
xor \U$12491 ( \12680 , \12675 , \12679 );
xor \U$12492 ( \12681 , \12666 , \12680 );
xor \U$12493 ( \12682 , \12657 , \12681 );
xor \U$12494 ( \12683 , \12604 , \12682 );
and \U$12495 ( \12684 , \12573 , \12594 );
nor \U$12496 ( \12685 , \12683 , \12684 );
nor \U$12497 ( \12686 , \12600 , \12685 );
nand \U$12498 ( \12687 , \12519 , \12686 );
and \U$12499 ( \12688 , \12608 , \12656 );
and \U$12500 ( \12689 , \12656 , \12681 );
and \U$12501 ( \12690 , \12608 , \12681 );
or \U$12502 ( \12691 , \12688 , \12689 , \12690 );
and \U$12503 ( \12692 , \7163 , \12612 );
and \U$12504 ( \12693 , \12612 , \12617 );
and \U$12505 ( \12694 , \7163 , \12617 );
or \U$12506 ( \12695 , \12692 , \12693 , \12694 );
and \U$12507 ( \12696 , \12670 , \12674 );
and \U$12508 ( \12697 , \12674 , \12679 );
and \U$12509 ( \12698 , \12670 , \12679 );
or \U$12510 ( \12699 , \12696 , \12697 , \12698 );
xor \U$12511 ( \12700 , \12695 , \12699 );
and \U$12512 ( \12701 , \12629 , \12633 );
and \U$12513 ( \12702 , \12633 , \12638 );
and \U$12514 ( \12703 , \12629 , \12638 );
or \U$12515 ( \12704 , \12701 , \12702 , \12703 );
xor \U$12516 ( \12705 , \12700 , \12704 );
and \U$12517 ( \12706 , \12645 , \12649 );
and \U$12518 ( \12707 , \12649 , \12654 );
and \U$12519 ( \12708 , \12645 , \12654 );
or \U$12520 ( \12709 , \12706 , \12707 , \12708 );
and \U$12521 ( \12710 , \12622 , \12624 );
and \U$12522 ( \12711 , \12624 , \12639 );
and \U$12523 ( \12712 , \12622 , \12639 );
or \U$12524 ( \12713 , \12710 , \12711 , \12712 );
xor \U$12525 ( \12714 , \12709 , \12713 );
and \U$12526 ( \12715 , \5893 , \6991 );
and \U$12527 ( \12716 , \5861 , \6988 );
nor \U$12528 ( \12717 , \12715 , \12716 );
xnor \U$12529 ( \12718 , \12717 , \6985 );
and \U$12530 ( \12719 , \5918 , \7006 );
and \U$12531 ( \12720 , \5881 , \7004 );
nor \U$12532 ( \12721 , \12719 , \12720 );
xnor \U$12533 ( \12722 , \12721 , \7012 );
xor \U$12534 ( \12723 , \12718 , \12722 );
and \U$12535 ( \12724 , \5937 , \7026 );
and \U$12536 ( \12725 , \5906 , \7024 );
nor \U$12537 ( \12726 , \12724 , \12725 );
xnor \U$12538 ( \12727 , \12726 , \7032 );
xor \U$12539 ( \12728 , \12723 , \12727 );
xor \U$12540 ( \12729 , \12714 , \12728 );
xor \U$12541 ( \12730 , \12705 , \12729 );
xor \U$12542 ( \12731 , \12691 , \12730 );
and \U$12543 ( \12732 , \12661 , \12665 );
and \U$12544 ( \12733 , \12665 , \12680 );
and \U$12545 ( \12734 , \12661 , \12680 );
or \U$12546 ( \12735 , \12732 , \12733 , \12734 );
and \U$12547 ( \12736 , \12618 , \12640 );
and \U$12548 ( \12737 , \12640 , \12655 );
and \U$12549 ( \12738 , \12618 , \12655 );
or \U$12550 ( \12739 , \12736 , \12737 , \12738 );
xor \U$12551 ( \12740 , \12735 , \12739 );
and \U$12552 ( \12741 , \6065 , \7157 );
and \U$12553 ( \12742 , \6048 , \7155 );
nor \U$12554 ( \12743 , \12741 , \12742 );
xnor \U$12555 ( \12744 , \12743 , \7163 );
and \U$12556 ( \12745 , \6018 , \7099 );
and \U$12557 ( \12746 , \5986 , \7097 );
nor \U$12558 ( \12747 , \12745 , \12746 );
xnor \U$12559 ( \12748 , \12747 , \7105 );
and \U$12560 ( \12749 , \6041 , \7117 );
and \U$12561 ( \12750 , \6006 , \7115 );
nor \U$12562 ( \12751 , \12749 , \12750 );
xnor \U$12563 ( \12752 , \12751 , \7123 );
xor \U$12564 ( \12753 , \12748 , \12752 );
and \U$12565 ( \12754 , \6057 , \7140 );
and \U$12566 ( \12755 , \6029 , \7138 );
nor \U$12567 ( \12756 , \12754 , \12755 );
xnor \U$12568 ( \12757 , \12756 , \7146 );
xor \U$12569 ( \12758 , \12753 , \12757 );
xor \U$12570 ( \12759 , \12744 , \12758 );
and \U$12571 ( \12760 , \5957 , \7043 );
and \U$12572 ( \12761 , \5925 , \7041 );
nor \U$12573 ( \12762 , \12760 , \12761 );
xnor \U$12574 ( \12763 , \12762 , \7049 );
and \U$12575 ( \12764 , \5979 , \7061 );
and \U$12576 ( \12765 , \5945 , \7059 );
nor \U$12577 ( \12766 , \12764 , \12765 );
xnor \U$12578 ( \12767 , \12766 , \7067 );
xor \U$12579 ( \12768 , \12763 , \12767 );
and \U$12580 ( \12769 , \5998 , \7082 );
and \U$12581 ( \12770 , \5967 , \7080 );
nor \U$12582 ( \12771 , \12769 , \12770 );
xnor \U$12583 ( \12772 , \12771 , \7088 );
xor \U$12584 ( \12773 , \12768 , \12772 );
xor \U$12585 ( \12774 , \12759 , \12773 );
xor \U$12586 ( \12775 , \12740 , \12774 );
xor \U$12587 ( \12776 , \12731 , \12775 );
and \U$12588 ( \12777 , \12604 , \12682 );
nor \U$12589 ( \12778 , \12776 , \12777 );
and \U$12590 ( \12779 , \12735 , \12739 );
and \U$12591 ( \12780 , \12739 , \12774 );
and \U$12592 ( \12781 , \12735 , \12774 );
or \U$12593 ( \12782 , \12779 , \12780 , \12781 );
and \U$12594 ( \12783 , \12705 , \12729 );
xor \U$12595 ( \12784 , \12782 , \12783 );
and \U$12596 ( \12785 , \12709 , \12713 );
and \U$12597 ( \12786 , \12713 , \12728 );
and \U$12598 ( \12787 , \12709 , \12728 );
or \U$12599 ( \12788 , \12785 , \12786 , \12787 );
and \U$12600 ( \12789 , \6029 , \7140 );
and \U$12601 ( \12790 , \6041 , \7138 );
nor \U$12602 ( \12791 , \12789 , \12790 );
xnor \U$12603 ( \12792 , \12791 , \7146 );
and \U$12604 ( \12793 , \6048 , \7157 );
and \U$12605 ( \12794 , \6057 , \7155 );
nor \U$12606 ( \12795 , \12793 , \12794 );
xnor \U$12607 ( \12796 , \12795 , \7163 );
xor \U$12608 ( \12797 , \12792 , \12796 );
nand \U$12609 ( \12798 , \6065 , \7173 );
xnor \U$12610 ( \12799 , \12798 , \7181 );
xor \U$12611 ( \12800 , \12797 , \12799 );
and \U$12612 ( \12801 , \5967 , \7082 );
and \U$12613 ( \12802 , \5979 , \7080 );
nor \U$12614 ( \12803 , \12801 , \12802 );
xnor \U$12615 ( \12804 , \12803 , \7088 );
and \U$12616 ( \12805 , \5986 , \7099 );
and \U$12617 ( \12806 , \5998 , \7097 );
nor \U$12618 ( \12807 , \12805 , \12806 );
xnor \U$12619 ( \12808 , \12807 , \7105 );
xor \U$12620 ( \12809 , \12804 , \12808 );
and \U$12621 ( \12810 , \6006 , \7117 );
and \U$12622 ( \12811 , \6018 , \7115 );
nor \U$12623 ( \12812 , \12810 , \12811 );
xnor \U$12624 ( \12813 , \12812 , \7123 );
xor \U$12625 ( \12814 , \12809 , \12813 );
xor \U$12626 ( \12815 , \12800 , \12814 );
and \U$12627 ( \12816 , \5906 , \7026 );
and \U$12628 ( \12817 , \5918 , \7024 );
nor \U$12629 ( \12818 , \12816 , \12817 );
xnor \U$12630 ( \12819 , \12818 , \7032 );
and \U$12631 ( \12820 , \5925 , \7043 );
and \U$12632 ( \12821 , \5937 , \7041 );
nor \U$12633 ( \12822 , \12820 , \12821 );
xnor \U$12634 ( \12823 , \12822 , \7049 );
xor \U$12635 ( \12824 , \12819 , \12823 );
and \U$12636 ( \12825 , \5945 , \7061 );
and \U$12637 ( \12826 , \5957 , \7059 );
nor \U$12638 ( \12827 , \12825 , \12826 );
xnor \U$12639 ( \12828 , \12827 , \7067 );
xor \U$12640 ( \12829 , \12824 , \12828 );
xor \U$12641 ( \12830 , \12815 , \12829 );
and \U$12642 ( \12831 , \12718 , \12722 );
and \U$12643 ( \12832 , \12722 , \12727 );
and \U$12644 ( \12833 , \12718 , \12727 );
or \U$12645 ( \12834 , \12831 , \12832 , \12833 );
and \U$12646 ( \12835 , \12763 , \12767 );
and \U$12647 ( \12836 , \12767 , \12772 );
and \U$12648 ( \12837 , \12763 , \12772 );
or \U$12649 ( \12838 , \12835 , \12836 , \12837 );
xor \U$12650 ( \12839 , \12834 , \12838 );
and \U$12651 ( \12840 , \12748 , \12752 );
and \U$12652 ( \12841 , \12752 , \12757 );
and \U$12653 ( \12842 , \12748 , \12757 );
or \U$12654 ( \12843 , \12840 , \12841 , \12842 );
xor \U$12655 ( \12844 , \12839 , \12843 );
xor \U$12656 ( \12845 , \12830 , \12844 );
xor \U$12657 ( \12846 , \12788 , \12845 );
and \U$12658 ( \12847 , \12695 , \12699 );
and \U$12659 ( \12848 , \12699 , \12704 );
and \U$12660 ( \12849 , \12695 , \12704 );
or \U$12661 ( \12850 , \12847 , \12848 , \12849 );
and \U$12662 ( \12851 , \12744 , \12758 );
and \U$12663 ( \12852 , \12758 , \12773 );
and \U$12664 ( \12853 , \12744 , \12773 );
or \U$12665 ( \12854 , \12851 , \12852 , \12853 );
xor \U$12666 ( \12855 , \12850 , \12854 );
and \U$12667 ( \12856 , \5861 , \6991 );
and \U$12668 ( \12857 , \5873 , \6988 );
nor \U$12669 ( \12858 , \12856 , \12857 );
xnor \U$12670 ( \12859 , \12858 , \6985 );
xor \U$12671 ( \12860 , \7181 , \12859 );
and \U$12672 ( \12861 , \5881 , \7006 );
and \U$12673 ( \12862 , \5893 , \7004 );
nor \U$12674 ( \12863 , \12861 , \12862 );
xnor \U$12675 ( \12864 , \12863 , \7012 );
xor \U$12676 ( \12865 , \12860 , \12864 );
xor \U$12677 ( \12866 , \12855 , \12865 );
xor \U$12678 ( \12867 , \12846 , \12866 );
xor \U$12679 ( \12868 , \12784 , \12867 );
and \U$12680 ( \12869 , \12691 , \12730 );
and \U$12681 ( \12870 , \12730 , \12775 );
and \U$12682 ( \12871 , \12691 , \12775 );
or \U$12683 ( \12872 , \12869 , \12870 , \12871 );
nor \U$12684 ( \12873 , \12868 , \12872 );
nor \U$12685 ( \12874 , \12778 , \12873 );
and \U$12686 ( \12875 , \12788 , \12845 );
and \U$12687 ( \12876 , \12845 , \12866 );
and \U$12688 ( \12877 , \12788 , \12866 );
or \U$12689 ( \12878 , \12875 , \12876 , \12877 );
and \U$12690 ( \12879 , \7181 , \12859 );
and \U$12691 ( \12880 , \12859 , \12864 );
and \U$12692 ( \12881 , \7181 , \12864 );
or \U$12693 ( \12882 , \12879 , \12880 , \12881 );
and \U$12694 ( \12883 , \12819 , \12823 );
and \U$12695 ( \12884 , \12823 , \12828 );
and \U$12696 ( \12885 , \12819 , \12828 );
or \U$12697 ( \12886 , \12883 , \12884 , \12885 );
xor \U$12698 ( \12887 , \12882 , \12886 );
and \U$12699 ( \12888 , \12804 , \12808 );
and \U$12700 ( \12889 , \12808 , \12813 );
and \U$12701 ( \12890 , \12804 , \12813 );
or \U$12702 ( \12891 , \12888 , \12889 , \12890 );
xor \U$12703 ( \12892 , \12887 , \12891 );
and \U$12704 ( \12893 , \12834 , \12838 );
and \U$12705 ( \12894 , \12838 , \12843 );
and \U$12706 ( \12895 , \12834 , \12843 );
or \U$12707 ( \12896 , \12893 , \12894 , \12895 );
and \U$12708 ( \12897 , \12800 , \12814 );
and \U$12709 ( \12898 , \12814 , \12829 );
and \U$12710 ( \12899 , \12800 , \12829 );
or \U$12711 ( \12900 , \12897 , \12898 , \12899 );
xor \U$12712 ( \12901 , \12896 , \12900 );
and \U$12713 ( \12902 , \5998 , \7099 );
and \U$12714 ( \12903 , \5967 , \7097 );
nor \U$12715 ( \12904 , \12902 , \12903 );
xnor \U$12716 ( \12905 , \12904 , \7105 );
and \U$12717 ( \12906 , \6018 , \7117 );
and \U$12718 ( \12907 , \5986 , \7115 );
nor \U$12719 ( \12908 , \12906 , \12907 );
xnor \U$12720 ( \12909 , \12908 , \7123 );
xor \U$12721 ( \12910 , \12905 , \12909 );
and \U$12722 ( \12911 , \6041 , \7140 );
and \U$12723 ( \12912 , \6006 , \7138 );
nor \U$12724 ( \12913 , \12911 , \12912 );
xnor \U$12725 ( \12914 , \12913 , \7146 );
xor \U$12726 ( \12915 , \12910 , \12914 );
and \U$12727 ( \12916 , \5937 , \7043 );
and \U$12728 ( \12917 , \5906 , \7041 );
nor \U$12729 ( \12918 , \12916 , \12917 );
xnor \U$12730 ( \12919 , \12918 , \7049 );
and \U$12731 ( \12920 , \5957 , \7061 );
and \U$12732 ( \12921 , \5925 , \7059 );
nor \U$12733 ( \12922 , \12920 , \12921 );
xnor \U$12734 ( \12923 , \12922 , \7067 );
xor \U$12735 ( \12924 , \12919 , \12923 );
and \U$12736 ( \12925 , \5979 , \7082 );
and \U$12737 ( \12926 , \5945 , \7080 );
nor \U$12738 ( \12927 , \12925 , \12926 );
xnor \U$12739 ( \12928 , \12927 , \7088 );
xor \U$12740 ( \12929 , \12924 , \12928 );
xor \U$12741 ( \12930 , \12915 , \12929 );
and \U$12742 ( \12931 , \5873 , \6991 );
and \U$12743 ( \12932 , \5842 , \6988 );
nor \U$12744 ( \12933 , \12931 , \12932 );
xnor \U$12745 ( \12934 , \12933 , \6985 );
and \U$12746 ( \12935 , \5893 , \7006 );
and \U$12747 ( \12936 , \5861 , \7004 );
nor \U$12748 ( \12937 , \12935 , \12936 );
xnor \U$12749 ( \12938 , \12937 , \7012 );
xor \U$12750 ( \12939 , \12934 , \12938 );
and \U$12751 ( \12940 , \5918 , \7026 );
and \U$12752 ( \12941 , \5881 , \7024 );
nor \U$12753 ( \12942 , \12940 , \12941 );
xnor \U$12754 ( \12943 , \12942 , \7032 );
xor \U$12755 ( \12944 , \12939 , \12943 );
xor \U$12756 ( \12945 , \12930 , \12944 );
xor \U$12757 ( \12946 , \12901 , \12945 );
xor \U$12758 ( \12947 , \12892 , \12946 );
xor \U$12759 ( \12948 , \12878 , \12947 );
and \U$12760 ( \12949 , \12850 , \12854 );
and \U$12761 ( \12950 , \12854 , \12865 );
and \U$12762 ( \12951 , \12850 , \12865 );
or \U$12763 ( \12952 , \12949 , \12950 , \12951 );
and \U$12764 ( \12953 , \12830 , \12844 );
xor \U$12765 ( \12954 , \12952 , \12953 );
and \U$12766 ( \12955 , \12792 , \12796 );
and \U$12767 ( \12956 , \12796 , \12799 );
and \U$12768 ( \12957 , \12792 , \12799 );
or \U$12769 ( \12958 , \12955 , \12956 , \12957 );
and \U$12770 ( \12959 , \6057 , \7157 );
and \U$12771 ( \12960 , \6029 , \7155 );
nor \U$12772 ( \12961 , \12959 , \12960 );
xnor \U$12773 ( \12962 , \12961 , \7163 );
xor \U$12774 ( \12963 , \12958 , \12962 );
and \U$12775 ( \12964 , \6065 , \7175 );
and \U$12776 ( \12965 , \6048 , \7173 );
nor \U$12777 ( \12966 , \12964 , \12965 );
xnor \U$12778 ( \12967 , \12966 , \7181 );
xor \U$12779 ( \12968 , \12963 , \12967 );
xor \U$12780 ( \12969 , \12954 , \12968 );
xor \U$12781 ( \12970 , \12948 , \12969 );
and \U$12782 ( \12971 , \12782 , \12783 );
and \U$12783 ( \12972 , \12783 , \12867 );
and \U$12784 ( \12973 , \12782 , \12867 );
or \U$12785 ( \12974 , \12971 , \12972 , \12973 );
nor \U$12786 ( \12975 , \12970 , \12974 );
and \U$12787 ( \12976 , \12952 , \12953 );
and \U$12788 ( \12977 , \12953 , \12968 );
and \U$12789 ( \12978 , \12952 , \12968 );
or \U$12790 ( \12979 , \12976 , \12977 , \12978 );
and \U$12791 ( \12980 , \12892 , \12946 );
xor \U$12792 ( \12981 , \12979 , \12980 );
and \U$12793 ( \12982 , \12896 , \12900 );
and \U$12794 ( \12983 , \12900 , \12945 );
and \U$12795 ( \12984 , \12896 , \12945 );
or \U$12796 ( \12985 , \12982 , \12983 , \12984 );
and \U$12797 ( \12986 , \5881 , \7026 );
and \U$12798 ( \12987 , \5893 , \7024 );
nor \U$12799 ( \12988 , \12986 , \12987 );
xnor \U$12800 ( \12989 , \12988 , \7032 );
and \U$12801 ( \12990 , \5906 , \7043 );
and \U$12802 ( \12991 , \5918 , \7041 );
nor \U$12803 ( \12992 , \12990 , \12991 );
xnor \U$12804 ( \12993 , \12992 , \7049 );
xor \U$12805 ( \12994 , \12989 , \12993 );
and \U$12806 ( \12995 , \5925 , \7061 );
and \U$12807 ( \12996 , \5937 , \7059 );
nor \U$12808 ( \12997 , \12995 , \12996 );
xnor \U$12809 ( \12998 , \12997 , \7067 );
xor \U$12810 ( \12999 , \12994 , \12998 );
and \U$12811 ( \13000 , \5842 , \6991 );
and \U$12812 ( \13001 , \5854 , \6988 );
nor \U$12813 ( \13002 , \13000 , \13001 );
xnor \U$12814 ( \13003 , \13002 , \6985 );
xor \U$12815 ( \13004 , \7198 , \13003 );
and \U$12816 ( \13005 , \5861 , \7006 );
and \U$12817 ( \13006 , \5873 , \7004 );
nor \U$12818 ( \13007 , \13005 , \13006 );
xnor \U$12819 ( \13008 , \13007 , \7012 );
xor \U$12820 ( \13009 , \13004 , \13008 );
xor \U$12821 ( \13010 , \12999 , \13009 );
nand \U$12822 ( \13011 , \6065 , \7190 );
xnor \U$12823 ( \13012 , \13011 , \7198 );
and \U$12824 ( \13013 , \6006 , \7140 );
and \U$12825 ( \13014 , \6018 , \7138 );
nor \U$12826 ( \13015 , \13013 , \13014 );
xnor \U$12827 ( \13016 , \13015 , \7146 );
and \U$12828 ( \13017 , \6029 , \7157 );
and \U$12829 ( \13018 , \6041 , \7155 );
nor \U$12830 ( \13019 , \13017 , \13018 );
xnor \U$12831 ( \13020 , \13019 , \7163 );
xor \U$12832 ( \13021 , \13016 , \13020 );
and \U$12833 ( \13022 , \6048 , \7175 );
and \U$12834 ( \13023 , \6057 , \7173 );
nor \U$12835 ( \13024 , \13022 , \13023 );
xnor \U$12836 ( \13025 , \13024 , \7181 );
xor \U$12837 ( \13026 , \13021 , \13025 );
xor \U$12838 ( \13027 , \13012 , \13026 );
and \U$12839 ( \13028 , \5945 , \7082 );
and \U$12840 ( \13029 , \5957 , \7080 );
nor \U$12841 ( \13030 , \13028 , \13029 );
xnor \U$12842 ( \13031 , \13030 , \7088 );
and \U$12843 ( \13032 , \5967 , \7099 );
and \U$12844 ( \13033 , \5979 , \7097 );
nor \U$12845 ( \13034 , \13032 , \13033 );
xnor \U$12846 ( \13035 , \13034 , \7105 );
xor \U$12847 ( \13036 , \13031 , \13035 );
and \U$12848 ( \13037 , \5986 , \7117 );
and \U$12849 ( \13038 , \5998 , \7115 );
nor \U$12850 ( \13039 , \13037 , \13038 );
xnor \U$12851 ( \13040 , \13039 , \7123 );
xor \U$12852 ( \13041 , \13036 , \13040 );
xor \U$12853 ( \13042 , \13027 , \13041 );
xor \U$12854 ( \13043 , \13010 , \13042 );
and \U$12855 ( \13044 , \12934 , \12938 );
and \U$12856 ( \13045 , \12938 , \12943 );
and \U$12857 ( \13046 , \12934 , \12943 );
or \U$12858 ( \13047 , \13044 , \13045 , \13046 );
and \U$12859 ( \13048 , \12919 , \12923 );
and \U$12860 ( \13049 , \12923 , \12928 );
and \U$12861 ( \13050 , \12919 , \12928 );
or \U$12862 ( \13051 , \13048 , \13049 , \13050 );
xor \U$12863 ( \13052 , \13047 , \13051 );
and \U$12864 ( \13053 , \12905 , \12909 );
and \U$12865 ( \13054 , \12909 , \12914 );
and \U$12866 ( \13055 , \12905 , \12914 );
or \U$12867 ( \13056 , \13053 , \13054 , \13055 );
xor \U$12868 ( \13057 , \13052 , \13056 );
xor \U$12869 ( \13058 , \13043 , \13057 );
xor \U$12870 ( \13059 , \12985 , \13058 );
and \U$12871 ( \13060 , \12882 , \12886 );
and \U$12872 ( \13061 , \12886 , \12891 );
and \U$12873 ( \13062 , \12882 , \12891 );
or \U$12874 ( \13063 , \13060 , \13061 , \13062 );
and \U$12875 ( \13064 , \12958 , \12962 );
and \U$12876 ( \13065 , \12962 , \12967 );
and \U$12877 ( \13066 , \12958 , \12967 );
or \U$12878 ( \13067 , \13064 , \13065 , \13066 );
xor \U$12879 ( \13068 , \13063 , \13067 );
and \U$12880 ( \13069 , \12915 , \12929 );
and \U$12881 ( \13070 , \12929 , \12944 );
and \U$12882 ( \13071 , \12915 , \12944 );
or \U$12883 ( \13072 , \13069 , \13070 , \13071 );
xor \U$12884 ( \13073 , \13068 , \13072 );
xor \U$12885 ( \13074 , \13059 , \13073 );
xor \U$12886 ( \13075 , \12981 , \13074 );
and \U$12887 ( \13076 , \12878 , \12947 );
and \U$12888 ( \13077 , \12947 , \12969 );
and \U$12889 ( \13078 , \12878 , \12969 );
or \U$12890 ( \13079 , \13076 , \13077 , \13078 );
nor \U$12891 ( \13080 , \13075 , \13079 );
nor \U$12892 ( \13081 , \12975 , \13080 );
nand \U$12893 ( \13082 , \12874 , \13081 );
nor \U$12894 ( \13083 , \12687 , \13082 );
and \U$12895 ( \13084 , \12985 , \13058 );
and \U$12896 ( \13085 , \13058 , \13073 );
and \U$12897 ( \13086 , \12985 , \13073 );
or \U$12898 ( \13087 , \13084 , \13085 , \13086 );
and \U$12899 ( \13088 , \13047 , \13051 );
and \U$12900 ( \13089 , \13051 , \13056 );
and \U$12901 ( \13090 , \13047 , \13056 );
or \U$12902 ( \13091 , \13088 , \13089 , \13090 );
and \U$12903 ( \13092 , \13012 , \13026 );
and \U$12904 ( \13093 , \13026 , \13041 );
and \U$12905 ( \13094 , \13012 , \13041 );
or \U$12906 ( \13095 , \13092 , \13093 , \13094 );
xor \U$12907 ( \13096 , \13091 , \13095 );
and \U$12908 ( \13097 , \12999 , \13009 );
xor \U$12909 ( \13098 , \13096 , \13097 );
xor \U$12910 ( \13099 , \13087 , \13098 );
and \U$12911 ( \13100 , \13063 , \13067 );
and \U$12912 ( \13101 , \13067 , \13072 );
and \U$12913 ( \13102 , \13063 , \13072 );
or \U$12914 ( \13103 , \13100 , \13101 , \13102 );
and \U$12915 ( \13104 , \13010 , \13042 );
and \U$12916 ( \13105 , \13042 , \13057 );
and \U$12917 ( \13106 , \13010 , \13057 );
or \U$12918 ( \13107 , \13104 , \13105 , \13106 );
xor \U$12919 ( \13108 , \13103 , \13107 );
and \U$12920 ( \13109 , \5918 , \7043 );
and \U$12921 ( \13110 , \5881 , \7041 );
nor \U$12922 ( \13111 , \13109 , \13110 );
xnor \U$12923 ( \13112 , \13111 , \7049 );
and \U$12924 ( \13113 , \5937 , \7061 );
and \U$12925 ( \13114 , \5906 , \7059 );
nor \U$12926 ( \13115 , \13113 , \13114 );
xnor \U$12927 ( \13116 , \13115 , \7067 );
xor \U$12928 ( \13117 , \13112 , \13116 );
and \U$12929 ( \13118 , \5957 , \7082 );
and \U$12930 ( \13119 , \5925 , \7080 );
nor \U$12931 ( \13120 , \13118 , \13119 );
xnor \U$12932 ( \13121 , \13120 , \7088 );
xor \U$12933 ( \13122 , \13117 , \13121 );
and \U$12934 ( \13123 , \5854 , \6991 );
and \U$12935 ( \13124 , \5819 , \6988 );
nor \U$12936 ( \13125 , \13123 , \13124 );
xnor \U$12937 ( \13126 , \13125 , \6985 );
and \U$12938 ( \13127 , \5873 , \7006 );
and \U$12939 ( \13128 , \5842 , \7004 );
nor \U$12940 ( \13129 , \13127 , \13128 );
xnor \U$12941 ( \13130 , \13129 , \7012 );
xor \U$12942 ( \13131 , \13126 , \13130 );
and \U$12943 ( \13132 , \5893 , \7026 );
and \U$12944 ( \13133 , \5861 , \7024 );
nor \U$12945 ( \13134 , \13132 , \13133 );
xnor \U$12946 ( \13135 , \13134 , \7032 );
xor \U$12947 ( \13136 , \13131 , \13135 );
xor \U$12948 ( \13137 , \13122 , \13136 );
and \U$12949 ( \13138 , \13016 , \13020 );
and \U$12950 ( \13139 , \13020 , \13025 );
and \U$12951 ( \13140 , \13016 , \13025 );
or \U$12952 ( \13141 , \13138 , \13139 , \13140 );
and \U$12953 ( \13142 , \6041 , \7157 );
and \U$12954 ( \13143 , \6006 , \7155 );
nor \U$12955 ( \13144 , \13142 , \13143 );
xnor \U$12956 ( \13145 , \13144 , \7163 );
and \U$12957 ( \13146 , \6057 , \7175 );
and \U$12958 ( \13147 , \6029 , \7173 );
nor \U$12959 ( \13148 , \13146 , \13147 );
xnor \U$12960 ( \13149 , \13148 , \7181 );
xor \U$12961 ( \13150 , \13145 , \13149 );
and \U$12962 ( \13151 , \6065 , \7192 );
and \U$12963 ( \13152 , \6048 , \7190 );
nor \U$12964 ( \13153 , \13151 , \13152 );
xnor \U$12965 ( \13154 , \13153 , \7198 );
xor \U$12966 ( \13155 , \13150 , \13154 );
xor \U$12967 ( \13156 , \13141 , \13155 );
and \U$12968 ( \13157 , \5979 , \7099 );
and \U$12969 ( \13158 , \5945 , \7097 );
nor \U$12970 ( \13159 , \13157 , \13158 );
xnor \U$12971 ( \13160 , \13159 , \7105 );
and \U$12972 ( \13161 , \5998 , \7117 );
and \U$12973 ( \13162 , \5967 , \7115 );
nor \U$12974 ( \13163 , \13161 , \13162 );
xnor \U$12975 ( \13164 , \13163 , \7123 );
xor \U$12976 ( \13165 , \13160 , \13164 );
and \U$12977 ( \13166 , \6018 , \7140 );
and \U$12978 ( \13167 , \5986 , \7138 );
nor \U$12979 ( \13168 , \13166 , \13167 );
xnor \U$12980 ( \13169 , \13168 , \7146 );
xor \U$12981 ( \13170 , \13165 , \13169 );
xor \U$12982 ( \13171 , \13156 , \13170 );
xor \U$12983 ( \13172 , \13137 , \13171 );
and \U$12984 ( \13173 , \7198 , \13003 );
and \U$12985 ( \13174 , \13003 , \13008 );
and \U$12986 ( \13175 , \7198 , \13008 );
or \U$12987 ( \13176 , \13173 , \13174 , \13175 );
and \U$12988 ( \13177 , \12989 , \12993 );
and \U$12989 ( \13178 , \12993 , \12998 );
and \U$12990 ( \13179 , \12989 , \12998 );
or \U$12991 ( \13180 , \13177 , \13178 , \13179 );
xor \U$12992 ( \13181 , \13176 , \13180 );
and \U$12993 ( \13182 , \13031 , \13035 );
and \U$12994 ( \13183 , \13035 , \13040 );
and \U$12995 ( \13184 , \13031 , \13040 );
or \U$12996 ( \13185 , \13182 , \13183 , \13184 );
xor \U$12997 ( \13186 , \13181 , \13185 );
xor \U$12998 ( \13187 , \13172 , \13186 );
xor \U$12999 ( \13188 , \13108 , \13187 );
xor \U$13000 ( \13189 , \13099 , \13188 );
and \U$13001 ( \13190 , \12979 , \12980 );
and \U$13002 ( \13191 , \12980 , \13074 );
and \U$13003 ( \13192 , \12979 , \13074 );
or \U$13004 ( \13193 , \13190 , \13191 , \13192 );
nor \U$13005 ( \13194 , \13189 , \13193 );
and \U$13006 ( \13195 , \13103 , \13107 );
and \U$13007 ( \13196 , \13107 , \13187 );
and \U$13008 ( \13197 , \13103 , \13187 );
or \U$13009 ( \13198 , \13195 , \13196 , \13197 );
and \U$13010 ( \13199 , \13176 , \13180 );
and \U$13011 ( \13200 , \13180 , \13185 );
and \U$13012 ( \13201 , \13176 , \13185 );
or \U$13013 ( \13202 , \13199 , \13200 , \13201 );
and \U$13014 ( \13203 , \13141 , \13155 );
and \U$13015 ( \13204 , \13155 , \13170 );
and \U$13016 ( \13205 , \13141 , \13170 );
or \U$13017 ( \13206 , \13203 , \13204 , \13205 );
xor \U$13018 ( \13207 , \13202 , \13206 );
and \U$13019 ( \13208 , \13122 , \13136 );
xor \U$13020 ( \13209 , \13207 , \13208 );
xor \U$13021 ( \13210 , \13198 , \13209 );
and \U$13022 ( \13211 , \13091 , \13095 );
and \U$13023 ( \13212 , \13095 , \13097 );
and \U$13024 ( \13213 , \13091 , \13097 );
or \U$13025 ( \13214 , \13211 , \13212 , \13213 );
and \U$13026 ( \13215 , \13137 , \13171 );
and \U$13027 ( \13216 , \13171 , \13186 );
and \U$13028 ( \13217 , \13137 , \13186 );
or \U$13029 ( \13218 , \13215 , \13216 , \13217 );
xor \U$13030 ( \13219 , \13214 , \13218 );
and \U$13031 ( \13220 , \5925 , \7082 );
and \U$13032 ( \13221 , \5937 , \7080 );
nor \U$13033 ( \13222 , \13220 , \13221 );
xnor \U$13034 ( \13223 , \13222 , \7088 );
and \U$13035 ( \13224 , \5945 , \7099 );
and \U$13036 ( \13225 , \5957 , \7097 );
nor \U$13037 ( \13226 , \13224 , \13225 );
xnor \U$13038 ( \13227 , \13226 , \7105 );
xor \U$13039 ( \13228 , \13223 , \13227 );
and \U$13040 ( \13229 , \5967 , \7117 );
and \U$13041 ( \13230 , \5979 , \7115 );
nor \U$13042 ( \13231 , \13229 , \13230 );
xnor \U$13043 ( \13232 , \13231 , \7123 );
xor \U$13044 ( \13233 , \13228 , \13232 );
and \U$13045 ( \13234 , \5861 , \7026 );
and \U$13046 ( \13235 , \5873 , \7024 );
nor \U$13047 ( \13236 , \13234 , \13235 );
xnor \U$13048 ( \13237 , \13236 , \7032 );
and \U$13049 ( \13238 , \5881 , \7043 );
and \U$13050 ( \13239 , \5893 , \7041 );
nor \U$13051 ( \13240 , \13238 , \13239 );
xnor \U$13052 ( \13241 , \13240 , \7049 );
xor \U$13053 ( \13242 , \13237 , \13241 );
and \U$13054 ( \13243 , \5906 , \7061 );
and \U$13055 ( \13244 , \5918 , \7059 );
nor \U$13056 ( \13245 , \13243 , \13244 );
xnor \U$13057 ( \13246 , \13245 , \7067 );
xor \U$13058 ( \13247 , \13242 , \13246 );
xor \U$13059 ( \13248 , \13233 , \13247 );
and \U$13060 ( \13249 , \5819 , \6991 );
and \U$13061 ( \13250 , \5831 , \6988 );
nor \U$13062 ( \13251 , \13249 , \13250 );
xnor \U$13063 ( \13252 , \13251 , \6985 );
xor \U$13064 ( \13253 , \6824 , \13252 );
and \U$13065 ( \13254 , \5842 , \7006 );
and \U$13066 ( \13255 , \5854 , \7004 );
nor \U$13067 ( \13256 , \13254 , \13255 );
xnor \U$13068 ( \13257 , \13256 , \7012 );
xor \U$13069 ( \13258 , \13253 , \13257 );
xor \U$13070 ( \13259 , \13248 , \13258 );
and \U$13071 ( \13260 , \13145 , \13149 );
and \U$13072 ( \13261 , \13149 , \13154 );
and \U$13073 ( \13262 , \13145 , \13154 );
or \U$13074 ( \13263 , \13260 , \13261 , \13262 );
and \U$13075 ( \13264 , \6048 , \7192 );
and \U$13076 ( \13265 , \6057 , \7190 );
nor \U$13077 ( \13266 , \13264 , \13265 );
xnor \U$13078 ( \13267 , \13266 , \7198 );
nand \U$13079 ( \13268 , \6065 , \7201 );
xnor \U$13080 ( \13269 , \13268 , \6824 );
xor \U$13081 ( \13270 , \13267 , \13269 );
xor \U$13082 ( \13271 , \13263 , \13270 );
and \U$13083 ( \13272 , \5986 , \7140 );
and \U$13084 ( \13273 , \5998 , \7138 );
nor \U$13085 ( \13274 , \13272 , \13273 );
xnor \U$13086 ( \13275 , \13274 , \7146 );
and \U$13087 ( \13276 , \6006 , \7157 );
and \U$13088 ( \13277 , \6018 , \7155 );
nor \U$13089 ( \13278 , \13276 , \13277 );
xnor \U$13090 ( \13279 , \13278 , \7163 );
xor \U$13091 ( \13280 , \13275 , \13279 );
and \U$13092 ( \13281 , \6029 , \7175 );
and \U$13093 ( \13282 , \6041 , \7173 );
nor \U$13094 ( \13283 , \13281 , \13282 );
xnor \U$13095 ( \13284 , \13283 , \7181 );
xor \U$13096 ( \13285 , \13280 , \13284 );
xor \U$13097 ( \13286 , \13271 , \13285 );
xor \U$13098 ( \13287 , \13259 , \13286 );
and \U$13099 ( \13288 , \13126 , \13130 );
and \U$13100 ( \13289 , \13130 , \13135 );
and \U$13101 ( \13290 , \13126 , \13135 );
or \U$13102 ( \13291 , \13288 , \13289 , \13290 );
and \U$13103 ( \13292 , \13112 , \13116 );
and \U$13104 ( \13293 , \13116 , \13121 );
and \U$13105 ( \13294 , \13112 , \13121 );
or \U$13106 ( \13295 , \13292 , \13293 , \13294 );
xor \U$13107 ( \13296 , \13291 , \13295 );
and \U$13108 ( \13297 , \13160 , \13164 );
and \U$13109 ( \13298 , \13164 , \13169 );
and \U$13110 ( \13299 , \13160 , \13169 );
or \U$13111 ( \13300 , \13297 , \13298 , \13299 );
xor \U$13112 ( \13301 , \13296 , \13300 );
xor \U$13113 ( \13302 , \13287 , \13301 );
xor \U$13114 ( \13303 , \13219 , \13302 );
xor \U$13115 ( \13304 , \13210 , \13303 );
and \U$13116 ( \13305 , \13087 , \13098 );
and \U$13117 ( \13306 , \13098 , \13188 );
and \U$13118 ( \13307 , \13087 , \13188 );
or \U$13119 ( \13308 , \13305 , \13306 , \13307 );
nor \U$13120 ( \13309 , \13304 , \13308 );
nor \U$13121 ( \13310 , \13194 , \13309 );
and \U$13122 ( \13311 , \13214 , \13218 );
and \U$13123 ( \13312 , \13218 , \13302 );
and \U$13124 ( \13313 , \13214 , \13302 );
or \U$13125 ( \13314 , \13311 , \13312 , \13313 );
xor \U$13126 ( \13315 , \7770 , \7774 );
xor \U$13127 ( \13316 , \13315 , \7779 );
xor \U$13128 ( \13317 , \7822 , \7826 );
xor \U$13129 ( \13318 , \13317 , \7831 );
xor \U$13130 ( \13319 , \7803 , \7807 );
xor \U$13131 ( \13320 , \13319 , \7812 );
xor \U$13132 ( \13321 , \13318 , \13320 );
xor \U$13133 ( \13322 , \7786 , \7790 );
xor \U$13134 ( \13323 , \13322 , \7795 );
xor \U$13135 ( \13324 , \13321 , \13323 );
xor \U$13136 ( \13325 , \13316 , \13324 );
and \U$13137 ( \13326 , \13275 , \13279 );
and \U$13138 ( \13327 , \13279 , \13284 );
and \U$13139 ( \13328 , \13275 , \13284 );
or \U$13140 ( \13329 , \13326 , \13327 , \13328 );
and \U$13141 ( \13330 , \13267 , \13269 );
xor \U$13142 ( \13331 , \13329 , \13330 );
and \U$13143 ( \13332 , \6065 , \7203 );
and \U$13144 ( \13333 , \6048 , \7201 );
nor \U$13145 ( \13334 , \13332 , \13333 );
xnor \U$13146 ( \13335 , \13334 , \6824 );
xor \U$13147 ( \13336 , \13331 , \13335 );
xor \U$13148 ( \13337 , \13325 , \13336 );
and \U$13149 ( \13338 , \13291 , \13295 );
and \U$13150 ( \13339 , \13295 , \13300 );
and \U$13151 ( \13340 , \13291 , \13300 );
or \U$13152 ( \13341 , \13338 , \13339 , \13340 );
and \U$13153 ( \13342 , \13263 , \13270 );
and \U$13154 ( \13343 , \13270 , \13285 );
and \U$13155 ( \13344 , \13263 , \13285 );
or \U$13156 ( \13345 , \13342 , \13343 , \13344 );
xor \U$13157 ( \13346 , \13341 , \13345 );
and \U$13158 ( \13347 , \13233 , \13247 );
and \U$13159 ( \13348 , \13247 , \13258 );
and \U$13160 ( \13349 , \13233 , \13258 );
or \U$13161 ( \13350 , \13347 , \13348 , \13349 );
xor \U$13162 ( \13351 , \13346 , \13350 );
xor \U$13163 ( \13352 , \13337 , \13351 );
xor \U$13164 ( \13353 , \13314 , \13352 );
and \U$13165 ( \13354 , \13202 , \13206 );
and \U$13166 ( \13355 , \13206 , \13208 );
and \U$13167 ( \13356 , \13202 , \13208 );
or \U$13168 ( \13357 , \13354 , \13355 , \13356 );
and \U$13169 ( \13358 , \13259 , \13286 );
and \U$13170 ( \13359 , \13286 , \13301 );
and \U$13171 ( \13360 , \13259 , \13301 );
or \U$13172 ( \13361 , \13358 , \13359 , \13360 );
xor \U$13173 ( \13362 , \13357 , \13361 );
and \U$13174 ( \13363 , \6824 , \13252 );
and \U$13175 ( \13364 , \13252 , \13257 );
and \U$13176 ( \13365 , \6824 , \13257 );
or \U$13177 ( \13366 , \13363 , \13364 , \13365 );
and \U$13178 ( \13367 , \13237 , \13241 );
and \U$13179 ( \13368 , \13241 , \13246 );
and \U$13180 ( \13369 , \13237 , \13246 );
or \U$13181 ( \13370 , \13367 , \13368 , \13369 );
xor \U$13182 ( \13371 , \13366 , \13370 );
and \U$13183 ( \13372 , \13223 , \13227 );
and \U$13184 ( \13373 , \13227 , \13232 );
and \U$13185 ( \13374 , \13223 , \13232 );
or \U$13186 ( \13375 , \13372 , \13373 , \13374 );
xor \U$13187 ( \13376 , \13371 , \13375 );
xor \U$13188 ( \13377 , \13362 , \13376 );
xor \U$13189 ( \13378 , \13353 , \13377 );
and \U$13190 ( \13379 , \13198 , \13209 );
and \U$13191 ( \13380 , \13209 , \13303 );
and \U$13192 ( \13381 , \13198 , \13303 );
or \U$13193 ( \13382 , \13379 , \13380 , \13381 );
nor \U$13194 ( \13383 , \13378 , \13382 );
and \U$13195 ( \13384 , \13341 , \13345 );
and \U$13196 ( \13385 , \13345 , \13350 );
and \U$13197 ( \13386 , \13341 , \13350 );
or \U$13198 ( \13387 , \13384 , \13385 , \13386 );
and \U$13199 ( \13388 , \13316 , \13324 );
and \U$13200 ( \13389 , \13324 , \13336 );
and \U$13201 ( \13390 , \13316 , \13336 );
or \U$13202 ( \13391 , \13388 , \13389 , \13390 );
xor \U$13203 ( \13392 , \13387 , \13391 );
xor \U$13204 ( \13393 , \7845 , \7847 );
xor \U$13205 ( \13394 , \13393 , \7850 );
xor \U$13206 ( \13395 , \7834 , \7836 );
xor \U$13207 ( \13396 , \13395 , \7839 );
xor \U$13208 ( \13397 , \13394 , \13396 );
xor \U$13209 ( \13398 , \7782 , \7798 );
xor \U$13210 ( \13399 , \13398 , \7815 );
xor \U$13211 ( \13400 , \13397 , \13399 );
xor \U$13212 ( \13401 , \13392 , \13400 );
and \U$13213 ( \13402 , \13357 , \13361 );
and \U$13214 ( \13403 , \13361 , \13376 );
and \U$13215 ( \13404 , \13357 , \13376 );
or \U$13216 ( \13405 , \13402 , \13403 , \13404 );
and \U$13217 ( \13406 , \13337 , \13351 );
xor \U$13218 ( \13407 , \13405 , \13406 );
and \U$13219 ( \13408 , \13366 , \13370 );
and \U$13220 ( \13409 , \13370 , \13375 );
and \U$13221 ( \13410 , \13366 , \13375 );
or \U$13222 ( \13411 , \13408 , \13409 , \13410 );
and \U$13223 ( \13412 , \13329 , \13330 );
and \U$13224 ( \13413 , \13330 , \13335 );
and \U$13225 ( \13414 , \13329 , \13335 );
or \U$13226 ( \13415 , \13412 , \13413 , \13414 );
xor \U$13227 ( \13416 , \13411 , \13415 );
and \U$13228 ( \13417 , \13318 , \13320 );
and \U$13229 ( \13418 , \13320 , \13323 );
and \U$13230 ( \13419 , \13318 , \13323 );
or \U$13231 ( \13420 , \13417 , \13418 , \13419 );
xor \U$13232 ( \13421 , \13416 , \13420 );
xor \U$13233 ( \13422 , \13407 , \13421 );
xor \U$13234 ( \13423 , \13401 , \13422 );
and \U$13235 ( \13424 , \13314 , \13352 );
and \U$13236 ( \13425 , \13352 , \13377 );
and \U$13237 ( \13426 , \13314 , \13377 );
or \U$13238 ( \13427 , \13424 , \13425 , \13426 );
nor \U$13239 ( \13428 , \13423 , \13427 );
nor \U$13240 ( \13429 , \13383 , \13428 );
nand \U$13241 ( \13430 , \13310 , \13429 );
and \U$13242 ( \13431 , \13405 , \13406 );
and \U$13243 ( \13432 , \13406 , \13421 );
and \U$13244 ( \13433 , \13405 , \13421 );
or \U$13245 ( \13434 , \13431 , \13432 , \13433 );
and \U$13246 ( \13435 , \13387 , \13391 );
and \U$13247 ( \13436 , \13391 , \13400 );
and \U$13248 ( \13437 , \13387 , \13400 );
or \U$13249 ( \13438 , \13435 , \13436 , \13437 );
xor \U$13250 ( \13439 , \7016 , \7071 );
xor \U$13251 ( \13440 , \13439 , \7127 );
xor \U$13252 ( \13441 , \7858 , \7860 );
xor \U$13253 ( \13442 , \13441 , \7863 );
xor \U$13254 ( \13443 , \13440 , \13442 );
xor \U$13255 ( \13444 , \7818 , \7842 );
xor \U$13256 ( \13445 , \13444 , \7853 );
xor \U$13257 ( \13446 , \13443 , \13445 );
xor \U$13258 ( \13447 , \13438 , \13446 );
and \U$13259 ( \13448 , \13411 , \13415 );
and \U$13260 ( \13449 , \13415 , \13420 );
and \U$13261 ( \13450 , \13411 , \13420 );
or \U$13262 ( \13451 , \13448 , \13449 , \13450 );
and \U$13263 ( \13452 , \13394 , \13396 );
and \U$13264 ( \13453 , \13396 , \13399 );
and \U$13265 ( \13454 , \13394 , \13399 );
or \U$13266 ( \13455 , \13452 , \13453 , \13454 );
xor \U$13267 ( \13456 , \13451 , \13455 );
xor \U$13268 ( \13457 , \7185 , \7213 );
xor \U$13269 ( \13458 , \13457 , \7218 );
xor \U$13270 ( \13459 , \13456 , \13458 );
xor \U$13271 ( \13460 , \13447 , \13459 );
xor \U$13272 ( \13461 , \13434 , \13460 );
and \U$13273 ( \13462 , \13401 , \13422 );
nor \U$13274 ( \13463 , \13461 , \13462 );
and \U$13275 ( \13464 , \13438 , \13446 );
and \U$13276 ( \13465 , \13446 , \13459 );
and \U$13277 ( \13466 , \13438 , \13459 );
or \U$13278 ( \13467 , \13464 , \13465 , \13466 );
xor \U$13279 ( \13468 , \7130 , \7221 );
xor \U$13280 ( \13469 , \13468 , \7258 );
xor \U$13281 ( \13470 , \7856 , \7866 );
xor \U$13282 ( \13471 , \13470 , \7869 );
xor \U$13283 ( \13472 , \13469 , \13471 );
xor \U$13284 ( \13473 , \13467 , \13472 );
and \U$13285 ( \13474 , \13451 , \13455 );
and \U$13286 ( \13475 , \13455 , \13458 );
and \U$13287 ( \13476 , \13451 , \13458 );
or \U$13288 ( \13477 , \13474 , \13475 , \13476 );
and \U$13289 ( \13478 , \13440 , \13442 );
and \U$13290 ( \13479 , \13442 , \13445 );
and \U$13291 ( \13480 , \13440 , \13445 );
or \U$13292 ( \13481 , \13478 , \13479 , \13480 );
xor \U$13293 ( \13482 , \13477 , \13481 );
xor \U$13294 ( \13483 , \7271 , \7315 );
xor \U$13295 ( \13484 , \13483 , \7338 );
xor \U$13296 ( \13485 , \13482 , \13484 );
xor \U$13297 ( \13486 , \13473 , \13485 );
and \U$13298 ( \13487 , \13434 , \13460 );
nor \U$13299 ( \13488 , \13486 , \13487 );
nor \U$13300 ( \13489 , \13463 , \13488 );
and \U$13301 ( \13490 , \13477 , \13481 );
and \U$13302 ( \13491 , \13481 , \13484 );
and \U$13303 ( \13492 , \13477 , \13484 );
or \U$13304 ( \13493 , \13490 , \13491 , \13492 );
and \U$13305 ( \13494 , \13469 , \13471 );
xor \U$13306 ( \13495 , \13493 , \13494 );
xor \U$13307 ( \13496 , \7872 , \7873 );
xor \U$13308 ( \13497 , \13496 , \7876 );
xor \U$13309 ( \13498 , \13495 , \13497 );
and \U$13310 ( \13499 , \13467 , \13472 );
and \U$13311 ( \13500 , \13472 , \13485 );
and \U$13312 ( \13501 , \13467 , \13485 );
or \U$13313 ( \13502 , \13499 , \13500 , \13501 );
nor \U$13314 ( \13503 , \13498 , \13502 );
xor \U$13315 ( \13504 , \7879 , \7880 );
xor \U$13316 ( \13505 , \13504 , \7883 );
and \U$13317 ( \13506 , \13493 , \13494 );
and \U$13318 ( \13507 , \13494 , \13497 );
and \U$13319 ( \13508 , \13493 , \13497 );
or \U$13320 ( \13509 , \13506 , \13507 , \13508 );
nor \U$13321 ( \13510 , \13505 , \13509 );
nor \U$13322 ( \13511 , \13503 , \13510 );
nand \U$13323 ( \13512 , \13489 , \13511 );
nor \U$13324 ( \13513 , \13430 , \13512 );
nand \U$13325 ( \13514 , \13083 , \13513 );
and \U$13326 ( \13515 , \6018 , \6991 );
and \U$13327 ( \13516 , \5986 , \6988 );
nor \U$13328 ( \13517 , \13515 , \13516 );
xnor \U$13329 ( \13518 , \13517 , \6985 );
and \U$13330 ( \13519 , \6041 , \7006 );
and \U$13331 ( \13520 , \6006 , \7004 );
nor \U$13332 ( \13521 , \13519 , \13520 );
xnor \U$13333 ( \13522 , \13521 , \7012 );
xor \U$13334 ( \13523 , \13518 , \13522 );
and \U$13335 ( \13524 , \6057 , \7026 );
and \U$13336 ( \13525 , \6029 , \7024 );
nor \U$13337 ( \13526 , \13524 , \13525 );
xnor \U$13338 ( \13527 , \13526 , \7032 );
xor \U$13339 ( \13528 , \13523 , \13527 );
and \U$13340 ( \13529 , \6006 , \6991 );
and \U$13341 ( \13530 , \6018 , \6988 );
nor \U$13342 ( \13531 , \13529 , \13530 );
xnor \U$13343 ( \13532 , \13531 , \6985 );
and \U$13344 ( \13533 , \7049 , \13532 );
and \U$13345 ( \13534 , \6029 , \7006 );
and \U$13346 ( \13535 , \6041 , \7004 );
nor \U$13347 ( \13536 , \13534 , \13535 );
xnor \U$13348 ( \13537 , \13536 , \7012 );
and \U$13349 ( \13538 , \13532 , \13537 );
and \U$13350 ( \13539 , \7049 , \13537 );
or \U$13351 ( \13540 , \13533 , \13538 , \13539 );
and \U$13352 ( \13541 , \6048 , \7026 );
and \U$13353 ( \13542 , \6057 , \7024 );
nor \U$13354 ( \13543 , \13541 , \13542 );
xnor \U$13355 ( \13544 , \13543 , \7032 );
nand \U$13356 ( \13545 , \6065 , \7041 );
xnor \U$13357 ( \13546 , \13545 , \7049 );
and \U$13358 ( \13547 , \13544 , \13546 );
xor \U$13359 ( \13548 , \13540 , \13547 );
and \U$13360 ( \13549 , \6065 , \7043 );
and \U$13361 ( \13550 , \6048 , \7041 );
nor \U$13362 ( \13551 , \13549 , \13550 );
xnor \U$13363 ( \13552 , \13551 , \7049 );
xor \U$13364 ( \13553 , \13548 , \13552 );
xor \U$13365 ( \13554 , \13528 , \13553 );
and \U$13366 ( \13555 , \6041 , \6991 );
and \U$13367 ( \13556 , \6006 , \6988 );
nor \U$13368 ( \13557 , \13555 , \13556 );
xnor \U$13369 ( \13558 , \13557 , \6985 );
and \U$13370 ( \13559 , \6057 , \7006 );
and \U$13371 ( \13560 , \6029 , \7004 );
nor \U$13372 ( \13561 , \13559 , \13560 );
xnor \U$13373 ( \13562 , \13561 , \7012 );
and \U$13374 ( \13563 , \13558 , \13562 );
and \U$13375 ( \13564 , \6065 , \7026 );
and \U$13376 ( \13565 , \6048 , \7024 );
nor \U$13377 ( \13566 , \13564 , \13565 );
xnor \U$13378 ( \13567 , \13566 , \7032 );
and \U$13379 ( \13568 , \13562 , \13567 );
and \U$13380 ( \13569 , \13558 , \13567 );
or \U$13381 ( \13570 , \13563 , \13568 , \13569 );
xor \U$13382 ( \13571 , \13544 , \13546 );
and \U$13383 ( \13572 , \13570 , \13571 );
xor \U$13384 ( \13573 , \7049 , \13532 );
xor \U$13385 ( \13574 , \13573 , \13537 );
and \U$13386 ( \13575 , \13571 , \13574 );
and \U$13387 ( \13576 , \13570 , \13574 );
or \U$13388 ( \13577 , \13572 , \13575 , \13576 );
nor \U$13389 ( \13578 , \13554 , \13577 );
and \U$13390 ( \13579 , \13540 , \13547 );
and \U$13391 ( \13580 , \13547 , \13552 );
and \U$13392 ( \13581 , \13540 , \13552 );
or \U$13393 ( \13582 , \13579 , \13580 , \13581 );
and \U$13394 ( \13583 , \13518 , \13522 );
and \U$13395 ( \13584 , \13522 , \13527 );
and \U$13396 ( \13585 , \13518 , \13527 );
or \U$13397 ( \13586 , \13583 , \13584 , \13585 );
and \U$13398 ( \13587 , \6029 , \7026 );
and \U$13399 ( \13588 , \6041 , \7024 );
nor \U$13400 ( \13589 , \13587 , \13588 );
xnor \U$13401 ( \13590 , \13589 , \7032 );
and \U$13402 ( \13591 , \6048 , \7043 );
and \U$13403 ( \13592 , \6057 , \7041 );
nor \U$13404 ( \13593 , \13591 , \13592 );
xnor \U$13405 ( \13594 , \13593 , \7049 );
xor \U$13406 ( \13595 , \13590 , \13594 );
nand \U$13407 ( \13596 , \6065 , \7059 );
xnor \U$13408 ( \13597 , \13596 , \7067 );
xor \U$13409 ( \13598 , \13595 , \13597 );
xor \U$13410 ( \13599 , \13586 , \13598 );
and \U$13411 ( \13600 , \5986 , \6991 );
and \U$13412 ( \13601 , \5998 , \6988 );
nor \U$13413 ( \13602 , \13600 , \13601 );
xnor \U$13414 ( \13603 , \13602 , \6985 );
xor \U$13415 ( \13604 , \7067 , \13603 );
and \U$13416 ( \13605 , \6006 , \7006 );
and \U$13417 ( \13606 , \6018 , \7004 );
nor \U$13418 ( \13607 , \13605 , \13606 );
xnor \U$13419 ( \13608 , \13607 , \7012 );
xor \U$13420 ( \13609 , \13604 , \13608 );
xor \U$13421 ( \13610 , \13599 , \13609 );
xor \U$13422 ( \13611 , \13582 , \13610 );
and \U$13423 ( \13612 , \13528 , \13553 );
nor \U$13424 ( \13613 , \13611 , \13612 );
nor \U$13425 ( \13614 , \13578 , \13613 );
and \U$13426 ( \13615 , \13586 , \13598 );
and \U$13427 ( \13616 , \13598 , \13609 );
and \U$13428 ( \13617 , \13586 , \13609 );
or \U$13429 ( \13618 , \13615 , \13616 , \13617 );
and \U$13430 ( \13619 , \6065 , \7061 );
and \U$13431 ( \13620 , \6048 , \7059 );
nor \U$13432 ( \13621 , \13619 , \13620 );
xnor \U$13433 ( \13622 , \13621 , \7067 );
and \U$13434 ( \13623 , \5998 , \6991 );
and \U$13435 ( \13624 , \5967 , \6988 );
nor \U$13436 ( \13625 , \13623 , \13624 );
xnor \U$13437 ( \13626 , \13625 , \6985 );
and \U$13438 ( \13627 , \6018 , \7006 );
and \U$13439 ( \13628 , \5986 , \7004 );
nor \U$13440 ( \13629 , \13627 , \13628 );
xnor \U$13441 ( \13630 , \13629 , \7012 );
xor \U$13442 ( \13631 , \13626 , \13630 );
and \U$13443 ( \13632 , \6041 , \7026 );
and \U$13444 ( \13633 , \6006 , \7024 );
nor \U$13445 ( \13634 , \13632 , \13633 );
xnor \U$13446 ( \13635 , \13634 , \7032 );
xor \U$13447 ( \13636 , \13631 , \13635 );
xor \U$13448 ( \13637 , \13622 , \13636 );
xor \U$13449 ( \13638 , \13618 , \13637 );
and \U$13450 ( \13639 , \7067 , \13603 );
and \U$13451 ( \13640 , \13603 , \13608 );
and \U$13452 ( \13641 , \7067 , \13608 );
or \U$13453 ( \13642 , \13639 , \13640 , \13641 );
and \U$13454 ( \13643 , \13590 , \13594 );
and \U$13455 ( \13644 , \13594 , \13597 );
and \U$13456 ( \13645 , \13590 , \13597 );
or \U$13457 ( \13646 , \13643 , \13644 , \13645 );
xor \U$13458 ( \13647 , \13642 , \13646 );
and \U$13459 ( \13648 , \6057 , \7043 );
and \U$13460 ( \13649 , \6029 , \7041 );
nor \U$13461 ( \13650 , \13648 , \13649 );
xnor \U$13462 ( \13651 , \13650 , \7049 );
xor \U$13463 ( \13652 , \13647 , \13651 );
xor \U$13464 ( \13653 , \13638 , \13652 );
and \U$13465 ( \13654 , \13582 , \13610 );
nor \U$13466 ( \13655 , \13653 , \13654 );
and \U$13467 ( \13656 , \13626 , \13630 );
and \U$13468 ( \13657 , \13630 , \13635 );
and \U$13469 ( \13658 , \13626 , \13635 );
or \U$13470 ( \13659 , \13656 , \13657 , \13658 );
nand \U$13471 ( \13660 , \6065 , \7080 );
xnor \U$13472 ( \13661 , \13660 , \7088 );
xor \U$13473 ( \13662 , \13659 , \13661 );
and \U$13474 ( \13663 , \6006 , \7026 );
and \U$13475 ( \13664 , \6018 , \7024 );
nor \U$13476 ( \13665 , \13663 , \13664 );
xnor \U$13477 ( \13666 , \13665 , \7032 );
and \U$13478 ( \13667 , \6029 , \7043 );
and \U$13479 ( \13668 , \6041 , \7041 );
nor \U$13480 ( \13669 , \13667 , \13668 );
xnor \U$13481 ( \13670 , \13669 , \7049 );
xor \U$13482 ( \13671 , \13666 , \13670 );
and \U$13483 ( \13672 , \6048 , \7061 );
and \U$13484 ( \13673 , \6057 , \7059 );
nor \U$13485 ( \13674 , \13672 , \13673 );
xnor \U$13486 ( \13675 , \13674 , \7067 );
xor \U$13487 ( \13676 , \13671 , \13675 );
xor \U$13488 ( \13677 , \13662 , \13676 );
and \U$13489 ( \13678 , \13642 , \13646 );
and \U$13490 ( \13679 , \13646 , \13651 );
and \U$13491 ( \13680 , \13642 , \13651 );
or \U$13492 ( \13681 , \13678 , \13679 , \13680 );
and \U$13493 ( \13682 , \13622 , \13636 );
xor \U$13494 ( \13683 , \13681 , \13682 );
and \U$13495 ( \13684 , \5967 , \6991 );
and \U$13496 ( \13685 , \5979 , \6988 );
nor \U$13497 ( \13686 , \13684 , \13685 );
xnor \U$13498 ( \13687 , \13686 , \6985 );
xor \U$13499 ( \13688 , \7088 , \13687 );
and \U$13500 ( \13689 , \5986 , \7006 );
and \U$13501 ( \13690 , \5998 , \7004 );
nor \U$13502 ( \13691 , \13689 , \13690 );
xnor \U$13503 ( \13692 , \13691 , \7012 );
xor \U$13504 ( \13693 , \13688 , \13692 );
xor \U$13505 ( \13694 , \13683 , \13693 );
xor \U$13506 ( \13695 , \13677 , \13694 );
and \U$13507 ( \13696 , \13618 , \13637 );
and \U$13508 ( \13697 , \13637 , \13652 );
and \U$13509 ( \13698 , \13618 , \13652 );
or \U$13510 ( \13699 , \13696 , \13697 , \13698 );
nor \U$13511 ( \13700 , \13695 , \13699 );
nor \U$13512 ( \13701 , \13655 , \13700 );
nand \U$13513 ( \13702 , \13614 , \13701 );
and \U$13514 ( \13703 , \13681 , \13682 );
and \U$13515 ( \13704 , \13682 , \13693 );
and \U$13516 ( \13705 , \13681 , \13693 );
or \U$13517 ( \13706 , \13703 , \13704 , \13705 );
and \U$13518 ( \13707 , \13659 , \13661 );
and \U$13519 ( \13708 , \13661 , \13676 );
and \U$13520 ( \13709 , \13659 , \13676 );
or \U$13521 ( \13710 , \13707 , \13708 , \13709 );
xor \U$13522 ( \13711 , \12379 , \12383 );
xor \U$13523 ( \13712 , \13711 , \12388 );
xor \U$13524 ( \13713 , \13710 , \13712 );
and \U$13525 ( \13714 , \7088 , \13687 );
and \U$13526 ( \13715 , \13687 , \13692 );
and \U$13527 ( \13716 , \7088 , \13692 );
or \U$13528 ( \13717 , \13714 , \13715 , \13716 );
and \U$13529 ( \13718 , \13666 , \13670 );
and \U$13530 ( \13719 , \13670 , \13675 );
and \U$13531 ( \13720 , \13666 , \13675 );
or \U$13532 ( \13721 , \13718 , \13719 , \13720 );
xor \U$13533 ( \13722 , \13717 , \13721 );
xor \U$13534 ( \13723 , \12395 , \12399 );
xor \U$13535 ( \13724 , \13723 , \12404 );
xor \U$13536 ( \13725 , \13722 , \13724 );
xor \U$13537 ( \13726 , \13713 , \13725 );
xor \U$13538 ( \13727 , \13706 , \13726 );
and \U$13539 ( \13728 , \13677 , \13694 );
nor \U$13540 ( \13729 , \13727 , \13728 );
and \U$13541 ( \13730 , \13710 , \13712 );
and \U$13542 ( \13731 , \13712 , \13725 );
and \U$13543 ( \13732 , \13710 , \13725 );
or \U$13544 ( \13733 , \13730 , \13731 , \13732 );
and \U$13545 ( \13734 , \13717 , \13721 );
and \U$13546 ( \13735 , \13721 , \13724 );
and \U$13547 ( \13736 , \13717 , \13724 );
or \U$13548 ( \13737 , \13734 , \13735 , \13736 );
xor \U$13549 ( \13738 , \12417 , \12419 );
xor \U$13550 ( \13739 , \13738 , \12422 );
xor \U$13551 ( \13740 , \13737 , \13739 );
xor \U$13552 ( \13741 , \12391 , \12407 );
xor \U$13553 ( \13742 , \13741 , \12412 );
xor \U$13554 ( \13743 , \13740 , \13742 );
xor \U$13555 ( \13744 , \13733 , \13743 );
and \U$13556 ( \13745 , \13706 , \13726 );
nor \U$13557 ( \13746 , \13744 , \13745 );
nor \U$13558 ( \13747 , \13729 , \13746 );
and \U$13559 ( \13748 , \13737 , \13739 );
and \U$13560 ( \13749 , \13739 , \13742 );
and \U$13561 ( \13750 , \13737 , \13742 );
or \U$13562 ( \13751 , \13748 , \13749 , \13750 );
xor \U$13563 ( \13752 , \12433 , \12435 );
xor \U$13564 ( \13753 , \13751 , \13752 );
xor \U$13565 ( \13754 , \12415 , \12425 );
xor \U$13566 ( \13755 , \13754 , \12428 );
xor \U$13567 ( \13756 , \13753 , \13755 );
and \U$13568 ( \13757 , \13733 , \13743 );
nor \U$13569 ( \13758 , \13756 , \13757 );
xor \U$13570 ( \13759 , \12431 , \12436 );
xor \U$13571 ( \13760 , \13759 , \12439 );
and \U$13572 ( \13761 , \13751 , \13752 );
and \U$13573 ( \13762 , \13752 , \13755 );
and \U$13574 ( \13763 , \13751 , \13755 );
or \U$13575 ( \13764 , \13761 , \13762 , \13763 );
nor \U$13576 ( \13765 , \13760 , \13764 );
nor \U$13577 ( \13766 , \13758 , \13765 );
nand \U$13578 ( \13767 , \13747 , \13766 );
nor \U$13579 ( \13768 , \13702 , \13767 );
and \U$13580 ( \13769 , \6057 , \6991 );
and \U$13581 ( \13770 , \6029 , \6988 );
nor \U$13582 ( \13771 , \13769 , \13770 );
xnor \U$13583 ( \13772 , \13771 , \6985 );
and \U$13584 ( \13773 , \6065 , \7006 );
and \U$13585 ( \13774 , \6048 , \7004 );
nor \U$13586 ( \13775 , \13773 , \13774 );
xnor \U$13587 ( \13776 , \13775 , \7012 );
xor \U$13588 ( \13777 , \13772 , \13776 );
and \U$13589 ( \13778 , \6048 , \6991 );
and \U$13590 ( \13779 , \6057 , \6988 );
nor \U$13591 ( \13780 , \13778 , \13779 );
xnor \U$13592 ( \13781 , \13780 , \6985 );
and \U$13593 ( \13782 , \13781 , \7012 );
nor \U$13594 ( \13783 , \13777 , \13782 );
nand \U$13595 ( \13784 , \6065 , \7024 );
xnor \U$13596 ( \13785 , \13784 , \7032 );
and \U$13597 ( \13786 , \6029 , \6991 );
and \U$13598 ( \13787 , \6041 , \6988 );
nor \U$13599 ( \13788 , \13786 , \13787 );
xnor \U$13600 ( \13789 , \13788 , \6985 );
xor \U$13601 ( \13790 , \7032 , \13789 );
and \U$13602 ( \13791 , \6048 , \7006 );
and \U$13603 ( \13792 , \6057 , \7004 );
nor \U$13604 ( \13793 , \13791 , \13792 );
xnor \U$13605 ( \13794 , \13793 , \7012 );
xor \U$13606 ( \13795 , \13790 , \13794 );
xor \U$13607 ( \13796 , \13785 , \13795 );
and \U$13608 ( \13797 , \13772 , \13776 );
nor \U$13609 ( \13798 , \13796 , \13797 );
nor \U$13610 ( \13799 , \13783 , \13798 );
and \U$13611 ( \13800 , \7032 , \13789 );
and \U$13612 ( \13801 , \13789 , \13794 );
and \U$13613 ( \13802 , \7032 , \13794 );
or \U$13614 ( \13803 , \13800 , \13801 , \13802 );
xor \U$13615 ( \13804 , \13558 , \13562 );
xor \U$13616 ( \13805 , \13804 , \13567 );
xor \U$13617 ( \13806 , \13803 , \13805 );
and \U$13618 ( \13807 , \13785 , \13795 );
nor \U$13619 ( \13808 , \13806 , \13807 );
xor \U$13620 ( \13809 , \13570 , \13571 );
xor \U$13621 ( \13810 , \13809 , \13574 );
and \U$13622 ( \13811 , \13803 , \13805 );
nor \U$13623 ( \13812 , \13810 , \13811 );
nor \U$13624 ( \13813 , \13808 , \13812 );
nand \U$13625 ( \13814 , \13799 , \13813 );
xor \U$13626 ( \13815 , \13781 , \7012 );
nand \U$13627 ( \13816 , \6065 , \7004 );
xnor \U$13628 ( \13817 , \13816 , \7012 );
nor \U$13629 ( \13818 , \13815 , \13817 );
and \U$13630 ( \13819 , \6065 , \6991 );
and \U$13631 ( \13820 , \6048 , \6988 );
nor \U$13632 ( \13821 , \13819 , \13820 );
xnor \U$13633 ( \13822 , \13821 , \6985 );
nand \U$13634 ( \13823 , \6065 , \6988 );
xnor \U$13635 ( \13824 , \13823 , \6985 );
and \U$13636 ( \13825 , \13824 , \6985 );
nand \U$13637 ( \13826 , \13822 , \13825 );
or \U$13638 ( \13827 , \13818 , \13826 );
nand \U$13639 ( \13828 , \13815 , \13817 );
nand \U$13640 ( \13829 , \13827 , \13828 );
not \U$13641 ( \13830 , \13829 );
or \U$13642 ( \13831 , \13814 , \13830 );
nand \U$13643 ( \13832 , \13777 , \13782 );
or \U$13644 ( \13833 , \13798 , \13832 );
nand \U$13645 ( \13834 , \13796 , \13797 );
nand \U$13646 ( \13835 , \13833 , \13834 );
and \U$13647 ( \13836 , \13813 , \13835 );
nand \U$13648 ( \13837 , \13806 , \13807 );
or \U$13649 ( \13838 , \13812 , \13837 );
nand \U$13650 ( \13839 , \13810 , \13811 );
nand \U$13651 ( \13840 , \13838 , \13839 );
nor \U$13652 ( \13841 , \13836 , \13840 );
nand \U$13653 ( \13842 , \13831 , \13841 );
and \U$13654 ( \13843 , \13768 , \13842 );
nand \U$13655 ( \13844 , \13554 , \13577 );
or \U$13656 ( \13845 , \13613 , \13844 );
nand \U$13657 ( \13846 , \13611 , \13612 );
nand \U$13658 ( \13847 , \13845 , \13846 );
and \U$13659 ( \13848 , \13701 , \13847 );
nand \U$13660 ( \13849 , \13653 , \13654 );
or \U$13661 ( \13850 , \13700 , \13849 );
nand \U$13662 ( \13851 , \13695 , \13699 );
nand \U$13663 ( \13852 , \13850 , \13851 );
nor \U$13664 ( \13853 , \13848 , \13852 );
or \U$13665 ( \13854 , \13767 , \13853 );
nand \U$13666 ( \13855 , \13727 , \13728 );
or \U$13667 ( \13856 , \13746 , \13855 );
nand \U$13668 ( \13857 , \13744 , \13745 );
nand \U$13669 ( \13858 , \13856 , \13857 );
and \U$13670 ( \13859 , \13766 , \13858 );
nand \U$13671 ( \13860 , \13756 , \13757 );
or \U$13672 ( \13861 , \13765 , \13860 );
nand \U$13673 ( \13862 , \13760 , \13764 );
nand \U$13674 ( \13863 , \13861 , \13862 );
nor \U$13675 ( \13864 , \13859 , \13863 );
nand \U$13676 ( \13865 , \13854 , \13864 );
nor \U$13677 ( \13866 , \13843 , \13865 );
or \U$13678 ( \13867 , \13514 , \13866 );
nand \U$13679 ( \13868 , \12375 , \12442 );
or \U$13680 ( \13869 , \12518 , \13868 );
nand \U$13681 ( \13870 , \12513 , \12517 );
nand \U$13682 ( \13871 , \13869 , \13870 );
and \U$13683 ( \13872 , \12686 , \13871 );
nand \U$13684 ( \13873 , \12595 , \12599 );
or \U$13685 ( \13874 , \12685 , \13873 );
nand \U$13686 ( \13875 , \12683 , \12684 );
nand \U$13687 ( \13876 , \13874 , \13875 );
nor \U$13688 ( \13877 , \13872 , \13876 );
or \U$13689 ( \13878 , \13082 , \13877 );
nand \U$13690 ( \13879 , \12776 , \12777 );
or \U$13691 ( \13880 , \12873 , \13879 );
nand \U$13692 ( \13881 , \12868 , \12872 );
nand \U$13693 ( \13882 , \13880 , \13881 );
and \U$13694 ( \13883 , \13081 , \13882 );
nand \U$13695 ( \13884 , \12970 , \12974 );
or \U$13696 ( \13885 , \13080 , \13884 );
nand \U$13697 ( \13886 , \13075 , \13079 );
nand \U$13698 ( \13887 , \13885 , \13886 );
nor \U$13699 ( \13888 , \13883 , \13887 );
nand \U$13700 ( \13889 , \13878 , \13888 );
and \U$13701 ( \13890 , \13513 , \13889 );
nand \U$13702 ( \13891 , \13189 , \13193 );
or \U$13703 ( \13892 , \13309 , \13891 );
nand \U$13704 ( \13893 , \13304 , \13308 );
nand \U$13705 ( \13894 , \13892 , \13893 );
and \U$13706 ( \13895 , \13429 , \13894 );
nand \U$13707 ( \13896 , \13378 , \13382 );
or \U$13708 ( \13897 , \13428 , \13896 );
nand \U$13709 ( \13898 , \13423 , \13427 );
nand \U$13710 ( \13899 , \13897 , \13898 );
nor \U$13711 ( \13900 , \13895 , \13899 );
or \U$13712 ( \13901 , \13512 , \13900 );
nand \U$13713 ( \13902 , \13461 , \13462 );
or \U$13714 ( \13903 , \13488 , \13902 );
nand \U$13715 ( \13904 , \13486 , \13487 );
nand \U$13716 ( \13905 , \13903 , \13904 );
and \U$13717 ( \13906 , \13511 , \13905 );
nand \U$13718 ( \13907 , \13498 , \13502 );
or \U$13719 ( \13908 , \13510 , \13907 );
nand \U$13720 ( \13909 , \13505 , \13509 );
nand \U$13721 ( \13910 , \13908 , \13909 );
nor \U$13722 ( \13911 , \13906 , \13910 );
nand \U$13723 ( \13912 , \13901 , \13911 );
nor \U$13724 ( \13913 , \13890 , \13912 );
nand \U$13725 ( \13914 , \13867 , \13913 );
and \U$13726 ( \13915 , \12202 , \13914 );
nand \U$13727 ( \13916 , \7766 , \7886 );
or \U$13728 ( \13917 , \8041 , \13916 );
nand \U$13729 ( \13918 , \8036 , \8040 );
nand \U$13730 ( \13919 , \13917 , \13918 );
and \U$13731 ( \13920 , \8360 , \13919 );
nand \U$13732 ( \13921 , \8195 , \8199 );
or \U$13733 ( \13922 , \8359 , \13921 );
nand \U$13734 ( \13923 , \8354 , \8358 );
nand \U$13735 ( \13924 , \13922 , \13923 );
nor \U$13736 ( \13925 , \13920 , \13924 );
or \U$13737 ( \13926 , \9009 , \13925 );
nand \U$13738 ( \13927 , \8516 , \8520 );
or \U$13739 ( \13928 , \8682 , \13927 );
nand \U$13740 ( \13929 , \8677 , \8681 );
nand \U$13741 ( \13930 , \13928 , \13929 );
and \U$13742 ( \13931 , \9008 , \13930 );
nand \U$13743 ( \13932 , \8841 , \8845 );
or \U$13744 ( \13933 , \9007 , \13932 );
nand \U$13745 ( \13934 , \9002 , \9006 );
nand \U$13746 ( \13935 , \13933 , \13934 );
nor \U$13747 ( \13936 , \13931 , \13935 );
nand \U$13748 ( \13937 , \13926 , \13936 );
and \U$13749 ( \13938 , \10313 , \13937 );
nand \U$13750 ( \13939 , \9168 , \9172 );
or \U$13751 ( \13940 , \9334 , \13939 );
nand \U$13752 ( \13941 , \9329 , \9333 );
nand \U$13753 ( \13942 , \13940 , \13941 );
and \U$13754 ( \13943 , \9660 , \13942 );
nand \U$13755 ( \13944 , \9493 , \9497 );
or \U$13756 ( \13945 , \9659 , \13944 );
nand \U$13757 ( \13946 , \9654 , \9658 );
nand \U$13758 ( \13947 , \13945 , \13946 );
nor \U$13759 ( \13948 , \13943 , \13947 );
or \U$13760 ( \13949 , \10312 , \13948 );
nand \U$13761 ( \13950 , \9819 , \9823 );
or \U$13762 ( \13951 , \9985 , \13950 );
nand \U$13763 ( \13952 , \9980 , \9984 );
nand \U$13764 ( \13953 , \13951 , \13952 );
and \U$13765 ( \13954 , \10311 , \13953 );
nand \U$13766 ( \13955 , \10144 , \10148 );
or \U$13767 ( \13956 , \10310 , \13955 );
nand \U$13768 ( \13957 , \10305 , \10309 );
nand \U$13769 ( \13958 , \13956 , \13957 );
nor \U$13770 ( \13959 , \13954 , \13958 );
nand \U$13771 ( \13960 , \13949 , \13959 );
nor \U$13772 ( \13961 , \13938 , \13960 );
or \U$13773 ( \13962 , \12201 , \13961 );
nand \U$13774 ( \13963 , \10472 , \10476 );
or \U$13775 ( \13964 , \10638 , \13963 );
nand \U$13776 ( \13965 , \10633 , \10637 );
nand \U$13777 ( \13966 , \13964 , \13965 );
and \U$13778 ( \13967 , \10964 , \13966 );
nand \U$13779 ( \13968 , \10797 , \10801 );
or \U$13780 ( \13969 , \10963 , \13968 );
nand \U$13781 ( \13970 , \10958 , \10962 );
nand \U$13782 ( \13971 , \13969 , \13970 );
nor \U$13783 ( \13972 , \13967 , \13971 );
or \U$13784 ( \13973 , \11616 , \13972 );
nand \U$13785 ( \13974 , \11123 , \11127 );
or \U$13786 ( \13975 , \11289 , \13974 );
nand \U$13787 ( \13976 , \11284 , \11288 );
nand \U$13788 ( \13977 , \13975 , \13976 );
and \U$13789 ( \13978 , \11615 , \13977 );
nand \U$13790 ( \13979 , \11448 , \11452 );
or \U$13791 ( \13980 , \11614 , \13979 );
nand \U$13792 ( \13981 , \11609 , \11613 );
nand \U$13793 ( \13982 , \13980 , \13981 );
nor \U$13794 ( \13983 , \13978 , \13982 );
nand \U$13795 ( \13984 , \13973 , \13983 );
and \U$13796 ( \13985 , \12200 , \13984 );
nand \U$13797 ( \13986 , \11775 , \11779 );
or \U$13798 ( \13987 , \11941 , \13986 );
nand \U$13799 ( \13988 , \11936 , \11940 );
nand \U$13800 ( \13989 , \13987 , \13988 );
and \U$13801 ( \13990 , \12106 , \13989 );
nand \U$13802 ( \13991 , \12035 , \12039 );
or \U$13803 ( \13992 , \12105 , \13991 );
nand \U$13804 ( \13993 , \12100 , \12104 );
nand \U$13805 ( \13994 , \13992 , \13993 );
nor \U$13806 ( \13995 , \13990 , \13994 );
or \U$13807 ( \13996 , \12199 , \13995 );
nand \U$13808 ( \13997 , \12144 , \12148 );
or \U$13809 ( \13998 , \12174 , \13997 );
nand \U$13810 ( \13999 , \12169 , \12173 );
nand \U$13811 ( \14000 , \13998 , \13999 );
and \U$13812 ( \14001 , \12198 , \14000 );
nand \U$13813 ( \14002 , \12185 , \12189 );
or \U$13814 ( \14003 , \12197 , \14002 );
nand \U$13815 ( \14004 , \12192 , \12196 );
nand \U$13816 ( \14005 , \14003 , \14004 );
nor \U$13817 ( \14006 , \14001 , \14005 );
nand \U$13818 ( \14007 , \13996 , \14006 );
nor \U$13819 ( \14008 , \13985 , \14007 );
nand \U$13820 ( \14009 , \13962 , \14008 );
nor \U$13821 ( \14010 , \13915 , \14009 );
not \U$13822 ( \14011 , \14010 );
xnor \U$13823 ( \14012 , \6982 , \14011 );
buf \U$13824 ( \14013 , \14012 );
buf \U$13825 ( \14014 , \14013 );
not \U$13826 ( \14015 , \12197 );
nand \U$13827 ( \14016 , \14004 , \14015 );
nor \U$13828 ( \14017 , \13510 , \7887 );
nor \U$13829 ( \14018 , \8041 , \8200 );
nand \U$13830 ( \14019 , \14017 , \14018 );
nor \U$13831 ( \14020 , \8359 , \8521 );
nor \U$13832 ( \14021 , \8682 , \8846 );
nand \U$13833 ( \14022 , \14020 , \14021 );
nor \U$13834 ( \14023 , \14019 , \14022 );
nor \U$13835 ( \14024 , \9007 , \9173 );
nor \U$13836 ( \14025 , \9334 , \9498 );
nand \U$13837 ( \14026 , \14024 , \14025 );
nor \U$13838 ( \14027 , \9659 , \9824 );
nor \U$13839 ( \14028 , \9985 , \10149 );
nand \U$13840 ( \14029 , \14027 , \14028 );
nor \U$13841 ( \14030 , \14026 , \14029 );
nand \U$13842 ( \14031 , \14023 , \14030 );
nor \U$13843 ( \14032 , \10310 , \10477 );
nor \U$13844 ( \14033 , \10638 , \10802 );
nand \U$13845 ( \14034 , \14032 , \14033 );
nor \U$13846 ( \14035 , \10963 , \11128 );
nor \U$13847 ( \14036 , \11289 , \11453 );
nand \U$13848 ( \14037 , \14035 , \14036 );
nor \U$13849 ( \14038 , \14034 , \14037 );
nor \U$13850 ( \14039 , \11614 , \11780 );
nor \U$13851 ( \14040 , \11941 , \12040 );
nand \U$13852 ( \14041 , \14039 , \14040 );
nor \U$13853 ( \14042 , \12105 , \12149 );
nor \U$13854 ( \14043 , \12174 , \12190 );
nand \U$13855 ( \14044 , \14042 , \14043 );
nor \U$13856 ( \14045 , \14041 , \14044 );
nand \U$13857 ( \14046 , \14038 , \14045 );
nor \U$13858 ( \14047 , \14031 , \14046 );
nor \U$13859 ( \14048 , \13765 , \12443 );
nor \U$13860 ( \14049 , \12518 , \12600 );
nand \U$13861 ( \14050 , \14048 , \14049 );
nor \U$13862 ( \14051 , \12685 , \12778 );
nor \U$13863 ( \14052 , \12873 , \12975 );
nand \U$13864 ( \14053 , \14051 , \14052 );
nor \U$13865 ( \14054 , \14050 , \14053 );
nor \U$13866 ( \14055 , \13080 , \13194 );
nor \U$13867 ( \14056 , \13309 , \13383 );
nand \U$13868 ( \14057 , \14055 , \14056 );
nor \U$13869 ( \14058 , \13428 , \13463 );
nor \U$13870 ( \14059 , \13488 , \13503 );
nand \U$13871 ( \14060 , \14058 , \14059 );
nor \U$13872 ( \14061 , \14057 , \14060 );
nand \U$13873 ( \14062 , \14054 , \14061 );
nor \U$13874 ( \14063 , \13812 , \13578 );
nor \U$13875 ( \14064 , \13613 , \13655 );
nand \U$13876 ( \14065 , \14063 , \14064 );
nor \U$13877 ( \14066 , \13700 , \13729 );
nor \U$13878 ( \14067 , \13746 , \13758 );
nand \U$13879 ( \14068 , \14066 , \14067 );
nor \U$13880 ( \14069 , \14065 , \14068 );
nor \U$13881 ( \14070 , \13818 , \13783 );
nor \U$13882 ( \14071 , \13798 , \13808 );
nand \U$13883 ( \14072 , \14070 , \14071 );
or \U$13884 ( \14073 , \14072 , \13826 );
or \U$13885 ( \14074 , \13783 , \13828 );
nand \U$13886 ( \14075 , \14074 , \13832 );
and \U$13887 ( \14076 , \14071 , \14075 );
or \U$13888 ( \14077 , \13808 , \13834 );
nand \U$13889 ( \14078 , \14077 , \13837 );
nor \U$13890 ( \14079 , \14076 , \14078 );
nand \U$13891 ( \14080 , \14073 , \14079 );
and \U$13892 ( \14081 , \14069 , \14080 );
or \U$13893 ( \14082 , \13578 , \13839 );
nand \U$13894 ( \14083 , \14082 , \13844 );
and \U$13895 ( \14084 , \14064 , \14083 );
or \U$13896 ( \14085 , \13655 , \13846 );
nand \U$13897 ( \14086 , \14085 , \13849 );
nor \U$13898 ( \14087 , \14084 , \14086 );
or \U$13899 ( \14088 , \14068 , \14087 );
or \U$13900 ( \14089 , \13729 , \13851 );
nand \U$13901 ( \14090 , \14089 , \13855 );
and \U$13902 ( \14091 , \14067 , \14090 );
or \U$13903 ( \14092 , \13758 , \13857 );
nand \U$13904 ( \14093 , \14092 , \13860 );
nor \U$13905 ( \14094 , \14091 , \14093 );
nand \U$13906 ( \14095 , \14088 , \14094 );
nor \U$13907 ( \14096 , \14081 , \14095 );
or \U$13908 ( \14097 , \14062 , \14096 );
or \U$13909 ( \14098 , \12443 , \13862 );
nand \U$13910 ( \14099 , \14098 , \13868 );
and \U$13911 ( \14100 , \14049 , \14099 );
or \U$13912 ( \14101 , \12600 , \13870 );
nand \U$13913 ( \14102 , \14101 , \13873 );
nor \U$13914 ( \14103 , \14100 , \14102 );
or \U$13915 ( \14104 , \14053 , \14103 );
or \U$13916 ( \14105 , \12778 , \13875 );
nand \U$13917 ( \14106 , \14105 , \13879 );
and \U$13918 ( \14107 , \14052 , \14106 );
or \U$13919 ( \14108 , \12975 , \13881 );
nand \U$13920 ( \14109 , \14108 , \13884 );
nor \U$13921 ( \14110 , \14107 , \14109 );
nand \U$13922 ( \14111 , \14104 , \14110 );
and \U$13923 ( \14112 , \14061 , \14111 );
or \U$13924 ( \14113 , \13194 , \13886 );
nand \U$13925 ( \14114 , \14113 , \13891 );
and \U$13926 ( \14115 , \14056 , \14114 );
or \U$13927 ( \14116 , \13383 , \13893 );
nand \U$13928 ( \14117 , \14116 , \13896 );
nor \U$13929 ( \14118 , \14115 , \14117 );
or \U$13930 ( \14119 , \14060 , \14118 );
or \U$13931 ( \14120 , \13463 , \13898 );
nand \U$13932 ( \14121 , \14120 , \13902 );
and \U$13933 ( \14122 , \14059 , \14121 );
or \U$13934 ( \14123 , \13503 , \13904 );
nand \U$13935 ( \14124 , \14123 , \13907 );
nor \U$13936 ( \14125 , \14122 , \14124 );
nand \U$13937 ( \14126 , \14119 , \14125 );
nor \U$13938 ( \14127 , \14112 , \14126 );
nand \U$13939 ( \14128 , \14097 , \14127 );
and \U$13940 ( \14129 , \14047 , \14128 );
or \U$13941 ( \14130 , \7887 , \13909 );
nand \U$13942 ( \14131 , \14130 , \13916 );
and \U$13943 ( \14132 , \14018 , \14131 );
or \U$13944 ( \14133 , \8200 , \13918 );
nand \U$13945 ( \14134 , \14133 , \13921 );
nor \U$13946 ( \14135 , \14132 , \14134 );
or \U$13947 ( \14136 , \14022 , \14135 );
or \U$13948 ( \14137 , \8521 , \13923 );
nand \U$13949 ( \14138 , \14137 , \13927 );
and \U$13950 ( \14139 , \14021 , \14138 );
or \U$13951 ( \14140 , \8846 , \13929 );
nand \U$13952 ( \14141 , \14140 , \13932 );
nor \U$13953 ( \14142 , \14139 , \14141 );
nand \U$13954 ( \14143 , \14136 , \14142 );
and \U$13955 ( \14144 , \14030 , \14143 );
or \U$13956 ( \14145 , \9173 , \13934 );
nand \U$13957 ( \14146 , \14145 , \13939 );
and \U$13958 ( \14147 , \14025 , \14146 );
or \U$13959 ( \14148 , \9498 , \13941 );
nand \U$13960 ( \14149 , \14148 , \13944 );
nor \U$13961 ( \14150 , \14147 , \14149 );
or \U$13962 ( \14151 , \14029 , \14150 );
or \U$13963 ( \14152 , \9824 , \13946 );
nand \U$13964 ( \14153 , \14152 , \13950 );
and \U$13965 ( \14154 , \14028 , \14153 );
or \U$13966 ( \14155 , \10149 , \13952 );
nand \U$13967 ( \14156 , \14155 , \13955 );
nor \U$13968 ( \14157 , \14154 , \14156 );
nand \U$13969 ( \14158 , \14151 , \14157 );
nor \U$13970 ( \14159 , \14144 , \14158 );
or \U$13971 ( \14160 , \14046 , \14159 );
or \U$13972 ( \14161 , \10477 , \13957 );
nand \U$13973 ( \14162 , \14161 , \13963 );
and \U$13974 ( \14163 , \14033 , \14162 );
or \U$13975 ( \14164 , \10802 , \13965 );
nand \U$13976 ( \14165 , \14164 , \13968 );
nor \U$13977 ( \14166 , \14163 , \14165 );
or \U$13978 ( \14167 , \14037 , \14166 );
or \U$13979 ( \14168 , \11128 , \13970 );
nand \U$13980 ( \14169 , \14168 , \13974 );
and \U$13981 ( \14170 , \14036 , \14169 );
or \U$13982 ( \14171 , \11453 , \13976 );
nand \U$13983 ( \14172 , \14171 , \13979 );
nor \U$13984 ( \14173 , \14170 , \14172 );
nand \U$13985 ( \14174 , \14167 , \14173 );
and \U$13986 ( \14175 , \14045 , \14174 );
or \U$13987 ( \14176 , \11780 , \13981 );
nand \U$13988 ( \14177 , \14176 , \13986 );
and \U$13989 ( \14178 , \14040 , \14177 );
or \U$13990 ( \14179 , \12040 , \13988 );
nand \U$13991 ( \14180 , \14179 , \13991 );
nor \U$13992 ( \14181 , \14178 , \14180 );
or \U$13993 ( \14182 , \14044 , \14181 );
or \U$13994 ( \14183 , \12149 , \13993 );
nand \U$13995 ( \14184 , \14183 , \13997 );
and \U$13996 ( \14185 , \14043 , \14184 );
or \U$13997 ( \14186 , \12190 , \13999 );
nand \U$13998 ( \14187 , \14186 , \14002 );
nor \U$13999 ( \14188 , \14185 , \14187 );
nand \U$14000 ( \14189 , \14182 , \14188 );
nor \U$14001 ( \14190 , \14175 , \14189 );
nand \U$14002 ( \14191 , \14160 , \14190 );
nor \U$14003 ( \14192 , \14129 , \14191 );
not \U$14004 ( \14193 , \14192 );
xnor \U$14005 ( \14194 , \14016 , \14193 );
buf \U$14006 ( \14195 , \14194 );
buf \U$14007 ( \14196 , \14195 );
not \U$14008 ( \14197 , \12190 );
nand \U$14009 ( \14198 , \14002 , \14197 );
nand \U$14010 ( \14199 , \13511 , \8042 );
nand \U$14011 ( \14200 , \8360 , \8683 );
nor \U$14012 ( \14201 , \14199 , \14200 );
nand \U$14013 ( \14202 , \9008 , \9335 );
nand \U$14014 ( \14203 , \9660 , \9986 );
nor \U$14015 ( \14204 , \14202 , \14203 );
nand \U$14016 ( \14205 , \14201 , \14204 );
nand \U$14017 ( \14206 , \10311 , \10639 );
nand \U$14018 ( \14207 , \10964 , \11290 );
nor \U$14019 ( \14208 , \14206 , \14207 );
nand \U$14020 ( \14209 , \11615 , \11942 );
nand \U$14021 ( \14210 , \12106 , \12175 );
nor \U$14022 ( \14211 , \14209 , \14210 );
nand \U$14023 ( \14212 , \14208 , \14211 );
nor \U$14024 ( \14213 , \14205 , \14212 );
nand \U$14025 ( \14214 , \13766 , \12519 );
nand \U$14026 ( \14215 , \12686 , \12874 );
nor \U$14027 ( \14216 , \14214 , \14215 );
nand \U$14028 ( \14217 , \13081 , \13310 );
nand \U$14029 ( \14218 , \13429 , \13489 );
nor \U$14030 ( \14219 , \14217 , \14218 );
nand \U$14031 ( \14220 , \14216 , \14219 );
nand \U$14032 ( \14221 , \13813 , \13614 );
nand \U$14033 ( \14222 , \13701 , \13747 );
nor \U$14034 ( \14223 , \14221 , \14222 );
and \U$14035 ( \14224 , \13799 , \13829 );
nor \U$14036 ( \14225 , \14224 , \13835 );
not \U$14037 ( \14226 , \14225 );
and \U$14038 ( \14227 , \14223 , \14226 );
and \U$14039 ( \14228 , \13614 , \13840 );
nor \U$14040 ( \14229 , \14228 , \13847 );
or \U$14041 ( \14230 , \14222 , \14229 );
and \U$14042 ( \14231 , \13747 , \13852 );
nor \U$14043 ( \14232 , \14231 , \13858 );
nand \U$14044 ( \14233 , \14230 , \14232 );
nor \U$14045 ( \14234 , \14227 , \14233 );
or \U$14046 ( \14235 , \14220 , \14234 );
and \U$14047 ( \14236 , \12519 , \13863 );
nor \U$14048 ( \14237 , \14236 , \13871 );
or \U$14049 ( \14238 , \14215 , \14237 );
and \U$14050 ( \14239 , \12874 , \13876 );
nor \U$14051 ( \14240 , \14239 , \13882 );
nand \U$14052 ( \14241 , \14238 , \14240 );
and \U$14053 ( \14242 , \14219 , \14241 );
and \U$14054 ( \14243 , \13310 , \13887 );
nor \U$14055 ( \14244 , \14243 , \13894 );
or \U$14056 ( \14245 , \14218 , \14244 );
and \U$14057 ( \14246 , \13489 , \13899 );
nor \U$14058 ( \14247 , \14246 , \13905 );
nand \U$14059 ( \14248 , \14245 , \14247 );
nor \U$14060 ( \14249 , \14242 , \14248 );
nand \U$14061 ( \14250 , \14235 , \14249 );
and \U$14062 ( \14251 , \14213 , \14250 );
and \U$14063 ( \14252 , \8042 , \13910 );
nor \U$14064 ( \14253 , \14252 , \13919 );
or \U$14065 ( \14254 , \14200 , \14253 );
and \U$14066 ( \14255 , \8683 , \13924 );
nor \U$14067 ( \14256 , \14255 , \13930 );
nand \U$14068 ( \14257 , \14254 , \14256 );
and \U$14069 ( \14258 , \14204 , \14257 );
and \U$14070 ( \14259 , \9335 , \13935 );
nor \U$14071 ( \14260 , \14259 , \13942 );
or \U$14072 ( \14261 , \14203 , \14260 );
and \U$14073 ( \14262 , \9986 , \13947 );
nor \U$14074 ( \14263 , \14262 , \13953 );
nand \U$14075 ( \14264 , \14261 , \14263 );
nor \U$14076 ( \14265 , \14258 , \14264 );
or \U$14077 ( \14266 , \14212 , \14265 );
and \U$14078 ( \14267 , \10639 , \13958 );
nor \U$14079 ( \14268 , \14267 , \13966 );
or \U$14080 ( \14269 , \14207 , \14268 );
and \U$14081 ( \14270 , \11290 , \13971 );
nor \U$14082 ( \14271 , \14270 , \13977 );
nand \U$14083 ( \14272 , \14269 , \14271 );
and \U$14084 ( \14273 , \14211 , \14272 );
and \U$14085 ( \14274 , \11942 , \13982 );
nor \U$14086 ( \14275 , \14274 , \13989 );
or \U$14087 ( \14276 , \14210 , \14275 );
and \U$14088 ( \14277 , \12175 , \13994 );
nor \U$14089 ( \14278 , \14277 , \14000 );
nand \U$14090 ( \14279 , \14276 , \14278 );
nor \U$14091 ( \14280 , \14273 , \14279 );
nand \U$14092 ( \14281 , \14266 , \14280 );
nor \U$14093 ( \14282 , \14251 , \14281 );
not \U$14094 ( \14283 , \14282 );
xnor \U$14095 ( \14284 , \14198 , \14283 );
buf \U$14096 ( \14285 , \14284 );
buf \U$14097 ( \14286 , \14285 );
not \U$14098 ( \14287 , \12174 );
nand \U$14099 ( \14288 , \13999 , \14287 );
nand \U$14100 ( \14289 , \14059 , \14017 );
nand \U$14101 ( \14290 , \14018 , \14020 );
nor \U$14102 ( \14291 , \14289 , \14290 );
nand \U$14103 ( \14292 , \14021 , \14024 );
nand \U$14104 ( \14293 , \14025 , \14027 );
nor \U$14105 ( \14294 , \14292 , \14293 );
nand \U$14106 ( \14295 , \14291 , \14294 );
nand \U$14107 ( \14296 , \14028 , \14032 );
nand \U$14108 ( \14297 , \14033 , \14035 );
nor \U$14109 ( \14298 , \14296 , \14297 );
nand \U$14110 ( \14299 , \14036 , \14039 );
nand \U$14111 ( \14300 , \14040 , \14042 );
nor \U$14112 ( \14301 , \14299 , \14300 );
nand \U$14113 ( \14302 , \14298 , \14301 );
nor \U$14114 ( \14303 , \14295 , \14302 );
nand \U$14115 ( \14304 , \14067 , \14048 );
nand \U$14116 ( \14305 , \14049 , \14051 );
nor \U$14117 ( \14306 , \14304 , \14305 );
nand \U$14118 ( \14307 , \14052 , \14055 );
nand \U$14119 ( \14308 , \14056 , \14058 );
nor \U$14120 ( \14309 , \14307 , \14308 );
nand \U$14121 ( \14310 , \14306 , \14309 );
nand \U$14122 ( \14311 , \14071 , \14063 );
nand \U$14123 ( \14312 , \14064 , \14066 );
nor \U$14124 ( \14313 , \14311 , \14312 );
not \U$14125 ( \14314 , \13826 );
and \U$14126 ( \14315 , \14070 , \14314 );
nor \U$14127 ( \14316 , \14315 , \14075 );
not \U$14128 ( \14317 , \14316 );
and \U$14129 ( \14318 , \14313 , \14317 );
and \U$14130 ( \14319 , \14063 , \14078 );
nor \U$14131 ( \14320 , \14319 , \14083 );
or \U$14132 ( \14321 , \14312 , \14320 );
and \U$14133 ( \14322 , \14066 , \14086 );
nor \U$14134 ( \14323 , \14322 , \14090 );
nand \U$14135 ( \14324 , \14321 , \14323 );
nor \U$14136 ( \14325 , \14318 , \14324 );
or \U$14137 ( \14326 , \14310 , \14325 );
and \U$14138 ( \14327 , \14048 , \14093 );
nor \U$14139 ( \14328 , \14327 , \14099 );
or \U$14140 ( \14329 , \14305 , \14328 );
and \U$14141 ( \14330 , \14051 , \14102 );
nor \U$14142 ( \14331 , \14330 , \14106 );
nand \U$14143 ( \14332 , \14329 , \14331 );
and \U$14144 ( \14333 , \14309 , \14332 );
and \U$14145 ( \14334 , \14055 , \14109 );
nor \U$14146 ( \14335 , \14334 , \14114 );
or \U$14147 ( \14336 , \14308 , \14335 );
and \U$14148 ( \14337 , \14058 , \14117 );
nor \U$14149 ( \14338 , \14337 , \14121 );
nand \U$14150 ( \14339 , \14336 , \14338 );
nor \U$14151 ( \14340 , \14333 , \14339 );
nand \U$14152 ( \14341 , \14326 , \14340 );
and \U$14153 ( \14342 , \14303 , \14341 );
and \U$14154 ( \14343 , \14017 , \14124 );
nor \U$14155 ( \14344 , \14343 , \14131 );
or \U$14156 ( \14345 , \14290 , \14344 );
and \U$14157 ( \14346 , \14020 , \14134 );
nor \U$14158 ( \14347 , \14346 , \14138 );
nand \U$14159 ( \14348 , \14345 , \14347 );
and \U$14160 ( \14349 , \14294 , \14348 );
and \U$14161 ( \14350 , \14024 , \14141 );
nor \U$14162 ( \14351 , \14350 , \14146 );
or \U$14163 ( \14352 , \14293 , \14351 );
and \U$14164 ( \14353 , \14027 , \14149 );
nor \U$14165 ( \14354 , \14353 , \14153 );
nand \U$14166 ( \14355 , \14352 , \14354 );
nor \U$14167 ( \14356 , \14349 , \14355 );
or \U$14168 ( \14357 , \14302 , \14356 );
and \U$14169 ( \14358 , \14032 , \14156 );
nor \U$14170 ( \14359 , \14358 , \14162 );
or \U$14171 ( \14360 , \14297 , \14359 );
and \U$14172 ( \14361 , \14035 , \14165 );
nor \U$14173 ( \14362 , \14361 , \14169 );
nand \U$14174 ( \14363 , \14360 , \14362 );
and \U$14175 ( \14364 , \14301 , \14363 );
and \U$14176 ( \14365 , \14039 , \14172 );
nor \U$14177 ( \14366 , \14365 , \14177 );
or \U$14178 ( \14367 , \14300 , \14366 );
and \U$14179 ( \14368 , \14042 , \14180 );
nor \U$14180 ( \14369 , \14368 , \14184 );
nand \U$14181 ( \14370 , \14367 , \14369 );
nor \U$14182 ( \14371 , \14364 , \14370 );
nand \U$14183 ( \14372 , \14357 , \14371 );
nor \U$14184 ( \14373 , \14342 , \14372 );
not \U$14185 ( \14374 , \14373 );
xnor \U$14186 ( \14375 , \14288 , \14374 );
buf \U$14187 ( \14376 , \14375 );
buf \U$14188 ( \14377 , \14376 );
not \U$14189 ( \14378 , \12149 );
nand \U$14190 ( \14379 , \13997 , \14378 );
nor \U$14191 ( \14380 , \13512 , \8361 );
nor \U$14192 ( \14381 , \9009 , \9661 );
nand \U$14193 ( \14382 , \14380 , \14381 );
nor \U$14194 ( \14383 , \10312 , \10965 );
nor \U$14195 ( \14384 , \11616 , \12107 );
nand \U$14196 ( \14385 , \14383 , \14384 );
nor \U$14197 ( \14386 , \14382 , \14385 );
nor \U$14198 ( \14387 , \13767 , \12687 );
nor \U$14199 ( \14388 , \13082 , \13430 );
nand \U$14200 ( \14389 , \14387 , \14388 );
nor \U$14201 ( \14390 , \13814 , \13702 );
and \U$14202 ( \14391 , \14390 , \13829 );
or \U$14203 ( \14392 , \13702 , \13841 );
nand \U$14204 ( \14393 , \14392 , \13853 );
nor \U$14205 ( \14394 , \14391 , \14393 );
or \U$14206 ( \14395 , \14389 , \14394 );
or \U$14207 ( \14396 , \12687 , \13864 );
nand \U$14208 ( \14397 , \14396 , \13877 );
and \U$14209 ( \14398 , \14388 , \14397 );
or \U$14210 ( \14399 , \13430 , \13888 );
nand \U$14211 ( \14400 , \14399 , \13900 );
nor \U$14212 ( \14401 , \14398 , \14400 );
nand \U$14213 ( \14402 , \14395 , \14401 );
and \U$14214 ( \14403 , \14386 , \14402 );
or \U$14215 ( \14404 , \8361 , \13911 );
nand \U$14216 ( \14405 , \14404 , \13925 );
and \U$14217 ( \14406 , \14381 , \14405 );
or \U$14218 ( \14407 , \9661 , \13936 );
nand \U$14219 ( \14408 , \14407 , \13948 );
nor \U$14220 ( \14409 , \14406 , \14408 );
or \U$14221 ( \14410 , \14385 , \14409 );
or \U$14222 ( \14411 , \10965 , \13959 );
nand \U$14223 ( \14412 , \14411 , \13972 );
and \U$14224 ( \14413 , \14384 , \14412 );
or \U$14225 ( \14414 , \12107 , \13983 );
nand \U$14226 ( \14415 , \14414 , \13995 );
nor \U$14227 ( \14416 , \14413 , \14415 );
nand \U$14228 ( \14417 , \14410 , \14416 );
nor \U$14229 ( \14418 , \14403 , \14417 );
not \U$14230 ( \14419 , \14418 );
xnor \U$14231 ( \14420 , \14379 , \14419 );
buf \U$14232 ( \14421 , \14420 );
buf \U$14233 ( \14422 , \14421 );
not \U$14234 ( \14423 , \12105 );
nand \U$14235 ( \14424 , \13993 , \14423 );
nor \U$14236 ( \14425 , \14060 , \14019 );
nor \U$14237 ( \14426 , \14022 , \14026 );
nand \U$14238 ( \14427 , \14425 , \14426 );
nor \U$14239 ( \14428 , \14029 , \14034 );
nor \U$14240 ( \14429 , \14037 , \14041 );
nand \U$14241 ( \14430 , \14428 , \14429 );
nor \U$14242 ( \14431 , \14427 , \14430 );
nor \U$14243 ( \14432 , \14068 , \14050 );
nor \U$14244 ( \14433 , \14053 , \14057 );
nand \U$14245 ( \14434 , \14432 , \14433 );
nor \U$14246 ( \14435 , \14072 , \14065 );
and \U$14247 ( \14436 , \14435 , \14314 );
or \U$14248 ( \14437 , \14065 , \14079 );
nand \U$14249 ( \14438 , \14437 , \14087 );
nor \U$14250 ( \14439 , \14436 , \14438 );
or \U$14251 ( \14440 , \14434 , \14439 );
or \U$14252 ( \14441 , \14050 , \14094 );
nand \U$14253 ( \14442 , \14441 , \14103 );
and \U$14254 ( \14443 , \14433 , \14442 );
or \U$14255 ( \14444 , \14057 , \14110 );
nand \U$14256 ( \14445 , \14444 , \14118 );
nor \U$14257 ( \14446 , \14443 , \14445 );
nand \U$14258 ( \14447 , \14440 , \14446 );
and \U$14259 ( \14448 , \14431 , \14447 );
or \U$14260 ( \14449 , \14019 , \14125 );
nand \U$14261 ( \14450 , \14449 , \14135 );
and \U$14262 ( \14451 , \14426 , \14450 );
or \U$14263 ( \14452 , \14026 , \14142 );
nand \U$14264 ( \14453 , \14452 , \14150 );
nor \U$14265 ( \14454 , \14451 , \14453 );
or \U$14266 ( \14455 , \14430 , \14454 );
or \U$14267 ( \14456 , \14034 , \14157 );
nand \U$14268 ( \14457 , \14456 , \14166 );
and \U$14269 ( \14458 , \14429 , \14457 );
or \U$14270 ( \14459 , \14041 , \14173 );
nand \U$14271 ( \14460 , \14459 , \14181 );
nor \U$14272 ( \14461 , \14458 , \14460 );
nand \U$14273 ( \14462 , \14455 , \14461 );
nor \U$14274 ( \14463 , \14448 , \14462 );
not \U$14275 ( \14464 , \14463 );
xnor \U$14276 ( \14465 , \14424 , \14464 );
buf \U$14277 ( \14466 , \14465 );
buf \U$14278 ( \14467 , \14466 );
not \U$14279 ( \14468 , \12040 );
nand \U$14280 ( \14469 , \13991 , \14468 );
nor \U$14281 ( \14470 , \14218 , \14199 );
nor \U$14282 ( \14471 , \14200 , \14202 );
nand \U$14283 ( \14472 , \14470 , \14471 );
nor \U$14284 ( \14473 , \14203 , \14206 );
nor \U$14285 ( \14474 , \14207 , \14209 );
nand \U$14286 ( \14475 , \14473 , \14474 );
nor \U$14287 ( \14476 , \14472 , \14475 );
nor \U$14288 ( \14477 , \14222 , \14214 );
nor \U$14289 ( \14478 , \14215 , \14217 );
nand \U$14290 ( \14479 , \14477 , \14478 );
or \U$14291 ( \14480 , \14221 , \14225 );
nand \U$14292 ( \14481 , \14480 , \14229 );
not \U$14293 ( \14482 , \14481 );
or \U$14294 ( \14483 , \14479 , \14482 );
or \U$14295 ( \14484 , \14214 , \14232 );
nand \U$14296 ( \14485 , \14484 , \14237 );
and \U$14297 ( \14486 , \14478 , \14485 );
or \U$14298 ( \14487 , \14217 , \14240 );
nand \U$14299 ( \14488 , \14487 , \14244 );
nor \U$14300 ( \14489 , \14486 , \14488 );
nand \U$14301 ( \14490 , \14483 , \14489 );
and \U$14302 ( \14491 , \14476 , \14490 );
or \U$14303 ( \14492 , \14199 , \14247 );
nand \U$14304 ( \14493 , \14492 , \14253 );
and \U$14305 ( \14494 , \14471 , \14493 );
or \U$14306 ( \14495 , \14202 , \14256 );
nand \U$14307 ( \14496 , \14495 , \14260 );
nor \U$14308 ( \14497 , \14494 , \14496 );
or \U$14309 ( \14498 , \14475 , \14497 );
or \U$14310 ( \14499 , \14206 , \14263 );
nand \U$14311 ( \14500 , \14499 , \14268 );
and \U$14312 ( \14501 , \14474 , \14500 );
or \U$14313 ( \14502 , \14209 , \14271 );
nand \U$14314 ( \14503 , \14502 , \14275 );
nor \U$14315 ( \14504 , \14501 , \14503 );
nand \U$14316 ( \14505 , \14498 , \14504 );
nor \U$14317 ( \14506 , \14491 , \14505 );
not \U$14318 ( \14507 , \14506 );
xnor \U$14319 ( \14508 , \14469 , \14507 );
buf \U$14320 ( \14509 , \14508 );
buf \U$14321 ( \14510 , \14509 );
not \U$14322 ( \14511 , \11941 );
nand \U$14323 ( \14512 , \13988 , \14511 );
nor \U$14324 ( \14513 , \14308 , \14289 );
nor \U$14325 ( \14514 , \14290 , \14292 );
nand \U$14326 ( \14515 , \14513 , \14514 );
nor \U$14327 ( \14516 , \14293 , \14296 );
nor \U$14328 ( \14517 , \14297 , \14299 );
nand \U$14329 ( \14518 , \14516 , \14517 );
nor \U$14330 ( \14519 , \14515 , \14518 );
nor \U$14331 ( \14520 , \14312 , \14304 );
nor \U$14332 ( \14521 , \14305 , \14307 );
nand \U$14333 ( \14522 , \14520 , \14521 );
or \U$14334 ( \14523 , \14311 , \14316 );
nand \U$14335 ( \14524 , \14523 , \14320 );
not \U$14336 ( \14525 , \14524 );
or \U$14337 ( \14526 , \14522 , \14525 );
or \U$14338 ( \14527 , \14304 , \14323 );
nand \U$14339 ( \14528 , \14527 , \14328 );
and \U$14340 ( \14529 , \14521 , \14528 );
or \U$14341 ( \14530 , \14307 , \14331 );
nand \U$14342 ( \14531 , \14530 , \14335 );
nor \U$14343 ( \14532 , \14529 , \14531 );
nand \U$14344 ( \14533 , \14526 , \14532 );
and \U$14345 ( \14534 , \14519 , \14533 );
or \U$14346 ( \14535 , \14289 , \14338 );
nand \U$14347 ( \14536 , \14535 , \14344 );
and \U$14348 ( \14537 , \14514 , \14536 );
or \U$14349 ( \14538 , \14292 , \14347 );
nand \U$14350 ( \14539 , \14538 , \14351 );
nor \U$14351 ( \14540 , \14537 , \14539 );
or \U$14352 ( \14541 , \14518 , \14540 );
or \U$14353 ( \14542 , \14296 , \14354 );
nand \U$14354 ( \14543 , \14542 , \14359 );
and \U$14355 ( \14544 , \14517 , \14543 );
or \U$14356 ( \14545 , \14299 , \14362 );
nand \U$14357 ( \14546 , \14545 , \14366 );
nor \U$14358 ( \14547 , \14544 , \14546 );
nand \U$14359 ( \14548 , \14541 , \14547 );
nor \U$14360 ( \14549 , \14534 , \14548 );
not \U$14361 ( \14550 , \14549 );
xnor \U$14362 ( \14551 , \14512 , \14550 );
buf \U$14363 ( \14552 , \14551 );
buf \U$14364 ( \14553 , \14552 );
not \U$14365 ( \14554 , \11780 );
nand \U$14366 ( \14555 , \13986 , \14554 );
nand \U$14367 ( \14556 , \13513 , \9010 );
nand \U$14368 ( \14557 , \10313 , \11617 );
nor \U$14369 ( \14558 , \14556 , \14557 );
nand \U$14370 ( \14559 , \13768 , \13083 );
not \U$14371 ( \14560 , \13842 );
or \U$14372 ( \14561 , \14559 , \14560 );
and \U$14373 ( \14562 , \13083 , \13865 );
nor \U$14374 ( \14563 , \14562 , \13889 );
nand \U$14375 ( \14564 , \14561 , \14563 );
and \U$14376 ( \14565 , \14558 , \14564 );
and \U$14377 ( \14566 , \9010 , \13912 );
nor \U$14378 ( \14567 , \14566 , \13937 );
or \U$14379 ( \14568 , \14557 , \14567 );
and \U$14380 ( \14569 , \11617 , \13960 );
nor \U$14381 ( \14570 , \14569 , \13984 );
nand \U$14382 ( \14571 , \14568 , \14570 );
nor \U$14383 ( \14572 , \14565 , \14571 );
not \U$14384 ( \14573 , \14572 );
xnor \U$14385 ( \14574 , \14555 , \14573 );
buf \U$14386 ( \14575 , \14574 );
buf \U$14387 ( \14576 , \14575 );
not \U$14388 ( \14577 , \11614 );
nand \U$14389 ( \14578 , \13981 , \14577 );
nand \U$14390 ( \14579 , \14061 , \14023 );
nand \U$14391 ( \14580 , \14030 , \14038 );
nor \U$14392 ( \14581 , \14579 , \14580 );
nand \U$14393 ( \14582 , \14069 , \14054 );
not \U$14394 ( \14583 , \14080 );
or \U$14395 ( \14584 , \14582 , \14583 );
and \U$14396 ( \14585 , \14054 , \14095 );
nor \U$14397 ( \14586 , \14585 , \14111 );
nand \U$14398 ( \14587 , \14584 , \14586 );
and \U$14399 ( \14588 , \14581 , \14587 );
and \U$14400 ( \14589 , \14023 , \14126 );
nor \U$14401 ( \14590 , \14589 , \14143 );
or \U$14402 ( \14591 , \14580 , \14590 );
and \U$14403 ( \14592 , \14038 , \14158 );
nor \U$14404 ( \14593 , \14592 , \14174 );
nand \U$14405 ( \14594 , \14591 , \14593 );
nor \U$14406 ( \14595 , \14588 , \14594 );
not \U$14407 ( \14596 , \14595 );
xnor \U$14408 ( \14597 , \14578 , \14596 );
buf \U$14409 ( \14598 , \14597 );
buf \U$14410 ( \14599 , \14598 );
not \U$14411 ( \14600 , \11453 );
nand \U$14412 ( \14601 , \13979 , \14600 );
nand \U$14413 ( \14602 , \14219 , \14201 );
nand \U$14414 ( \14603 , \14204 , \14208 );
nor \U$14415 ( \14604 , \14602 , \14603 );
nand \U$14416 ( \14605 , \14223 , \14216 );
or \U$14417 ( \14606 , \14605 , \14225 );
and \U$14418 ( \14607 , \14216 , \14233 );
nor \U$14419 ( \14608 , \14607 , \14241 );
nand \U$14420 ( \14609 , \14606 , \14608 );
and \U$14421 ( \14610 , \14604 , \14609 );
and \U$14422 ( \14611 , \14201 , \14248 );
nor \U$14423 ( \14612 , \14611 , \14257 );
or \U$14424 ( \14613 , \14603 , \14612 );
and \U$14425 ( \14614 , \14208 , \14264 );
nor \U$14426 ( \14615 , \14614 , \14272 );
nand \U$14427 ( \14616 , \14613 , \14615 );
nor \U$14428 ( \14617 , \14610 , \14616 );
not \U$14429 ( \14618 , \14617 );
xnor \U$14430 ( \14619 , \14601 , \14618 );
buf \U$14431 ( \14620 , \14619 );
buf \U$14432 ( \14621 , \14620 );
not \U$14433 ( \14622 , \11289 );
nand \U$14434 ( \14623 , \13976 , \14622 );
nand \U$14435 ( \14624 , \14309 , \14291 );
nand \U$14436 ( \14625 , \14294 , \14298 );
nor \U$14437 ( \14626 , \14624 , \14625 );
nand \U$14438 ( \14627 , \14313 , \14306 );
or \U$14439 ( \14628 , \14627 , \14316 );
and \U$14440 ( \14629 , \14306 , \14324 );
nor \U$14441 ( \14630 , \14629 , \14332 );
nand \U$14442 ( \14631 , \14628 , \14630 );
and \U$14443 ( \14632 , \14626 , \14631 );
and \U$14444 ( \14633 , \14291 , \14339 );
nor \U$14445 ( \14634 , \14633 , \14348 );
or \U$14446 ( \14635 , \14625 , \14634 );
and \U$14447 ( \14636 , \14298 , \14355 );
nor \U$14448 ( \14637 , \14636 , \14363 );
nand \U$14449 ( \14638 , \14635 , \14637 );
nor \U$14450 ( \14639 , \14632 , \14638 );
not \U$14451 ( \14640 , \14639 );
xnor \U$14452 ( \14641 , \14623 , \14640 );
buf \U$14453 ( \14642 , \14641 );
buf \U$14454 ( \14643 , \14642 );
not \U$14455 ( \14644 , \11128 );
nand \U$14456 ( \14645 , \13974 , \14644 );
nand \U$14457 ( \14646 , \14388 , \14380 );
nand \U$14458 ( \14647 , \14381 , \14383 );
nor \U$14459 ( \14648 , \14646 , \14647 );
nand \U$14460 ( \14649 , \14390 , \14387 );
or \U$14461 ( \14650 , \14649 , \13830 );
and \U$14462 ( \14651 , \14387 , \14393 );
nor \U$14463 ( \14652 , \14651 , \14397 );
nand \U$14464 ( \14653 , \14650 , \14652 );
and \U$14465 ( \14654 , \14648 , \14653 );
and \U$14466 ( \14655 , \14380 , \14400 );
nor \U$14467 ( \14656 , \14655 , \14405 );
or \U$14468 ( \14657 , \14647 , \14656 );
and \U$14469 ( \14658 , \14383 , \14408 );
nor \U$14470 ( \14659 , \14658 , \14412 );
nand \U$14471 ( \14660 , \14657 , \14659 );
nor \U$14472 ( \14661 , \14654 , \14660 );
not \U$14473 ( \14662 , \14661 );
xnor \U$14474 ( \14663 , \14645 , \14662 );
buf \U$14475 ( \14664 , \14663 );
buf \U$14476 ( \14665 , \14664 );
not \U$14477 ( \14666 , \10963 );
nand \U$14478 ( \14667 , \13970 , \14666 );
nand \U$14479 ( \14668 , \14433 , \14425 );
nand \U$14480 ( \14669 , \14426 , \14428 );
nor \U$14481 ( \14670 , \14668 , \14669 );
nand \U$14482 ( \14671 , \14435 , \14432 );
or \U$14483 ( \14672 , \14671 , \13826 );
and \U$14484 ( \14673 , \14432 , \14438 );
nor \U$14485 ( \14674 , \14673 , \14442 );
nand \U$14486 ( \14675 , \14672 , \14674 );
and \U$14487 ( \14676 , \14670 , \14675 );
and \U$14488 ( \14677 , \14425 , \14445 );
nor \U$14489 ( \14678 , \14677 , \14450 );
or \U$14490 ( \14679 , \14669 , \14678 );
and \U$14491 ( \14680 , \14428 , \14453 );
nor \U$14492 ( \14681 , \14680 , \14457 );
nand \U$14493 ( \14682 , \14679 , \14681 );
nor \U$14494 ( \14683 , \14676 , \14682 );
not \U$14495 ( \14684 , \14683 );
xnor \U$14496 ( \14685 , \14667 , \14684 );
buf \U$14497 ( \14686 , \14685 );
buf \U$14498 ( \14687 , \14686 );
not \U$14499 ( \14688 , \10802 );
nand \U$14500 ( \14689 , \13968 , \14688 );
nand \U$14501 ( \14690 , \14478 , \14470 );
nand \U$14502 ( \14691 , \14471 , \14473 );
nor \U$14503 ( \14692 , \14690 , \14691 );
and \U$14504 ( \14693 , \14477 , \14481 );
nor \U$14505 ( \14694 , \14693 , \14485 );
not \U$14506 ( \14695 , \14694 );
and \U$14507 ( \14696 , \14692 , \14695 );
and \U$14508 ( \14697 , \14470 , \14488 );
nor \U$14509 ( \14698 , \14697 , \14493 );
or \U$14510 ( \14699 , \14691 , \14698 );
and \U$14511 ( \14700 , \14473 , \14496 );
nor \U$14512 ( \14701 , \14700 , \14500 );
nand \U$14513 ( \14702 , \14699 , \14701 );
nor \U$14514 ( \14703 , \14696 , \14702 );
not \U$14515 ( \14704 , \14703 );
xnor \U$14516 ( \14705 , \14689 , \14704 );
buf \U$14517 ( \14706 , \14705 );
buf \U$14518 ( \14707 , \14706 );
not \U$14519 ( \14708 , \10638 );
nand \U$14520 ( \14709 , \13965 , \14708 );
nand \U$14521 ( \14710 , \14521 , \14513 );
nand \U$14522 ( \14711 , \14514 , \14516 );
nor \U$14523 ( \14712 , \14710 , \14711 );
and \U$14524 ( \14713 , \14520 , \14524 );
nor \U$14525 ( \14714 , \14713 , \14528 );
not \U$14526 ( \14715 , \14714 );
and \U$14527 ( \14716 , \14712 , \14715 );
and \U$14528 ( \14717 , \14513 , \14531 );
nor \U$14529 ( \14718 , \14717 , \14536 );
or \U$14530 ( \14719 , \14711 , \14718 );
and \U$14531 ( \14720 , \14516 , \14539 );
nor \U$14532 ( \14721 , \14720 , \14543 );
nand \U$14533 ( \14722 , \14719 , \14721 );
nor \U$14534 ( \14723 , \14716 , \14722 );
not \U$14535 ( \14724 , \14723 );
xnor \U$14536 ( \14725 , \14709 , \14724 );
buf \U$14537 ( \14726 , \14725 );
buf \U$14538 ( \14727 , \14726 );
not \U$14539 ( \14728 , \10477 );
nand \U$14540 ( \14729 , \13963 , \14728 );
nor \U$14541 ( \14730 , \13514 , \10314 );
not \U$14542 ( \14731 , \13866 );
and \U$14543 ( \14732 , \14730 , \14731 );
or \U$14544 ( \14733 , \10314 , \13913 );
nand \U$14545 ( \14734 , \14733 , \13961 );
nor \U$14546 ( \14735 , \14732 , \14734 );
not \U$14547 ( \14736 , \14735 );
xnor \U$14548 ( \14737 , \14729 , \14736 );
buf \U$14549 ( \14738 , \14737 );
buf \U$14550 ( \14739 , \14738 );
not \U$14551 ( \14740 , \10310 );
nand \U$14552 ( \14741 , \13957 , \14740 );
nor \U$14553 ( \14742 , \14062 , \14031 );
not \U$14554 ( \14743 , \14096 );
and \U$14555 ( \14744 , \14742 , \14743 );
or \U$14556 ( \14745 , \14031 , \14127 );
nand \U$14557 ( \14746 , \14745 , \14159 );
nor \U$14558 ( \14747 , \14744 , \14746 );
not \U$14559 ( \14748 , \14747 );
xnor \U$14560 ( \14749 , \14741 , \14748 );
buf \U$14561 ( \14750 , \14749 );
buf \U$14562 ( \14751 , \14750 );
not \U$14563 ( \14752 , \10149 );
nand \U$14564 ( \14753 , \13955 , \14752 );
nor \U$14565 ( \14754 , \14220 , \14205 );
not \U$14566 ( \14755 , \14234 );
and \U$14567 ( \14756 , \14754 , \14755 );
or \U$14568 ( \14757 , \14205 , \14249 );
nand \U$14569 ( \14758 , \14757 , \14265 );
nor \U$14570 ( \14759 , \14756 , \14758 );
not \U$14571 ( \14760 , \14759 );
xnor \U$14572 ( \14761 , \14753 , \14760 );
buf \U$14573 ( \14762 , \14761 );
buf \U$14574 ( \14763 , \14762 );
not \U$14575 ( \14764 , \9985 );
nand \U$14576 ( \14765 , \13952 , \14764 );
nor \U$14577 ( \14766 , \14310 , \14295 );
not \U$14578 ( \14767 , \14325 );
and \U$14579 ( \14768 , \14766 , \14767 );
or \U$14580 ( \14769 , \14295 , \14340 );
nand \U$14581 ( \14770 , \14769 , \14356 );
nor \U$14582 ( \14771 , \14768 , \14770 );
not \U$14583 ( \14772 , \14771 );
xnor \U$14584 ( \14773 , \14765 , \14772 );
buf \U$14585 ( \14774 , \14773 );
buf \U$14586 ( \14775 , \14774 );
not \U$14587 ( \14776 , \9824 );
nand \U$14588 ( \14777 , \13950 , \14776 );
nor \U$14589 ( \14778 , \14389 , \14382 );
not \U$14590 ( \14779 , \14394 );
and \U$14591 ( \14780 , \14778 , \14779 );
or \U$14592 ( \14781 , \14382 , \14401 );
nand \U$14593 ( \14782 , \14781 , \14409 );
nor \U$14594 ( \14783 , \14780 , \14782 );
not \U$14595 ( \14784 , \14783 );
xnor \U$14596 ( \14785 , \14777 , \14784 );
buf \U$14597 ( \14786 , \14785 );
buf \U$14598 ( \14787 , \14786 );
not \U$14599 ( \14788 , \9659 );
nand \U$14600 ( \14789 , \13946 , \14788 );
nor \U$14601 ( \14790 , \14434 , \14427 );
not \U$14602 ( \14791 , \14439 );
and \U$14603 ( \14792 , \14790 , \14791 );
or \U$14604 ( \14793 , \14427 , \14446 );
nand \U$14605 ( \14794 , \14793 , \14454 );
nor \U$14606 ( \14795 , \14792 , \14794 );
not \U$14607 ( \14796 , \14795 );
xnor \U$14608 ( \14797 , \14789 , \14796 );
buf \U$14609 ( \14798 , \14797 );
buf \U$14610 ( \14799 , \14798 );
not \U$14611 ( \14800 , \9498 );
nand \U$14612 ( \14801 , \13944 , \14800 );
nor \U$14613 ( \14802 , \14479 , \14472 );
and \U$14614 ( \14803 , \14802 , \14481 );
or \U$14615 ( \14804 , \14472 , \14489 );
nand \U$14616 ( \14805 , \14804 , \14497 );
nor \U$14617 ( \14806 , \14803 , \14805 );
not \U$14618 ( \14807 , \14806 );
xnor \U$14619 ( \14808 , \14801 , \14807 );
buf \U$14620 ( \14809 , \14808 );
buf \U$14621 ( \14810 , \14809 );
not \U$14622 ( \14811 , \9334 );
nand \U$14623 ( \14812 , \13941 , \14811 );
nor \U$14624 ( \14813 , \14522 , \14515 );
and \U$14625 ( \14814 , \14813 , \14524 );
or \U$14626 ( \14815 , \14515 , \14532 );
nand \U$14627 ( \14816 , \14815 , \14540 );
nor \U$14628 ( \14817 , \14814 , \14816 );
not \U$14629 ( \14818 , \14817 );
xnor \U$14630 ( \14819 , \14812 , \14818 );
buf \U$14631 ( \14820 , \14819 );
buf \U$14632 ( \14821 , \14820 );
not \U$14633 ( \14822 , \9173 );
nand \U$14634 ( \14823 , \13939 , \14822 );
nor \U$14635 ( \14824 , \14559 , \14556 );
and \U$14636 ( \14825 , \14824 , \13842 );
or \U$14637 ( \14826 , \14556 , \14563 );
nand \U$14638 ( \14827 , \14826 , \14567 );
nor \U$14639 ( \14828 , \14825 , \14827 );
not \U$14640 ( \14829 , \14828 );
xnor \U$14641 ( \14830 , \14823 , \14829 );
buf \U$14642 ( \14831 , \14830 );
buf \U$14643 ( \14832 , \14831 );
not \U$14644 ( \14833 , \9007 );
nand \U$14645 ( \14834 , \13934 , \14833 );
nor \U$14646 ( \14835 , \14582 , \14579 );
and \U$14647 ( \14836 , \14835 , \14080 );
or \U$14648 ( \14837 , \14579 , \14586 );
nand \U$14649 ( \14838 , \14837 , \14590 );
nor \U$14650 ( \14839 , \14836 , \14838 );
not \U$14651 ( \14840 , \14839 );
xnor \U$14652 ( \14841 , \14834 , \14840 );
buf \U$14653 ( \14842 , \14841 );
buf \U$14654 ( \14843 , \14842 );
not \U$14655 ( \14844 , \8846 );
nand \U$14656 ( \14845 , \13932 , \14844 );
nor \U$14657 ( \14846 , \14605 , \14602 );
and \U$14658 ( \14847 , \14846 , \14226 );
or \U$14659 ( \14848 , \14602 , \14608 );
nand \U$14660 ( \14849 , \14848 , \14612 );
nor \U$14661 ( \14850 , \14847 , \14849 );
not \U$14662 ( \14851 , \14850 );
xnor \U$14663 ( \14852 , \14845 , \14851 );
buf \U$14664 ( \14853 , \14852 );
buf \U$14665 ( \14854 , \14853 );
not \U$14666 ( \14855 , \8682 );
nand \U$14667 ( \14856 , \13929 , \14855 );
nor \U$14668 ( \14857 , \14627 , \14624 );
and \U$14669 ( \14858 , \14857 , \14317 );
or \U$14670 ( \14859 , \14624 , \14630 );
nand \U$14671 ( \14860 , \14859 , \14634 );
nor \U$14672 ( \14861 , \14858 , \14860 );
not \U$14673 ( \14862 , \14861 );
xnor \U$14674 ( \14863 , \14856 , \14862 );
buf \U$14675 ( \14864 , \14863 );
buf \U$14676 ( \14865 , \14864 );
not \U$14677 ( \14866 , \8521 );
nand \U$14678 ( \14867 , \13927 , \14866 );
nor \U$14679 ( \14868 , \14649 , \14646 );
and \U$14680 ( \14869 , \14868 , \13829 );
or \U$14681 ( \14870 , \14646 , \14652 );
nand \U$14682 ( \14871 , \14870 , \14656 );
nor \U$14683 ( \14872 , \14869 , \14871 );
not \U$14684 ( \14873 , \14872 );
xnor \U$14685 ( \14874 , \14867 , \14873 );
buf \U$14686 ( \14875 , \14874 );
buf \U$14687 ( \14876 , \14875 );
not \U$14688 ( \14877 , \8359 );
nand \U$14689 ( \14878 , \13923 , \14877 );
nor \U$14690 ( \14879 , \14671 , \14668 );
and \U$14691 ( \14880 , \14879 , \14314 );
or \U$14692 ( \14881 , \14668 , \14674 );
nand \U$14693 ( \14882 , \14881 , \14678 );
nor \U$14694 ( \14883 , \14880 , \14882 );
not \U$14695 ( \14884 , \14883 );
xnor \U$14696 ( \14885 , \14878 , \14884 );
buf \U$14697 ( \14886 , \14885 );
buf \U$14698 ( \14887 , \14886 );
not \U$14699 ( \14888 , \8200 );
nand \U$14700 ( \14889 , \13921 , \14888 );
or \U$14701 ( \14890 , \14690 , \14694 );
nand \U$14702 ( \14891 , \14890 , \14698 );
xnor \U$14703 ( \14892 , \14889 , \14891 );
buf \U$14704 ( \14893 , \14892 );
buf \U$14705 ( \14894 , \14893 );
not \U$14706 ( \14895 , \8041 );
nand \U$14707 ( \14896 , \13918 , \14895 );
or \U$14708 ( \14897 , \14710 , \14714 );
nand \U$14709 ( \14898 , \14897 , \14718 );
xnor \U$14710 ( \14899 , \14896 , \14898 );
buf \U$14711 ( \14900 , \14899 );
buf \U$14712 ( \14901 , \14900 );
not \U$14713 ( \14902 , \7887 );
nand \U$14714 ( \14903 , \13916 , \14902 );
xnor \U$14715 ( \14904 , \14903 , \13914 );
buf \U$14716 ( \14905 , \14904 );
buf \U$14717 ( \14906 , \14905 );
not \U$14718 ( \14907 , \13510 );
nand \U$14719 ( \14908 , \13909 , \14907 );
xnor \U$14720 ( \14909 , \14908 , \14128 );
buf \U$14721 ( \14910 , \14909 );
buf \U$14722 ( \14911 , \14910 );
not \U$14723 ( \14912 , \13503 );
nand \U$14724 ( \14913 , \13907 , \14912 );
xnor \U$14725 ( \14914 , \14913 , \14250 );
buf \U$14726 ( \14915 , \14914 );
buf \U$14727 ( \14916 , \14915 );
not \U$14728 ( \14917 , \13488 );
nand \U$14729 ( \14918 , \13904 , \14917 );
xnor \U$14730 ( \14919 , \14918 , \14341 );
buf \U$14731 ( \14920 , \14919 );
buf \U$14732 ( \14921 , \14920 );
not \U$14733 ( \14922 , \13463 );
nand \U$14734 ( \14923 , \13902 , \14922 );
xnor \U$14735 ( \14924 , \14923 , \14402 );
buf \U$14736 ( \14925 , \14924 );
buf \U$14737 ( \14926 , \14925 );
not \U$14738 ( \14927 , \13428 );
nand \U$14739 ( \14928 , \13898 , \14927 );
xnor \U$14740 ( \14929 , \14928 , \14447 );
buf \U$14741 ( \14930 , \14929 );
buf \U$14742 ( \14931 , \14930 );
not \U$14743 ( \14932 , \13383 );
nand \U$14744 ( \14933 , \13896 , \14932 );
xnor \U$14745 ( \14934 , \14933 , \14490 );
buf \U$14746 ( \14935 , \14934 );
buf \U$14747 ( \14936 , \14935 );
not \U$14748 ( \14937 , \13309 );
nand \U$14749 ( \14938 , \13893 , \14937 );
xnor \U$14750 ( \14939 , \14938 , \14533 );
buf \U$14751 ( \14940 , \14939 );
buf \U$14752 ( \14941 , \14940 );
not \U$14753 ( \14942 , \13194 );
nand \U$14754 ( \14943 , \13891 , \14942 );
xnor \U$14755 ( \14944 , \14943 , \14564 );
buf \U$14756 ( \14945 , \14944 );
buf \U$14757 ( \14946 , \14945 );
not \U$14758 ( \14947 , \13080 );
nand \U$14759 ( \14948 , \13886 , \14947 );
xnor \U$14760 ( \14949 , \14948 , \14587 );
buf \U$14761 ( \14950 , \14949 );
buf \U$14762 ( \14951 , \14950 );
not \U$14763 ( \14952 , \12975 );
nand \U$14764 ( \14953 , \13884 , \14952 );
xnor \U$14765 ( \14954 , \14953 , \14609 );
buf \U$14766 ( \14955 , \14954 );
buf \U$14767 ( \14956 , \14955 );
not \U$14768 ( \14957 , \12873 );
nand \U$14769 ( \14958 , \13881 , \14957 );
xnor \U$14770 ( \14959 , \14958 , \14631 );
buf \U$14771 ( \14960 , \14959 );
buf \U$14772 ( \14961 , \14960 );
not \U$14773 ( \14962 , \12778 );
nand \U$14774 ( \14963 , \13879 , \14962 );
xnor \U$14775 ( \14964 , \14963 , \14653 );
buf \U$14776 ( \14965 , \14964 );
buf \U$14777 ( \14966 , \14965 );
not \U$14778 ( \14967 , \12685 );
nand \U$14779 ( \14968 , \13875 , \14967 );
xnor \U$14780 ( \14969 , \14968 , \14675 );
buf \U$14781 ( \14970 , \14969 );
buf \U$14782 ( \14971 , \14970 );
not \U$14783 ( \14972 , \12600 );
nand \U$14784 ( \14973 , \13873 , \14972 );
xnor \U$14785 ( \14974 , \14973 , \14695 );
buf \U$14786 ( \14975 , \14974 );
buf \U$14787 ( \14976 , \14975 );
not \U$14788 ( \14977 , \12518 );
nand \U$14789 ( \14978 , \13870 , \14977 );
xnor \U$14790 ( \14979 , \14978 , \14715 );
buf \U$14791 ( \14980 , \14979 );
buf \U$14792 ( \14981 , \14980 );
not \U$14793 ( \14982 , \12443 );
nand \U$14794 ( \14983 , \13868 , \14982 );
xnor \U$14795 ( \14984 , \14983 , \14731 );
buf \U$14796 ( \14985 , \14984 );
buf \U$14797 ( \14986 , \14985 );
not \U$14798 ( \14987 , \13765 );
nand \U$14799 ( \14988 , \13862 , \14987 );
xnor \U$14800 ( \14989 , \14988 , \14743 );
buf \U$14801 ( \14990 , \14989 );
buf \U$14802 ( \14991 , \14990 );
not \U$14803 ( \14992 , \13758 );
nand \U$14804 ( \14993 , \13860 , \14992 );
xnor \U$14805 ( \14994 , \14993 , \14755 );
buf \U$14806 ( \14995 , \14994 );
buf \U$14807 ( \14996 , \14995 );
not \U$14808 ( \14997 , \13746 );
nand \U$14809 ( \14998 , \13857 , \14997 );
xnor \U$14810 ( \14999 , \14998 , \14767 );
buf \U$14811 ( \15000 , \14999 );
buf \U$14812 ( \15001 , \15000 );
not \U$14813 ( \15002 , \13729 );
nand \U$14814 ( \15003 , \13855 , \15002 );
xnor \U$14815 ( \15004 , \15003 , \14779 );
buf \U$14816 ( \15005 , \15004 );
buf \U$14817 ( \15006 , \15005 );
not \U$14818 ( \15007 , \13700 );
nand \U$14819 ( \15008 , \13851 , \15007 );
xnor \U$14820 ( \15009 , \15008 , \14791 );
buf \U$14821 ( \15010 , \15009 );
buf \U$14822 ( \15011 , \15010 );
not \U$14823 ( \15012 , \13655 );
nand \U$14824 ( \15013 , \13849 , \15012 );
xnor \U$14825 ( \15014 , \15013 , \14481 );
buf \U$14826 ( \15015 , \15014 );
buf \U$14827 ( \15016 , \15015 );
not \U$14828 ( \15017 , \13613 );
nand \U$14829 ( \15018 , \13846 , \15017 );
xnor \U$14830 ( \15019 , \15018 , \14524 );
buf \U$14831 ( \15020 , \15019 );
buf \U$14832 ( \15021 , \15020 );
not \U$14833 ( \15022 , \13578 );
nand \U$14834 ( \15023 , \13844 , \15022 );
xnor \U$14835 ( \15024 , \15023 , \13842 );
buf \U$14836 ( \15025 , \15024 );
buf \U$14837 ( \15026 , \15025 );
not \U$14838 ( \15027 , \13812 );
nand \U$14839 ( \15028 , \13839 , \15027 );
xnor \U$14840 ( \15029 , \15028 , \14080 );
buf \U$14841 ( \15030 , \15029 );
buf \U$14842 ( \15031 , \15030 );
endmodule

