//
// Conformal-LEC Version 20.10-d005 (29-Apr-2020)
//
module top(RI2b1c4342d4e0_65,RI2b1c4342b6e0_1,RI2b1c4342c5e0_33,RI2b1c4342b758_2,RI2b1c4342c658_34,RI2b1c4342b7d0_3,RI2b1c4342c6d0_35,RI2b1c4342b848_4,RI2b1c4342c748_36,
        RI2b1c4342b8c0_5,RI2b1c4342c7c0_37,RI2b1c4342b938_6,RI2b1c4342c838_38,RI2b1c4342b9b0_7,RI2b1c4342c8b0_39,RI2b1c4342ba28_8,RI2b1c4342c928_40,RI2b1c4342baa0_9,RI2b1c4342c9a0_41,
        RI2b1c4342bb18_10,RI2b1c4342ca18_42,RI2b1c4342bb90_11,RI2b1c4342ca90_43,RI2b1c4342bc08_12,RI2b1c4342cb08_44,RI2b1c4342bc80_13,RI2b1c4342cb80_45,RI2b1c4342bcf8_14,RI2b1c4342cbf8_46,
        RI2b1c4342bd70_15,RI2b1c4342cc70_47,RI2b1c4342bde8_16,RI2b1c4342cce8_48,RI2b1c4342be60_17,RI2b1c4342cd60_49,RI2b1c4342bed8_18,RI2b1c4342cdd8_50,RI2b1c4342bf50_19,RI2b1c4342ce50_51,
        RI2b1c4342bfc8_20,RI2b1c4342cec8_52,RI2b1c4342c040_21,RI2b1c4342cf40_53,RI2b1c4342c0b8_22,RI2b1c4342cfb8_54,RI2b1c4342c130_23,RI2b1c4342d030_55,RI2b1c4342c1a8_24,RI2b1c4342d0a8_56,
        RI2b1c4342c220_25,RI2b1c4342d120_57,RI2b1c4342c298_26,RI2b1c4342d198_58,RI2b1c4342c310_27,RI2b1c4342d210_59,RI2b1c4342c388_28,RI2b1c4342d288_60,RI2b1c4342c400_29,RI2b1c4342d300_61,
        RI2b1c4342c478_30,RI2b1c4342d378_62,RI2b1c4342c4f0_31,RI2b1c4342d3f0_63,RI2b1c4342c568_32,RI2b1c4342d468_64,RI2b1c4342d558_66,RI2b1c4342d5d0_67,RI2b1c4342d648_68,RI2b1c4342d6c0_69,
        RI2b1c4342d738_70,RI2b1c4342d7b0_71,RI2b1c4342d828_72,RI2b1c4342d8a0_73,RI2b1c4342d918_74,RI2b1c4342d990_75,RI2b1c4342da08_76,RI2b1c4342da80_77,RI2b1c4342daf8_78,RI2b1c4342db70_79,
        RI2b1c4342dbe8_80,RI2b1c4342dc60_81,RI2b1c4342dcd8_82,RI2b1c4342dd50_83,RI2b1c4342ddc8_84,RI2b1c4342de40_85,RI2b1c4342deb8_86,RI2b1c4342df30_87,RI2b1c4342dfa8_88,RI2b1c4342e020_89,
        RI2b1c4342e098_90,RI2b1c4342e110_91,RI2b1c4342e188_92,RI2b1c4342e200_93,RI2b1c4342e278_94,RI2b1c4342e2f0_95,RI2b1c4342e368_96,R_61_7d2b4e8,R_62_7d2b590,R_63_7d2b638,
        R_64_7d2b6e0,R_65_7d2b788,R_66_7d2b830,R_67_7d2b8d8,R_68_7d2b980,R_69_7d2ba28,R_6a_7d2bad0,R_6b_7d2bb78,R_6c_7d2bc20,R_6d_7d2bcc8,
        R_6e_7d2bd70,R_6f_7d2be18,R_70_7d2bec0,R_71_7d2bf68,R_72_7d2c010,R_73_7d2c0b8,R_74_7d2c160,R_75_7d2c208,R_76_7d2c2b0,R_77_7d2c358,
        R_78_7d2c400,R_79_7d2c4a8,R_7a_7d2c550,R_7b_7d2c5f8,R_7c_7d2c6a0,R_7d_7d2c748,R_7e_7d2c7f0,R_7f_7d2c898,R_80_7d2c940,R_81_7d2c9e8,
        R_82_7d2ca90,R_83_7d2cb38,R_84_7d2cbe0,R_85_7d2cc88,R_86_7d2cd30,R_87_7d2cdd8,R_88_7d2ce80,R_89_7d2cf28,R_8a_7d2cfd0,R_8b_7d2d078,
        R_8c_7d2d120,R_8d_7d2d1c8,R_8e_7d2d270,R_8f_7d2d318,R_90_7d2d3c0,R_91_7d2d468,R_92_7d2d510,R_93_7d2d5b8,R_94_7d2d660,R_95_7d2d708,
        R_96_7d2d7b0,R_97_7d2d858,R_98_7d2d900,R_99_7d2d9a8,R_9a_7d2da50,R_9b_7d2daf8);
input RI2b1c4342d4e0_65,RI2b1c4342b6e0_1,RI2b1c4342c5e0_33,RI2b1c4342b758_2,RI2b1c4342c658_34,RI2b1c4342b7d0_3,RI2b1c4342c6d0_35,RI2b1c4342b848_4,RI2b1c4342c748_36,
        RI2b1c4342b8c0_5,RI2b1c4342c7c0_37,RI2b1c4342b938_6,RI2b1c4342c838_38,RI2b1c4342b9b0_7,RI2b1c4342c8b0_39,RI2b1c4342ba28_8,RI2b1c4342c928_40,RI2b1c4342baa0_9,RI2b1c4342c9a0_41,
        RI2b1c4342bb18_10,RI2b1c4342ca18_42,RI2b1c4342bb90_11,RI2b1c4342ca90_43,RI2b1c4342bc08_12,RI2b1c4342cb08_44,RI2b1c4342bc80_13,RI2b1c4342cb80_45,RI2b1c4342bcf8_14,RI2b1c4342cbf8_46,
        RI2b1c4342bd70_15,RI2b1c4342cc70_47,RI2b1c4342bde8_16,RI2b1c4342cce8_48,RI2b1c4342be60_17,RI2b1c4342cd60_49,RI2b1c4342bed8_18,RI2b1c4342cdd8_50,RI2b1c4342bf50_19,RI2b1c4342ce50_51,
        RI2b1c4342bfc8_20,RI2b1c4342cec8_52,RI2b1c4342c040_21,RI2b1c4342cf40_53,RI2b1c4342c0b8_22,RI2b1c4342cfb8_54,RI2b1c4342c130_23,RI2b1c4342d030_55,RI2b1c4342c1a8_24,RI2b1c4342d0a8_56,
        RI2b1c4342c220_25,RI2b1c4342d120_57,RI2b1c4342c298_26,RI2b1c4342d198_58,RI2b1c4342c310_27,RI2b1c4342d210_59,RI2b1c4342c388_28,RI2b1c4342d288_60,RI2b1c4342c400_29,RI2b1c4342d300_61,
        RI2b1c4342c478_30,RI2b1c4342d378_62,RI2b1c4342c4f0_31,RI2b1c4342d3f0_63,RI2b1c4342c568_32,RI2b1c4342d468_64,RI2b1c4342d558_66,RI2b1c4342d5d0_67,RI2b1c4342d648_68,RI2b1c4342d6c0_69,
        RI2b1c4342d738_70,RI2b1c4342d7b0_71,RI2b1c4342d828_72,RI2b1c4342d8a0_73,RI2b1c4342d918_74,RI2b1c4342d990_75,RI2b1c4342da08_76,RI2b1c4342da80_77,RI2b1c4342daf8_78,RI2b1c4342db70_79,
        RI2b1c4342dbe8_80,RI2b1c4342dc60_81,RI2b1c4342dcd8_82,RI2b1c4342dd50_83,RI2b1c4342ddc8_84,RI2b1c4342de40_85,RI2b1c4342deb8_86,RI2b1c4342df30_87,RI2b1c4342dfa8_88,RI2b1c4342e020_89,
        RI2b1c4342e098_90,RI2b1c4342e110_91,RI2b1c4342e188_92,RI2b1c4342e200_93,RI2b1c4342e278_94,RI2b1c4342e2f0_95,RI2b1c4342e368_96;
output R_61_7d2b4e8,R_62_7d2b590,R_63_7d2b638,R_64_7d2b6e0,R_65_7d2b788,R_66_7d2b830,R_67_7d2b8d8,R_68_7d2b980,R_69_7d2ba28,
        R_6a_7d2bad0,R_6b_7d2bb78,R_6c_7d2bc20,R_6d_7d2bcc8,R_6e_7d2bd70,R_6f_7d2be18,R_70_7d2bec0,R_71_7d2bf68,R_72_7d2c010,R_73_7d2c0b8,
        R_74_7d2c160,R_75_7d2c208,R_76_7d2c2b0,R_77_7d2c358,R_78_7d2c400,R_79_7d2c4a8,R_7a_7d2c550,R_7b_7d2c5f8,R_7c_7d2c6a0,R_7d_7d2c748,
        R_7e_7d2c7f0,R_7f_7d2c898,R_80_7d2c940,R_81_7d2c9e8,R_82_7d2ca90,R_83_7d2cb38,R_84_7d2cbe0,R_85_7d2cc88,R_86_7d2cd30,R_87_7d2cdd8,
        R_88_7d2ce80,R_89_7d2cf28,R_8a_7d2cfd0,R_8b_7d2d078,R_8c_7d2d120,R_8d_7d2d1c8,R_8e_7d2d270,R_8f_7d2d318,R_90_7d2d3c0,R_91_7d2d468,
        R_92_7d2d510,R_93_7d2d5b8,R_94_7d2d660,R_95_7d2d708,R_96_7d2d7b0,R_97_7d2d858,R_98_7d2d900,R_99_7d2d9a8,R_9a_7d2da50,R_9b_7d2daf8;

wire \156 , \157 , \158 , \159 , \160 , \161 , \162 , \163 , \164 ,
         \165 , \166 , \167 , \168 , \169 , \170 , \171 , \172 , \173 , \174 ,
         \175 , \176 , \177 , \178 , \179 , \180 , \181 , \182 , \183 , \184 ,
         \185 , \186 , \187 , \188 , \189_N$1 , \190_N$2 , \191_N$3 , \192_N$4 , \193_N$5 , \194_N$6 ,
         \195_N$7 , \196_N$8 , \197_N$9 , \198_N$10 , \199_N$11 , \200_N$12 , \201_N$13 , \202_N$14 , \203_N$15 , \204_N$16 ,
         \205_N$17 , \206_N$18 , \207_N$19 , \208_N$20 , \209_N$21 , \210_N$22 , \211_N$23 , \212_N$24 , \213_N$25 , \214_N$26 ,
         \215_N$27 , \216_N$28 , \217_N$29 , \218_N$30 , \219_N$31 , \220_N$32 , \221_ZERO , \222_ONE , \223 , \224 ,
         \225 , \226 , \227 , \228 , \229 , \230 , \231 , \232 , \233 , \234 ,
         \235 , \236 , \237 , \238 , \239 , \240 , \241 , \242 , \243 , \244 ,
         \245 , \246 , \247 , \248 , \249 , \250 , \251 , \252 , \253 , \254 ,
         \255 , \256 , \257 , \258 , \259 , \260 , \261 , \262 , \263 , \264 ,
         \265 , \266 , \267 , \268 , \269 , \270 , \271 , \272 , \273 , \274 ,
         \275 , \276 , \277 , \278 , \279 , \280 , \281 , \282 , \283 , \284 ,
         \285 , \286 , \287 , \288 , \289 , \290 , \291 , \292 , \293 , \294 ,
         \295 , \296 , \297 , \298 , \299 , \300 , \301 , \302 , \303 , \304 ,
         \305 , \306 , \307 , \308 , \309 , \310 , \311 , \312 , \313 , \314 ,
         \315 , \316 , \317 , \318 , \319 , \320 , \321 , \322 , \323 , \324 ,
         \325 , \326 , \327 , \328 , \329 , \330 , \331 , \332 , \333 , \334 ,
         \335 , \336 , \337 , \338 , \339 , \340 , \341 , \342 , \343 , \344 ,
         \345 , \346 , \347 , \348 , \349 , \350 , \351 , \352 , \353 , \354 ,
         \355 , \356 , \357 , \358 , \359 , \360 , \361 , \362 , \363 , \364 ,
         \365 , \366 , \367 , \368 , \369 , \370 , \371 , \372 , \373 , \374 ,
         \375 , \376 , \377 , \378 , \379 , \380 , \381 , \382 , \383 , \384 ,
         \385 , \386 , \387 , \388 , \389 , \390 , \391 , \392 , \393 , \394 ,
         \395 , \396 , \397 , \398 , \399 , \400 , \401 , \402 , \403 , \404 ,
         \405 , \406 , \407 , \408 , \409 , \410 , \411 , \412 , \413 , \414 ,
         \415 , \416 , \417 , \418 , \419 , \420 , \421 , \422 , \423 , \424 ,
         \425 , \426 , \427 , \428 , \429 , \430 , \431 , \432 , \433 , \434 ,
         \435 , \436 , \437 , \438 , \439 , \440 , \441 , \442 , \443 , \444 ,
         \445 , \446 , \447 , \448 , \449 , \450 , \451 , \452 , \453 , \454 ,
         \455 , \456 , \457 , \458 , \459 , \460 , \461 , \462 , \463 , \464 ,
         \465 , \466 , \467 , \468 , \469 , \470 , \471 , \472 , \473 , \474 ,
         \475 , \476_nR2b9 , \477 , \478 , \479 , \480 , \481 , \482 , \483_nR2ad , \484 ,
         \485 , \486 , \487 , \488 , \489 , \490 , \491_nR2a1 , \492 , \493 , \494 ,
         \495 , \496 , \497 , \498 , \499 , \500 , \501 , \502 , \503 , \504 ,
         \505 , \506 , \507 , \508 , \509 , \510 , \511 , \512 , \513 , \514 ,
         \515 , \516 , \517 , \518 , \519_nR295 , \520 , \521 , \522 , \523 , \524 ,
         \525 , \526_nR289 , \527 , \528 , \529 , \530 , \531 , \532 , \533 , \534 ,
         \535 , \536 , \537 , \538 , \539 , \540 , \541 , \542 , \543 , \544 ,
         \545 , \546 , \547 , \548 , \549 , \550 , \551 , \552 , \553 , \554 ,
         \555_nR27d , \556 , \557 , \558 , \559 , \560 , \561 , \562_nR271 , \563 , \564 ,
         \565 , \566 , \567 , \568 , \569 , \570 , \571 , \572 , \573_nR151 , \574 ,
         \575 , \576 , \577 , \578 , \579_nR129 , \580 , \581 , \582 , \583 , \584 ,
         \585 , \586 , \587 , \588 , \589 , \590 , \591 , \592 , \593 , \594 ,
         \595 , \596 , \597 , \598 , \599 , \600 , \601 , \602 , \603 , \604 ,
         \605 , \606 , \607 , \608 , \609 , \610 , \611 , \612 , \613 , \614 ,
         \615 , \616 , \617 , \618 , \619 , \620 , \621 , \622 , \623 , \624 ,
         \625 , \626 , \627_nR169 , \628 , \629 , \630 , \631 , \632 , \633 , \634_nR15d ,
         \635 , \636 , \637 , \638 , \639 , \640 , \641 , \642 , \643 , \644 ,
         \645 , \646 , \647 , \648 , \649 , \650 , \651 , \652 , \653 , \654 ,
         \655 , \656 , \657_nR181 , \658 , \659 , \660 , \661 , \662 , \663 , \664_nR175 ,
         \665 , \666 , \667 , \668 , \669 , \670 , \671 , \672 , \673 , \674 ,
         \675 , \676 , \677 , \678 , \679 , \680 , \681 , \682 , \683 , \684_nR199 ,
         \685 , \686 , \687 , \688 , \689 , \690 , \691_nR18d , \692 , \693 , \694 ,
         \695 , \696 , \697 , \698 , \699 , \700 , \701 , \702 , \703 , \704 ,
         \705 , \706 , \707 , \708 , \709 , \710 , \711 , \712_nR1b1 , \713 , \714 ,
         \715 , \716 , \717 , \718 , \719_nR1a5 , \720 , \721 , \722 , \723 , \724 ,
         \725 , \726 , \727 , \728 , \729 , \730 , \731 , \732 , \733 , \734 ,
         \735 , \736 , \737 , \738 , \739 , \740 , \741 , \742 , \743_nR1c9 , \744 ,
         \745 , \746 , \747 , \748 , \749 , \750_nR1bd , \751 , \752 , \753 , \754 ,
         \755 , \756 , \757 , \758 , \759 , \760 , \761 , \762 , \763 , \764 ,
         \765 , \766 , \767 , \768 , \769 , \770_nR1e1 , \771 , \772 , \773 , \774 ,
         \775 , \776 , \777_nR1d5 , \778 , \779 , \780 , \781 , \782 , \783 , \784 ,
         \785 , \786 , \787 , \788 , \789 , \790 , \791 , \792 , \793 , \794 ,
         \795 , \796 , \797 , \798_nR1f9 , \799 , \800 , \801 , \802 , \803 , \804 ,
         \805_nR1ed , \806 , \807 , \808 , \809 , \810 , \811 , \812 , \813 , \814 ,
         \815 , \816 , \817 , \818 , \819 , \820 , \821 , \822 , \823 , \824 ,
         \825 , \826 , \827 , \828 , \829 , \830 , \831_nR211 , \832 , \833 , \834 ,
         \835 , \836 , \837 , \838_nR205 , \839 , \840 , \841 , \842 , \843 , \844 ,
         \845 , \846 , \847 , \848 , \849 , \850 , \851 , \852 , \853 , \854 ,
         \855 , \856 , \857 , \858_nR229 , \859 , \860 , \861 , \862 , \863 , \864 ,
         \865_nR21d , \866 , \867 , \868 , \869 , \870 , \871 , \872 , \873 , \874 ,
         \875 , \876 , \877 , \878 , \879 , \880 , \881 , \882 , \883 , \884 ,
         \885 , \886_nR241 , \887 , \888 , \889 , \890 , \891 , \892 , \893_nR235 , \894 ,
         \895 , \896 , \897 , \898 , \899 , \900 , \901 , \902 , \903 , \904 ,
         \905 , \906 , \907 , \908 , \909 , \910 , \911 , \912 , \913 , \914 ,
         \915 , \916_nR259 , \917 , \918 , \919 , \920 , \921 , \922 , \923_nR24d , \924 ,
         \925 , \926 , \927 , \928 , \929 , \930 , \931 , \932 , \933 , \934 ,
         \935 , \936 , \937 , \938 , \939 , \940 , \941 , \942 , \943_nR265 , \944 ,
         \945 , \946 , \947 , \948 , \949 , \950 , \951 , \952 , \953 , \954 ,
         \955 , \956 , \957 , \958 , \959 , \960 , \961 , \962 , \963 , \964 ,
         \965 , \966 , \967 , \968 , \969 , \970 , \971 , \972 , \973 , \974 ,
         \975 , \976 , \977 , \978 , \979 , \980 , \981 , \982 , \983 , \984 ,
         \985 , \986 , \987 , \988 , \989 , \990 , \991 , \992 , \993 , \994 ,
         \995 , \996 , \997 , \998 , \999 , \1000 , \1001 , \1002 , \1003 , \1004 ,
         \1005 , \1006 , \1007 , \1008 , \1009 , \1010 , \1011 , \1012 , \1013 , \1014 ,
         \1015 , \1016 , \1017 , \1018 , \1019 , \1020 , \1021 , \1022 , \1023 , \1024 ,
         \1025 , \1026 , \1027 , \1028 , \1029 , \1030 , \1031 , \1032 , \1033 , \1034 ,
         \1035 , \1036 , \1037 , \1038 , \1039 , \1040 , \1041 , \1042 , \1043 , \1044 ,
         \1045 , \1046 , \1047 , \1048 , \1049 , \1050 , \1051 , \1052 , \1053 , \1054 ,
         \1055 , \1056 , \1057 , \1058 , \1059 , \1060 , \1061 , \1062 , \1063 , \1064 ,
         \1065 , \1066 , \1067 , \1068 , \1069 , \1070 , \1071 , \1072 , \1073 , \1074 ,
         \1075 , \1076 , \1077 , \1078 , \1079 , \1080 , \1081 , \1082 , \1083 , \1084 ,
         \1085 , \1086 , \1087 , \1088 , \1089 , \1090 , \1091 , \1092 , \1093 , \1094 ,
         \1095 , \1096 , \1097 , \1098 , \1099 , \1100 , \1101 , \1102 , \1103 , \1104 ,
         \1105 , \1106 , \1107 , \1108 , \1109 , \1110 , \1111 , \1112 , \1113 , \1114 ,
         \1115 , \1116 , \1117 , \1118 , \1119 , \1120 , \1121 , \1122 , \1123 , \1124 ,
         \1125 , \1126 , \1127 , \1128 , \1129 , \1130 , \1131 , \1132 , \1133 , \1134 ,
         \1135 , \1136 , \1137 , \1138 , \1139 , \1140 , \1141 , \1142 , \1143 , \1144 ,
         \1145 , \1146 , \1147 , \1148 , \1149 , \1150 , \1151 , \1152 , \1153 , \1154 ,
         \1155 , \1156 , \1157 , \1158 , \1159 , \1160 , \1161 , \1162 , \1163 , \1164 ,
         \1165 , \1166 , \1167 , \1168 , \1169 , \1170 , \1171 , \1172 , \1173 , \1174 ,
         \1175 , \1176 , \1177 , \1178 , \1179 , \1180 , \1181 , \1182 , \1183 , \1184 ,
         \1185 , \1186 , \1187 , \1188 , \1189 , \1190 , \1191 , \1192 , \1193 , \1194 ,
         \1195 , \1196 , \1197 , \1198 , \1199 , \1200 , \1201 , \1202 , \1203 , \1204 ,
         \1205 , \1206 , \1207 , \1208 , \1209 , \1210 , \1211 , \1212 , \1213 , \1214 ,
         \1215 , \1216 , \1217 , \1218 , \1219 , \1220 , \1221 , \1222 , \1223 , \1224 ,
         \1225 , \1226 , \1227 , \1228 , \1229 , \1230 , \1231 , \1232 , \1233 , \1234 ,
         \1235 , \1236 , \1237 , \1238 , \1239 , \1240 , \1241 , \1242 , \1243 , \1244 ,
         \1245 , \1246 , \1247 , \1248 , \1249 , \1250 , \1251 , \1252 , \1253 , \1254 ,
         \1255 , \1256 , \1257 , \1258 , \1259 , \1260 , \1261 , \1262 , \1263 , \1264 ,
         \1265 , \1266 , \1267 , \1268 , \1269 , \1270 , \1271 , \1272 , \1273 , \1274 ,
         \1275 , \1276 , \1277 , \1278 , \1279 , \1280 , \1281 , \1282 , \1283 , \1284 ,
         \1285 , \1286 , \1287 , \1288 , \1289 , \1290 , \1291 , \1292 , \1293 , \1294 ,
         \1295 , \1296 , \1297 , \1298 , \1299 , \1300 , \1301 , \1302 , \1303 , \1304 ,
         \1305 , \1306 , \1307 , \1308 , \1309 , \1310 , \1311 , \1312 , \1313 , \1314 ,
         \1315 , \1316 , \1317 , \1318 , \1319 , \1320 , \1321 , \1322 , \1323 , \1324 ,
         \1325 , \1326 , \1327 , \1328 , \1329 , \1330 , \1331 , \1332 , \1333 , \1334 ,
         \1335 , \1336 , \1337 , \1338 , \1339 , \1340 , \1341 , \1342 , \1343 , \1344 ,
         \1345 , \1346 , \1347 , \1348 , \1349 , \1350 , \1351 , \1352 , \1353 , \1354 ,
         \1355 , \1356 , \1357 , \1358 , \1359 , \1360 , \1361 , \1362 , \1363 , \1364 ,
         \1365 , \1366 , \1367 , \1368 , \1369 , \1370 , \1371 , \1372 , \1373 , \1374 ,
         \1375 , \1376 , \1377 , \1378 , \1379 , \1380 , \1381 , \1382 , \1383 , \1384 ,
         \1385 , \1386 , \1387 , \1388 , \1389 , \1390 , \1391 , \1392 , \1393 , \1394 ,
         \1395 , \1396 , \1397 , \1398 , \1399 , \1400 , \1401 , \1402 , \1403 , \1404 ,
         \1405 , \1406 , \1407 , \1408 , \1409 , \1410 , \1411 , \1412 , \1413 , \1414 ,
         \1415 , \1416 , \1417 , \1418 , \1419 , \1420 , \1421 , \1422 , \1423 , \1424 ,
         \1425 , \1426 , \1427 , \1428 , \1429 , \1430 , \1431 , \1432 , \1433 , \1434 ,
         \1435 , \1436 , \1437 , \1438 , \1439 , \1440 , \1441 , \1442 , \1443 , \1444 ,
         \1445 , \1446 , \1447 , \1448 , \1449 , \1450 , \1451 , \1452 , \1453 , \1454 ,
         \1455 , \1456 , \1457 , \1458 , \1459 , \1460 , \1461 , \1462 , \1463 , \1464 ,
         \1465 , \1466 , \1467 , \1468 , \1469 , \1470 , \1471 , \1472 , \1473 , \1474 ,
         \1475 , \1476 , \1477 , \1478 , \1479 , \1480 , \1481 , \1482 , \1483 , \1484 ,
         \1485 , \1486 , \1487 , \1488 , \1489 , \1490 , \1491 , \1492 , \1493 , \1494 ,
         \1495 , \1496 , \1497 , \1498 , \1499 , \1500 , \1501 , \1502 , \1503 , \1504 ,
         \1505 , \1506 , \1507 , \1508 , \1509 , \1510 , \1511 , \1512 , \1513 , \1514 ,
         \1515 , \1516 , \1517 , \1518 , \1519 , \1520 , \1521 , \1522 , \1523 , \1524 ,
         \1525 , \1526 , \1527 , \1528 , \1529 , \1530 , \1531 , \1532 , \1533 , \1534 ,
         \1535 , \1536 , \1537 , \1538 , \1539 , \1540 , \1541 , \1542 , \1543 , \1544 ,
         \1545 , \1546 , \1547 , \1548 , \1549 , \1550 , \1551 , \1552 , \1553 , \1554 ,
         \1555 , \1556 , \1557 , \1558 , \1559 , \1560 , \1561 , \1562 , \1563 , \1564 ,
         \1565 , \1566 , \1567 , \1568 , \1569 , \1570 , \1571 , \1572 , \1573 , \1574 ,
         \1575 , \1576 , \1577 , \1578 , \1579 , \1580 , \1581 , \1582 , \1583 , \1584 ,
         \1585 , \1586 , \1587 , \1588 , \1589 , \1590 , \1591 , \1592 , \1593 , \1594 ,
         \1595 , \1596 , \1597 , \1598 , \1599 , \1600 , \1601 , \1602 , \1603 , \1604 ,
         \1605 , \1606 , \1607 , \1608 , \1609 , \1610 , \1611 , \1612 , \1613 , \1614 ,
         \1615 , \1616 , \1617 , \1618 , \1619 , \1620 , \1621 , \1622 , \1623 , \1624 ,
         \1625 , \1626 , \1627 , \1628 , \1629 , \1630 , \1631 , \1632 , \1633 , \1634 ,
         \1635 , \1636 , \1637 , \1638 , \1639 , \1640 , \1641 , \1642 , \1643 , \1644 ,
         \1645 , \1646 , \1647 , \1648 , \1649 , \1650 , \1651 , \1652 , \1653 , \1654 ,
         \1655 , \1656 , \1657 , \1658 , \1659 , \1660 , \1661 , \1662 , \1663 , \1664 ,
         \1665 , \1666 , \1667 , \1668 , \1669 , \1670 , \1671 , \1672 , \1673 , \1674 ,
         \1675 , \1676 , \1677 , \1678 , \1679 , \1680 , \1681 , \1682 , \1683 , \1684 ,
         \1685 , \1686 , \1687 , \1688 , \1689 , \1690 , \1691 , \1692 , \1693 , \1694 ,
         \1695 , \1696 , \1697 , \1698 , \1699 , \1700 , \1701 , \1702 , \1703 , \1704 ,
         \1705 , \1706 , \1707 , \1708 , \1709 , \1710 , \1711 , \1712 , \1713 , \1714 ,
         \1715 , \1716 , \1717 , \1718 , \1719 , \1720 , \1721 , \1722 , \1723 , \1724 ,
         \1725 , \1726 , \1727 , \1728 , \1729 , \1730 , \1731 , \1732 , \1733 , \1734 ,
         \1735 , \1736 , \1737 , \1738 , \1739 , \1740 , \1741 , \1742 , \1743 , \1744 ,
         \1745 , \1746 , \1747 , \1748 , \1749 , \1750 , \1751 , \1752 , \1753 , \1754 ,
         \1755 , \1756 , \1757 , \1758 , \1759 , \1760 , \1761 , \1762 , \1763 , \1764 ,
         \1765 , \1766 , \1767 , \1768 , \1769 , \1770 , \1771 , \1772 , \1773 , \1774 ,
         \1775 , \1776 , \1777 , \1778 , \1779 , \1780 , \1781 , \1782 , \1783 , \1784 ,
         \1785 , \1786 , \1787 , \1788 , \1789 , \1790 , \1791 , \1792 , \1793 , \1794 ,
         \1795 , \1796 , \1797 , \1798 , \1799 , \1800 , \1801 , \1802 , \1803 , \1804 ,
         \1805 , \1806 , \1807 , \1808 , \1809 , \1810 , \1811 , \1812 , \1813 , \1814 ,
         \1815 , \1816 , \1817 , \1818 , \1819 , \1820 , \1821 , \1822 , \1823 , \1824 ,
         \1825 , \1826 , \1827 , \1828 , \1829 , \1830 , \1831 , \1832 , \1833 , \1834 ,
         \1835 , \1836 , \1837 , \1838 , \1839 , \1840 , \1841 , \1842 , \1843 , \1844 ,
         \1845 , \1846 , \1847 , \1848 , \1849 , \1850 , \1851 , \1852 , \1853 , \1854 ,
         \1855 , \1856 , \1857 , \1858 , \1859 , \1860 , \1861 , \1862 , \1863 , \1864 ,
         \1865 , \1866 , \1867 , \1868 , \1869 , \1870 , \1871 , \1872 , \1873 , \1874 ,
         \1875 , \1876 , \1877 , \1878 , \1879 , \1880 , \1881 , \1882 , \1883 , \1884 ,
         \1885 , \1886 , \1887 , \1888 , \1889 , \1890 , \1891 , \1892 , \1893 , \1894 ,
         \1895 , \1896 , \1897 , \1898 , \1899 , \1900 , \1901 , \1902 , \1903 , \1904 ,
         \1905 , \1906 , \1907 , \1908 , \1909 , \1910 , \1911 , \1912 , \1913 , \1914 ,
         \1915 , \1916 , \1917 , \1918 , \1919 , \1920 , \1921 , \1922 , \1923 , \1924 ,
         \1925 , \1926 , \1927 , \1928 , \1929 , \1930 , \1931 , \1932 , \1933 , \1934 ,
         \1935 , \1936 , \1937 , \1938 , \1939 , \1940 , \1941 , \1942 , \1943 , \1944 ,
         \1945 , \1946 , \1947 , \1948 , \1949 , \1950 , \1951 , \1952 , \1953 , \1954 ,
         \1955 , \1956 , \1957 , \1958 , \1959 , \1960 , \1961 , \1962 , \1963 , \1964 ,
         \1965 , \1966 , \1967 , \1968 , \1969 , \1970 , \1971 , \1972 , \1973 , \1974 ,
         \1975 , \1976 , \1977 , \1978 , \1979 , \1980 , \1981 , \1982 , \1983 , \1984 ,
         \1985 , \1986 , \1987 , \1988 , \1989 , \1990 , \1991 , \1992 , \1993 , \1994 ,
         \1995 , \1996 , \1997 , \1998 , \1999 , \2000 , \2001 , \2002 , \2003 , \2004 ,
         \2005 , \2006 , \2007 , \2008 , \2009 , \2010 , \2011 , \2012 , \2013 , \2014 ,
         \2015 , \2016 , \2017 , \2018 , \2019 , \2020 , \2021 , \2022 , \2023 , \2024 ,
         \2025 , \2026 , \2027 , \2028 , \2029 , \2030 , \2031 , \2032 , \2033 , \2034 ,
         \2035 , \2036 , \2037 , \2038 , \2039 , \2040 , \2041 , \2042 , \2043 , \2044 ,
         \2045 , \2046 , \2047 , \2048 , \2049 , \2050 , \2051 , \2052 , \2053 , \2054 ,
         \2055 , \2056 , \2057 , \2058 , \2059 , \2060 , \2061 , \2062 , \2063 , \2064 ,
         \2065 , \2066 , \2067 , \2068 , \2069 , \2070 , \2071 , \2072 , \2073 , \2074 ,
         \2075 , \2076 , \2077 , \2078 , \2079 , \2080 , \2081 , \2082 , \2083 , \2084 ,
         \2085 , \2086 , \2087 , \2088 , \2089 , \2090 , \2091 , \2092 , \2093 , \2094 ,
         \2095 , \2096 , \2097 , \2098 , \2099 , \2100 , \2101 , \2102 , \2103 , \2104 ,
         \2105 , \2106 , \2107 , \2108 , \2109 , \2110 , \2111 , \2112 , \2113 , \2114 ,
         \2115 , \2116 , \2117 , \2118 , \2119 , \2120 , \2121 , \2122 , \2123 , \2124 ,
         \2125 , \2126 , \2127 , \2128 , \2129 , \2130 , \2131 , \2132 , \2133 , \2134 ,
         \2135 , \2136 , \2137 , \2138 , \2139 , \2140 , \2141 , \2142 , \2143 , \2144 ,
         \2145 , \2146 , \2147 , \2148 , \2149 , \2150 , \2151 , \2152 , \2153 , \2154 ,
         \2155 , \2156 , \2157 , \2158 , \2159 , \2160 , \2161 , \2162 , \2163 , \2164 ,
         \2165 , \2166 , \2167 , \2168 , \2169 , \2170 , \2171 , \2172 , \2173 , \2174 ,
         \2175 , \2176 , \2177 , \2178 , \2179 , \2180 , \2181 , \2182 , \2183 , \2184 ,
         \2185 , \2186 , \2187 , \2188 , \2189 , \2190 , \2191 , \2192 , \2193 , \2194 ,
         \2195 , \2196 , \2197 , \2198 , \2199 , \2200 , \2201 , \2202 , \2203 , \2204 ,
         \2205 , \2206 , \2207 , \2208 , \2209 , \2210 , \2211 , \2212 , \2213 , \2214 ,
         \2215 , \2216 , \2217 , \2218 , \2219 , \2220 , \2221 , \2222 , \2223 , \2224 ,
         \2225 , \2226 , \2227 , \2228 , \2229 , \2230 , \2231 , \2232 , \2233 , \2234 ,
         \2235 , \2236 , \2237 , \2238 , \2239 , \2240 , \2241 , \2242 , \2243 , \2244 ,
         \2245 , \2246 , \2247 , \2248 , \2249 , \2250 , \2251 , \2252 , \2253 , \2254 ,
         \2255 , \2256 , \2257 , \2258 , \2259 , \2260 , \2261 , \2262 , \2263 , \2264 ,
         \2265 , \2266 , \2267 , \2268 , \2269 , \2270 , \2271 , \2272 , \2273 , \2274 ,
         \2275 , \2276 , \2277 , \2278 , \2279 , \2280 , \2281 , \2282 , \2283 , \2284 ,
         \2285 , \2286 , \2287 , \2288 , \2289 , \2290 , \2291 , \2292 , \2293 , \2294 ,
         \2295 , \2296 , \2297 , \2298 , \2299 , \2300 , \2301 , \2302 , \2303 , \2304 ,
         \2305 , \2306 , \2307 , \2308 , \2309 , \2310 , \2311 , \2312 , \2313 , \2314 ,
         \2315 , \2316 , \2317 , \2318 , \2319 , \2320 , \2321 , \2322 , \2323 , \2324 ,
         \2325 , \2326 , \2327 , \2328 , \2329 , \2330 , \2331 , \2332 , \2333 , \2334 ,
         \2335 , \2336 , \2337 , \2338 , \2339 , \2340 , \2341 , \2342 , \2343 , \2344 ,
         \2345 , \2346 , \2347 , \2348 , \2349 , \2350 , \2351 , \2352 , \2353 , \2354 ,
         \2355 , \2356 , \2357 , \2358 , \2359 , \2360 , \2361 , \2362 , \2363 , \2364 ,
         \2365 , \2366 , \2367 , \2368 , \2369 , \2370 , \2371 , \2372 , \2373 , \2374 ,
         \2375 , \2376 , \2377 , \2378 , \2379 , \2380 , \2381 , \2382 , \2383 , \2384 ,
         \2385 , \2386 , \2387 , \2388 , \2389 , \2390 , \2391 , \2392 , \2393 , \2394 ,
         \2395 , \2396 , \2397 , \2398 , \2399 , \2400 , \2401 , \2402 , \2403 , \2404 ,
         \2405 , \2406 , \2407 , \2408 , \2409 , \2410 , \2411 , \2412 , \2413 , \2414 ,
         \2415 , \2416 , \2417 , \2418 , \2419 , \2420 , \2421 , \2422 , \2423 , \2424 ,
         \2425 , \2426 , \2427 , \2428 , \2429 , \2430 , \2431 , \2432 , \2433 , \2434 ,
         \2435 , \2436 , \2437 , \2438 , \2439 , \2440 , \2441 , \2442 , \2443 , \2444 ,
         \2445 , \2446 , \2447 , \2448 , \2449 , \2450 , \2451 , \2452 , \2453 , \2454 ,
         \2455 , \2456 , \2457 , \2458 , \2459 , \2460 , \2461 , \2462 , \2463 , \2464 ,
         \2465 , \2466 , \2467 , \2468 , \2469 , \2470 , \2471 , \2472 , \2473 , \2474 ,
         \2475 , \2476 , \2477 , \2478 , \2479 , \2480 , \2481 , \2482 , \2483 , \2484 ,
         \2485 , \2486 , \2487 , \2488 , \2489 , \2490 , \2491 , \2492 , \2493 , \2494 ,
         \2495 , \2496 , \2497 , \2498 , \2499 , \2500 , \2501 , \2502 , \2503 , \2504 ,
         \2505 , \2506 , \2507 , \2508 , \2509 , \2510 , \2511 , \2512 , \2513 , \2514 ,
         \2515 , \2516 , \2517 , \2518 , \2519 , \2520 , \2521 , \2522 , \2523 , \2524 ,
         \2525 , \2526 , \2527 , \2528 , \2529 , \2530 , \2531 , \2532 , \2533 , \2534 ,
         \2535 , \2536 , \2537 , \2538 , \2539 , \2540 , \2541 , \2542 , \2543 , \2544 ,
         \2545 , \2546 , \2547 , \2548 , \2549 , \2550 , \2551 , \2552 , \2553 , \2554 ,
         \2555 , \2556 , \2557 , \2558 , \2559 , \2560 , \2561 , \2562 , \2563 , \2564 ,
         \2565 , \2566 , \2567 , \2568 , \2569 , \2570 , \2571 , \2572 , \2573 , \2574 ,
         \2575 , \2576 , \2577 , \2578 , \2579 , \2580 , \2581 , \2582 , \2583 , \2584 ,
         \2585 , \2586 , \2587 , \2588 , \2589 , \2590 , \2591 , \2592 , \2593 , \2594 ,
         \2595 , \2596 , \2597 , \2598 , \2599 , \2600 , \2601 , \2602 , \2603 , \2604 ,
         \2605 , \2606 , \2607 , \2608 , \2609 , \2610 , \2611 , \2612 , \2613 , \2614 ,
         \2615 , \2616 , \2617 , \2618 , \2619 , \2620 , \2621 , \2622 , \2623 , \2624 ,
         \2625 , \2626 , \2627 , \2628 , \2629 , \2630 , \2631 , \2632 , \2633 , \2634 ,
         \2635 , \2636 , \2637 , \2638 , \2639 , \2640 , \2641 , \2642 , \2643 , \2644 ,
         \2645 , \2646 , \2647 , \2648 , \2649 , \2650 , \2651 , \2652 , \2653 , \2654 ,
         \2655 , \2656 , \2657 , \2658 , \2659 , \2660 , \2661 , \2662 , \2663 , \2664 ,
         \2665 , \2666 , \2667 , \2668 , \2669 , \2670 , \2671 , \2672 , \2673 , \2674 ,
         \2675 , \2676 , \2677 , \2678 , \2679 , \2680 , \2681 , \2682 , \2683 , \2684 ,
         \2685 , \2686 , \2687 , \2688 , \2689 , \2690 , \2691 , \2692 , \2693 , \2694 ,
         \2695 , \2696 , \2697 , \2698 , \2699 , \2700 , \2701 , \2702 , \2703 , \2704 ,
         \2705 , \2706 , \2707 , \2708 , \2709 , \2710 , \2711 , \2712 , \2713 , \2714 ,
         \2715 , \2716 , \2717 , \2718 , \2719 , \2720 , \2721 , \2722 , \2723 , \2724 ,
         \2725 , \2726 , \2727 , \2728 , \2729 , \2730 , \2731 , \2732 , \2733 , \2734 ,
         \2735 , \2736 , \2737 , \2738 , \2739 , \2740 , \2741 , \2742 , \2743 , \2744 ,
         \2745 , \2746 , \2747 , \2748 , \2749 , \2750 , \2751 , \2752 , \2753 , \2754 ,
         \2755 , \2756 , \2757 , \2758 , \2759 , \2760 , \2761 , \2762 , \2763 , \2764 ,
         \2765 , \2766 , \2767 , \2768 , \2769 , \2770 , \2771 , \2772 , \2773 , \2774 ,
         \2775 , \2776 , \2777 , \2778 , \2779 , \2780 , \2781 , \2782 , \2783 , \2784 ,
         \2785 , \2786 , \2787 , \2788 , \2789 , \2790 , \2791 , \2792 , \2793 , \2794 ,
         \2795 , \2796 , \2797 , \2798 , \2799 , \2800 , \2801 , \2802 , \2803 , \2804 ,
         \2805 , \2806 , \2807 , \2808 , \2809 , \2810 , \2811 , \2812 , \2813 , \2814 ,
         \2815 , \2816 , \2817 , \2818 , \2819 , \2820 , \2821 , \2822 , \2823 , \2824 ,
         \2825 , \2826 , \2827 , \2828 , \2829 , \2830 , \2831 , \2832 , \2833 , \2834 ,
         \2835 , \2836 , \2837 , \2838 , \2839 , \2840 , \2841 , \2842 , \2843 , \2844 ,
         \2845 , \2846 , \2847 , \2848 , \2849 , \2850 , \2851 , \2852 , \2853 , \2854 ,
         \2855 , \2856 , \2857 , \2858 , \2859 , \2860 , \2861 , \2862 , \2863 , \2864 ,
         \2865 , \2866 , \2867 , \2868 , \2869 , \2870 , \2871 , \2872 , \2873 , \2874 ,
         \2875 , \2876 , \2877 , \2878 , \2879 , \2880 , \2881 , \2882 , \2883 , \2884 ,
         \2885 , \2886 , \2887 , \2888 , \2889 , \2890 , \2891 , \2892 , \2893 , \2894 ,
         \2895 , \2896 , \2897 , \2898 , \2899 , \2900 , \2901 , \2902 , \2903 , \2904 ,
         \2905 , \2906 , \2907 , \2908 , \2909 , \2910 , \2911 , \2912 , \2913 , \2914 ,
         \2915 , \2916 , \2917 , \2918 , \2919 , \2920 , \2921 , \2922 , \2923 , \2924 ,
         \2925 , \2926 , \2927 , \2928 , \2929 , \2930 , \2931 , \2932 , \2933 , \2934 ,
         \2935 , \2936 , \2937 , \2938 , \2939 , \2940 , \2941 , \2942 , \2943 , \2944 ,
         \2945 , \2946 , \2947 , \2948 , \2949 , \2950 , \2951 , \2952 , \2953 , \2954 ,
         \2955 , \2956 , \2957 , \2958 , \2959 , \2960 , \2961 , \2962 , \2963 , \2964 ,
         \2965 , \2966 , \2967 , \2968 , \2969 , \2970 , \2971 , \2972 , \2973 , \2974 ,
         \2975 , \2976 , \2977 , \2978 , \2979 , \2980 , \2981 , \2982 , \2983 , \2984 ,
         \2985 , \2986 , \2987 , \2988 , \2989 , \2990 , \2991 , \2992 , \2993 , \2994 ,
         \2995 , \2996 , \2997 , \2998 , \2999 , \3000 , \3001 , \3002 , \3003 , \3004 ,
         \3005 , \3006 , \3007 , \3008 , \3009 , \3010 , \3011 , \3012 , \3013 , \3014 ,
         \3015 , \3016 , \3017 , \3018 , \3019 , \3020 , \3021 , \3022 , \3023 , \3024 ,
         \3025 , \3026 , \3027 , \3028 , \3029 , \3030 , \3031 , \3032 , \3033 , \3034 ,
         \3035 , \3036 , \3037 , \3038 , \3039 , \3040 , \3041 , \3042 , \3043 , \3044 ,
         \3045 , \3046 , \3047 , \3048 , \3049 , \3050 , \3051 , \3052 , \3053 , \3054 ,
         \3055 , \3056 , \3057 , \3058 , \3059 , \3060 , \3061 , \3062 , \3063 , \3064 ,
         \3065 , \3066 , \3067 , \3068 , \3069 , \3070 , \3071 , \3072 , \3073 , \3074 ,
         \3075 , \3076 , \3077 , \3078 , \3079 , \3080 , \3081 , \3082 , \3083 , \3084 ,
         \3085 , \3086 , \3087 , \3088 , \3089 , \3090 , \3091 , \3092 , \3093 , \3094 ,
         \3095 , \3096 , \3097 , \3098 , \3099 , \3100 , \3101 , \3102 , \3103 , \3104 ,
         \3105 , \3106 , \3107 , \3108 , \3109 , \3110 , \3111 , \3112 , \3113 , \3114 ,
         \3115 , \3116 , \3117 , \3118 , \3119 , \3120 , \3121 , \3122 , \3123 , \3124 ,
         \3125 , \3126 , \3127 , \3128 , \3129 , \3130 , \3131 , \3132 , \3133 , \3134 ,
         \3135 , \3136 , \3137 , \3138 , \3139 , \3140 , \3141 , \3142 , \3143 , \3144 ,
         \3145 , \3146 , \3147 , \3148 , \3149 , \3150 , \3151 , \3152 , \3153 , \3154 ,
         \3155 , \3156 , \3157 , \3158 , \3159 , \3160 , \3161 , \3162 , \3163 , \3164 ,
         \3165 , \3166 , \3167 , \3168 , \3169 , \3170 , \3171 , \3172 , \3173 , \3174 ,
         \3175 , \3176 , \3177 , \3178 , \3179 , \3180 , \3181 , \3182 , \3183 , \3184 ,
         \3185 , \3186 , \3187 , \3188 , \3189 , \3190 , \3191 , \3192 , \3193 , \3194 ,
         \3195 , \3196 , \3197 , \3198 , \3199 , \3200 , \3201 , \3202 , \3203 , \3204 ,
         \3205 , \3206 , \3207 , \3208 , \3209 , \3210 , \3211 , \3212 , \3213 , \3214 ,
         \3215 , \3216 , \3217 , \3218 , \3219 , \3220 , \3221 , \3222 , \3223 , \3224 ,
         \3225 , \3226 , \3227 , \3228 , \3229 , \3230 , \3231 , \3232 , \3233 , \3234 ,
         \3235 , \3236 , \3237 , \3238 , \3239 , \3240 , \3241 , \3242 , \3243 , \3244 ,
         \3245 , \3246 , \3247 , \3248 , \3249 , \3250 , \3251 , \3252 , \3253 , \3254 ,
         \3255 , \3256 , \3257 , \3258 , \3259 , \3260 , \3261 , \3262 , \3263 , \3264 ,
         \3265 , \3266 , \3267 , \3268 , \3269 , \3270 , \3271 , \3272 , \3273 , \3274 ,
         \3275 , \3276 , \3277 , \3278 , \3279 , \3280 , \3281 , \3282 , \3283 , \3284 ,
         \3285 , \3286 , \3287 , \3288 , \3289 , \3290 , \3291 , \3292 , \3293 , \3294 ,
         \3295 , \3296 , \3297 , \3298 , \3299 , \3300 , \3301 , \3302 , \3303 , \3304 ,
         \3305 , \3306 , \3307 , \3308 , \3309 , \3310 , \3311 , \3312 , \3313 , \3314 ,
         \3315 , \3316 , \3317 , \3318 , \3319 , \3320 , \3321 , \3322 , \3323 , \3324 ,
         \3325 , \3326 , \3327 , \3328 , \3329 , \3330 , \3331 , \3332 , \3333 , \3334 ,
         \3335 , \3336 , \3337 , \3338 , \3339 , \3340 , \3341 , \3342 , \3343 , \3344 ,
         \3345 , \3346 , \3347 , \3348 , \3349 , \3350 , \3351 , \3352 , \3353 , \3354 ,
         \3355 , \3356 , \3357 , \3358 , \3359 , \3360 , \3361 , \3362 , \3363 , \3364 ,
         \3365 , \3366 , \3367 , \3368 , \3369 , \3370 , \3371 , \3372 , \3373 , \3374 ,
         \3375 , \3376 , \3377 , \3378 , \3379 , \3380 , \3381 , \3382 , \3383 , \3384 ,
         \3385 , \3386 , \3387 , \3388 , \3389 , \3390 , \3391 , \3392 , \3393 , \3394 ,
         \3395 , \3396 , \3397 , \3398 , \3399 , \3400 , \3401 , \3402 , \3403 , \3404 ,
         \3405 , \3406 , \3407 , \3408 , \3409 , \3410 , \3411 , \3412 , \3413 , \3414 ,
         \3415 , \3416 , \3417 , \3418 , \3419 , \3420 , \3421 , \3422 , \3423 , \3424 ,
         \3425 , \3426 , \3427 , \3428 , \3429 , \3430 , \3431 , \3432 , \3433 , \3434 ,
         \3435 , \3436 , \3437 , \3438 , \3439 , \3440 , \3441 , \3442 , \3443 , \3444 ,
         \3445 , \3446 , \3447 , \3448 , \3449 , \3450 , \3451 , \3452 , \3453 , \3454 ,
         \3455 , \3456 , \3457 , \3458 , \3459 , \3460 , \3461 , \3462 , \3463 , \3464 ,
         \3465 , \3466 , \3467 , \3468 , \3469 , \3470 , \3471 , \3472 , \3473 , \3474 ,
         \3475 , \3476 , \3477 , \3478 , \3479 , \3480 , \3481 , \3482 , \3483 , \3484 ,
         \3485 , \3486 , \3487 , \3488 , \3489 , \3490 , \3491 , \3492 , \3493 , \3494 ,
         \3495 , \3496 , \3497 , \3498 , \3499 , \3500 , \3501 , \3502 , \3503 , \3504 ,
         \3505 , \3506 , \3507 , \3508 , \3509 , \3510 , \3511 , \3512 , \3513 , \3514 ,
         \3515 , \3516 , \3517 , \3518 , \3519 , \3520 , \3521 , \3522 , \3523 , \3524 ,
         \3525 , \3526 , \3527 , \3528 , \3529 , \3530 , \3531 , \3532 , \3533 , \3534 ,
         \3535 , \3536 , \3537 , \3538 , \3539 , \3540 , \3541 , \3542 , \3543 , \3544 ,
         \3545 , \3546 , \3547 , \3548 , \3549 , \3550 , \3551 , \3552 , \3553 , \3554 ,
         \3555 , \3556 , \3557 , \3558 , \3559 , \3560 , \3561 , \3562 , \3563 , \3564 ,
         \3565 , \3566 , \3567 , \3568 , \3569 , \3570 , \3571 , \3572 , \3573 , \3574 ,
         \3575 , \3576 , \3577 , \3578 , \3579 , \3580 , \3581 , \3582 , \3583 , \3584 ,
         \3585 , \3586 , \3587 , \3588 , \3589 , \3590 , \3591 , \3592 , \3593 , \3594 ,
         \3595 , \3596 , \3597 , \3598 , \3599 , \3600 , \3601 , \3602 , \3603 , \3604 ,
         \3605 , \3606 , \3607 , \3608 , \3609 , \3610 , \3611 , \3612 , \3613 , \3614 ,
         \3615 , \3616 , \3617 , \3618 , \3619 , \3620 , \3621 , \3622 , \3623 , \3624 ,
         \3625 , \3626 , \3627 , \3628 , \3629 , \3630 , \3631 , \3632 , \3633 , \3634 ,
         \3635 , \3636 , \3637 , \3638 , \3639 , \3640 , \3641 , \3642 , \3643 , \3644 ,
         \3645 , \3646 , \3647 , \3648 , \3649 , \3650 , \3651 , \3652 , \3653 , \3654 ,
         \3655 , \3656 , \3657 , \3658 , \3659 , \3660 , \3661 , \3662 , \3663 , \3664 ,
         \3665 , \3666 , \3667 , \3668 , \3669 , \3670 , \3671 , \3672 , \3673 , \3674 ,
         \3675 , \3676 , \3677 , \3678 , \3679 , \3680 , \3681 , \3682 , \3683 , \3684 ,
         \3685 , \3686 , \3687 , \3688 , \3689 , \3690 , \3691 , \3692 , \3693 , \3694 ,
         \3695 , \3696 , \3697 , \3698 , \3699 , \3700 , \3701 , \3702 , \3703 , \3704 ,
         \3705 , \3706 , \3707 , \3708 , \3709 , \3710 , \3711 , \3712 , \3713 , \3714 ,
         \3715 , \3716 , \3717 , \3718 , \3719 , \3720 , \3721 , \3722 , \3723 , \3724 ,
         \3725 , \3726 , \3727 , \3728 , \3729 , \3730 , \3731 , \3732 , \3733 , \3734 ,
         \3735 , \3736 , \3737 , \3738 , \3739 , \3740 , \3741 , \3742 , \3743 , \3744 ,
         \3745 , \3746 , \3747 , \3748 , \3749 , \3750 , \3751 , \3752 , \3753 , \3754 ,
         \3755 , \3756 , \3757 , \3758 , \3759 , \3760 , \3761 , \3762 , \3763 , \3764 ,
         \3765 , \3766 , \3767 , \3768 , \3769 , \3770 , \3771 , \3772 , \3773 , \3774 ,
         \3775 , \3776 , \3777 , \3778 , \3779 , \3780 , \3781 , \3782 , \3783 , \3784 ,
         \3785 , \3786 , \3787 , \3788 , \3789 , \3790 , \3791 , \3792 , \3793 , \3794 ,
         \3795 , \3796 , \3797 , \3798 , \3799 , \3800 , \3801 , \3802 , \3803 , \3804 ,
         \3805 , \3806 , \3807 , \3808 , \3809 , \3810 , \3811 , \3812 , \3813 , \3814 ,
         \3815 , \3816 , \3817 , \3818 , \3819 , \3820 , \3821 , \3822 , \3823 , \3824 ,
         \3825 , \3826 , \3827 , \3828 , \3829 , \3830 , \3831 , \3832 , \3833 , \3834 ,
         \3835 , \3836 , \3837 , \3838 , \3839 , \3840 , \3841 , \3842 , \3843 , \3844 ,
         \3845 , \3846 , \3847 , \3848 , \3849 , \3850 , \3851 , \3852 , \3853 , \3854 ,
         \3855 , \3856 , \3857 , \3858 , \3859 , \3860 , \3861 , \3862 , \3863 , \3864 ,
         \3865 , \3866 , \3867 , \3868 , \3869 , \3870 , \3871 , \3872 , \3873 , \3874 ,
         \3875 , \3876 , \3877 , \3878 , \3879 , \3880 , \3881 , \3882 , \3883 , \3884 ,
         \3885 , \3886 , \3887 , \3888 , \3889 , \3890 , \3891 , \3892 , \3893 , \3894 ,
         \3895 , \3896 , \3897 , \3898 , \3899 , \3900 , \3901 , \3902 , \3903 , \3904 ,
         \3905 , \3906 , \3907 , \3908 , \3909 , \3910 , \3911 , \3912 , \3913 , \3914 ,
         \3915 , \3916 , \3917 , \3918 , \3919 , \3920 , \3921 , \3922 , \3923 , \3924 ,
         \3925 , \3926 , \3927 , \3928 , \3929 , \3930 , \3931 , \3932 , \3933 , \3934 ,
         \3935 , \3936 , \3937 , \3938 , \3939 , \3940 , \3941 , \3942 , \3943 , \3944 ,
         \3945 , \3946 , \3947 , \3948 , \3949 , \3950 , \3951 , \3952 , \3953 , \3954 ,
         \3955 , \3956 , \3957 , \3958 , \3959 , \3960 , \3961 , \3962 , \3963 , \3964 ,
         \3965 , \3966 , \3967 , \3968 , \3969 , \3970 , \3971 , \3972 , \3973 , \3974 ,
         \3975 , \3976 , \3977 , \3978 , \3979 , \3980 , \3981 , \3982 , \3983 , \3984 ,
         \3985 , \3986 , \3987 , \3988 , \3989 , \3990 , \3991 , \3992 , \3993 , \3994 ,
         \3995 , \3996 , \3997 , \3998 , \3999 , \4000 , \4001 , \4002 , \4003 , \4004 ,
         \4005 , \4006 , \4007 , \4008 , \4009 , \4010 , \4011 , \4012 , \4013 , \4014 ,
         \4015 , \4016 , \4017 , \4018 , \4019 , \4020 , \4021 , \4022 , \4023 , \4024 ,
         \4025 , \4026 , \4027 , \4028 , \4029 , \4030 , \4031 , \4032 , \4033 , \4034 ,
         \4035 , \4036 , \4037 , \4038 , \4039 , \4040 , \4041 , \4042 , \4043 , \4044 ,
         \4045 , \4046 , \4047 , \4048 , \4049 , \4050 , \4051 , \4052 , \4053 , \4054 ,
         \4055 , \4056 , \4057 , \4058 , \4059 , \4060 , \4061 , \4062 , \4063 , \4064 ,
         \4065 , \4066 , \4067 , \4068 , \4069 , \4070 , \4071 , \4072 , \4073 , \4074 ,
         \4075 , \4076 , \4077 , \4078 , \4079 , \4080 , \4081 , \4082 , \4083 , \4084 ,
         \4085 , \4086 , \4087 , \4088 , \4089 , \4090 , \4091 , \4092 , \4093 , \4094 ,
         \4095 , \4096 , \4097 , \4098 , \4099 , \4100 , \4101 , \4102 , \4103 , \4104 ,
         \4105 , \4106 , \4107 , \4108 , \4109 , \4110 , \4111 , \4112 , \4113 , \4114 ,
         \4115 , \4116 , \4117 , \4118 , \4119 , \4120 , \4121 , \4122 , \4123 , \4124 ,
         \4125 , \4126 , \4127 , \4128 , \4129 , \4130 , \4131 , \4132 , \4133 , \4134 ,
         \4135 , \4136 , \4137 , \4138 , \4139 , \4140 , \4141 , \4142 , \4143 , \4144 ,
         \4145 , \4146 , \4147 , \4148 , \4149 , \4150 , \4151 , \4152 , \4153 , \4154 ,
         \4155 , \4156 , \4157 , \4158 , \4159 , \4160 , \4161 , \4162 , \4163 , \4164 ,
         \4165 , \4166 , \4167 , \4168 , \4169 , \4170 , \4171 , \4172 , \4173 , \4174 ,
         \4175 , \4176 , \4177 , \4178 , \4179 , \4180 , \4181 , \4182 , \4183 , \4184 ,
         \4185 , \4186 , \4187 , \4188 , \4189 , \4190 , \4191 , \4192 , \4193 , \4194 ,
         \4195 , \4196 , \4197 , \4198 , \4199 , \4200 , \4201 , \4202 , \4203 , \4204 ,
         \4205 , \4206 , \4207 , \4208 , \4209 , \4210 , \4211 , \4212 , \4213 , \4214 ,
         \4215 , \4216 , \4217 , \4218 , \4219 , \4220 , \4221 , \4222 , \4223 , \4224 ,
         \4225 , \4226 , \4227 , \4228 , \4229 , \4230 , \4231 , \4232 , \4233 , \4234 ,
         \4235 , \4236 , \4237 , \4238 , \4239 , \4240 , \4241 , \4242 , \4243 , \4244 ,
         \4245 , \4246 , \4247 , \4248 , \4249 , \4250 , \4251 , \4252 , \4253 , \4254 ,
         \4255 , \4256 , \4257 , \4258 , \4259 , \4260 , \4261 , \4262 , \4263 , \4264 ,
         \4265 , \4266 , \4267 , \4268 , \4269 , \4270 , \4271 , \4272 , \4273 , \4274 ,
         \4275 , \4276 , \4277 , \4278 , \4279 , \4280 , \4281 , \4282 , \4283 , \4284 ,
         \4285 , \4286 , \4287 , \4288 , \4289 , \4290 , \4291 , \4292 , \4293 , \4294 ,
         \4295 , \4296 , \4297 , \4298 , \4299 , \4300 , \4301 , \4302 , \4303 , \4304 ,
         \4305 , \4306 , \4307 , \4308 , \4309 , \4310 , \4311 , \4312 , \4313 , \4314 ,
         \4315 , \4316 , \4317 , \4318 , \4319 , \4320 , \4321 , \4322 , \4323 , \4324 ,
         \4325 , \4326 , \4327 , \4328 , \4329 , \4330 , \4331 , \4332 , \4333 , \4334 ,
         \4335 , \4336 , \4337 , \4338 , \4339 , \4340 , \4341 , \4342 , \4343 , \4344 ,
         \4345 , \4346 , \4347 , \4348 , \4349 , \4350 , \4351 , \4352 , \4353 , \4354 ,
         \4355 , \4356 , \4357 , \4358 , \4359 , \4360 , \4361 , \4362 , \4363 , \4364 ,
         \4365 , \4366 , \4367 , \4368 , \4369 , \4370 , \4371 , \4372 , \4373 , \4374 ,
         \4375 , \4376 , \4377 , \4378 , \4379 , \4380 , \4381 , \4382 , \4383 , \4384 ,
         \4385 , \4386 , \4387 , \4388 , \4389 , \4390 , \4391 , \4392 , \4393 , \4394 ,
         \4395 , \4396 , \4397 , \4398 , \4399 , \4400 , \4401 , \4402 , \4403 , \4404 ,
         \4405 , \4406 , \4407 , \4408 , \4409 , \4410 , \4411 , \4412 , \4413 , \4414 ,
         \4415 , \4416 , \4417 , \4418 , \4419 , \4420 , \4421 , \4422 , \4423 , \4424 ,
         \4425 , \4426 , \4427 , \4428 , \4429 , \4430 , \4431 , \4432 , \4433 , \4434 ,
         \4435 , \4436 , \4437 , \4438 , \4439 , \4440 , \4441 , \4442 , \4443 , \4444 ,
         \4445 , \4446 , \4447 , \4448 , \4449 , \4450 , \4451 , \4452 , \4453 , \4454 ,
         \4455 , \4456 , \4457 , \4458 , \4459 , \4460 , \4461 , \4462 , \4463 , \4464 ,
         \4465 , \4466 , \4467 , \4468 , \4469 , \4470 , \4471 , \4472 , \4473 , \4474 ,
         \4475 , \4476 , \4477 , \4478 , \4479 , \4480 , \4481 , \4482 , \4483 , \4484 ,
         \4485 , \4486 , \4487 , \4488 , \4489 , \4490 , \4491 , \4492 , \4493 , \4494 ,
         \4495 , \4496 , \4497 , \4498 , \4499 , \4500 , \4501 , \4502 , \4503 , \4504 ,
         \4505 , \4506 , \4507 , \4508 , \4509 , \4510 , \4511 , \4512 , \4513 , \4514 ,
         \4515 , \4516 , \4517 , \4518 , \4519 , \4520 , \4521 , \4522 , \4523 , \4524 ,
         \4525 , \4526 , \4527 , \4528 , \4529 , \4530 , \4531 , \4532 , \4533 , \4534 ,
         \4535 , \4536 , \4537 , \4538 , \4539 , \4540 , \4541 , \4542 , \4543 , \4544 ,
         \4545 , \4546 , \4547 , \4548 , \4549 , \4550 , \4551 , \4552 , \4553 , \4554 ,
         \4555 , \4556 , \4557 , \4558 , \4559 , \4560 , \4561 , \4562 , \4563 , \4564 ,
         \4565 , \4566 , \4567 , \4568 , \4569 , \4570 , \4571 , \4572 , \4573 , \4574 ,
         \4575 , \4576 , \4577 , \4578 , \4579 , \4580 , \4581 , \4582 , \4583 , \4584 ,
         \4585 , \4586 , \4587 , \4588 , \4589 , \4590 , \4591 , \4592 , \4593 , \4594 ,
         \4595 , \4596 , \4597 , \4598 , \4599 , \4600 , \4601 , \4602 , \4603 , \4604 ,
         \4605 , \4606 , \4607 , \4608 , \4609 , \4610 , \4611 , \4612 , \4613 , \4614 ,
         \4615 , \4616 , \4617 , \4618 , \4619 , \4620 , \4621 , \4622 , \4623 , \4624 ,
         \4625 , \4626 , \4627 , \4628 , \4629 , \4630 , \4631 , \4632 , \4633 , \4634 ,
         \4635 , \4636 , \4637 , \4638 , \4639 , \4640 , \4641 , \4642 , \4643 , \4644 ,
         \4645 , \4646 , \4647 , \4648 , \4649 , \4650 , \4651 , \4652 , \4653 , \4654 ,
         \4655 , \4656 , \4657 , \4658 , \4659 , \4660 , \4661 , \4662 , \4663 , \4664 ,
         \4665 , \4666 , \4667 , \4668 , \4669 , \4670 , \4671 , \4672 , \4673 , \4674 ,
         \4675 , \4676 , \4677 , \4678 , \4679 , \4680 , \4681 , \4682 , \4683 , \4684 ,
         \4685 , \4686 , \4687 , \4688 , \4689 , \4690 , \4691 , \4692 , \4693 , \4694 ,
         \4695 , \4696 , \4697 , \4698 , \4699 , \4700 , \4701 , \4702 , \4703 , \4704 ,
         \4705 , \4706 , \4707 , \4708 , \4709 , \4710 , \4711 , \4712 , \4713 , \4714 ,
         \4715 , \4716 , \4717 , \4718 , \4719 , \4720 , \4721 , \4722 , \4723 , \4724 ,
         \4725 , \4726 , \4727 , \4728 , \4729 , \4730 , \4731 , \4732 , \4733 , \4734 ,
         \4735 , \4736 , \4737 , \4738 , \4739 , \4740 , \4741 , \4742 , \4743 , \4744 ,
         \4745 , \4746 , \4747 , \4748 , \4749 , \4750 , \4751 , \4752 , \4753 , \4754 ,
         \4755 , \4756 , \4757 , \4758 , \4759 , \4760 , \4761 , \4762 , \4763 , \4764 ,
         \4765 , \4766 , \4767 , \4768 , \4769 , \4770 , \4771 , \4772 , \4773 , \4774 ,
         \4775 , \4776 , \4777 , \4778 , \4779 , \4780 , \4781 , \4782 , \4783 , \4784 ,
         \4785 , \4786 , \4787 , \4788 , \4789 , \4790 , \4791 , \4792 , \4793 , \4794 ,
         \4795 , \4796 , \4797 , \4798 , \4799 , \4800 , \4801 , \4802 , \4803 , \4804 ,
         \4805 , \4806 , \4807 , \4808 , \4809 , \4810 , \4811 , \4812 , \4813 , \4814 ,
         \4815 , \4816 , \4817 , \4818 , \4819 , \4820 , \4821 , \4822 , \4823 , \4824 ,
         \4825 , \4826 , \4827 , \4828 , \4829 , \4830 , \4831 , \4832 , \4833 , \4834 ,
         \4835 , \4836 , \4837 , \4838 , \4839 , \4840 , \4841 , \4842 , \4843 , \4844 ,
         \4845 , \4846 , \4847 , \4848 , \4849 , \4850 , \4851 , \4852 , \4853 , \4854 ,
         \4855 , \4856 , \4857 , \4858 , \4859 , \4860 , \4861 , \4862 , \4863 , \4864 ,
         \4865 , \4866 , \4867 , \4868 , \4869 , \4870 , \4871 , \4872 , \4873 , \4874 ,
         \4875 , \4876 , \4877 , \4878 , \4879 , \4880 , \4881 , \4882 , \4883 , \4884 ,
         \4885 , \4886 , \4887 , \4888 , \4889 , \4890 , \4891 , \4892 , \4893 , \4894 ,
         \4895 , \4896 , \4897 , \4898 , \4899 , \4900 , \4901 , \4902 , \4903 , \4904 ,
         \4905 , \4906 , \4907 , \4908 , \4909 , \4910 , \4911 , \4912 , \4913 , \4914 ,
         \4915 , \4916 , \4917 , \4918 , \4919 , \4920 , \4921 , \4922 , \4923 , \4924 ,
         \4925 , \4926 , \4927 , \4928 , \4929 , \4930 , \4931 , \4932 , \4933 , \4934 ,
         \4935 , \4936 , \4937 , \4938 , \4939 , \4940 , \4941 , \4942 , \4943 , \4944 ,
         \4945 , \4946 , \4947 , \4948 , \4949 , \4950 , \4951 , \4952 , \4953 , \4954 ,
         \4955 , \4956 , \4957 , \4958 , \4959 , \4960 , \4961 , \4962 , \4963 , \4964 ,
         \4965 , \4966 , \4967 , \4968 , \4969 , \4970 , \4971 , \4972 , \4973 , \4974 ,
         \4975 , \4976 , \4977 , \4978 , \4979 , \4980 , \4981 , \4982 , \4983 , \4984 ,
         \4985 , \4986 , \4987 , \4988 , \4989 , \4990 , \4991 , \4992 , \4993 , \4994 ,
         \4995 , \4996 , \4997 , \4998 , \4999 , \5000 , \5001 , \5002 , \5003 , \5004 ,
         \5005 , \5006 , \5007 , \5008 , \5009 , \5010 , \5011 , \5012 , \5013 , \5014 ,
         \5015 , \5016 , \5017 , \5018 , \5019 , \5020 , \5021 , \5022 , \5023 , \5024 ,
         \5025 , \5026 , \5027 , \5028 , \5029 , \5030 , \5031 , \5032 , \5033 , \5034 ,
         \5035 , \5036 , \5037 , \5038 , \5039 , \5040 , \5041 , \5042 , \5043 , \5044 ,
         \5045 , \5046 , \5047 , \5048 , \5049 , \5050 , \5051 , \5052 , \5053 , \5054 ,
         \5055 , \5056 , \5057 , \5058 , \5059 , \5060 , \5061 , \5062 , \5063 , \5064 ,
         \5065 , \5066 , \5067 , \5068 , \5069 , \5070 , \5071 , \5072 , \5073 , \5074 ,
         \5075 , \5076 , \5077 , \5078 , \5079 , \5080 , \5081 , \5082 , \5083 , \5084 ,
         \5085 , \5086 , \5087 , \5088 , \5089 , \5090 , \5091 , \5092 , \5093 , \5094 ,
         \5095 , \5096 , \5097 , \5098 , \5099 , \5100 , \5101 , \5102 , \5103 , \5104 ,
         \5105 , \5106 , \5107 , \5108 , \5109 , \5110 , \5111 , \5112 , \5113 , \5114 ,
         \5115 , \5116 , \5117 , \5118 , \5119 , \5120 , \5121 , \5122 , \5123 , \5124 ,
         \5125 , \5126 , \5127 , \5128 , \5129 , \5130 , \5131 , \5132 , \5133 , \5134 ,
         \5135 , \5136 , \5137 , \5138 , \5139 , \5140 , \5141 , \5142 , \5143 , \5144 ,
         \5145 , \5146 , \5147 , \5148 , \5149 , \5150 , \5151 , \5152 , \5153 , \5154 ,
         \5155 , \5156 , \5157 , \5158 , \5159 , \5160 , \5161 , \5162 , \5163 , \5164 ,
         \5165 , \5166 , \5167 , \5168 , \5169 , \5170 , \5171 , \5172 , \5173 , \5174 ,
         \5175 , \5176 , \5177 , \5178 , \5179 , \5180 , \5181 , \5182 , \5183 , \5184 ,
         \5185 , \5186 , \5187 , \5188 , \5189 , \5190 , \5191 , \5192 , \5193 , \5194 ,
         \5195 , \5196 , \5197 , \5198 , \5199 , \5200 , \5201 , \5202 , \5203 , \5204 ,
         \5205 , \5206 , \5207 , \5208 , \5209 , \5210 , \5211 , \5212 , \5213 , \5214 ,
         \5215 , \5216 , \5217 , \5218 , \5219 , \5220 , \5221 , \5222 , \5223 , \5224 ,
         \5225 , \5226 , \5227 , \5228 , \5229 , \5230 , \5231 , \5232 , \5233 , \5234 ,
         \5235 , \5236 , \5237 , \5238 , \5239 , \5240 , \5241 , \5242 , \5243 , \5244 ,
         \5245 , \5246 , \5247 , \5248 , \5249 , \5250 , \5251 , \5252 , \5253 , \5254 ,
         \5255 , \5256 , \5257 , \5258 , \5259 , \5260 , \5261 , \5262 , \5263 , \5264 ,
         \5265 , \5266 , \5267 , \5268 , \5269 , \5270 , \5271 , \5272 , \5273 , \5274 ,
         \5275 , \5276 , \5277 , \5278 , \5279 , \5280 , \5281 , \5282 , \5283 , \5284 ,
         \5285 , \5286 , \5287 , \5288 , \5289 , \5290 , \5291 , \5292 , \5293 , \5294 ,
         \5295 , \5296 , \5297 , \5298 , \5299 , \5300 , \5301 , \5302 , \5303 , \5304 ,
         \5305 , \5306 , \5307 , \5308 , \5309 , \5310 , \5311 , \5312 , \5313 , \5314 ,
         \5315 , \5316 , \5317 , \5318 , \5319 , \5320 , \5321 , \5322 , \5323 , \5324 ,
         \5325 , \5326 , \5327 , \5328 , \5329 , \5330 , \5331 , \5332 , \5333 , \5334 ,
         \5335 , \5336 , \5337 , \5338 , \5339 , \5340 , \5341 , \5342 , \5343 , \5344 ,
         \5345 , \5346 , \5347 , \5348 , \5349 , \5350 , \5351 , \5352 , \5353 , \5354 ,
         \5355 , \5356 , \5357 , \5358 , \5359 , \5360 , \5361 , \5362 , \5363 , \5364 ,
         \5365 , \5366 , \5367 , \5368 , \5369 , \5370 , \5371 , \5372 , \5373 , \5374 ,
         \5375 , \5376 , \5377 , \5378 , \5379 , \5380 , \5381 , \5382 , \5383 , \5384 ,
         \5385 , \5386 , \5387 , \5388 , \5389 , \5390 , \5391 , \5392 , \5393 , \5394 ,
         \5395 , \5396 , \5397 , \5398 , \5399 , \5400 , \5401 , \5402 , \5403 , \5404 ,
         \5405 , \5406 , \5407 , \5408 , \5409 , \5410 , \5411 , \5412 , \5413 , \5414 ,
         \5415 , \5416 , \5417 , \5418 , \5419 , \5420 , \5421 , \5422 , \5423 , \5424 ,
         \5425 , \5426 , \5427 , \5428 , \5429 , \5430 , \5431 , \5432 , \5433 , \5434 ,
         \5435 , \5436 , \5437 , \5438 , \5439 , \5440 , \5441 , \5442 , \5443 , \5444 ,
         \5445 , \5446 , \5447 , \5448 , \5449 , \5450 , \5451 , \5452 , \5453 , \5454 ,
         \5455 , \5456 , \5457 , \5458 , \5459 , \5460 , \5461 , \5462 , \5463 , \5464 ,
         \5465 , \5466 , \5467 , \5468 , \5469 , \5470 , \5471 , \5472 , \5473 , \5474 ,
         \5475 , \5476 , \5477 , \5478 , \5479 , \5480 , \5481 , \5482 , \5483 , \5484 ,
         \5485 , \5486 , \5487 , \5488 , \5489 , \5490 , \5491 , \5492 , \5493 , \5494 ,
         \5495 , \5496 , \5497 , \5498 , \5499 , \5500 , \5501 , \5502 , \5503 , \5504 ,
         \5505 , \5506 , \5507 , \5508 , \5509 , \5510 , \5511 , \5512 , \5513 , \5514 ,
         \5515 , \5516 , \5517 , \5518 , \5519 , \5520 , \5521 , \5522 , \5523 , \5524 ,
         \5525 , \5526 , \5527 , \5528 , \5529 , \5530 , \5531 , \5532 , \5533 , \5534 ,
         \5535 , \5536 , \5537 , \5538 , \5539 , \5540 , \5541 , \5542 , \5543 , \5544 ,
         \5545 , \5546 , \5547 , \5548 , \5549 , \5550 , \5551 , \5552 , \5553 , \5554 ,
         \5555 , \5556 , \5557 , \5558 , \5559 , \5560 , \5561 , \5562 , \5563 , \5564 ,
         \5565 , \5566 , \5567 , \5568 , \5569 , \5570 , \5571 , \5572 , \5573 , \5574 ,
         \5575 , \5576 , \5577 , \5578 , \5579 , \5580 , \5581 , \5582 , \5583 , \5584 ,
         \5585 , \5586 , \5587 , \5588 , \5589 , \5590 , \5591 , \5592 , \5593 , \5594 ,
         \5595 , \5596 , \5597 , \5598 , \5599 , \5600 , \5601 , \5602 , \5603 , \5604 ,
         \5605 , \5606 , \5607 , \5608 , \5609 , \5610 , \5611 , \5612 , \5613 , \5614 ,
         \5615 , \5616 , \5617 , \5618 , \5619 , \5620 , \5621 , \5622 , \5623 , \5624 ,
         \5625 , \5626 , \5627 , \5628 , \5629 , \5630 , \5631 , \5632 , \5633 , \5634 ,
         \5635 , \5636 , \5637 , \5638 , \5639 , \5640 , \5641 , \5642 , \5643 , \5644 ,
         \5645 , \5646 , \5647 , \5648 , \5649 , \5650 , \5651 , \5652 , \5653 , \5654 ,
         \5655 , \5656 , \5657 , \5658 , \5659 , \5660 , \5661 , \5662 , \5663 , \5664 ,
         \5665 , \5666 , \5667 , \5668 , \5669 , \5670 , \5671 , \5672 , \5673 , \5674 ,
         \5675 , \5676 , \5677 , \5678 , \5679 , \5680 , \5681 , \5682 , \5683 , \5684 ,
         \5685 , \5686 , \5687 , \5688 , \5689 , \5690 , \5691 , \5692 , \5693 , \5694 ,
         \5695 , \5696 , \5697 , \5698 , \5699 , \5700 , \5701 , \5702 , \5703 , \5704 ,
         \5705 , \5706 , \5707 , \5708 , \5709 , \5710 , \5711 , \5712 , \5713 , \5714 ,
         \5715 , \5716 , \5717 , \5718 , \5719 , \5720 , \5721 , \5722 , \5723 , \5724 ,
         \5725 , \5726 , \5727 , \5728 , \5729 , \5730 , \5731 , \5732 , \5733 , \5734 ,
         \5735 , \5736 , \5737 , \5738 , \5739 , \5740 , \5741 , \5742 , \5743 , \5744 ,
         \5745 , \5746 , \5747 , \5748 , \5749 , \5750 , \5751 , \5752 , \5753 , \5754 ,
         \5755 , \5756 , \5757 , \5758 , \5759 , \5760 , \5761 , \5762 , \5763 , \5764 ,
         \5765 , \5766 , \5767 , \5768 , \5769 , \5770 , \5771 , \5772 , \5773 , \5774 ,
         \5775 , \5776 , \5777 , \5778 , \5779 , \5780 , \5781 , \5782 , \5783 , \5784 ,
         \5785 , \5786 , \5787 , \5788 , \5789 , \5790 , \5791 , \5792 , \5793 , \5794 ,
         \5795 , \5796 , \5797 , \5798 , \5799 , \5800 , \5801 , \5802 , \5803 , \5804 ,
         \5805 , \5806 , \5807 , \5808 , \5809 , \5810 , \5811 , \5812 , \5813 , \5814 ,
         \5815 , \5816 , \5817 , \5818 , \5819 , \5820 , \5821 , \5822 , \5823 , \5824 ,
         \5825 , \5826 , \5827 , \5828 , \5829 , \5830 , \5831 , \5832 , \5833 , \5834 ,
         \5835 , \5836 , \5837 , \5838 , \5839 , \5840 , \5841 , \5842 , \5843 , \5844 ,
         \5845 , \5846 , \5847 , \5848 , \5849 , \5850 , \5851 , \5852 , \5853 , \5854 ,
         \5855 , \5856 , \5857 , \5858 , \5859 , \5860 , \5861 , \5862 , \5863 , \5864 ,
         \5865 , \5866 , \5867 , \5868 , \5869 , \5870 , \5871 , \5872 , \5873 , \5874 ,
         \5875 , \5876 , \5877 , \5878 , \5879 , \5880 , \5881 , \5882 , \5883 , \5884 ,
         \5885 , \5886 , \5887 , \5888 , \5889 , \5890 , \5891 , \5892 , \5893 , \5894 ,
         \5895 , \5896 , \5897 , \5898 , \5899 , \5900 , \5901 , \5902 , \5903 , \5904 ,
         \5905 , \5906 , \5907 , \5908 , \5909 , \5910 , \5911 , \5912 , \5913 , \5914 ,
         \5915 , \5916 , \5917 , \5918 , \5919 , \5920 , \5921 , \5922 , \5923 , \5924 ,
         \5925 , \5926 , \5927 , \5928 , \5929 , \5930 , \5931 , \5932 , \5933 , \5934 ,
         \5935 , \5936 , \5937 , \5938 , \5939 , \5940 , \5941 , \5942 , \5943 , \5944 ,
         \5945 , \5946 , \5947 , \5948 , \5949 , \5950 , \5951 , \5952 , \5953 , \5954 ,
         \5955 , \5956 , \5957 , \5958 , \5959 , \5960 , \5961 , \5962 , \5963 , \5964 ,
         \5965 , \5966 , \5967 , \5968 , \5969 , \5970 , \5971 , \5972 , \5973 , \5974 ,
         \5975 , \5976 , \5977 , \5978 , \5979 , \5980 , \5981 , \5982 , \5983 , \5984 ,
         \5985 , \5986 , \5987 , \5988 , \5989 , \5990 , \5991 , \5992 , \5993 , \5994 ,
         \5995 , \5996 , \5997 , \5998 , \5999 , \6000 , \6001 , \6002 , \6003 , \6004 ,
         \6005 , \6006 , \6007 , \6008 , \6009 , \6010 , \6011 , \6012 , \6013 , \6014 ,
         \6015 , \6016 , \6017 , \6018 , \6019 , \6020 , \6021 , \6022 , \6023 , \6024 ,
         \6025 , \6026 , \6027 , \6028 , \6029 , \6030 , \6031 , \6032 , \6033 , \6034 ,
         \6035 , \6036 , \6037 , \6038 , \6039 , \6040 , \6041 , \6042 , \6043 , \6044 ,
         \6045 , \6046 , \6047 , \6048 , \6049 , \6050 , \6051 , \6052 , \6053 , \6054 ,
         \6055 , \6056 , \6057 , \6058 , \6059 , \6060 , \6061 , \6062 , \6063 , \6064 ,
         \6065 , \6066 , \6067 , \6068 , \6069 , \6070 , \6071 , \6072 , \6073 , \6074 ,
         \6075 , \6076 , \6077 , \6078 , \6079 , \6080 , \6081 , \6082 , \6083 , \6084 ,
         \6085 , \6086 , \6087 , \6088 , \6089 , \6090 , \6091 , \6092 , \6093 , \6094 ,
         \6095 , \6096 , \6097 , \6098 , \6099 , \6100 , \6101 , \6102 , \6103 , \6104 ,
         \6105 , \6106 , \6107 , \6108 , \6109 , \6110 , \6111 , \6112 , \6113 , \6114 ,
         \6115 , \6116 , \6117 , \6118 , \6119 , \6120 , \6121 , \6122 , \6123 , \6124 ,
         \6125 , \6126 , \6127 , \6128 , \6129 , \6130 , \6131 , \6132 , \6133 , \6134 ,
         \6135 , \6136 , \6137 , \6138 , \6139 , \6140 , \6141 , \6142 , \6143 , \6144 ,
         \6145 , \6146 , \6147 , \6148 , \6149 , \6150 , \6151 , \6152 , \6153 , \6154 ,
         \6155 , \6156 , \6157 , \6158 , \6159 , \6160 , \6161 , \6162 , \6163 , \6164 ,
         \6165 , \6166 , \6167 , \6168 , \6169 , \6170 , \6171 , \6172 , \6173 , \6174 ,
         \6175 , \6176 , \6177 , \6178 , \6179 , \6180 , \6181 , \6182 , \6183 , \6184 ,
         \6185 , \6186 , \6187 , \6188 , \6189 , \6190 , \6191 , \6192 , \6193 , \6194 ,
         \6195 , \6196 , \6197 , \6198 , \6199 , \6200 , \6201 , \6202 , \6203 , \6204 ,
         \6205 , \6206 , \6207 , \6208 , \6209 , \6210 , \6211 , \6212 , \6213 , \6214 ,
         \6215 , \6216 , \6217 , \6218 , \6219 , \6220 , \6221 , \6222 , \6223 , \6224 ,
         \6225 , \6226 , \6227 , \6228 , \6229 , \6230 , \6231 , \6232 , \6233 , \6234 ,
         \6235 , \6236 , \6237 , \6238 , \6239 , \6240 , \6241 , \6242 , \6243 , \6244 ,
         \6245 , \6246 , \6247 , \6248 , \6249 , \6250 , \6251 , \6252 , \6253 , \6254 ,
         \6255 , \6256 , \6257 , \6258 , \6259 , \6260 , \6261 , \6262 , \6263 , \6264 ,
         \6265 , \6266 , \6267 , \6268 , \6269 , \6270 , \6271 , \6272 , \6273 , \6274 ,
         \6275 , \6276 , \6277 , \6278 , \6279 , \6280 , \6281 , \6282 , \6283 , \6284 ,
         \6285 , \6286 , \6287 , \6288 , \6289 , \6290 , \6291 , \6292 , \6293 , \6294 ,
         \6295 , \6296 , \6297 , \6298 , \6299 , \6300 , \6301 , \6302 , \6303 , \6304 ,
         \6305 , \6306 , \6307 , \6308 , \6309 , \6310 , \6311 , \6312 , \6313 , \6314 ,
         \6315 , \6316 , \6317 , \6318 , \6319 , \6320 , \6321 , \6322 , \6323 , \6324 ,
         \6325 , \6326 , \6327 , \6328 , \6329 , \6330 , \6331 , \6332 , \6333 , \6334 ,
         \6335 , \6336 , \6337 , \6338 , \6339 , \6340 , \6341 , \6342 , \6343 , \6344 ,
         \6345 , \6346 , \6347 , \6348 , \6349 , \6350 , \6351 , \6352 , \6353 , \6354 ,
         \6355 , \6356 , \6357 , \6358 , \6359 , \6360 , \6361 , \6362 , \6363 , \6364 ,
         \6365 , \6366 , \6367 , \6368 , \6369 , \6370 , \6371 , \6372 , \6373 , \6374 ,
         \6375 , \6376 , \6377 , \6378 , \6379 , \6380 , \6381 , \6382 , \6383 , \6384 ,
         \6385 , \6386 , \6387 , \6388 , \6389 , \6390 , \6391 , \6392 , \6393 , \6394 ,
         \6395 , \6396 , \6397 , \6398 , \6399 , \6400 , \6401 , \6402 , \6403 , \6404 ,
         \6405 , \6406 , \6407 , \6408 , \6409 , \6410 , \6411 , \6412 , \6413 , \6414 ,
         \6415 , \6416 , \6417 , \6418 , \6419 , \6420 , \6421 , \6422 , \6423 , \6424 ,
         \6425 , \6426 , \6427 , \6428 , \6429 , \6430 , \6431 , \6432 , \6433 , \6434 ,
         \6435 , \6436 , \6437 , \6438 , \6439 , \6440 , \6441 , \6442 , \6443 , \6444 ,
         \6445 , \6446 , \6447 , \6448 , \6449 , \6450 , \6451 , \6452 , \6453 , \6454 ,
         \6455 , \6456 , \6457 , \6458 , \6459 , \6460 , \6461 , \6462 , \6463 , \6464 ,
         \6465 , \6466 , \6467 , \6468 , \6469 , \6470 , \6471 , \6472 , \6473 , \6474 ,
         \6475 , \6476 , \6477 , \6478 , \6479 , \6480 , \6481 , \6482 , \6483 , \6484 ,
         \6485 , \6486 , \6487 , \6488 , \6489 , \6490 , \6491 , \6492 , \6493 , \6494 ,
         \6495 , \6496 , \6497 , \6498 , \6499 , \6500 , \6501 , \6502 , \6503 , \6504 ,
         \6505 , \6506 , \6507 , \6508 , \6509 , \6510 , \6511 , \6512 , \6513 , \6514 ,
         \6515 , \6516 , \6517 , \6518 , \6519 , \6520 , \6521 , \6522 , \6523 , \6524 ,
         \6525 , \6526 , \6527 , \6528 , \6529 , \6530 , \6531 , \6532 , \6533 , \6534 ,
         \6535 , \6536 , \6537 , \6538 , \6539 , \6540 , \6541 , \6542 , \6543 , \6544 ,
         \6545 , \6546 , \6547 , \6548 , \6549 , \6550 , \6551 , \6552 , \6553 , \6554 ,
         \6555 , \6556 , \6557 , \6558 , \6559 , \6560 , \6561 , \6562 , \6563 , \6564 ,
         \6565 , \6566 , \6567 , \6568 , \6569 , \6570 , \6571 , \6572 , \6573 , \6574 ,
         \6575 , \6576 , \6577 , \6578 , \6579 , \6580 , \6581 , \6582 , \6583 , \6584 ,
         \6585 , \6586 , \6587 , \6588 , \6589 , \6590 , \6591 , \6592 , \6593 , \6594 ,
         \6595 , \6596 , \6597 , \6598 , \6599 , \6600 , \6601 , \6602 , \6603 , \6604 ,
         \6605 , \6606 , \6607 , \6608 , \6609 , \6610 , \6611 , \6612 , \6613 , \6614 ,
         \6615 , \6616 , \6617 , \6618 , \6619 , \6620 , \6621 , \6622 , \6623 , \6624 ,
         \6625 , \6626 , \6627 , \6628 , \6629 , \6630 , \6631 , \6632 , \6633 , \6634 ,
         \6635 , \6636 , \6637 , \6638 , \6639 , \6640 , \6641 , \6642 , \6643 , \6644 ,
         \6645 , \6646 , \6647 , \6648 , \6649 , \6650 , \6651 , \6652 , \6653 , \6654 ,
         \6655 , \6656 , \6657 , \6658 , \6659 , \6660 , \6661 , \6662 , \6663 , \6664 ,
         \6665 , \6666 , \6667 , \6668 , \6669 , \6670 , \6671 , \6672 , \6673 , \6674 ,
         \6675 , \6676 , \6677 , \6678 , \6679 , \6680 , \6681 , \6682 , \6683 , \6684 ,
         \6685 , \6686 , \6687 , \6688 , \6689 , \6690 , \6691 , \6692 , \6693 , \6694 ,
         \6695 , \6696 , \6697 , \6698 , \6699 , \6700 , \6701 , \6702 , \6703 , \6704 ,
         \6705 , \6706 , \6707 , \6708 , \6709 , \6710 , \6711 , \6712 , \6713 , \6714 ,
         \6715 , \6716 , \6717 , \6718 , \6719 , \6720 , \6721 , \6722 , \6723 , \6724 ,
         \6725 , \6726 , \6727 , \6728 , \6729 , \6730 , \6731 , \6732 , \6733 , \6734 ,
         \6735 , \6736 , \6737 , \6738 , \6739 , \6740 , \6741 , \6742 , \6743 , \6744 ,
         \6745 , \6746 , \6747 , \6748 , \6749 , \6750 , \6751 , \6752 , \6753 , \6754 ,
         \6755 , \6756 , \6757 , \6758 , \6759 , \6760 , \6761 , \6762 , \6763 , \6764 ,
         \6765 , \6766 , \6767 , \6768 , \6769 , \6770 , \6771 , \6772 , \6773 , \6774 ,
         \6775 , \6776 , \6777 , \6778 , \6779 , \6780 , \6781 , \6782 , \6783 , \6784 ,
         \6785 , \6786 , \6787 , \6788 , \6789 , \6790 , \6791 , \6792 , \6793 , \6794 ,
         \6795 , \6796 , \6797 , \6798 , \6799 , \6800 , \6801 , \6802 , \6803 , \6804 ,
         \6805 , \6806 , \6807 , \6808 , \6809 , \6810 , \6811 , \6812 , \6813 , \6814 ,
         \6815 , \6816 , \6817 , \6818 , \6819 , \6820 , \6821 , \6822 , \6823 , \6824 ,
         \6825 , \6826 , \6827 , \6828 , \6829 , \6830 , \6831 , \6832 , \6833 , \6834 ,
         \6835 , \6836 , \6837 , \6838 , \6839 , \6840 , \6841 , \6842 , \6843 , \6844 ,
         \6845 , \6846 , \6847 , \6848 , \6849 , \6850 , \6851 , \6852 , \6853 , \6854 ,
         \6855 , \6856 , \6857 , \6858 , \6859 , \6860 , \6861 , \6862 , \6863 , \6864 ,
         \6865 , \6866 , \6867 , \6868 , \6869 , \6870 , \6871 , \6872 , \6873 , \6874 ,
         \6875 , \6876 , \6877 , \6878 , \6879 , \6880 , \6881 , \6882 , \6883 , \6884 ,
         \6885 , \6886 , \6887 , \6888 , \6889 , \6890 , \6891 , \6892 , \6893 , \6894 ,
         \6895 , \6896 , \6897 , \6898 , \6899 , \6900 , \6901 , \6902 , \6903 , \6904 ,
         \6905 , \6906 , \6907 , \6908 , \6909 , \6910 , \6911 , \6912 , \6913 , \6914 ,
         \6915 , \6916 , \6917 , \6918 , \6919 , \6920 , \6921 , \6922 , \6923 , \6924 ,
         \6925 , \6926 , \6927 , \6928 , \6929 , \6930 , \6931 , \6932 , \6933 , \6934 ,
         \6935 , \6936 , \6937 , \6938 , \6939 , \6940 , \6941 , \6942 , \6943 , \6944 ,
         \6945 , \6946 , \6947 , \6948 , \6949 , \6950 , \6951 , \6952 , \6953 , \6954 ,
         \6955 , \6956 , \6957 , \6958 , \6959 , \6960 , \6961 , \6962 , \6963 , \6964 ,
         \6965 , \6966 , \6967 , \6968 , \6969 , \6970 , \6971 , \6972 , \6973 , \6974 ,
         \6975 , \6976 , \6977 , \6978 , \6979 , \6980 , \6981 , \6982 , \6983 , \6984 ,
         \6985 , \6986 , \6987 , \6988 , \6989 , \6990 , \6991 , \6992 , \6993 , \6994 ,
         \6995 , \6996 , \6997 , \6998 , \6999 , \7000 , \7001 , \7002 , \7003 , \7004 ,
         \7005 , \7006 , \7007 , \7008 , \7009 , \7010 , \7011 , \7012 , \7013 , \7014 ,
         \7015 , \7016 , \7017 , \7018 , \7019 , \7020 , \7021 , \7022 , \7023 , \7024 ,
         \7025 , \7026 , \7027 , \7028 , \7029 , \7030 , \7031 , \7032 , \7033 , \7034 ,
         \7035 , \7036 , \7037 , \7038 , \7039 , \7040 , \7041 , \7042 , \7043 , \7044 ,
         \7045 , \7046 , \7047 , \7048 , \7049 , \7050 , \7051 , \7052 , \7053 , \7054 ,
         \7055 , \7056 , \7057 , \7058 , \7059 , \7060 , \7061 , \7062 , \7063 , \7064 ,
         \7065 , \7066 , \7067 , \7068 , \7069 , \7070 , \7071 , \7072 , \7073 , \7074 ,
         \7075 , \7076 , \7077 , \7078 , \7079 , \7080 , \7081 , \7082 , \7083 , \7084 ,
         \7085 , \7086 , \7087 , \7088 , \7089 , \7090 , \7091 , \7092 , \7093 , \7094 ,
         \7095 , \7096 , \7097 , \7098 , \7099 , \7100 , \7101 , \7102 , \7103 , \7104 ,
         \7105 , \7106 , \7107 , \7108 , \7109 , \7110 , \7111 , \7112 , \7113 , \7114 ,
         \7115 , \7116 , \7117 , \7118 , \7119 , \7120 , \7121 , \7122 , \7123 , \7124 ,
         \7125 , \7126 , \7127 , \7128 , \7129 , \7130 , \7131 , \7132 , \7133 , \7134 ,
         \7135 , \7136 , \7137 , \7138 , \7139 , \7140 , \7141 , \7142 , \7143 , \7144 ,
         \7145 , \7146 , \7147 , \7148 , \7149 , \7150 , \7151 , \7152 , \7153 , \7154 ,
         \7155 , \7156 , \7157 , \7158 , \7159 , \7160 , \7161 , \7162 , \7163 , \7164 ,
         \7165 , \7166 , \7167 , \7168 , \7169 , \7170 , \7171 , \7172 , \7173 , \7174 ,
         \7175 , \7176 , \7177 , \7178 , \7179 , \7180 , \7181 , \7182 , \7183 , \7184 ,
         \7185 , \7186 , \7187 , \7188 , \7189 , \7190 , \7191 , \7192 , \7193 , \7194 ,
         \7195 , \7196 , \7197 , \7198 , \7199 , \7200 , \7201 , \7202 , \7203 , \7204 ,
         \7205 , \7206 , \7207 , \7208 , \7209 , \7210 , \7211 , \7212 , \7213 , \7214 ,
         \7215 , \7216 , \7217 , \7218 , \7219 , \7220 , \7221 , \7222 , \7223 , \7224 ,
         \7225 , \7226 , \7227 , \7228 , \7229 , \7230 , \7231 , \7232 , \7233 , \7234 ,
         \7235 , \7236 , \7237 , \7238 , \7239 , \7240 , \7241 , \7242 , \7243 , \7244 ,
         \7245 , \7246 , \7247 , \7248 , \7249 , \7250 , \7251 , \7252 , \7253 , \7254 ,
         \7255 , \7256 , \7257 , \7258 , \7259 , \7260 , \7261 , \7262 , \7263 , \7264 ,
         \7265 , \7266 , \7267 , \7268 , \7269 , \7270 , \7271 , \7272 , \7273 , \7274 ,
         \7275 , \7276 , \7277 , \7278 , \7279 , \7280 , \7281 , \7282 , \7283 , \7284 ,
         \7285 , \7286 , \7287 , \7288 , \7289 , \7290 , \7291 , \7292 , \7293 , \7294 ,
         \7295 , \7296 , \7297 , \7298 , \7299 , \7300 , \7301 , \7302 , \7303 , \7304 ,
         \7305 , \7306 , \7307 , \7308 , \7309 , \7310 , \7311 , \7312 , \7313 , \7314 ,
         \7315 , \7316 , \7317 , \7318 , \7319 , \7320 ;
buf \U$labaj754 ( R_61_7d2b4e8, \6298 );
buf \U$labaj755 ( R_62_7d2b590, \6480 );
buf \U$labaj756 ( R_63_7d2b638, \6570 );
buf \U$labaj757 ( R_64_7d2b6e0, \6661 );
buf \U$labaj758 ( R_65_7d2b788, \6706 );
buf \U$labaj759 ( R_66_7d2b830, \6751 );
buf \U$labaj760 ( R_67_7d2b8d8, \6794 );
buf \U$labaj761 ( R_68_7d2b980, \6837 );
buf \U$labaj762 ( R_69_7d2ba28, \6860 );
buf \U$labaj763 ( R_6a_7d2bad0, \6883 );
buf \U$labaj764 ( R_6b_7d2bb78, \6905 );
buf \U$labaj765 ( R_6c_7d2bc20, \6927 );
buf \U$labaj766 ( R_6d_7d2bcc8, \6949 );
buf \U$labaj767 ( R_6e_7d2bd70, \6971 );
buf \U$labaj768 ( R_6f_7d2be18, \6991 );
buf \U$labaj769 ( R_70_7d2bec0, \7011 );
buf \U$labaj770 ( R_71_7d2bf68, \7023 );
buf \U$labaj771 ( R_72_7d2c010, \7035 );
buf \U$labaj772 ( R_73_7d2c0b8, \7047 );
buf \U$labaj773 ( R_74_7d2c160, \7059 );
buf \U$labaj774 ( R_75_7d2c208, \7071 );
buf \U$labaj775 ( R_76_7d2c2b0, \7083 );
buf \U$labaj776 ( R_77_7d2c358, \7094 );
buf \U$labaj777 ( R_78_7d2c400, \7105 );
buf \U$labaj778 ( R_79_7d2c4a8, \7116 );
buf \U$labaj779 ( R_7a_7d2c550, \7127 );
buf \U$labaj780 ( R_7b_7d2c5f8, \7138 );
buf \U$labaj781 ( R_7c_7d2c6a0, \7149 );
buf \U$labaj782 ( R_7d_7d2c748, \7160 );
buf \U$labaj783 ( R_7e_7d2c7f0, \7171 );
buf \U$labaj784 ( R_7f_7d2c898, \7178 );
buf \U$labaj785 ( R_80_7d2c940, \7185 );
buf \U$labaj786 ( R_81_7d2c9e8, \7190 );
buf \U$labaj787 ( R_82_7d2ca90, \7195 );
buf \U$labaj788 ( R_83_7d2cb38, \7200 );
buf \U$labaj789 ( R_84_7d2cbe0, \7205 );
buf \U$labaj790 ( R_85_7d2cc88, \7210 );
buf \U$labaj791 ( R_86_7d2cd30, \7215 );
buf \U$labaj792 ( R_87_7d2cdd8, \7220 );
buf \U$labaj793 ( R_88_7d2ce80, \7225 );
buf \U$labaj794 ( R_89_7d2cf28, \7230 );
buf \U$labaj795 ( R_8a_7d2cfd0, \7235 );
buf \U$labaj796 ( R_8b_7d2d078, \7240 );
buf \U$labaj797 ( R_8c_7d2d120, \7245 );
buf \U$labaj798 ( R_8d_7d2d1c8, \7250 );
buf \U$labaj799 ( R_8e_7d2d270, \7255 );
buf \U$labaj800 ( R_8f_7d2d318, \7260 );
buf \U$labaj801 ( R_90_7d2d3c0, \7265 );
buf \U$labaj802 ( R_91_7d2d468, \7270 );
buf \U$labaj803 ( R_92_7d2d510, \7275 );
buf \U$labaj804 ( R_93_7d2d5b8, \7280 );
buf \U$labaj805 ( R_94_7d2d660, \7285 );
buf \U$labaj806 ( R_95_7d2d708, \7290 );
buf \U$labaj807 ( R_96_7d2d7b0, \7295 );
buf \U$labaj808 ( R_97_7d2d858, \7300 );
buf \U$labaj809 ( R_98_7d2d900, \7305 );
buf \U$labaj810 ( R_99_7d2d9a8, \7310 );
buf \U$labaj811 ( R_9a_7d2da50, \7315 );
buf \U$labaj812 ( R_9b_7d2daf8, \7320 );
buf \U$1 ( \223 , RI2b1c4342d4e0_65);
buf \U$2 ( \224 , RI2b1c4342b6e0_1);
buf \U$3 ( \225 , RI2b1c4342c5e0_33);
xor \U$4 ( \226 , \224 , \225 );
buf \U$5 ( \227 , RI2b1c4342b758_2);
buf \U$6 ( \228 , RI2b1c4342c658_34);
and \U$7 ( \229 , \227 , \228 );
buf \U$8 ( \230 , RI2b1c4342b7d0_3);
buf \U$9 ( \231 , RI2b1c4342c6d0_35);
and \U$10 ( \232 , \230 , \231 );
buf \U$11 ( \233 , RI2b1c4342b848_4);
buf \U$12 ( \234 , RI2b1c4342c748_36);
and \U$13 ( \235 , \233 , \234 );
buf \U$14 ( \236 , RI2b1c4342b8c0_5);
buf \U$15 ( \237 , RI2b1c4342c7c0_37);
and \U$16 ( \238 , \236 , \237 );
buf \U$17 ( \239 , RI2b1c4342b938_6);
buf \U$18 ( \240 , RI2b1c4342c838_38);
and \U$19 ( \241 , \239 , \240 );
buf \U$20 ( \242 , RI2b1c4342b9b0_7);
buf \U$21 ( \243 , RI2b1c4342c8b0_39);
and \U$22 ( \244 , \242 , \243 );
buf \U$23 ( \245 , RI2b1c4342ba28_8);
buf \U$24 ( \246 , RI2b1c4342c928_40);
and \U$25 ( \247 , \245 , \246 );
buf \U$26 ( \248 , RI2b1c4342baa0_9);
buf \U$27 ( \249 , RI2b1c4342c9a0_41);
and \U$28 ( \250 , \248 , \249 );
buf \U$29 ( \251 , RI2b1c4342bb18_10);
buf \U$30 ( \252 , RI2b1c4342ca18_42);
and \U$31 ( \253 , \251 , \252 );
buf \U$32 ( \254 , RI2b1c4342bb90_11);
buf \U$33 ( \255 , RI2b1c4342ca90_43);
and \U$34 ( \256 , \254 , \255 );
buf \U$35 ( \257 , RI2b1c4342bc08_12);
buf \U$36 ( \258 , RI2b1c4342cb08_44);
and \U$37 ( \259 , \257 , \258 );
buf \U$38 ( \260 , RI2b1c4342bc80_13);
buf \U$39 ( \261 , RI2b1c4342cb80_45);
and \U$40 ( \262 , \260 , \261 );
buf \U$41 ( \263 , RI2b1c4342bcf8_14);
buf \U$42 ( \264 , RI2b1c4342cbf8_46);
and \U$43 ( \265 , \263 , \264 );
buf \U$44 ( \266 , RI2b1c4342bd70_15);
buf \U$45 ( \267 , RI2b1c4342cc70_47);
and \U$46 ( \268 , \266 , \267 );
buf \U$47 ( \269 , RI2b1c4342bde8_16);
buf \U$48 ( \270 , RI2b1c4342cce8_48);
and \U$49 ( \271 , \269 , \270 );
buf \U$50 ( \272 , RI2b1c4342be60_17);
buf \U$51 ( \273 , RI2b1c4342cd60_49);
and \U$52 ( \274 , \272 , \273 );
buf \U$53 ( \275 , RI2b1c4342bed8_18);
buf \U$54 ( \276 , RI2b1c4342cdd8_50);
and \U$55 ( \277 , \275 , \276 );
buf \U$56 ( \278 , RI2b1c4342bf50_19);
buf \U$57 ( \279 , RI2b1c4342ce50_51);
and \U$58 ( \280 , \278 , \279 );
buf \U$59 ( \281 , RI2b1c4342bfc8_20);
buf \U$60 ( \282 , RI2b1c4342cec8_52);
and \U$61 ( \283 , \281 , \282 );
buf \U$62 ( \284 , RI2b1c4342c040_21);
buf \U$63 ( \285 , RI2b1c4342cf40_53);
and \U$64 ( \286 , \284 , \285 );
buf \U$65 ( \287 , RI2b1c4342c0b8_22);
buf \U$66 ( \288 , RI2b1c4342cfb8_54);
and \U$67 ( \289 , \287 , \288 );
buf \U$68 ( \290 , RI2b1c4342c130_23);
buf \U$69 ( \291 , RI2b1c4342d030_55);
and \U$70 ( \292 , \290 , \291 );
buf \U$71 ( \293 , RI2b1c4342c1a8_24);
buf \U$72 ( \294 , RI2b1c4342d0a8_56);
and \U$73 ( \295 , \293 , \294 );
buf \U$74 ( \296 , RI2b1c4342c220_25);
buf \U$75 ( \297 , RI2b1c4342d120_57);
and \U$76 ( \298 , \296 , \297 );
buf \U$77 ( \299 , RI2b1c4342c298_26);
buf \U$78 ( \300 , RI2b1c4342d198_58);
and \U$79 ( \301 , \299 , \300 );
buf \U$80 ( \302 , RI2b1c4342c310_27);
buf \U$81 ( \303 , RI2b1c4342d210_59);
and \U$82 ( \304 , \302 , \303 );
buf \U$83 ( \305 , RI2b1c4342c388_28);
buf \U$84 ( \306 , RI2b1c4342d288_60);
and \U$85 ( \307 , \305 , \306 );
buf \U$86 ( \308 , RI2b1c4342c400_29);
buf \U$87 ( \309 , RI2b1c4342d300_61);
and \U$88 ( \310 , \308 , \309 );
buf \U$89 ( \311 , RI2b1c4342c478_30);
buf \U$90 ( \312 , RI2b1c4342d378_62);
and \U$91 ( \313 , \311 , \312 );
buf \U$92 ( \314 , RI2b1c4342c4f0_31);
buf \U$93 ( \315 , RI2b1c4342d3f0_63);
and \U$94 ( \316 , \314 , \315 );
buf \U$95 ( \317 , RI2b1c4342c568_32);
buf \U$96 ( \318 , RI2b1c4342d468_64);
and \U$97 ( \319 , \317 , \318 );
and \U$98 ( \320 , \315 , \319 );
and \U$99 ( \321 , \314 , \319 );
or \U$100 ( \322 , \316 , \320 , \321 );
and \U$101 ( \323 , \312 , \322 );
and \U$102 ( \324 , \311 , \322 );
or \U$103 ( \325 , \313 , \323 , \324 );
and \U$104 ( \326 , \309 , \325 );
and \U$105 ( \327 , \308 , \325 );
or \U$106 ( \328 , \310 , \326 , \327 );
and \U$107 ( \329 , \306 , \328 );
and \U$108 ( \330 , \305 , \328 );
or \U$109 ( \331 , \307 , \329 , \330 );
and \U$110 ( \332 , \303 , \331 );
and \U$111 ( \333 , \302 , \331 );
or \U$112 ( \334 , \304 , \332 , \333 );
and \U$113 ( \335 , \300 , \334 );
and \U$114 ( \336 , \299 , \334 );
or \U$115 ( \337 , \301 , \335 , \336 );
and \U$116 ( \338 , \297 , \337 );
and \U$117 ( \339 , \296 , \337 );
or \U$118 ( \340 , \298 , \338 , \339 );
and \U$119 ( \341 , \294 , \340 );
and \U$120 ( \342 , \293 , \340 );
or \U$121 ( \343 , \295 , \341 , \342 );
and \U$122 ( \344 , \291 , \343 );
and \U$123 ( \345 , \290 , \343 );
or \U$124 ( \346 , \292 , \344 , \345 );
and \U$125 ( \347 , \288 , \346 );
and \U$126 ( \348 , \287 , \346 );
or \U$127 ( \349 , \289 , \347 , \348 );
and \U$128 ( \350 , \285 , \349 );
and \U$129 ( \351 , \284 , \349 );
or \U$130 ( \352 , \286 , \350 , \351 );
and \U$131 ( \353 , \282 , \352 );
and \U$132 ( \354 , \281 , \352 );
or \U$133 ( \355 , \283 , \353 , \354 );
and \U$134 ( \356 , \279 , \355 );
and \U$135 ( \357 , \278 , \355 );
or \U$136 ( \358 , \280 , \356 , \357 );
and \U$137 ( \359 , \276 , \358 );
and \U$138 ( \360 , \275 , \358 );
or \U$139 ( \361 , \277 , \359 , \360 );
and \U$140 ( \362 , \273 , \361 );
and \U$141 ( \363 , \272 , \361 );
or \U$142 ( \364 , \274 , \362 , \363 );
and \U$143 ( \365 , \270 , \364 );
and \U$144 ( \366 , \269 , \364 );
or \U$145 ( \367 , \271 , \365 , \366 );
and \U$146 ( \368 , \267 , \367 );
and \U$147 ( \369 , \266 , \367 );
or \U$148 ( \370 , \268 , \368 , \369 );
and \U$149 ( \371 , \264 , \370 );
and \U$150 ( \372 , \263 , \370 );
or \U$151 ( \373 , \265 , \371 , \372 );
and \U$152 ( \374 , \261 , \373 );
and \U$153 ( \375 , \260 , \373 );
or \U$154 ( \376 , \262 , \374 , \375 );
and \U$155 ( \377 , \258 , \376 );
and \U$156 ( \378 , \257 , \376 );
or \U$157 ( \379 , \259 , \377 , \378 );
and \U$158 ( \380 , \255 , \379 );
and \U$159 ( \381 , \254 , \379 );
or \U$160 ( \382 , \256 , \380 , \381 );
and \U$161 ( \383 , \252 , \382 );
and \U$162 ( \384 , \251 , \382 );
or \U$163 ( \385 , \253 , \383 , \384 );
and \U$164 ( \386 , \249 , \385 );
and \U$165 ( \387 , \248 , \385 );
or \U$166 ( \388 , \250 , \386 , \387 );
and \U$167 ( \389 , \246 , \388 );
and \U$168 ( \390 , \245 , \388 );
or \U$169 ( \391 , \247 , \389 , \390 );
and \U$170 ( \392 , \243 , \391 );
and \U$171 ( \393 , \242 , \391 );
or \U$172 ( \394 , \244 , \392 , \393 );
and \U$173 ( \395 , \240 , \394 );
and \U$174 ( \396 , \239 , \394 );
or \U$175 ( \397 , \241 , \395 , \396 );
and \U$176 ( \398 , \237 , \397 );
and \U$177 ( \399 , \236 , \397 );
or \U$178 ( \400 , \238 , \398 , \399 );
and \U$179 ( \401 , \234 , \400 );
and \U$180 ( \402 , \233 , \400 );
or \U$181 ( \403 , \235 , \401 , \402 );
and \U$182 ( \404 , \231 , \403 );
and \U$183 ( \405 , \230 , \403 );
or \U$184 ( \406 , \232 , \404 , \405 );
and \U$185 ( \407 , \228 , \406 );
and \U$186 ( \408 , \227 , \406 );
or \U$187 ( \409 , \229 , \407 , \408 );
xor \U$188 ( \410 , \226 , \409 );
buf \U$189 ( \411 , \410 );
not \U$190 ( \412 , RI2b1c4342d4e0_65);
not \U$191 ( \413 , RI2b1c4342d558_66);
xor \U$192 ( \414 , \412 , \413 );
not \U$193 ( \415 , RI2b1c4342d5d0_67);
not \U$194 ( \416 , RI2b1c4342d648_68);
xor \U$195 ( \417 , \415 , \416 );
xor \U$196 ( \418 , \414 , \417 );
not \U$197 ( \419 , RI2b1c4342d6c0_69);
not \U$198 ( \420 , RI2b1c4342d738_70);
xor \U$199 ( \421 , \419 , \420 );
not \U$200 ( \422 , RI2b1c4342d7b0_71);
not \U$201 ( \423 , RI2b1c4342d828_72);
xor \U$202 ( \424 , \422 , \423 );
xor \U$203 ( \425 , \421 , \424 );
xor \U$204 ( \426 , \418 , \425 );
not \U$205 ( \427 , RI2b1c4342d8a0_73);
not \U$206 ( \428 , RI2b1c4342d918_74);
xor \U$207 ( \429 , \427 , \428 );
not \U$208 ( \430 , RI2b1c4342d990_75);
not \U$209 ( \431 , RI2b1c4342da08_76);
xor \U$210 ( \432 , \430 , \431 );
xor \U$211 ( \433 , \429 , \432 );
not \U$212 ( \434 , RI2b1c4342da80_77);
not \U$213 ( \435 , RI2b1c4342daf8_78);
xor \U$214 ( \436 , \434 , \435 );
not \U$215 ( \437 , RI2b1c4342db70_79);
not \U$216 ( \438 , RI2b1c4342dbe8_80);
xor \U$217 ( \439 , \437 , \438 );
xor \U$218 ( \440 , \436 , \439 );
xor \U$219 ( \441 , \433 , \440 );
xor \U$220 ( \442 , \426 , \441 );
not \U$221 ( \443 , RI2b1c4342dc60_81);
not \U$222 ( \444 , RI2b1c4342dcd8_82);
xor \U$223 ( \445 , \443 , \444 );
not \U$224 ( \446 , RI2b1c4342dd50_83);
not \U$225 ( \447 , RI2b1c4342ddc8_84);
xor \U$226 ( \448 , \446 , \447 );
xor \U$227 ( \449 , \445 , \448 );
not \U$228 ( \450 , RI2b1c4342de40_85);
not \U$229 ( \451 , RI2b1c4342deb8_86);
xor \U$230 ( \452 , \450 , \451 );
not \U$231 ( \453 , RI2b1c4342df30_87);
not \U$232 ( \454 , RI2b1c4342dfa8_88);
xor \U$233 ( \455 , \453 , \454 );
xor \U$234 ( \456 , \452 , \455 );
xor \U$235 ( \457 , \449 , \456 );
not \U$236 ( \458 , RI2b1c4342e020_89);
not \U$237 ( \459 , RI2b1c4342e098_90);
xor \U$238 ( \460 , \458 , \459 );
not \U$239 ( \461 , RI2b1c4342e110_91);
not \U$240 ( \462 , RI2b1c4342e188_92);
xor \U$241 ( \463 , \461 , \462 );
xor \U$242 ( \464 , \460 , \463 );
not \U$243 ( \465 , RI2b1c4342e200_93);
not \U$244 ( \466 , RI2b1c4342e278_94);
xor \U$245 ( \467 , \465 , \466 );
not \U$246 ( \468 , RI2b1c4342e2f0_95);
not \U$247 ( \469 , RI2b1c4342e368_96);
xor \U$248 ( \470 , \468 , \469 );
xor \U$249 ( \471 , \467 , \470 );
xor \U$250 ( \472 , \464 , \471 );
xor \U$251 ( \473 , \457 , \472 );
xor \U$252 ( \474 , \442 , \473 );
not \U$253 ( \475 , \474 );
_DC r2b9 ( \476_nR2b9 , \411 , \475 );
buf \U$254 ( \477 , RI2b1c4342b6e0_1);
and \U$255 ( \478 , \476_nR2b9 , \477 );
buf \U$256 ( \479 , \478 );
xor \U$257 ( \480 , \227 , \228 );
xor \U$258 ( \481 , \480 , \406 );
buf \U$259 ( \482 , \481 );
_DC r2ad ( \483_nR2ad , \482 , \475 );
buf \U$260 ( \484 , RI2b1c4342b758_2);
and \U$261 ( \485 , \483_nR2ad , \484 );
buf \U$262 ( \486 , \485 );
xor \U$263 ( \487 , \479 , \486 );
xor \U$264 ( \488 , \230 , \231 );
xor \U$265 ( \489 , \488 , \403 );
buf \U$266 ( \490 , \489 );
_DC r2a1 ( \491_nR2a1 , \490 , \475 );
buf \U$267 ( \492 , RI2b1c4342b7d0_3);
and \U$268 ( \493 , \491_nR2a1 , \492 );
buf \U$269 ( \494 , \493 );
xor \U$270 ( \495 , \486 , \494 );
not \U$271 ( \496 , \495 );
and \U$272 ( \497 , \487 , \496 );
and \U$273 ( \498 , \223 , \497 );
not \U$274 ( \499 , \498 );
and \U$275 ( \500 , \486 , \494 );
not \U$276 ( \501 , \500 );
and \U$277 ( \502 , \479 , \501 );
xnor \U$278 ( \503 , \499 , \502 );
buf \U$280 ( \504 , RI2b1c4342d558_66);
xor \U$283 ( \505 , 1'b0 , \479 );
and \U$284 ( \506 , \504 , \505 );
nor \U$285 ( \507 , 1'b0 , \506 );
not \U$286 ( \508 , \507 );
or \U$287 ( \509 , \503 , \508 );
not \U$288 ( \510 , \502 );
xor \U$289 ( \511 , \509 , \510 );
and \U$291 ( \512 , \223 , \505 );
nor \U$292 ( \513 , 1'b0 , \512 );
not \U$293 ( \514 , \513 );
xor \U$294 ( \515 , \511 , \514 );
xor \U$295 ( \516 , \233 , \234 );
xor \U$296 ( \517 , \516 , \400 );
buf \U$297 ( \518 , \517 );
_DC r295 ( \519_nR295 , \518 , \475 );
buf \U$298 ( \520 , RI2b1c4342b848_4);
and \U$299 ( \521 , \519_nR295 , \520 );
buf \U$300 ( \522 , \521 );
xor \U$301 ( \523 , \236 , \237 );
xor \U$302 ( \524 , \523 , \397 );
buf \U$303 ( \525 , \524 );
_DC r289 ( \526_nR289 , \525 , \475 );
buf \U$304 ( \527 , RI2b1c4342b8c0_5);
and \U$305 ( \528 , \526_nR289 , \527 );
buf \U$306 ( \529 , \528 );
and \U$307 ( \530 , \522 , \529 );
not \U$308 ( \531 , \530 );
and \U$309 ( \532 , \494 , \531 );
not \U$310 ( \533 , \532 );
and \U$311 ( \534 , \504 , \497 );
and \U$312 ( \535 , \223 , \495 );
nor \U$313 ( \536 , \534 , \535 );
xnor \U$314 ( \537 , \536 , \502 );
and \U$315 ( \538 , \533 , \537 );
buf \U$317 ( \539 , RI2b1c4342d5d0_67);
and \U$318 ( \540 , \539 , \505 );
nor \U$319 ( \541 , 1'b0 , \540 );
not \U$320 ( \542 , \541 );
and \U$321 ( \543 , \537 , \542 );
and \U$322 ( \544 , \533 , \542 );
or \U$323 ( \545 , \538 , \543 , \544 );
xnor \U$324 ( \546 , \503 , \508 );
and \U$325 ( \547 , \545 , \546 );
nand \U$326 ( \548 , \515 , \547 );
nor \U$327 ( \549 , \515 , \547 );
not \U$328 ( \550 , \549 );
nand \U$329 ( \551 , \548 , \550 );
xor \U$330 ( \552 , \239 , \240 );
xor \U$331 ( \553 , \552 , \394 );
buf \U$332 ( \554 , \553 );
_DC r27d ( \555_nR27d , \554 , \475 );
buf \U$333 ( \556 , RI2b1c4342b938_6);
and \U$334 ( \557 , \555_nR27d , \556 );
buf \U$335 ( \558 , \557 );
xor \U$336 ( \559 , \242 , \243 );
xor \U$337 ( \560 , \559 , \391 );
buf \U$338 ( \561 , \560 );
_DC r271 ( \562_nR271 , \561 , \475 );
buf \U$339 ( \563 , RI2b1c4342b9b0_7);
and \U$340 ( \564 , \562_nR271 , \563 );
buf \U$341 ( \565 , \564 );
and \U$342 ( \566 , \558 , \565 );
not \U$343 ( \567 , \566 );
and \U$344 ( \568 , \529 , \567 );
buf \U$345 ( \569 , RI2b1c4342d7b0_71);
xor \U$346 ( \570 , \314 , \315 );
xor \U$347 ( \571 , \570 , \319 );
buf \U$348 ( \572 , \571 );
_DC r151 ( \573_nR151 , \572 , \475 );
buf \U$349 ( \574 , RI2b1c4342c4f0_31);
and \U$350 ( \575 , \573_nR151 , \574 );
buf \U$351 ( \576 , \575 );
xor \U$352 ( \577 , \317 , \318 );
buf \U$353 ( \578 , \577 );
_DC r129 ( \579_nR129 , \578 , \475 );
xor \U$354 ( \580 , RI2b1c4342c5e0_33, RI2b1c4342c658_34);
xor \U$355 ( \581 , RI2b1c4342c6d0_35, RI2b1c4342c748_36);
xor \U$356 ( \582 , \580 , \581 );
xor \U$357 ( \583 , RI2b1c4342c7c0_37, RI2b1c4342c838_38);
xor \U$358 ( \584 , RI2b1c4342c8b0_39, RI2b1c4342c928_40);
xor \U$359 ( \585 , \583 , \584 );
xor \U$360 ( \586 , \582 , \585 );
xor \U$361 ( \587 , RI2b1c4342c9a0_41, RI2b1c4342ca18_42);
xor \U$362 ( \588 , RI2b1c4342ca90_43, RI2b1c4342cb08_44);
xor \U$363 ( \589 , \587 , \588 );
xor \U$364 ( \590 , RI2b1c4342cb80_45, RI2b1c4342cbf8_46);
xor \U$365 ( \591 , RI2b1c4342cc70_47, RI2b1c4342cce8_48);
xor \U$366 ( \592 , \590 , \591 );
xor \U$367 ( \593 , \589 , \592 );
xor \U$368 ( \594 , \586 , \593 );
xor \U$369 ( \595 , RI2b1c4342cd60_49, RI2b1c4342cdd8_50);
xor \U$370 ( \596 , RI2b1c4342ce50_51, RI2b1c4342cec8_52);
xor \U$371 ( \597 , \595 , \596 );
xor \U$372 ( \598 , RI2b1c4342cf40_53, RI2b1c4342cfb8_54);
xor \U$373 ( \599 , RI2b1c4342d030_55, RI2b1c4342d0a8_56);
xor \U$374 ( \600 , \598 , \599 );
xor \U$375 ( \601 , \597 , \600 );
xor \U$376 ( \602 , RI2b1c4342d120_57, RI2b1c4342d198_58);
xor \U$377 ( \603 , RI2b1c4342d210_59, RI2b1c4342d288_60);
xor \U$378 ( \604 , \602 , \603 );
xor \U$379 ( \605 , RI2b1c4342d300_61, RI2b1c4342d378_62);
xor \U$380 ( \606 , RI2b1c4342d3f0_63, RI2b1c4342d468_64);
xor \U$381 ( \607 , \605 , \606 );
xor \U$382 ( \608 , \604 , \607 );
xor \U$383 ( \609 , \601 , \608 );
xor \U$384 ( \610 , \594 , \609 );
xor \U$385 ( \611 , \610 , RI2b1c4342c568_32);
and \U$386 ( \612 , \579_nR129 , \611 );
buf \U$387 ( \613 , \612 );
xor \U$388 ( \614 , \576 , \613 );
not \U$389 ( \615 , \613 );
and \U$390 ( \616 , \614 , \615 );
and \U$391 ( \617 , \569 , \616 );
buf \U$392 ( \618 , RI2b1c4342d738_70);
and \U$393 ( \619 , \618 , \613 );
nor \U$394 ( \620 , \617 , \619 );
xnor \U$395 ( \621 , \620 , \576 );
and \U$396 ( \622 , \568 , \621 );
buf \U$397 ( \623 , RI2b1c4342d8a0_73);
xor \U$398 ( \624 , \308 , \309 );
xor \U$399 ( \625 , \624 , \325 );
buf \U$400 ( \626 , \625 );
_DC r169 ( \627_nR169 , \626 , \475 );
buf \U$401 ( \628 , RI2b1c4342c400_29);
and \U$402 ( \629 , \627_nR169 , \628 );
buf \U$403 ( \630 , \629 );
xor \U$404 ( \631 , \311 , \312 );
xor \U$405 ( \632 , \631 , \322 );
buf \U$406 ( \633 , \632 );
_DC r15d ( \634_nR15d , \633 , \475 );
buf \U$407 ( \635 , RI2b1c4342c478_30);
and \U$408 ( \636 , \634_nR15d , \635 );
buf \U$409 ( \637 , \636 );
xor \U$410 ( \638 , \630 , \637 );
xor \U$411 ( \639 , \637 , \576 );
not \U$412 ( \640 , \639 );
and \U$413 ( \641 , \638 , \640 );
and \U$414 ( \642 , \623 , \641 );
buf \U$415 ( \643 , RI2b1c4342d828_72);
and \U$416 ( \644 , \643 , \639 );
nor \U$417 ( \645 , \642 , \644 );
and \U$418 ( \646 , \637 , \576 );
not \U$419 ( \647 , \646 );
and \U$420 ( \648 , \630 , \647 );
xnor \U$421 ( \649 , \645 , \648 );
and \U$422 ( \650 , \621 , \649 );
and \U$423 ( \651 , \568 , \649 );
or \U$424 ( \652 , \622 , \650 , \651 );
buf \U$425 ( \653 , RI2b1c4342d990_75);
xor \U$426 ( \654 , \302 , \303 );
xor \U$427 ( \655 , \654 , \331 );
buf \U$428 ( \656 , \655 );
_DC r181 ( \657_nR181 , \656 , \475 );
buf \U$429 ( \658 , RI2b1c4342c310_27);
and \U$430 ( \659 , \657_nR181 , \658 );
buf \U$431 ( \660 , \659 );
xor \U$432 ( \661 , \305 , \306 );
xor \U$433 ( \662 , \661 , \328 );
buf \U$434 ( \663 , \662 );
_DC r175 ( \664_nR175 , \663 , \475 );
buf \U$435 ( \665 , RI2b1c4342c388_28);
and \U$436 ( \666 , \664_nR175 , \665 );
buf \U$437 ( \667 , \666 );
xor \U$438 ( \668 , \660 , \667 );
xor \U$439 ( \669 , \667 , \630 );
not \U$440 ( \670 , \669 );
and \U$441 ( \671 , \668 , \670 );
and \U$442 ( \672 , \653 , \671 );
buf \U$443 ( \673 , RI2b1c4342d918_74);
and \U$444 ( \674 , \673 , \669 );
nor \U$445 ( \675 , \672 , \674 );
and \U$446 ( \676 , \667 , \630 );
not \U$447 ( \677 , \676 );
and \U$448 ( \678 , \660 , \677 );
xnor \U$449 ( \679 , \675 , \678 );
buf \U$450 ( \680 , RI2b1c4342da80_77);
xor \U$451 ( \681 , \296 , \297 );
xor \U$452 ( \682 , \681 , \337 );
buf \U$453 ( \683 , \682 );
_DC r199 ( \684_nR199 , \683 , \475 );
buf \U$454 ( \685 , RI2b1c4342c220_25);
and \U$455 ( \686 , \684_nR199 , \685 );
buf \U$456 ( \687 , \686 );
xor \U$457 ( \688 , \299 , \300 );
xor \U$458 ( \689 , \688 , \334 );
buf \U$459 ( \690 , \689 );
_DC r18d ( \691_nR18d , \690 , \475 );
buf \U$460 ( \692 , RI2b1c4342c298_26);
and \U$461 ( \693 , \691_nR18d , \692 );
buf \U$462 ( \694 , \693 );
xor \U$463 ( \695 , \687 , \694 );
xor \U$464 ( \696 , \694 , \660 );
not \U$465 ( \697 , \696 );
and \U$466 ( \698 , \695 , \697 );
and \U$467 ( \699 , \680 , \698 );
buf \U$468 ( \700 , RI2b1c4342da08_76);
and \U$469 ( \701 , \700 , \696 );
nor \U$470 ( \702 , \699 , \701 );
and \U$471 ( \703 , \694 , \660 );
not \U$472 ( \704 , \703 );
and \U$473 ( \705 , \687 , \704 );
xnor \U$474 ( \706 , \702 , \705 );
and \U$475 ( \707 , \679 , \706 );
buf \U$476 ( \708 , RI2b1c4342db70_79);
xor \U$477 ( \709 , \290 , \291 );
xor \U$478 ( \710 , \709 , \343 );
buf \U$479 ( \711 , \710 );
_DC r1b1 ( \712_nR1b1 , \711 , \475 );
buf \U$480 ( \713 , RI2b1c4342c130_23);
and \U$481 ( \714 , \712_nR1b1 , \713 );
buf \U$482 ( \715 , \714 );
xor \U$483 ( \716 , \293 , \294 );
xor \U$484 ( \717 , \716 , \340 );
buf \U$485 ( \718 , \717 );
_DC r1a5 ( \719_nR1a5 , \718 , \475 );
buf \U$486 ( \720 , RI2b1c4342c1a8_24);
and \U$487 ( \721 , \719_nR1a5 , \720 );
buf \U$488 ( \722 , \721 );
xor \U$489 ( \723 , \715 , \722 );
xor \U$490 ( \724 , \722 , \687 );
not \U$491 ( \725 , \724 );
and \U$492 ( \726 , \723 , \725 );
and \U$493 ( \727 , \708 , \726 );
buf \U$494 ( \728 , RI2b1c4342daf8_78);
and \U$495 ( \729 , \728 , \724 );
nor \U$496 ( \730 , \727 , \729 );
and \U$497 ( \731 , \722 , \687 );
not \U$498 ( \732 , \731 );
and \U$499 ( \733 , \715 , \732 );
xnor \U$500 ( \734 , \730 , \733 );
and \U$501 ( \735 , \706 , \734 );
and \U$502 ( \736 , \679 , \734 );
or \U$503 ( \737 , \707 , \735 , \736 );
and \U$504 ( \738 , \652 , \737 );
buf \U$505 ( \739 , RI2b1c4342dc60_81);
xor \U$506 ( \740 , \284 , \285 );
xor \U$507 ( \741 , \740 , \349 );
buf \U$508 ( \742 , \741 );
_DC r1c9 ( \743_nR1c9 , \742 , \475 );
buf \U$509 ( \744 , RI2b1c4342c040_21);
and \U$510 ( \745 , \743_nR1c9 , \744 );
buf \U$511 ( \746 , \745 );
xor \U$512 ( \747 , \287 , \288 );
xor \U$513 ( \748 , \747 , \346 );
buf \U$514 ( \749 , \748 );
_DC r1bd ( \750_nR1bd , \749 , \475 );
buf \U$515 ( \751 , RI2b1c4342c0b8_22);
and \U$516 ( \752 , \750_nR1bd , \751 );
buf \U$517 ( \753 , \752 );
xor \U$518 ( \754 , \746 , \753 );
xor \U$519 ( \755 , \753 , \715 );
not \U$520 ( \756 , \755 );
and \U$521 ( \757 , \754 , \756 );
and \U$522 ( \758 , \739 , \757 );
buf \U$523 ( \759 , RI2b1c4342dbe8_80);
and \U$524 ( \760 , \759 , \755 );
nor \U$525 ( \761 , \758 , \760 );
and \U$526 ( \762 , \753 , \715 );
not \U$527 ( \763 , \762 );
and \U$528 ( \764 , \746 , \763 );
xnor \U$529 ( \765 , \761 , \764 );
buf \U$530 ( \766 , RI2b1c4342dd50_83);
xor \U$531 ( \767 , \278 , \279 );
xor \U$532 ( \768 , \767 , \355 );
buf \U$533 ( \769 , \768 );
_DC r1e1 ( \770_nR1e1 , \769 , \475 );
buf \U$534 ( \771 , RI2b1c4342bf50_19);
and \U$535 ( \772 , \770_nR1e1 , \771 );
buf \U$536 ( \773 , \772 );
xor \U$537 ( \774 , \281 , \282 );
xor \U$538 ( \775 , \774 , \352 );
buf \U$539 ( \776 , \775 );
_DC r1d5 ( \777_nR1d5 , \776 , \475 );
buf \U$540 ( \778 , RI2b1c4342bfc8_20);
and \U$541 ( \779 , \777_nR1d5 , \778 );
buf \U$542 ( \780 , \779 );
xor \U$543 ( \781 , \773 , \780 );
xor \U$544 ( \782 , \780 , \746 );
not \U$545 ( \783 , \782 );
and \U$546 ( \784 , \781 , \783 );
and \U$547 ( \785 , \766 , \784 );
buf \U$548 ( \786 , RI2b1c4342dcd8_82);
and \U$549 ( \787 , \786 , \782 );
nor \U$550 ( \788 , \785 , \787 );
and \U$551 ( \789 , \780 , \746 );
not \U$552 ( \790 , \789 );
and \U$553 ( \791 , \773 , \790 );
xnor \U$554 ( \792 , \788 , \791 );
and \U$555 ( \793 , \765 , \792 );
buf \U$556 ( \794 , RI2b1c4342de40_85);
xor \U$557 ( \795 , \272 , \273 );
xor \U$558 ( \796 , \795 , \361 );
buf \U$559 ( \797 , \796 );
_DC r1f9 ( \798_nR1f9 , \797 , \475 );
buf \U$560 ( \799 , RI2b1c4342be60_17);
and \U$561 ( \800 , \798_nR1f9 , \799 );
buf \U$562 ( \801 , \800 );
xor \U$563 ( \802 , \275 , \276 );
xor \U$564 ( \803 , \802 , \358 );
buf \U$565 ( \804 , \803 );
_DC r1ed ( \805_nR1ed , \804 , \475 );
buf \U$566 ( \806 , RI2b1c4342bed8_18);
and \U$567 ( \807 , \805_nR1ed , \806 );
buf \U$568 ( \808 , \807 );
xor \U$569 ( \809 , \801 , \808 );
xor \U$570 ( \810 , \808 , \773 );
not \U$571 ( \811 , \810 );
and \U$572 ( \812 , \809 , \811 );
and \U$573 ( \813 , \794 , \812 );
buf \U$574 ( \814 , RI2b1c4342ddc8_84);
and \U$575 ( \815 , \814 , \810 );
nor \U$576 ( \816 , \813 , \815 );
and \U$577 ( \817 , \808 , \773 );
not \U$578 ( \818 , \817 );
and \U$579 ( \819 , \801 , \818 );
xnor \U$580 ( \820 , \816 , \819 );
and \U$581 ( \821 , \792 , \820 );
and \U$582 ( \822 , \765 , \820 );
or \U$583 ( \823 , \793 , \821 , \822 );
and \U$584 ( \824 , \737 , \823 );
and \U$585 ( \825 , \652 , \823 );
or \U$586 ( \826 , \738 , \824 , \825 );
buf \U$587 ( \827 , RI2b1c4342df30_87);
xor \U$588 ( \828 , \266 , \267 );
xor \U$589 ( \829 , \828 , \367 );
buf \U$590 ( \830 , \829 );
_DC r211 ( \831_nR211 , \830 , \475 );
buf \U$591 ( \832 , RI2b1c4342bd70_15);
and \U$592 ( \833 , \831_nR211 , \832 );
buf \U$593 ( \834 , \833 );
xor \U$594 ( \835 , \269 , \270 );
xor \U$595 ( \836 , \835 , \364 );
buf \U$596 ( \837 , \836 );
_DC r205 ( \838_nR205 , \837 , \475 );
buf \U$597 ( \839 , RI2b1c4342bde8_16);
and \U$598 ( \840 , \838_nR205 , \839 );
buf \U$599 ( \841 , \840 );
xor \U$600 ( \842 , \834 , \841 );
xor \U$601 ( \843 , \841 , \801 );
not \U$602 ( \844 , \843 );
and \U$603 ( \845 , \842 , \844 );
and \U$604 ( \846 , \827 , \845 );
buf \U$605 ( \847 , RI2b1c4342deb8_86);
and \U$606 ( \848 , \847 , \843 );
nor \U$607 ( \849 , \846 , \848 );
and \U$608 ( \850 , \841 , \801 );
not \U$609 ( \851 , \850 );
and \U$610 ( \852 , \834 , \851 );
xnor \U$611 ( \853 , \849 , \852 );
buf \U$612 ( \854 , RI2b1c4342e020_89);
xor \U$613 ( \855 , \260 , \261 );
xor \U$614 ( \856 , \855 , \373 );
buf \U$615 ( \857 , \856 );
_DC r229 ( \858_nR229 , \857 , \475 );
buf \U$616 ( \859 , RI2b1c4342bc80_13);
and \U$617 ( \860 , \858_nR229 , \859 );
buf \U$618 ( \861 , \860 );
xor \U$619 ( \862 , \263 , \264 );
xor \U$620 ( \863 , \862 , \370 );
buf \U$621 ( \864 , \863 );
_DC r21d ( \865_nR21d , \864 , \475 );
buf \U$622 ( \866 , RI2b1c4342bcf8_14);
and \U$623 ( \867 , \865_nR21d , \866 );
buf \U$624 ( \868 , \867 );
xor \U$625 ( \869 , \861 , \868 );
xor \U$626 ( \870 , \868 , \834 );
not \U$627 ( \871 , \870 );
and \U$628 ( \872 , \869 , \871 );
and \U$629 ( \873 , \854 , \872 );
buf \U$630 ( \874 , RI2b1c4342dfa8_88);
and \U$631 ( \875 , \874 , \870 );
nor \U$632 ( \876 , \873 , \875 );
and \U$633 ( \877 , \868 , \834 );
not \U$634 ( \878 , \877 );
and \U$635 ( \879 , \861 , \878 );
xnor \U$636 ( \880 , \876 , \879 );
and \U$637 ( \881 , \853 , \880 );
buf \U$638 ( \882 , RI2b1c4342e110_91);
xor \U$639 ( \883 , \254 , \255 );
xor \U$640 ( \884 , \883 , \379 );
buf \U$641 ( \885 , \884 );
_DC r241 ( \886_nR241 , \885 , \475 );
buf \U$642 ( \887 , RI2b1c4342bb90_11);
and \U$643 ( \888 , \886_nR241 , \887 );
buf \U$644 ( \889 , \888 );
xor \U$645 ( \890 , \257 , \258 );
xor \U$646 ( \891 , \890 , \376 );
buf \U$647 ( \892 , \891 );
_DC r235 ( \893_nR235 , \892 , \475 );
buf \U$648 ( \894 , RI2b1c4342bc08_12);
and \U$649 ( \895 , \893_nR235 , \894 );
buf \U$650 ( \896 , \895 );
xor \U$651 ( \897 , \889 , \896 );
xor \U$652 ( \898 , \896 , \861 );
not \U$653 ( \899 , \898 );
and \U$654 ( \900 , \897 , \899 );
and \U$655 ( \901 , \882 , \900 );
buf \U$656 ( \902 , RI2b1c4342e098_90);
and \U$657 ( \903 , \902 , \898 );
nor \U$658 ( \904 , \901 , \903 );
and \U$659 ( \905 , \896 , \861 );
not \U$660 ( \906 , \905 );
and \U$661 ( \907 , \889 , \906 );
xnor \U$662 ( \908 , \904 , \907 );
and \U$663 ( \909 , \880 , \908 );
and \U$664 ( \910 , \853 , \908 );
or \U$665 ( \911 , \881 , \909 , \910 );
buf \U$666 ( \912 , RI2b1c4342e200_93);
xor \U$667 ( \913 , \248 , \249 );
xor \U$668 ( \914 , \913 , \385 );
buf \U$669 ( \915 , \914 );
_DC r259 ( \916_nR259 , \915 , \475 );
buf \U$670 ( \917 , RI2b1c4342baa0_9);
and \U$671 ( \918 , \916_nR259 , \917 );
buf \U$672 ( \919 , \918 );
xor \U$673 ( \920 , \251 , \252 );
xor \U$674 ( \921 , \920 , \382 );
buf \U$675 ( \922 , \921 );
_DC r24d ( \923_nR24d , \922 , \475 );
buf \U$676 ( \924 , RI2b1c4342bb18_10);
and \U$677 ( \925 , \923_nR24d , \924 );
buf \U$678 ( \926 , \925 );
xor \U$679 ( \927 , \919 , \926 );
xor \U$680 ( \928 , \926 , \889 );
not \U$681 ( \929 , \928 );
and \U$682 ( \930 , \927 , \929 );
and \U$683 ( \931 , \912 , \930 );
buf \U$684 ( \932 , RI2b1c4342e188_92);
and \U$685 ( \933 , \932 , \928 );
nor \U$686 ( \934 , \931 , \933 );
and \U$687 ( \935 , \926 , \889 );
not \U$688 ( \936 , \935 );
and \U$689 ( \937 , \919 , \936 );
xnor \U$690 ( \938 , \934 , \937 );
buf \U$691 ( \939 , RI2b1c4342e2f0_95);
xor \U$692 ( \940 , \245 , \246 );
xor \U$693 ( \941 , \940 , \388 );
buf \U$694 ( \942 , \941 );
_DC r265 ( \943_nR265 , \942 , \475 );
buf \U$695 ( \944 , RI2b1c4342ba28_8);
and \U$696 ( \945 , \943_nR265 , \944 );
buf \U$697 ( \946 , \945 );
xor \U$698 ( \947 , \565 , \946 );
xor \U$699 ( \948 , \946 , \919 );
not \U$700 ( \949 , \948 );
and \U$701 ( \950 , \947 , \949 );
and \U$702 ( \951 , \939 , \950 );
buf \U$703 ( \952 , RI2b1c4342e278_94);
and \U$704 ( \953 , \952 , \948 );
nor \U$705 ( \954 , \951 , \953 );
and \U$706 ( \955 , \946 , \919 );
not \U$707 ( \956 , \955 );
and \U$708 ( \957 , \565 , \956 );
xnor \U$709 ( \958 , \954 , \957 );
and \U$710 ( \959 , \938 , \958 );
buf \U$711 ( \960 , RI2b1c4342e368_96);
xor \U$712 ( \961 , \558 , \565 );
nand \U$713 ( \962 , \960 , \961 );
xnor \U$714 ( \963 , \962 , \568 );
and \U$715 ( \964 , \958 , \963 );
and \U$716 ( \965 , \938 , \963 );
or \U$717 ( \966 , \959 , \964 , \965 );
and \U$718 ( \967 , \911 , \966 );
and \U$719 ( \968 , \952 , \950 );
and \U$720 ( \969 , \912 , \948 );
nor \U$721 ( \970 , \968 , \969 );
xnor \U$722 ( \971 , \970 , \957 );
and \U$723 ( \972 , \966 , \971 );
and \U$724 ( \973 , \911 , \971 );
or \U$725 ( \974 , \967 , \972 , \973 );
and \U$726 ( \975 , \826 , \974 );
xor \U$727 ( \976 , \529 , \558 );
not \U$728 ( \977 , \961 );
and \U$729 ( \978 , \976 , \977 );
and \U$730 ( \979 , \960 , \978 );
and \U$731 ( \980 , \939 , \961 );
nor \U$732 ( \981 , \979 , \980 );
xnor \U$733 ( \982 , \981 , \568 );
and \U$734 ( \983 , \874 , \872 );
and \U$735 ( \984 , \827 , \870 );
nor \U$736 ( \985 , \983 , \984 );
xnor \U$737 ( \986 , \985 , \879 );
and \U$738 ( \987 , \902 , \900 );
and \U$739 ( \988 , \854 , \898 );
nor \U$740 ( \989 , \987 , \988 );
xnor \U$741 ( \990 , \989 , \907 );
xor \U$742 ( \991 , \986 , \990 );
and \U$743 ( \992 , \932 , \930 );
and \U$744 ( \993 , \882 , \928 );
nor \U$745 ( \994 , \992 , \993 );
xnor \U$746 ( \995 , \994 , \937 );
xor \U$747 ( \996 , \991 , \995 );
and \U$748 ( \997 , \982 , \996 );
and \U$749 ( \998 , \786 , \784 );
and \U$750 ( \999 , \739 , \782 );
nor \U$751 ( \1000 , \998 , \999 );
xnor \U$752 ( \1001 , \1000 , \791 );
and \U$753 ( \1002 , \814 , \812 );
and \U$754 ( \1003 , \766 , \810 );
nor \U$755 ( \1004 , \1002 , \1003 );
xnor \U$756 ( \1005 , \1004 , \819 );
xor \U$757 ( \1006 , \1001 , \1005 );
and \U$758 ( \1007 , \847 , \845 );
and \U$759 ( \1008 , \794 , \843 );
nor \U$760 ( \1009 , \1007 , \1008 );
xnor \U$761 ( \1010 , \1009 , \852 );
xor \U$762 ( \1011 , \1006 , \1010 );
and \U$763 ( \1012 , \996 , \1011 );
and \U$764 ( \1013 , \982 , \1011 );
or \U$765 ( \1014 , \997 , \1012 , \1013 );
and \U$766 ( \1015 , \974 , \1014 );
and \U$767 ( \1016 , \826 , \1014 );
or \U$768 ( \1017 , \975 , \1015 , \1016 );
buf \U$769 ( \1018 , RI2b1c4342d6c0_69);
and \U$770 ( \1019 , \1018 , \616 );
buf \U$771 ( \1020 , RI2b1c4342d648_68);
and \U$772 ( \1021 , \1020 , \613 );
nor \U$773 ( \1022 , \1019 , \1021 );
xnor \U$774 ( \1023 , \1022 , \576 );
xor \U$775 ( \1024 , \532 , \1023 );
and \U$776 ( \1025 , \569 , \641 );
and \U$777 ( \1026 , \618 , \639 );
nor \U$778 ( \1027 , \1025 , \1026 );
xnor \U$779 ( \1028 , \1027 , \648 );
xor \U$780 ( \1029 , \1024 , \1028 );
and \U$781 ( \1030 , \794 , \845 );
and \U$782 ( \1031 , \814 , \843 );
nor \U$783 ( \1032 , \1030 , \1031 );
xnor \U$784 ( \1033 , \1032 , \852 );
and \U$785 ( \1034 , \827 , \872 );
and \U$786 ( \1035 , \847 , \870 );
nor \U$787 ( \1036 , \1034 , \1035 );
xnor \U$788 ( \1037 , \1036 , \879 );
xor \U$789 ( \1038 , \1033 , \1037 );
and \U$790 ( \1039 , \854 , \900 );
and \U$791 ( \1040 , \874 , \898 );
nor \U$792 ( \1041 , \1039 , \1040 );
xnor \U$793 ( \1042 , \1041 , \907 );
xor \U$794 ( \1043 , \1038 , \1042 );
and \U$795 ( \1044 , \708 , \757 );
and \U$796 ( \1045 , \728 , \755 );
nor \U$797 ( \1046 , \1044 , \1045 );
xnor \U$798 ( \1047 , \1046 , \764 );
and \U$799 ( \1048 , \739 , \784 );
and \U$800 ( \1049 , \759 , \782 );
nor \U$801 ( \1050 , \1048 , \1049 );
xnor \U$802 ( \1051 , \1050 , \791 );
xor \U$803 ( \1052 , \1047 , \1051 );
and \U$804 ( \1053 , \766 , \812 );
and \U$805 ( \1054 , \786 , \810 );
nor \U$806 ( \1055 , \1053 , \1054 );
xnor \U$807 ( \1056 , \1055 , \819 );
xor \U$808 ( \1057 , \1052 , \1056 );
xor \U$809 ( \1058 , \1043 , \1057 );
and \U$810 ( \1059 , \623 , \671 );
and \U$811 ( \1060 , \643 , \669 );
nor \U$812 ( \1061 , \1059 , \1060 );
xnor \U$813 ( \1062 , \1061 , \678 );
and \U$814 ( \1063 , \653 , \698 );
and \U$815 ( \1064 , \673 , \696 );
nor \U$816 ( \1065 , \1063 , \1064 );
xnor \U$817 ( \1066 , \1065 , \705 );
xor \U$818 ( \1067 , \1062 , \1066 );
and \U$819 ( \1068 , \680 , \726 );
and \U$820 ( \1069 , \700 , \724 );
nor \U$821 ( \1070 , \1068 , \1069 );
xnor \U$822 ( \1071 , \1070 , \733 );
xor \U$823 ( \1072 , \1067 , \1071 );
xor \U$824 ( \1073 , \1058 , \1072 );
and \U$825 ( \1074 , \1029 , \1073 );
and \U$826 ( \1075 , \986 , \990 );
and \U$827 ( \1076 , \990 , \995 );
and \U$828 ( \1077 , \986 , \995 );
or \U$829 ( \1078 , \1075 , \1076 , \1077 );
xor \U$830 ( \1079 , \522 , \529 );
nand \U$831 ( \1080 , \960 , \1079 );
xnor \U$832 ( \1081 , \1080 , \532 );
xor \U$833 ( \1082 , \1078 , \1081 );
and \U$834 ( \1083 , \882 , \930 );
and \U$835 ( \1084 , \902 , \928 );
nor \U$836 ( \1085 , \1083 , \1084 );
xnor \U$837 ( \1086 , \1085 , \937 );
and \U$838 ( \1087 , \912 , \950 );
and \U$839 ( \1088 , \932 , \948 );
nor \U$840 ( \1089 , \1087 , \1088 );
xnor \U$841 ( \1090 , \1089 , \957 );
xor \U$842 ( \1091 , \1086 , \1090 );
and \U$843 ( \1092 , \939 , \978 );
and \U$844 ( \1093 , \952 , \961 );
nor \U$845 ( \1094 , \1092 , \1093 );
xnor \U$846 ( \1095 , \1094 , \568 );
xor \U$847 ( \1096 , \1091 , \1095 );
xor \U$848 ( \1097 , \1082 , \1096 );
and \U$849 ( \1098 , \1073 , \1097 );
and \U$850 ( \1099 , \1029 , \1097 );
or \U$851 ( \1100 , \1074 , \1098 , \1099 );
and \U$852 ( \1101 , \1017 , \1100 );
and \U$853 ( \1102 , \532 , \1023 );
and \U$854 ( \1103 , \1023 , \1028 );
and \U$855 ( \1104 , \532 , \1028 );
or \U$856 ( \1105 , \1102 , \1103 , \1104 );
and \U$857 ( \1106 , \1062 , \1066 );
and \U$858 ( \1107 , \1066 , \1071 );
and \U$859 ( \1108 , \1062 , \1071 );
or \U$860 ( \1109 , \1106 , \1107 , \1108 );
xor \U$861 ( \1110 , \1105 , \1109 );
and \U$862 ( \1111 , \1047 , \1051 );
and \U$863 ( \1112 , \1051 , \1056 );
and \U$864 ( \1113 , \1047 , \1056 );
or \U$865 ( \1114 , \1111 , \1112 , \1113 );
xor \U$866 ( \1115 , \1110 , \1114 );
and \U$867 ( \1116 , \1100 , \1115 );
and \U$868 ( \1117 , \1017 , \1115 );
or \U$869 ( \1118 , \1101 , \1116 , \1117 );
and \U$870 ( \1119 , \1020 , \616 );
and \U$871 ( \1120 , \539 , \613 );
nor \U$872 ( \1121 , \1119 , \1120 );
xnor \U$873 ( \1122 , \1121 , \576 );
and \U$874 ( \1123 , \618 , \641 );
and \U$875 ( \1124 , \1018 , \639 );
nor \U$876 ( \1125 , \1123 , \1124 );
xnor \U$877 ( \1126 , \1125 , \648 );
xor \U$878 ( \1127 , \1122 , \1126 );
and \U$879 ( \1128 , \643 , \671 );
and \U$880 ( \1129 , \569 , \669 );
nor \U$881 ( \1130 , \1128 , \1129 );
xnor \U$882 ( \1131 , \1130 , \678 );
xor \U$883 ( \1132 , \1127 , \1131 );
and \U$884 ( \1133 , \847 , \872 );
and \U$885 ( \1134 , \794 , \870 );
nor \U$886 ( \1135 , \1133 , \1134 );
xnor \U$887 ( \1136 , \1135 , \879 );
and \U$888 ( \1137 , \874 , \900 );
and \U$889 ( \1138 , \827 , \898 );
nor \U$890 ( \1139 , \1137 , \1138 );
xnor \U$891 ( \1140 , \1139 , \907 );
xor \U$892 ( \1141 , \1136 , \1140 );
and \U$893 ( \1142 , \902 , \930 );
and \U$894 ( \1143 , \854 , \928 );
nor \U$895 ( \1144 , \1142 , \1143 );
xnor \U$896 ( \1145 , \1144 , \937 );
xor \U$897 ( \1146 , \1141 , \1145 );
and \U$898 ( \1147 , \759 , \784 );
and \U$899 ( \1148 , \708 , \782 );
nor \U$900 ( \1149 , \1147 , \1148 );
xnor \U$901 ( \1150 , \1149 , \791 );
and \U$902 ( \1151 , \786 , \812 );
and \U$903 ( \1152 , \739 , \810 );
nor \U$904 ( \1153 , \1151 , \1152 );
xnor \U$905 ( \1154 , \1153 , \819 );
xor \U$906 ( \1155 , \1150 , \1154 );
and \U$907 ( \1156 , \814 , \845 );
and \U$908 ( \1157 , \766 , \843 );
nor \U$909 ( \1158 , \1156 , \1157 );
xnor \U$910 ( \1159 , \1158 , \852 );
xor \U$911 ( \1160 , \1155 , \1159 );
xor \U$912 ( \1161 , \1146 , \1160 );
and \U$913 ( \1162 , \673 , \698 );
and \U$914 ( \1163 , \623 , \696 );
nor \U$915 ( \1164 , \1162 , \1163 );
xnor \U$916 ( \1165 , \1164 , \705 );
and \U$917 ( \1166 , \700 , \726 );
and \U$918 ( \1167 , \653 , \724 );
nor \U$919 ( \1168 , \1166 , \1167 );
xnor \U$920 ( \1169 , \1168 , \733 );
xor \U$921 ( \1170 , \1165 , \1169 );
and \U$922 ( \1171 , \728 , \757 );
and \U$923 ( \1172 , \680 , \755 );
nor \U$924 ( \1173 , \1171 , \1172 );
xnor \U$925 ( \1174 , \1173 , \764 );
xor \U$926 ( \1175 , \1170 , \1174 );
xor \U$927 ( \1176 , \1161 , \1175 );
xor \U$928 ( \1177 , \1132 , \1176 );
and \U$929 ( \1178 , \1033 , \1037 );
and \U$930 ( \1179 , \1037 , \1042 );
and \U$931 ( \1180 , \1033 , \1042 );
or \U$932 ( \1181 , \1178 , \1179 , \1180 );
and \U$933 ( \1182 , \1086 , \1090 );
and \U$934 ( \1183 , \1090 , \1095 );
and \U$935 ( \1184 , \1086 , \1095 );
or \U$936 ( \1185 , \1182 , \1183 , \1184 );
xor \U$937 ( \1186 , \1181 , \1185 );
and \U$938 ( \1187 , \932 , \950 );
and \U$939 ( \1188 , \882 , \948 );
nor \U$940 ( \1189 , \1187 , \1188 );
xnor \U$941 ( \1190 , \1189 , \957 );
and \U$942 ( \1191 , \952 , \978 );
and \U$943 ( \1192 , \912 , \961 );
nor \U$944 ( \1193 , \1191 , \1192 );
xnor \U$945 ( \1194 , \1193 , \568 );
xor \U$946 ( \1195 , \1190 , \1194 );
xor \U$947 ( \1196 , \494 , \522 );
not \U$948 ( \1197 , \1079 );
and \U$949 ( \1198 , \1196 , \1197 );
and \U$950 ( \1199 , \960 , \1198 );
and \U$951 ( \1200 , \939 , \1079 );
nor \U$952 ( \1201 , \1199 , \1200 );
xnor \U$953 ( \1202 , \1201 , \532 );
xor \U$954 ( \1203 , \1195 , \1202 );
xor \U$955 ( \1204 , \1186 , \1203 );
xor \U$956 ( \1205 , \1177 , \1204 );
and \U$957 ( \1206 , \618 , \616 );
and \U$958 ( \1207 , \1018 , \613 );
nor \U$959 ( \1208 , \1206 , \1207 );
xnor \U$960 ( \1209 , \1208 , \576 );
and \U$961 ( \1210 , \643 , \641 );
and \U$962 ( \1211 , \569 , \639 );
nor \U$963 ( \1212 , \1210 , \1211 );
xnor \U$964 ( \1213 , \1212 , \648 );
and \U$965 ( \1214 , \1209 , \1213 );
and \U$966 ( \1215 , \673 , \671 );
and \U$967 ( \1216 , \623 , \669 );
nor \U$968 ( \1217 , \1215 , \1216 );
xnor \U$969 ( \1218 , \1217 , \678 );
and \U$970 ( \1219 , \1213 , \1218 );
and \U$971 ( \1220 , \1209 , \1218 );
or \U$972 ( \1221 , \1214 , \1219 , \1220 );
and \U$973 ( \1222 , \700 , \698 );
and \U$974 ( \1223 , \653 , \696 );
nor \U$975 ( \1224 , \1222 , \1223 );
xnor \U$976 ( \1225 , \1224 , \705 );
and \U$977 ( \1226 , \728 , \726 );
and \U$978 ( \1227 , \680 , \724 );
nor \U$979 ( \1228 , \1226 , \1227 );
xnor \U$980 ( \1229 , \1228 , \733 );
and \U$981 ( \1230 , \1225 , \1229 );
and \U$982 ( \1231 , \759 , \757 );
and \U$983 ( \1232 , \708 , \755 );
nor \U$984 ( \1233 , \1231 , \1232 );
xnor \U$985 ( \1234 , \1233 , \764 );
and \U$986 ( \1235 , \1229 , \1234 );
and \U$987 ( \1236 , \1225 , \1234 );
or \U$988 ( \1237 , \1230 , \1235 , \1236 );
and \U$989 ( \1238 , \1221 , \1237 );
and \U$990 ( \1239 , \1001 , \1005 );
and \U$991 ( \1240 , \1005 , \1010 );
and \U$992 ( \1241 , \1001 , \1010 );
or \U$993 ( \1242 , \1239 , \1240 , \1241 );
and \U$994 ( \1243 , \1237 , \1242 );
and \U$995 ( \1244 , \1221 , \1242 );
or \U$996 ( \1245 , \1238 , \1243 , \1244 );
and \U$997 ( \1246 , \1078 , \1081 );
and \U$998 ( \1247 , \1081 , \1096 );
and \U$999 ( \1248 , \1078 , \1096 );
or \U$1000 ( \1249 , \1246 , \1247 , \1248 );
xor \U$1001 ( \1250 , \1245 , \1249 );
and \U$1002 ( \1251 , \1043 , \1057 );
and \U$1003 ( \1252 , \1057 , \1072 );
and \U$1004 ( \1253 , \1043 , \1072 );
or \U$1005 ( \1254 , \1251 , \1252 , \1253 );
xor \U$1006 ( \1255 , \1250 , \1254 );
and \U$1007 ( \1256 , \1205 , \1255 );
and \U$1008 ( \1257 , \1118 , \1256 );
and \U$1009 ( \1258 , \680 , \757 );
and \U$1010 ( \1259 , \700 , \755 );
nor \U$1011 ( \1260 , \1258 , \1259 );
xnor \U$1012 ( \1261 , \1260 , \764 );
and \U$1013 ( \1262 , \708 , \784 );
and \U$1014 ( \1263 , \728 , \782 );
nor \U$1015 ( \1264 , \1262 , \1263 );
xnor \U$1016 ( \1265 , \1264 , \791 );
xor \U$1017 ( \1266 , \1261 , \1265 );
and \U$1018 ( \1267 , \739 , \812 );
and \U$1019 ( \1268 , \759 , \810 );
nor \U$1020 ( \1269 , \1267 , \1268 );
xnor \U$1021 ( \1270 , \1269 , \819 );
xor \U$1022 ( \1271 , \1266 , \1270 );
and \U$1023 ( \1272 , \569 , \671 );
and \U$1024 ( \1273 , \618 , \669 );
nor \U$1025 ( \1274 , \1272 , \1273 );
xnor \U$1026 ( \1275 , \1274 , \678 );
and \U$1027 ( \1276 , \623 , \698 );
and \U$1028 ( \1277 , \643 , \696 );
nor \U$1029 ( \1278 , \1276 , \1277 );
xnor \U$1030 ( \1279 , \1278 , \705 );
xor \U$1031 ( \1280 , \1275 , \1279 );
and \U$1032 ( \1281 , \653 , \726 );
and \U$1033 ( \1282 , \673 , \724 );
nor \U$1034 ( \1283 , \1281 , \1282 );
xnor \U$1035 ( \1284 , \1283 , \733 );
xor \U$1036 ( \1285 , \1280 , \1284 );
xor \U$1037 ( \1286 , \1271 , \1285 );
and \U$1038 ( \1287 , \539 , \616 );
and \U$1039 ( \1288 , \504 , \613 );
nor \U$1040 ( \1289 , \1287 , \1288 );
xnor \U$1041 ( \1290 , \1289 , \576 );
xor \U$1042 ( \1291 , \502 , \1290 );
and \U$1043 ( \1292 , \1018 , \641 );
and \U$1044 ( \1293 , \1020 , \639 );
nor \U$1045 ( \1294 , \1292 , \1293 );
xnor \U$1046 ( \1295 , \1294 , \648 );
xor \U$1047 ( \1296 , \1291 , \1295 );
xor \U$1048 ( \1297 , \1286 , \1296 );
nand \U$1049 ( \1298 , \960 , \495 );
xnor \U$1050 ( \1299 , \1298 , \502 );
and \U$1051 ( \1300 , \854 , \930 );
and \U$1052 ( \1301 , \874 , \928 );
nor \U$1053 ( \1302 , \1300 , \1301 );
xnor \U$1054 ( \1303 , \1302 , \937 );
and \U$1055 ( \1304 , \882 , \950 );
and \U$1056 ( \1305 , \902 , \948 );
nor \U$1057 ( \1306 , \1304 , \1305 );
xnor \U$1058 ( \1307 , \1306 , \957 );
xor \U$1059 ( \1308 , \1303 , \1307 );
and \U$1060 ( \1309 , \912 , \978 );
and \U$1061 ( \1310 , \932 , \961 );
nor \U$1062 ( \1311 , \1309 , \1310 );
xnor \U$1063 ( \1312 , \1311 , \568 );
xor \U$1064 ( \1313 , \1308 , \1312 );
xor \U$1065 ( \1314 , \1299 , \1313 );
and \U$1066 ( \1315 , \766 , \845 );
and \U$1067 ( \1316 , \786 , \843 );
nor \U$1068 ( \1317 , \1315 , \1316 );
xnor \U$1069 ( \1318 , \1317 , \852 );
and \U$1070 ( \1319 , \794 , \872 );
and \U$1071 ( \1320 , \814 , \870 );
nor \U$1072 ( \1321 , \1319 , \1320 );
xnor \U$1073 ( \1322 , \1321 , \879 );
xor \U$1074 ( \1323 , \1318 , \1322 );
and \U$1075 ( \1324 , \827 , \900 );
and \U$1076 ( \1325 , \847 , \898 );
nor \U$1077 ( \1326 , \1324 , \1325 );
xnor \U$1078 ( \1327 , \1326 , \907 );
xor \U$1079 ( \1328 , \1323 , \1327 );
xor \U$1080 ( \1329 , \1314 , \1328 );
xor \U$1081 ( \1330 , \1297 , \1329 );
and \U$1082 ( \1331 , \1136 , \1140 );
and \U$1083 ( \1332 , \1140 , \1145 );
and \U$1084 ( \1333 , \1136 , \1145 );
or \U$1085 ( \1334 , \1331 , \1332 , \1333 );
and \U$1086 ( \1335 , \1190 , \1194 );
and \U$1087 ( \1336 , \1194 , \1202 );
and \U$1088 ( \1337 , \1190 , \1202 );
or \U$1089 ( \1338 , \1335 , \1336 , \1337 );
xor \U$1090 ( \1339 , \1334 , \1338 );
and \U$1091 ( \1340 , \939 , \1198 );
and \U$1092 ( \1341 , \952 , \1079 );
nor \U$1093 ( \1342 , \1340 , \1341 );
xnor \U$1094 ( \1343 , \1342 , \532 );
xor \U$1095 ( \1344 , \1339 , \1343 );
xor \U$1096 ( \1345 , \1330 , \1344 );
and \U$1097 ( \1346 , \1256 , \1345 );
and \U$1098 ( \1347 , \1118 , \1345 );
or \U$1099 ( \1348 , \1257 , \1346 , \1347 );
and \U$1100 ( \1349 , \1105 , \1109 );
and \U$1101 ( \1350 , \1109 , \1114 );
and \U$1102 ( \1351 , \1105 , \1114 );
or \U$1103 ( \1352 , \1349 , \1350 , \1351 );
and \U$1104 ( \1353 , \1181 , \1185 );
and \U$1105 ( \1354 , \1185 , \1203 );
and \U$1106 ( \1355 , \1181 , \1203 );
or \U$1107 ( \1356 , \1353 , \1354 , \1355 );
xor \U$1108 ( \1357 , \1352 , \1356 );
and \U$1109 ( \1358 , \1146 , \1160 );
and \U$1110 ( \1359 , \1160 , \1175 );
and \U$1111 ( \1360 , \1146 , \1175 );
or \U$1112 ( \1361 , \1358 , \1359 , \1360 );
xor \U$1113 ( \1362 , \1357 , \1361 );
and \U$1114 ( \1363 , \1245 , \1249 );
and \U$1115 ( \1364 , \1249 , \1254 );
and \U$1116 ( \1365 , \1245 , \1254 );
or \U$1117 ( \1366 , \1363 , \1364 , \1365 );
and \U$1118 ( \1367 , \1132 , \1176 );
and \U$1119 ( \1368 , \1176 , \1204 );
and \U$1120 ( \1369 , \1132 , \1204 );
or \U$1121 ( \1370 , \1367 , \1368 , \1369 );
xor \U$1122 ( \1371 , \1366 , \1370 );
and \U$1123 ( \1372 , \1122 , \1126 );
and \U$1124 ( \1373 , \1126 , \1131 );
and \U$1125 ( \1374 , \1122 , \1131 );
or \U$1126 ( \1375 , \1372 , \1373 , \1374 );
and \U$1127 ( \1376 , \1165 , \1169 );
and \U$1128 ( \1377 , \1169 , \1174 );
and \U$1129 ( \1378 , \1165 , \1174 );
or \U$1130 ( \1379 , \1376 , \1377 , \1378 );
xor \U$1131 ( \1380 , \1375 , \1379 );
and \U$1132 ( \1381 , \1150 , \1154 );
and \U$1133 ( \1382 , \1154 , \1159 );
and \U$1134 ( \1383 , \1150 , \1159 );
or \U$1135 ( \1384 , \1381 , \1382 , \1383 );
xor \U$1136 ( \1385 , \1380 , \1384 );
xor \U$1137 ( \1386 , \1371 , \1385 );
and \U$1138 ( \1387 , \1362 , \1386 );
xor \U$1139 ( \1388 , \1348 , \1387 );
and \U$1140 ( \1389 , \1366 , \1370 );
and \U$1141 ( \1390 , \1370 , \1385 );
and \U$1142 ( \1391 , \1366 , \1385 );
or \U$1143 ( \1392 , \1389 , \1390 , \1391 );
and \U$1144 ( \1393 , \1271 , \1285 );
and \U$1145 ( \1394 , \1285 , \1296 );
and \U$1146 ( \1395 , \1271 , \1296 );
or \U$1147 ( \1396 , \1393 , \1394 , \1395 );
and \U$1148 ( \1397 , \643 , \698 );
and \U$1149 ( \1398 , \569 , \696 );
nor \U$1150 ( \1399 , \1397 , \1398 );
xnor \U$1151 ( \1400 , \1399 , \705 );
and \U$1152 ( \1401 , \673 , \726 );
and \U$1153 ( \1402 , \623 , \724 );
nor \U$1154 ( \1403 , \1401 , \1402 );
xnor \U$1155 ( \1404 , \1403 , \733 );
xor \U$1156 ( \1405 , \1400 , \1404 );
and \U$1157 ( \1406 , \700 , \757 );
and \U$1158 ( \1407 , \653 , \755 );
nor \U$1159 ( \1408 , \1406 , \1407 );
xnor \U$1160 ( \1409 , \1408 , \764 );
xor \U$1161 ( \1410 , \1405 , \1409 );
xor \U$1162 ( \1411 , \1396 , \1410 );
and \U$1163 ( \1412 , \504 , \616 );
and \U$1164 ( \1413 , \223 , \613 );
nor \U$1165 ( \1414 , \1412 , \1413 );
xnor \U$1166 ( \1415 , \1414 , \576 );
and \U$1167 ( \1416 , \1020 , \641 );
and \U$1168 ( \1417 , \539 , \639 );
nor \U$1169 ( \1418 , \1416 , \1417 );
xnor \U$1170 ( \1419 , \1418 , \648 );
xor \U$1171 ( \1420 , \1415 , \1419 );
and \U$1172 ( \1421 , \618 , \671 );
and \U$1173 ( \1422 , \1018 , \669 );
nor \U$1174 ( \1423 , \1421 , \1422 );
xnor \U$1175 ( \1424 , \1423 , \678 );
xor \U$1176 ( \1425 , \1420 , \1424 );
xor \U$1177 ( \1426 , \1411 , \1425 );
and \U$1178 ( \1427 , \1375 , \1379 );
and \U$1179 ( \1428 , \1379 , \1384 );
and \U$1180 ( \1429 , \1375 , \1384 );
or \U$1181 ( \1430 , \1427 , \1428 , \1429 );
and \U$1182 ( \1431 , \1334 , \1338 );
and \U$1183 ( \1432 , \1338 , \1343 );
and \U$1184 ( \1433 , \1334 , \1343 );
or \U$1185 ( \1434 , \1431 , \1432 , \1433 );
xor \U$1186 ( \1435 , \1430 , \1434 );
and \U$1187 ( \1436 , \1299 , \1313 );
and \U$1188 ( \1437 , \1313 , \1328 );
and \U$1189 ( \1438 , \1299 , \1328 );
or \U$1190 ( \1439 , \1436 , \1437 , \1438 );
xor \U$1191 ( \1440 , \1435 , \1439 );
xor \U$1192 ( \1441 , \1426 , \1440 );
xor \U$1193 ( \1442 , \1392 , \1441 );
and \U$1194 ( \1443 , \1352 , \1356 );
and \U$1195 ( \1444 , \1356 , \1361 );
and \U$1196 ( \1445 , \1352 , \1361 );
or \U$1197 ( \1446 , \1443 , \1444 , \1445 );
and \U$1198 ( \1447 , \1297 , \1329 );
and \U$1199 ( \1448 , \1329 , \1344 );
and \U$1200 ( \1449 , \1297 , \1344 );
or \U$1201 ( \1450 , \1447 , \1448 , \1449 );
xor \U$1202 ( \1451 , \1446 , \1450 );
and \U$1203 ( \1452 , \902 , \950 );
and \U$1204 ( \1453 , \854 , \948 );
nor \U$1205 ( \1454 , \1452 , \1453 );
xnor \U$1206 ( \1455 , \1454 , \957 );
and \U$1207 ( \1456 , \932 , \978 );
and \U$1208 ( \1457 , \882 , \961 );
nor \U$1209 ( \1458 , \1456 , \1457 );
xnor \U$1210 ( \1459 , \1458 , \568 );
xor \U$1211 ( \1460 , \1455 , \1459 );
and \U$1212 ( \1461 , \952 , \1198 );
and \U$1213 ( \1462 , \912 , \1079 );
nor \U$1214 ( \1463 , \1461 , \1462 );
xnor \U$1215 ( \1464 , \1463 , \532 );
xor \U$1216 ( \1465 , \1460 , \1464 );
and \U$1217 ( \1466 , \814 , \872 );
and \U$1218 ( \1467 , \766 , \870 );
nor \U$1219 ( \1468 , \1466 , \1467 );
xnor \U$1220 ( \1469 , \1468 , \879 );
and \U$1221 ( \1470 , \847 , \900 );
and \U$1222 ( \1471 , \794 , \898 );
nor \U$1223 ( \1472 , \1470 , \1471 );
xnor \U$1224 ( \1473 , \1472 , \907 );
xor \U$1225 ( \1474 , \1469 , \1473 );
and \U$1226 ( \1475 , \874 , \930 );
and \U$1227 ( \1476 , \827 , \928 );
nor \U$1228 ( \1477 , \1475 , \1476 );
xnor \U$1229 ( \1478 , \1477 , \937 );
xor \U$1230 ( \1479 , \1474 , \1478 );
xor \U$1231 ( \1480 , \1465 , \1479 );
and \U$1232 ( \1481 , \728 , \784 );
and \U$1233 ( \1482 , \680 , \782 );
nor \U$1234 ( \1483 , \1481 , \1482 );
xnor \U$1235 ( \1484 , \1483 , \791 );
and \U$1236 ( \1485 , \759 , \812 );
and \U$1237 ( \1486 , \708 , \810 );
nor \U$1238 ( \1487 , \1485 , \1486 );
xnor \U$1239 ( \1488 , \1487 , \819 );
xor \U$1240 ( \1489 , \1484 , \1488 );
and \U$1241 ( \1490 , \786 , \845 );
and \U$1242 ( \1491 , \739 , \843 );
nor \U$1243 ( \1492 , \1490 , \1491 );
xnor \U$1244 ( \1493 , \1492 , \852 );
xor \U$1245 ( \1494 , \1489 , \1493 );
xor \U$1246 ( \1495 , \1480 , \1494 );
and \U$1247 ( \1496 , \1318 , \1322 );
and \U$1248 ( \1497 , \1322 , \1327 );
and \U$1249 ( \1498 , \1318 , \1327 );
or \U$1250 ( \1499 , \1496 , \1497 , \1498 );
and \U$1251 ( \1500 , \1303 , \1307 );
and \U$1252 ( \1501 , \1307 , \1312 );
and \U$1253 ( \1502 , \1303 , \1312 );
or \U$1254 ( \1503 , \1500 , \1501 , \1502 );
xor \U$1255 ( \1504 , \1499 , \1503 );
and \U$1256 ( \1505 , \960 , \497 );
and \U$1257 ( \1506 , \939 , \495 );
nor \U$1258 ( \1507 , \1505 , \1506 );
xnor \U$1259 ( \1508 , \1507 , \502 );
xor \U$1260 ( \1509 , \1504 , \1508 );
xor \U$1261 ( \1510 , \1495 , \1509 );
and \U$1262 ( \1511 , \502 , \1290 );
and \U$1263 ( \1512 , \1290 , \1295 );
and \U$1264 ( \1513 , \502 , \1295 );
or \U$1265 ( \1514 , \1511 , \1512 , \1513 );
and \U$1266 ( \1515 , \1275 , \1279 );
and \U$1267 ( \1516 , \1279 , \1284 );
and \U$1268 ( \1517 , \1275 , \1284 );
or \U$1269 ( \1518 , \1515 , \1516 , \1517 );
xor \U$1270 ( \1519 , \1514 , \1518 );
and \U$1271 ( \1520 , \1261 , \1265 );
and \U$1272 ( \1521 , \1265 , \1270 );
and \U$1273 ( \1522 , \1261 , \1270 );
or \U$1274 ( \1523 , \1520 , \1521 , \1522 );
xor \U$1275 ( \1524 , \1519 , \1523 );
xor \U$1276 ( \1525 , \1510 , \1524 );
xor \U$1277 ( \1526 , \1451 , \1525 );
xor \U$1278 ( \1527 , \1442 , \1526 );
xor \U$1279 ( \1528 , \1388 , \1527 );
and \U$1280 ( \1529 , \643 , \616 );
and \U$1281 ( \1530 , \569 , \613 );
nor \U$1282 ( \1531 , \1529 , \1530 );
xnor \U$1283 ( \1532 , \1531 , \576 );
and \U$1284 ( \1533 , \673 , \641 );
and \U$1285 ( \1534 , \623 , \639 );
nor \U$1286 ( \1535 , \1533 , \1534 );
xnor \U$1287 ( \1536 , \1535 , \648 );
and \U$1288 ( \1537 , \1532 , \1536 );
and \U$1289 ( \1538 , \700 , \671 );
and \U$1290 ( \1539 , \653 , \669 );
nor \U$1291 ( \1540 , \1538 , \1539 );
xnor \U$1292 ( \1541 , \1540 , \678 );
and \U$1293 ( \1542 , \1536 , \1541 );
and \U$1294 ( \1543 , \1532 , \1541 );
or \U$1295 ( \1544 , \1537 , \1542 , \1543 );
and \U$1296 ( \1545 , \728 , \698 );
and \U$1297 ( \1546 , \680 , \696 );
nor \U$1298 ( \1547 , \1545 , \1546 );
xnor \U$1299 ( \1548 , \1547 , \705 );
and \U$1300 ( \1549 , \759 , \726 );
and \U$1301 ( \1550 , \708 , \724 );
nor \U$1302 ( \1551 , \1549 , \1550 );
xnor \U$1303 ( \1552 , \1551 , \733 );
and \U$1304 ( \1553 , \1548 , \1552 );
and \U$1305 ( \1554 , \786 , \757 );
and \U$1306 ( \1555 , \739 , \755 );
nor \U$1307 ( \1556 , \1554 , \1555 );
xnor \U$1308 ( \1557 , \1556 , \764 );
and \U$1309 ( \1558 , \1552 , \1557 );
and \U$1310 ( \1559 , \1548 , \1557 );
or \U$1311 ( \1560 , \1553 , \1558 , \1559 );
and \U$1312 ( \1561 , \1544 , \1560 );
and \U$1313 ( \1562 , \814 , \784 );
and \U$1314 ( \1563 , \766 , \782 );
nor \U$1315 ( \1564 , \1562 , \1563 );
xnor \U$1316 ( \1565 , \1564 , \791 );
and \U$1317 ( \1566 , \847 , \812 );
and \U$1318 ( \1567 , \794 , \810 );
nor \U$1319 ( \1568 , \1566 , \1567 );
xnor \U$1320 ( \1569 , \1568 , \819 );
and \U$1321 ( \1570 , \1565 , \1569 );
and \U$1322 ( \1571 , \874 , \845 );
and \U$1323 ( \1572 , \827 , \843 );
nor \U$1324 ( \1573 , \1571 , \1572 );
xnor \U$1325 ( \1574 , \1573 , \852 );
and \U$1326 ( \1575 , \1569 , \1574 );
and \U$1327 ( \1576 , \1565 , \1574 );
or \U$1328 ( \1577 , \1570 , \1575 , \1576 );
and \U$1329 ( \1578 , \1560 , \1577 );
and \U$1330 ( \1579 , \1544 , \1577 );
or \U$1331 ( \1580 , \1561 , \1578 , \1579 );
and \U$1332 ( \1581 , \902 , \872 );
and \U$1333 ( \1582 , \854 , \870 );
nor \U$1334 ( \1583 , \1581 , \1582 );
xnor \U$1335 ( \1584 , \1583 , \879 );
and \U$1336 ( \1585 , \932 , \900 );
and \U$1337 ( \1586 , \882 , \898 );
nor \U$1338 ( \1587 , \1585 , \1586 );
xnor \U$1339 ( \1588 , \1587 , \907 );
and \U$1340 ( \1589 , \1584 , \1588 );
and \U$1341 ( \1590 , \952 , \930 );
and \U$1342 ( \1591 , \912 , \928 );
nor \U$1343 ( \1592 , \1590 , \1591 );
xnor \U$1344 ( \1593 , \1592 , \937 );
and \U$1345 ( \1594 , \1588 , \1593 );
and \U$1346 ( \1595 , \1584 , \1593 );
or \U$1347 ( \1596 , \1589 , \1594 , \1595 );
xor \U$1348 ( \1597 , \938 , \958 );
xor \U$1349 ( \1598 , \1597 , \963 );
and \U$1350 ( \1599 , \1596 , \1598 );
xor \U$1351 ( \1600 , \853 , \880 );
xor \U$1352 ( \1601 , \1600 , \908 );
and \U$1353 ( \1602 , \1598 , \1601 );
and \U$1354 ( \1603 , \1596 , \1601 );
or \U$1355 ( \1604 , \1599 , \1602 , \1603 );
and \U$1356 ( \1605 , \1580 , \1604 );
xor \U$1357 ( \1606 , \765 , \792 );
xor \U$1358 ( \1607 , \1606 , \820 );
xor \U$1359 ( \1608 , \679 , \706 );
xor \U$1360 ( \1609 , \1608 , \734 );
and \U$1361 ( \1610 , \1607 , \1609 );
xor \U$1362 ( \1611 , \568 , \621 );
xor \U$1363 ( \1612 , \1611 , \649 );
and \U$1364 ( \1613 , \1609 , \1612 );
and \U$1365 ( \1614 , \1607 , \1612 );
or \U$1366 ( \1615 , \1610 , \1613 , \1614 );
and \U$1367 ( \1616 , \1604 , \1615 );
and \U$1368 ( \1617 , \1580 , \1615 );
or \U$1369 ( \1618 , \1605 , \1616 , \1617 );
xor \U$1370 ( \1619 , \1225 , \1229 );
xor \U$1371 ( \1620 , \1619 , \1234 );
xor \U$1372 ( \1621 , \1209 , \1213 );
xor \U$1373 ( \1622 , \1621 , \1218 );
and \U$1374 ( \1623 , \1620 , \1622 );
xor \U$1375 ( \1624 , \982 , \996 );
xor \U$1376 ( \1625 , \1624 , \1011 );
and \U$1377 ( \1626 , \1622 , \1625 );
and \U$1378 ( \1627 , \1620 , \1625 );
or \U$1379 ( \1628 , \1623 , \1626 , \1627 );
and \U$1380 ( \1629 , \1618 , \1628 );
xor \U$1381 ( \1630 , \1221 , \1237 );
xor \U$1382 ( \1631 , \1630 , \1242 );
and \U$1383 ( \1632 , \1628 , \1631 );
and \U$1384 ( \1633 , \1618 , \1631 );
or \U$1385 ( \1634 , \1629 , \1632 , \1633 );
xor \U$1386 ( \1635 , \1205 , \1255 );
and \U$1387 ( \1636 , \1634 , \1635 );
xor \U$1388 ( \1637 , \1017 , \1100 );
xor \U$1389 ( \1638 , \1637 , \1115 );
and \U$1390 ( \1639 , \1635 , \1638 );
and \U$1391 ( \1640 , \1634 , \1638 );
or \U$1392 ( \1641 , \1636 , \1639 , \1640 );
xor \U$1393 ( \1642 , \1362 , \1386 );
and \U$1394 ( \1643 , \1641 , \1642 );
xor \U$1395 ( \1644 , \1118 , \1256 );
xor \U$1396 ( \1645 , \1644 , \1345 );
and \U$1397 ( \1646 , \1642 , \1645 );
and \U$1398 ( \1647 , \1641 , \1645 );
or \U$1399 ( \1648 , \1643 , \1646 , \1647 );
nor \U$1400 ( \1649 , \1528 , \1648 );
and \U$1401 ( \1650 , \1392 , \1441 );
and \U$1402 ( \1651 , \1441 , \1526 );
and \U$1403 ( \1652 , \1392 , \1526 );
or \U$1404 ( \1653 , \1650 , \1651 , \1652 );
and \U$1405 ( \1654 , \1430 , \1434 );
and \U$1406 ( \1655 , \1434 , \1439 );
and \U$1407 ( \1656 , \1430 , \1439 );
or \U$1408 ( \1657 , \1654 , \1655 , \1656 );
and \U$1409 ( \1658 , \1396 , \1410 );
and \U$1410 ( \1659 , \1410 , \1425 );
and \U$1411 ( \1660 , \1396 , \1425 );
or \U$1412 ( \1661 , \1658 , \1659 , \1660 );
xor \U$1413 ( \1662 , \1657 , \1661 );
and \U$1414 ( \1663 , \1495 , \1509 );
and \U$1415 ( \1664 , \1509 , \1524 );
and \U$1416 ( \1665 , \1495 , \1524 );
or \U$1417 ( \1666 , \1663 , \1664 , \1665 );
xor \U$1418 ( \1667 , \1662 , \1666 );
xor \U$1419 ( \1668 , \1653 , \1667 );
and \U$1420 ( \1669 , \1446 , \1450 );
and \U$1421 ( \1670 , \1450 , \1525 );
and \U$1422 ( \1671 , \1446 , \1525 );
or \U$1423 ( \1672 , \1669 , \1670 , \1671 );
and \U$1424 ( \1673 , \1426 , \1440 );
xor \U$1425 ( \1674 , \1672 , \1673 );
and \U$1426 ( \1675 , \1469 , \1473 );
and \U$1427 ( \1676 , \1473 , \1478 );
and \U$1428 ( \1677 , \1469 , \1478 );
or \U$1429 ( \1678 , \1675 , \1676 , \1677 );
and \U$1430 ( \1679 , \1455 , \1459 );
and \U$1431 ( \1680 , \1459 , \1464 );
and \U$1432 ( \1681 , \1455 , \1464 );
or \U$1433 ( \1682 , \1679 , \1680 , \1681 );
xor \U$1434 ( \1683 , \1678 , \1682 );
and \U$1435 ( \1684 , \912 , \1198 );
and \U$1436 ( \1685 , \932 , \1079 );
nor \U$1437 ( \1686 , \1684 , \1685 );
xnor \U$1438 ( \1687 , \1686 , \532 );
and \U$1439 ( \1688 , \939 , \497 );
and \U$1440 ( \1689 , \952 , \495 );
nor \U$1441 ( \1690 , \1688 , \1689 );
xnor \U$1442 ( \1691 , \1690 , \502 );
xor \U$1443 ( \1692 , \1687 , \1691 );
nand \U$1444 ( \1693 , \960 , \505 );
not \U$1445 ( \1694 , \1693 );
xor \U$1446 ( \1695 , \1692 , \1694 );
xor \U$1447 ( \1696 , \1683 , \1695 );
and \U$1448 ( \1697 , \1415 , \1419 );
and \U$1449 ( \1698 , \1419 , \1424 );
and \U$1450 ( \1699 , \1415 , \1424 );
or \U$1451 ( \1700 , \1697 , \1698 , \1699 );
and \U$1452 ( \1701 , \1400 , \1404 );
and \U$1453 ( \1702 , \1404 , \1409 );
and \U$1454 ( \1703 , \1400 , \1409 );
or \U$1455 ( \1704 , \1701 , \1702 , \1703 );
xor \U$1456 ( \1705 , \1700 , \1704 );
and \U$1457 ( \1706 , \1484 , \1488 );
and \U$1458 ( \1707 , \1488 , \1493 );
and \U$1459 ( \1708 , \1484 , \1493 );
or \U$1460 ( \1709 , \1706 , \1707 , \1708 );
xor \U$1461 ( \1710 , \1705 , \1709 );
xor \U$1462 ( \1711 , \1696 , \1710 );
and \U$1463 ( \1712 , \1018 , \671 );
and \U$1464 ( \1713 , \1020 , \669 );
nor \U$1465 ( \1714 , \1712 , \1713 );
xnor \U$1466 ( \1715 , \1714 , \678 );
and \U$1467 ( \1716 , \569 , \698 );
and \U$1468 ( \1717 , \618 , \696 );
nor \U$1469 ( \1718 , \1716 , \1717 );
xnor \U$1470 ( \1719 , \1718 , \705 );
xor \U$1471 ( \1720 , \1715 , \1719 );
and \U$1472 ( \1721 , \623 , \726 );
and \U$1473 ( \1722 , \643 , \724 );
nor \U$1474 ( \1723 , \1721 , \1722 );
xnor \U$1475 ( \1724 , \1723 , \733 );
xor \U$1476 ( \1725 , \1720 , \1724 );
and \U$1477 ( \1726 , \223 , \616 );
not \U$1478 ( \1727 , \1726 );
xnor \U$1479 ( \1728 , \1727 , \576 );
and \U$1480 ( \1729 , \539 , \641 );
and \U$1481 ( \1730 , \504 , \639 );
nor \U$1482 ( \1731 , \1729 , \1730 );
xnor \U$1483 ( \1732 , \1731 , \648 );
xor \U$1484 ( \1733 , \1728 , \1732 );
xor \U$1485 ( \1734 , \1725 , \1733 );
and \U$1486 ( \1735 , \827 , \930 );
and \U$1487 ( \1736 , \847 , \928 );
nor \U$1488 ( \1737 , \1735 , \1736 );
xnor \U$1489 ( \1738 , \1737 , \937 );
and \U$1490 ( \1739 , \854 , \950 );
and \U$1491 ( \1740 , \874 , \948 );
nor \U$1492 ( \1741 , \1739 , \1740 );
xnor \U$1493 ( \1742 , \1741 , \957 );
xor \U$1494 ( \1743 , \1738 , \1742 );
and \U$1495 ( \1744 , \882 , \978 );
and \U$1496 ( \1745 , \902 , \961 );
nor \U$1497 ( \1746 , \1744 , \1745 );
xnor \U$1498 ( \1747 , \1746 , \568 );
xor \U$1499 ( \1748 , \1743 , \1747 );
and \U$1500 ( \1749 , \739 , \845 );
and \U$1501 ( \1750 , \759 , \843 );
nor \U$1502 ( \1751 , \1749 , \1750 );
xnor \U$1503 ( \1752 , \1751 , \852 );
and \U$1504 ( \1753 , \766 , \872 );
and \U$1505 ( \1754 , \786 , \870 );
nor \U$1506 ( \1755 , \1753 , \1754 );
xnor \U$1507 ( \1756 , \1755 , \879 );
xor \U$1508 ( \1757 , \1752 , \1756 );
and \U$1509 ( \1758 , \794 , \900 );
and \U$1510 ( \1759 , \814 , \898 );
nor \U$1511 ( \1760 , \1758 , \1759 );
xnor \U$1512 ( \1761 , \1760 , \907 );
xor \U$1513 ( \1762 , \1757 , \1761 );
xor \U$1514 ( \1763 , \1748 , \1762 );
and \U$1515 ( \1764 , \653 , \757 );
and \U$1516 ( \1765 , \673 , \755 );
nor \U$1517 ( \1766 , \1764 , \1765 );
xnor \U$1518 ( \1767 , \1766 , \764 );
and \U$1519 ( \1768 , \680 , \784 );
and \U$1520 ( \1769 , \700 , \782 );
nor \U$1521 ( \1770 , \1768 , \1769 );
xnor \U$1522 ( \1771 , \1770 , \791 );
xor \U$1523 ( \1772 , \1767 , \1771 );
and \U$1524 ( \1773 , \708 , \812 );
and \U$1525 ( \1774 , \728 , \810 );
nor \U$1526 ( \1775 , \1773 , \1774 );
xnor \U$1527 ( \1776 , \1775 , \819 );
xor \U$1528 ( \1777 , \1772 , \1776 );
xor \U$1529 ( \1778 , \1763 , \1777 );
xor \U$1530 ( \1779 , \1734 , \1778 );
xor \U$1531 ( \1780 , \1711 , \1779 );
and \U$1532 ( \1781 , \1514 , \1518 );
and \U$1533 ( \1782 , \1518 , \1523 );
and \U$1534 ( \1783 , \1514 , \1523 );
or \U$1535 ( \1784 , \1781 , \1782 , \1783 );
and \U$1536 ( \1785 , \1499 , \1503 );
and \U$1537 ( \1786 , \1503 , \1508 );
and \U$1538 ( \1787 , \1499 , \1508 );
or \U$1539 ( \1788 , \1785 , \1786 , \1787 );
xor \U$1540 ( \1789 , \1784 , \1788 );
and \U$1541 ( \1790 , \1465 , \1479 );
and \U$1542 ( \1791 , \1479 , \1494 );
and \U$1543 ( \1792 , \1465 , \1494 );
or \U$1544 ( \1793 , \1790 , \1791 , \1792 );
xor \U$1545 ( \1794 , \1789 , \1793 );
xor \U$1546 ( \1795 , \1780 , \1794 );
xor \U$1547 ( \1796 , \1674 , \1795 );
xor \U$1548 ( \1797 , \1668 , \1796 );
and \U$1549 ( \1798 , \1348 , \1387 );
and \U$1550 ( \1799 , \1387 , \1527 );
and \U$1551 ( \1800 , \1348 , \1527 );
or \U$1552 ( \1801 , \1798 , \1799 , \1800 );
nor \U$1553 ( \1802 , \1797 , \1801 );
nor \U$1554 ( \1803 , \1649 , \1802 );
and \U$1555 ( \1804 , \1672 , \1673 );
and \U$1556 ( \1805 , \1673 , \1795 );
and \U$1557 ( \1806 , \1672 , \1795 );
or \U$1558 ( \1807 , \1804 , \1805 , \1806 );
and \U$1559 ( \1808 , \1784 , \1788 );
and \U$1560 ( \1809 , \1788 , \1793 );
and \U$1561 ( \1810 , \1784 , \1793 );
or \U$1562 ( \1811 , \1808 , \1809 , \1810 );
and \U$1563 ( \1812 , \1725 , \1733 );
and \U$1564 ( \1813 , \1733 , \1778 );
and \U$1565 ( \1814 , \1725 , \1778 );
or \U$1566 ( \1815 , \1812 , \1813 , \1814 );
xor \U$1567 ( \1816 , \1811 , \1815 );
and \U$1568 ( \1817 , \1696 , \1710 );
xor \U$1569 ( \1818 , \1816 , \1817 );
xor \U$1570 ( \1819 , \1807 , \1818 );
and \U$1571 ( \1820 , \1657 , \1661 );
and \U$1572 ( \1821 , \1661 , \1666 );
and \U$1573 ( \1822 , \1657 , \1666 );
or \U$1574 ( \1823 , \1820 , \1821 , \1822 );
and \U$1575 ( \1824 , \1711 , \1779 );
and \U$1576 ( \1825 , \1779 , \1794 );
and \U$1577 ( \1826 , \1711 , \1794 );
or \U$1578 ( \1827 , \1824 , \1825 , \1826 );
xor \U$1579 ( \1828 , \1823 , \1827 );
and \U$1580 ( \1829 , \1728 , \1732 );
and \U$1581 ( \1830 , \1715 , \1719 );
and \U$1582 ( \1831 , \1719 , \1724 );
and \U$1583 ( \1832 , \1715 , \1724 );
or \U$1584 ( \1833 , \1830 , \1831 , \1832 );
xor \U$1585 ( \1834 , \1829 , \1833 );
and \U$1586 ( \1835 , \1767 , \1771 );
and \U$1587 ( \1836 , \1771 , \1776 );
and \U$1588 ( \1837 , \1767 , \1776 );
or \U$1589 ( \1838 , \1835 , \1836 , \1837 );
xor \U$1590 ( \1839 , \1834 , \1838 );
and \U$1591 ( \1840 , \700 , \784 );
and \U$1592 ( \1841 , \653 , \782 );
nor \U$1593 ( \1842 , \1840 , \1841 );
xnor \U$1594 ( \1843 , \1842 , \791 );
and \U$1595 ( \1844 , \728 , \812 );
and \U$1596 ( \1845 , \680 , \810 );
nor \U$1597 ( \1846 , \1844 , \1845 );
xnor \U$1598 ( \1847 , \1846 , \819 );
xor \U$1599 ( \1848 , \1843 , \1847 );
and \U$1600 ( \1849 , \759 , \845 );
and \U$1601 ( \1850 , \708 , \843 );
nor \U$1602 ( \1851 , \1849 , \1850 );
xnor \U$1603 ( \1852 , \1851 , \852 );
xor \U$1604 ( \1853 , \1848 , \1852 );
and \U$1605 ( \1854 , \618 , \698 );
and \U$1606 ( \1855 , \1018 , \696 );
nor \U$1607 ( \1856 , \1854 , \1855 );
xnor \U$1608 ( \1857 , \1856 , \705 );
and \U$1609 ( \1858 , \643 , \726 );
and \U$1610 ( \1859 , \569 , \724 );
nor \U$1611 ( \1860 , \1858 , \1859 );
xnor \U$1612 ( \1861 , \1860 , \733 );
xor \U$1613 ( \1862 , \1857 , \1861 );
and \U$1614 ( \1863 , \673 , \757 );
and \U$1615 ( \1864 , \623 , \755 );
nor \U$1616 ( \1865 , \1863 , \1864 );
xnor \U$1617 ( \1866 , \1865 , \764 );
xor \U$1618 ( \1867 , \1862 , \1866 );
xor \U$1619 ( \1868 , \1853 , \1867 );
not \U$1620 ( \1869 , \576 );
and \U$1621 ( \1870 , \504 , \641 );
and \U$1622 ( \1871 , \223 , \639 );
nor \U$1623 ( \1872 , \1870 , \1871 );
xnor \U$1624 ( \1873 , \1872 , \648 );
xor \U$1625 ( \1874 , \1869 , \1873 );
and \U$1626 ( \1875 , \1020 , \671 );
and \U$1627 ( \1876 , \539 , \669 );
nor \U$1628 ( \1877 , \1875 , \1876 );
xnor \U$1629 ( \1878 , \1877 , \678 );
xor \U$1630 ( \1879 , \1874 , \1878 );
xor \U$1631 ( \1880 , \1868 , \1879 );
and \U$1632 ( \1881 , \952 , \497 );
and \U$1633 ( \1882 , \912 , \495 );
nor \U$1634 ( \1883 , \1881 , \1882 );
xnor \U$1635 ( \1884 , \1883 , \502 );
and \U$1637 ( \1885 , \939 , \505 );
nor \U$1638 ( \1886 , 1'b0 , \1885 );
not \U$1639 ( \1887 , \1886 );
xnor \U$1640 ( \1888 , \1884 , \1887 );
and \U$1641 ( \1889 , \874 , \950 );
and \U$1642 ( \1890 , \827 , \948 );
nor \U$1643 ( \1891 , \1889 , \1890 );
xnor \U$1644 ( \1892 , \1891 , \957 );
and \U$1645 ( \1893 , \902 , \978 );
and \U$1646 ( \1894 , \854 , \961 );
nor \U$1647 ( \1895 , \1893 , \1894 );
xnor \U$1648 ( \1896 , \1895 , \568 );
xor \U$1649 ( \1897 , \1892 , \1896 );
and \U$1650 ( \1898 , \932 , \1198 );
and \U$1651 ( \1899 , \882 , \1079 );
nor \U$1652 ( \1900 , \1898 , \1899 );
xnor \U$1653 ( \1901 , \1900 , \532 );
xor \U$1654 ( \1902 , \1897 , \1901 );
xor \U$1655 ( \1903 , \1888 , \1902 );
and \U$1656 ( \1904 , \786 , \872 );
and \U$1657 ( \1905 , \739 , \870 );
nor \U$1658 ( \1906 , \1904 , \1905 );
xnor \U$1659 ( \1907 , \1906 , \879 );
and \U$1660 ( \1908 , \814 , \900 );
and \U$1661 ( \1909 , \766 , \898 );
nor \U$1662 ( \1910 , \1908 , \1909 );
xnor \U$1663 ( \1911 , \1910 , \907 );
xor \U$1664 ( \1912 , \1907 , \1911 );
and \U$1665 ( \1913 , \847 , \930 );
and \U$1666 ( \1914 , \794 , \928 );
nor \U$1667 ( \1915 , \1913 , \1914 );
xnor \U$1668 ( \1916 , \1915 , \937 );
xor \U$1669 ( \1917 , \1912 , \1916 );
xor \U$1670 ( \1918 , \1903 , \1917 );
xor \U$1671 ( \1919 , \1880 , \1918 );
and \U$1672 ( \1920 , \1752 , \1756 );
and \U$1673 ( \1921 , \1756 , \1761 );
and \U$1674 ( \1922 , \1752 , \1761 );
or \U$1675 ( \1923 , \1920 , \1921 , \1922 );
and \U$1676 ( \1924 , \1738 , \1742 );
and \U$1677 ( \1925 , \1742 , \1747 );
and \U$1678 ( \1926 , \1738 , \1747 );
or \U$1679 ( \1927 , \1924 , \1925 , \1926 );
xor \U$1680 ( \1928 , \1923 , \1927 );
and \U$1681 ( \1929 , \1687 , \1691 );
and \U$1682 ( \1930 , \1691 , \1694 );
and \U$1683 ( \1931 , \1687 , \1694 );
or \U$1684 ( \1932 , \1929 , \1930 , \1931 );
xor \U$1685 ( \1933 , \1928 , \1932 );
xor \U$1686 ( \1934 , \1919 , \1933 );
xor \U$1687 ( \1935 , \1839 , \1934 );
and \U$1688 ( \1936 , \1700 , \1704 );
and \U$1689 ( \1937 , \1704 , \1709 );
and \U$1690 ( \1938 , \1700 , \1709 );
or \U$1691 ( \1939 , \1936 , \1937 , \1938 );
and \U$1692 ( \1940 , \1678 , \1682 );
and \U$1693 ( \1941 , \1682 , \1695 );
and \U$1694 ( \1942 , \1678 , \1695 );
or \U$1695 ( \1943 , \1940 , \1941 , \1942 );
xor \U$1696 ( \1944 , \1939 , \1943 );
and \U$1697 ( \1945 , \1748 , \1762 );
and \U$1698 ( \1946 , \1762 , \1777 );
and \U$1699 ( \1947 , \1748 , \1777 );
or \U$1700 ( \1948 , \1945 , \1946 , \1947 );
xor \U$1701 ( \1949 , \1944 , \1948 );
xor \U$1702 ( \1950 , \1935 , \1949 );
xor \U$1703 ( \1951 , \1828 , \1950 );
xor \U$1704 ( \1952 , \1819 , \1951 );
and \U$1705 ( \1953 , \1653 , \1667 );
and \U$1706 ( \1954 , \1667 , \1796 );
and \U$1707 ( \1955 , \1653 , \1796 );
or \U$1708 ( \1956 , \1953 , \1954 , \1955 );
nor \U$1709 ( \1957 , \1952 , \1956 );
and \U$1710 ( \1958 , \1823 , \1827 );
and \U$1711 ( \1959 , \1827 , \1950 );
and \U$1712 ( \1960 , \1823 , \1950 );
or \U$1713 ( \1961 , \1958 , \1959 , \1960 );
and \U$1714 ( \1962 , \1939 , \1943 );
and \U$1715 ( \1963 , \1943 , \1948 );
and \U$1716 ( \1964 , \1939 , \1948 );
or \U$1717 ( \1965 , \1962 , \1963 , \1964 );
and \U$1718 ( \1966 , \1880 , \1918 );
and \U$1719 ( \1967 , \1918 , \1933 );
and \U$1720 ( \1968 , \1880 , \1933 );
or \U$1721 ( \1969 , \1966 , \1967 , \1968 );
xor \U$1722 ( \1970 , \1965 , \1969 );
and \U$1723 ( \1971 , \1907 , \1911 );
and \U$1724 ( \1972 , \1911 , \1916 );
and \U$1725 ( \1973 , \1907 , \1916 );
or \U$1726 ( \1974 , \1971 , \1972 , \1973 );
and \U$1727 ( \1975 , \1892 , \1896 );
and \U$1728 ( \1976 , \1896 , \1901 );
and \U$1729 ( \1977 , \1892 , \1901 );
or \U$1730 ( \1978 , \1975 , \1976 , \1977 );
xor \U$1731 ( \1979 , \1974 , \1978 );
or \U$1732 ( \1980 , \1884 , \1887 );
xor \U$1733 ( \1981 , \1979 , \1980 );
xor \U$1734 ( \1982 , \1970 , \1981 );
xor \U$1735 ( \1983 , \1961 , \1982 );
and \U$1736 ( \1984 , \1811 , \1815 );
and \U$1737 ( \1985 , \1815 , \1817 );
and \U$1738 ( \1986 , \1811 , \1817 );
or \U$1739 ( \1987 , \1984 , \1985 , \1986 );
and \U$1740 ( \1988 , \1839 , \1934 );
and \U$1741 ( \1989 , \1934 , \1949 );
and \U$1742 ( \1990 , \1839 , \1949 );
or \U$1743 ( \1991 , \1988 , \1989 , \1990 );
xor \U$1744 ( \1992 , \1987 , \1991 );
and \U$1745 ( \1993 , \1869 , \1873 );
and \U$1746 ( \1994 , \1873 , \1878 );
and \U$1747 ( \1995 , \1869 , \1878 );
or \U$1748 ( \1996 , \1993 , \1994 , \1995 );
and \U$1749 ( \1997 , \1857 , \1861 );
and \U$1750 ( \1998 , \1861 , \1866 );
and \U$1751 ( \1999 , \1857 , \1866 );
or \U$1752 ( \2000 , \1997 , \1998 , \1999 );
xor \U$1753 ( \2001 , \1996 , \2000 );
and \U$1754 ( \2002 , \1843 , \1847 );
and \U$1755 ( \2003 , \1847 , \1852 );
and \U$1756 ( \2004 , \1843 , \1852 );
or \U$1757 ( \2005 , \2002 , \2003 , \2004 );
xor \U$1758 ( \2006 , \2001 , \2005 );
and \U$1759 ( \2007 , \1853 , \1867 );
and \U$1760 ( \2008 , \1867 , \1879 );
and \U$1761 ( \2009 , \1853 , \1879 );
or \U$1762 ( \2010 , \2007 , \2008 , \2009 );
and \U$1763 ( \2011 , \680 , \812 );
and \U$1764 ( \2012 , \700 , \810 );
nor \U$1765 ( \2013 , \2011 , \2012 );
xnor \U$1766 ( \2014 , \2013 , \819 );
and \U$1767 ( \2015 , \708 , \845 );
and \U$1768 ( \2016 , \728 , \843 );
nor \U$1769 ( \2017 , \2015 , \2016 );
xnor \U$1770 ( \2018 , \2017 , \852 );
xor \U$1771 ( \2019 , \2014 , \2018 );
and \U$1772 ( \2020 , \739 , \872 );
and \U$1773 ( \2021 , \759 , \870 );
nor \U$1774 ( \2022 , \2020 , \2021 );
xnor \U$1775 ( \2023 , \2022 , \879 );
xor \U$1776 ( \2024 , \2019 , \2023 );
and \U$1777 ( \2025 , \569 , \726 );
and \U$1778 ( \2026 , \618 , \724 );
nor \U$1779 ( \2027 , \2025 , \2026 );
xnor \U$1780 ( \2028 , \2027 , \733 );
and \U$1781 ( \2029 , \623 , \757 );
and \U$1782 ( \2030 , \643 , \755 );
nor \U$1783 ( \2031 , \2029 , \2030 );
xnor \U$1784 ( \2032 , \2031 , \764 );
xor \U$1785 ( \2033 , \2028 , \2032 );
and \U$1786 ( \2034 , \653 , \784 );
and \U$1787 ( \2035 , \673 , \782 );
nor \U$1788 ( \2036 , \2034 , \2035 );
xnor \U$1789 ( \2037 , \2036 , \791 );
xor \U$1790 ( \2038 , \2033 , \2037 );
xor \U$1791 ( \2039 , \2024 , \2038 );
and \U$1792 ( \2040 , \223 , \641 );
not \U$1793 ( \2041 , \2040 );
xnor \U$1794 ( \2042 , \2041 , \648 );
and \U$1795 ( \2043 , \539 , \671 );
and \U$1796 ( \2044 , \504 , \669 );
nor \U$1797 ( \2045 , \2043 , \2044 );
xnor \U$1798 ( \2046 , \2045 , \678 );
xor \U$1799 ( \2047 , \2042 , \2046 );
and \U$1800 ( \2048 , \1018 , \698 );
and \U$1801 ( \2049 , \1020 , \696 );
nor \U$1802 ( \2050 , \2048 , \2049 );
xnor \U$1803 ( \2051 , \2050 , \705 );
xor \U$1804 ( \2052 , \2047 , \2051 );
xor \U$1805 ( \2053 , \2039 , \2052 );
xor \U$1806 ( \2054 , \2010 , \2053 );
and \U$1808 ( \2055 , \952 , \505 );
nor \U$1809 ( \2056 , 1'b0 , \2055 );
and \U$1810 ( \2057 , \854 , \978 );
and \U$1811 ( \2058 , \874 , \961 );
nor \U$1812 ( \2059 , \2057 , \2058 );
xnor \U$1813 ( \2060 , \2059 , \568 );
and \U$1814 ( \2061 , \882 , \1198 );
and \U$1815 ( \2062 , \902 , \1079 );
nor \U$1816 ( \2063 , \2061 , \2062 );
xnor \U$1817 ( \2064 , \2063 , \532 );
xor \U$1818 ( \2065 , \2060 , \2064 );
and \U$1819 ( \2066 , \912 , \497 );
and \U$1820 ( \2067 , \932 , \495 );
nor \U$1821 ( \2068 , \2066 , \2067 );
xnor \U$1822 ( \2069 , \2068 , \502 );
xor \U$1823 ( \2070 , \2065 , \2069 );
xor \U$1824 ( \2071 , \2056 , \2070 );
and \U$1825 ( \2072 , \766 , \900 );
and \U$1826 ( \2073 , \786 , \898 );
nor \U$1827 ( \2074 , \2072 , \2073 );
xnor \U$1828 ( \2075 , \2074 , \907 );
and \U$1829 ( \2076 , \794 , \930 );
and \U$1830 ( \2077 , \814 , \928 );
nor \U$1831 ( \2078 , \2076 , \2077 );
xnor \U$1832 ( \2079 , \2078 , \937 );
xor \U$1833 ( \2080 , \2075 , \2079 );
and \U$1834 ( \2081 , \827 , \950 );
and \U$1835 ( \2082 , \847 , \948 );
nor \U$1836 ( \2083 , \2081 , \2082 );
xnor \U$1837 ( \2084 , \2083 , \957 );
xor \U$1838 ( \2085 , \2080 , \2084 );
xor \U$1839 ( \2086 , \2071 , \2085 );
xor \U$1840 ( \2087 , \2054 , \2086 );
xor \U$1841 ( \2088 , \2006 , \2087 );
and \U$1842 ( \2089 , \1829 , \1833 );
and \U$1843 ( \2090 , \1833 , \1838 );
and \U$1844 ( \2091 , \1829 , \1838 );
or \U$1845 ( \2092 , \2089 , \2090 , \2091 );
and \U$1846 ( \2093 , \1923 , \1927 );
and \U$1847 ( \2094 , \1927 , \1932 );
and \U$1848 ( \2095 , \1923 , \1932 );
or \U$1849 ( \2096 , \2093 , \2094 , \2095 );
xor \U$1850 ( \2097 , \2092 , \2096 );
and \U$1851 ( \2098 , \1888 , \1902 );
and \U$1852 ( \2099 , \1902 , \1917 );
and \U$1853 ( \2100 , \1888 , \1917 );
or \U$1854 ( \2101 , \2098 , \2099 , \2100 );
xor \U$1855 ( \2102 , \2097 , \2101 );
xor \U$1856 ( \2103 , \2088 , \2102 );
xor \U$1857 ( \2104 , \1992 , \2103 );
xor \U$1858 ( \2105 , \1983 , \2104 );
and \U$1859 ( \2106 , \1807 , \1818 );
and \U$1860 ( \2107 , \1818 , \1951 );
and \U$1861 ( \2108 , \1807 , \1951 );
or \U$1862 ( \2109 , \2106 , \2107 , \2108 );
nor \U$1863 ( \2110 , \2105 , \2109 );
nor \U$1864 ( \2111 , \1957 , \2110 );
nand \U$1865 ( \2112 , \1803 , \2111 );
and \U$1866 ( \2113 , \1987 , \1991 );
and \U$1867 ( \2114 , \1991 , \2103 );
and \U$1868 ( \2115 , \1987 , \2103 );
or \U$1869 ( \2116 , \2113 , \2114 , \2115 );
and \U$1870 ( \2117 , \2092 , \2096 );
and \U$1871 ( \2118 , \2096 , \2101 );
and \U$1872 ( \2119 , \2092 , \2101 );
or \U$1873 ( \2120 , \2117 , \2118 , \2119 );
and \U$1874 ( \2121 , \2010 , \2053 );
and \U$1875 ( \2122 , \2053 , \2086 );
and \U$1876 ( \2123 , \2010 , \2086 );
or \U$1877 ( \2124 , \2121 , \2122 , \2123 );
xor \U$1878 ( \2125 , \2120 , \2124 );
and \U$1879 ( \2126 , \2075 , \2079 );
and \U$1880 ( \2127 , \2079 , \2084 );
and \U$1881 ( \2128 , \2075 , \2084 );
or \U$1882 ( \2129 , \2126 , \2127 , \2128 );
and \U$1883 ( \2130 , \2060 , \2064 );
and \U$1884 ( \2131 , \2064 , \2069 );
and \U$1885 ( \2132 , \2060 , \2069 );
or \U$1886 ( \2133 , \2130 , \2131 , \2132 );
xor \U$1887 ( \2134 , \2129 , \2133 );
not \U$1888 ( \2135 , \2056 );
xor \U$1889 ( \2136 , \2134 , \2135 );
xor \U$1890 ( \2137 , \2125 , \2136 );
xor \U$1891 ( \2138 , \2116 , \2137 );
and \U$1892 ( \2139 , \1965 , \1969 );
and \U$1893 ( \2140 , \1969 , \1981 );
and \U$1894 ( \2141 , \1965 , \1981 );
or \U$1895 ( \2142 , \2139 , \2140 , \2141 );
and \U$1896 ( \2143 , \2006 , \2087 );
and \U$1897 ( \2144 , \2087 , \2102 );
and \U$1898 ( \2145 , \2006 , \2102 );
or \U$1899 ( \2146 , \2143 , \2144 , \2145 );
xor \U$1900 ( \2147 , \2142 , \2146 );
and \U$1901 ( \2148 , \2042 , \2046 );
and \U$1902 ( \2149 , \2046 , \2051 );
and \U$1903 ( \2150 , \2042 , \2051 );
or \U$1904 ( \2151 , \2148 , \2149 , \2150 );
and \U$1905 ( \2152 , \2028 , \2032 );
and \U$1906 ( \2153 , \2032 , \2037 );
and \U$1907 ( \2154 , \2028 , \2037 );
or \U$1908 ( \2155 , \2152 , \2153 , \2154 );
xor \U$1909 ( \2156 , \2151 , \2155 );
and \U$1910 ( \2157 , \2014 , \2018 );
and \U$1911 ( \2158 , \2018 , \2023 );
and \U$1912 ( \2159 , \2014 , \2023 );
or \U$1913 ( \2160 , \2157 , \2158 , \2159 );
xor \U$1914 ( \2161 , \2156 , \2160 );
and \U$1915 ( \2162 , \2024 , \2038 );
and \U$1916 ( \2163 , \2038 , \2052 );
and \U$1917 ( \2164 , \2024 , \2052 );
or \U$1918 ( \2165 , \2162 , \2163 , \2164 );
and \U$1919 ( \2166 , \700 , \812 );
and \U$1920 ( \2167 , \653 , \810 );
nor \U$1921 ( \2168 , \2166 , \2167 );
xnor \U$1922 ( \2169 , \2168 , \819 );
and \U$1923 ( \2170 , \728 , \845 );
and \U$1924 ( \2171 , \680 , \843 );
nor \U$1925 ( \2172 , \2170 , \2171 );
xnor \U$1926 ( \2173 , \2172 , \852 );
xor \U$1927 ( \2174 , \2169 , \2173 );
and \U$1928 ( \2175 , \759 , \872 );
and \U$1929 ( \2176 , \708 , \870 );
nor \U$1930 ( \2177 , \2175 , \2176 );
xnor \U$1931 ( \2178 , \2177 , \879 );
xor \U$1932 ( \2179 , \2174 , \2178 );
and \U$1933 ( \2180 , \618 , \726 );
and \U$1934 ( \2181 , \1018 , \724 );
nor \U$1935 ( \2182 , \2180 , \2181 );
xnor \U$1936 ( \2183 , \2182 , \733 );
and \U$1937 ( \2184 , \643 , \757 );
and \U$1938 ( \2185 , \569 , \755 );
nor \U$1939 ( \2186 , \2184 , \2185 );
xnor \U$1940 ( \2187 , \2186 , \764 );
xor \U$1941 ( \2188 , \2183 , \2187 );
and \U$1942 ( \2189 , \673 , \784 );
and \U$1943 ( \2190 , \623 , \782 );
nor \U$1944 ( \2191 , \2189 , \2190 );
xnor \U$1945 ( \2192 , \2191 , \791 );
xor \U$1946 ( \2193 , \2188 , \2192 );
xor \U$1947 ( \2194 , \2179 , \2193 );
not \U$1948 ( \2195 , \648 );
and \U$1949 ( \2196 , \504 , \671 );
and \U$1950 ( \2197 , \223 , \669 );
nor \U$1951 ( \2198 , \2196 , \2197 );
xnor \U$1952 ( \2199 , \2198 , \678 );
xor \U$1953 ( \2200 , \2195 , \2199 );
and \U$1954 ( \2201 , \1020 , \698 );
and \U$1955 ( \2202 , \539 , \696 );
nor \U$1956 ( \2203 , \2201 , \2202 );
xnor \U$1957 ( \2204 , \2203 , \705 );
xor \U$1958 ( \2205 , \2200 , \2204 );
xor \U$1959 ( \2206 , \2194 , \2205 );
xor \U$1960 ( \2207 , \2165 , \2206 );
and \U$1962 ( \2208 , \912 , \505 );
nor \U$1963 ( \2209 , 1'b0 , \2208 );
not \U$1964 ( \2210 , \2209 );
and \U$1965 ( \2211 , \874 , \978 );
and \U$1966 ( \2212 , \827 , \961 );
nor \U$1967 ( \2213 , \2211 , \2212 );
xnor \U$1968 ( \2214 , \2213 , \568 );
and \U$1969 ( \2215 , \902 , \1198 );
and \U$1970 ( \2216 , \854 , \1079 );
nor \U$1971 ( \2217 , \2215 , \2216 );
xnor \U$1972 ( \2218 , \2217 , \532 );
xor \U$1973 ( \2219 , \2214 , \2218 );
and \U$1974 ( \2220 , \932 , \497 );
and \U$1975 ( \2221 , \882 , \495 );
nor \U$1976 ( \2222 , \2220 , \2221 );
xnor \U$1977 ( \2223 , \2222 , \502 );
xor \U$1978 ( \2224 , \2219 , \2223 );
xor \U$1979 ( \2225 , \2210 , \2224 );
and \U$1980 ( \2226 , \786 , \900 );
and \U$1981 ( \2227 , \739 , \898 );
nor \U$1982 ( \2228 , \2226 , \2227 );
xnor \U$1983 ( \2229 , \2228 , \907 );
and \U$1984 ( \2230 , \814 , \930 );
and \U$1985 ( \2231 , \766 , \928 );
nor \U$1986 ( \2232 , \2230 , \2231 );
xnor \U$1987 ( \2233 , \2232 , \937 );
xor \U$1988 ( \2234 , \2229 , \2233 );
and \U$1989 ( \2235 , \847 , \950 );
and \U$1990 ( \2236 , \794 , \948 );
nor \U$1991 ( \2237 , \2235 , \2236 );
xnor \U$1992 ( \2238 , \2237 , \957 );
xor \U$1993 ( \2239 , \2234 , \2238 );
xor \U$1994 ( \2240 , \2225 , \2239 );
xor \U$1995 ( \2241 , \2207 , \2240 );
xor \U$1996 ( \2242 , \2161 , \2241 );
and \U$1997 ( \2243 , \1996 , \2000 );
and \U$1998 ( \2244 , \2000 , \2005 );
and \U$1999 ( \2245 , \1996 , \2005 );
or \U$2000 ( \2246 , \2243 , \2244 , \2245 );
and \U$2001 ( \2247 , \1974 , \1978 );
and \U$2002 ( \2248 , \1978 , \1980 );
and \U$2003 ( \2249 , \1974 , \1980 );
or \U$2004 ( \2250 , \2247 , \2248 , \2249 );
xor \U$2005 ( \2251 , \2246 , \2250 );
and \U$2006 ( \2252 , \2056 , \2070 );
and \U$2007 ( \2253 , \2070 , \2085 );
and \U$2008 ( \2254 , \2056 , \2085 );
or \U$2009 ( \2255 , \2252 , \2253 , \2254 );
xor \U$2010 ( \2256 , \2251 , \2255 );
xor \U$2011 ( \2257 , \2242 , \2256 );
xor \U$2012 ( \2258 , \2147 , \2257 );
xor \U$2013 ( \2259 , \2138 , \2258 );
and \U$2014 ( \2260 , \1961 , \1982 );
and \U$2015 ( \2261 , \1982 , \2104 );
and \U$2016 ( \2262 , \1961 , \2104 );
or \U$2017 ( \2263 , \2260 , \2261 , \2262 );
nor \U$2018 ( \2264 , \2259 , \2263 );
and \U$2019 ( \2265 , \2142 , \2146 );
and \U$2020 ( \2266 , \2146 , \2257 );
and \U$2021 ( \2267 , \2142 , \2257 );
or \U$2022 ( \2268 , \2265 , \2266 , \2267 );
and \U$2023 ( \2269 , \2151 , \2155 );
and \U$2024 ( \2270 , \2155 , \2160 );
and \U$2025 ( \2271 , \2151 , \2160 );
or \U$2026 ( \2272 , \2269 , \2270 , \2271 );
and \U$2027 ( \2273 , \2129 , \2133 );
and \U$2028 ( \2274 , \2133 , \2135 );
and \U$2029 ( \2275 , \2129 , \2135 );
or \U$2030 ( \2276 , \2273 , \2274 , \2275 );
xor \U$2031 ( \2277 , \2272 , \2276 );
and \U$2032 ( \2278 , \2210 , \2224 );
and \U$2033 ( \2279 , \2224 , \2239 );
and \U$2034 ( \2280 , \2210 , \2239 );
or \U$2035 ( \2281 , \2278 , \2279 , \2280 );
xor \U$2036 ( \2282 , \2277 , \2281 );
and \U$2037 ( \2283 , \2246 , \2250 );
and \U$2038 ( \2284 , \2250 , \2255 );
and \U$2039 ( \2285 , \2246 , \2255 );
or \U$2040 ( \2286 , \2283 , \2284 , \2285 );
and \U$2041 ( \2287 , \2165 , \2206 );
and \U$2042 ( \2288 , \2206 , \2240 );
and \U$2043 ( \2289 , \2165 , \2240 );
or \U$2044 ( \2290 , \2287 , \2288 , \2289 );
xor \U$2045 ( \2291 , \2286 , \2290 );
and \U$2046 ( \2292 , \854 , \1198 );
and \U$2047 ( \2293 , \874 , \1079 );
nor \U$2048 ( \2294 , \2292 , \2293 );
xnor \U$2049 ( \2295 , \2294 , \532 );
and \U$2050 ( \2296 , \882 , \497 );
and \U$2051 ( \2297 , \902 , \495 );
nor \U$2052 ( \2298 , \2296 , \2297 );
xnor \U$2053 ( \2299 , \2298 , \502 );
xor \U$2054 ( \2300 , \2295 , \2299 );
and \U$2056 ( \2301 , \932 , \505 );
nor \U$2057 ( \2302 , 1'b0 , \2301 );
not \U$2058 ( \2303 , \2302 );
xor \U$2059 ( \2304 , \2300 , \2303 );
and \U$2060 ( \2305 , \766 , \930 );
and \U$2061 ( \2306 , \786 , \928 );
nor \U$2062 ( \2307 , \2305 , \2306 );
xnor \U$2063 ( \2308 , \2307 , \937 );
and \U$2064 ( \2309 , \794 , \950 );
and \U$2065 ( \2310 , \814 , \948 );
nor \U$2066 ( \2311 , \2309 , \2310 );
xnor \U$2067 ( \2312 , \2311 , \957 );
xor \U$2068 ( \2313 , \2308 , \2312 );
and \U$2069 ( \2314 , \827 , \978 );
and \U$2070 ( \2315 , \847 , \961 );
nor \U$2071 ( \2316 , \2314 , \2315 );
xnor \U$2072 ( \2317 , \2316 , \568 );
xor \U$2073 ( \2318 , \2313 , \2317 );
xor \U$2074 ( \2319 , \2304 , \2318 );
and \U$2075 ( \2320 , \680 , \845 );
and \U$2076 ( \2321 , \700 , \843 );
nor \U$2077 ( \2322 , \2320 , \2321 );
xnor \U$2078 ( \2323 , \2322 , \852 );
and \U$2079 ( \2324 , \708 , \872 );
and \U$2080 ( \2325 , \728 , \870 );
nor \U$2081 ( \2326 , \2324 , \2325 );
xnor \U$2082 ( \2327 , \2326 , \879 );
xor \U$2083 ( \2328 , \2323 , \2327 );
and \U$2084 ( \2329 , \739 , \900 );
and \U$2085 ( \2330 , \759 , \898 );
nor \U$2086 ( \2331 , \2329 , \2330 );
xnor \U$2087 ( \2332 , \2331 , \907 );
xor \U$2088 ( \2333 , \2328 , \2332 );
xor \U$2089 ( \2334 , \2319 , \2333 );
and \U$2090 ( \2335 , \2229 , \2233 );
and \U$2091 ( \2336 , \2233 , \2238 );
and \U$2092 ( \2337 , \2229 , \2238 );
or \U$2093 ( \2338 , \2335 , \2336 , \2337 );
and \U$2094 ( \2339 , \2214 , \2218 );
and \U$2095 ( \2340 , \2218 , \2223 );
and \U$2096 ( \2341 , \2214 , \2223 );
or \U$2097 ( \2342 , \2339 , \2340 , \2341 );
xnor \U$2098 ( \2343 , \2338 , \2342 );
xor \U$2099 ( \2344 , \2334 , \2343 );
and \U$2100 ( \2345 , \2195 , \2199 );
and \U$2101 ( \2346 , \2199 , \2204 );
and \U$2102 ( \2347 , \2195 , \2204 );
or \U$2103 ( \2348 , \2345 , \2346 , \2347 );
and \U$2104 ( \2349 , \2183 , \2187 );
and \U$2105 ( \2350 , \2187 , \2192 );
and \U$2106 ( \2351 , \2183 , \2192 );
or \U$2107 ( \2352 , \2349 , \2350 , \2351 );
xor \U$2108 ( \2353 , \2348 , \2352 );
and \U$2109 ( \2354 , \2169 , \2173 );
and \U$2110 ( \2355 , \2173 , \2178 );
and \U$2111 ( \2356 , \2169 , \2178 );
or \U$2112 ( \2357 , \2354 , \2355 , \2356 );
xor \U$2113 ( \2358 , \2353 , \2357 );
xor \U$2114 ( \2359 , \2344 , \2358 );
xor \U$2115 ( \2360 , \2291 , \2359 );
xor \U$2116 ( \2361 , \2282 , \2360 );
xor \U$2117 ( \2362 , \2268 , \2361 );
and \U$2118 ( \2363 , \2120 , \2124 );
and \U$2119 ( \2364 , \2124 , \2136 );
and \U$2120 ( \2365 , \2120 , \2136 );
or \U$2121 ( \2366 , \2363 , \2364 , \2365 );
and \U$2122 ( \2367 , \2161 , \2241 );
and \U$2123 ( \2368 , \2241 , \2256 );
and \U$2124 ( \2369 , \2161 , \2256 );
or \U$2125 ( \2370 , \2367 , \2368 , \2369 );
xor \U$2126 ( \2371 , \2366 , \2370 );
and \U$2127 ( \2372 , \2179 , \2193 );
and \U$2128 ( \2373 , \2193 , \2205 );
and \U$2129 ( \2374 , \2179 , \2205 );
or \U$2130 ( \2375 , \2372 , \2373 , \2374 );
and \U$2131 ( \2376 , \569 , \757 );
and \U$2132 ( \2377 , \618 , \755 );
nor \U$2133 ( \2378 , \2376 , \2377 );
xnor \U$2134 ( \2379 , \2378 , \764 );
and \U$2135 ( \2380 , \623 , \784 );
and \U$2136 ( \2381 , \643 , \782 );
nor \U$2137 ( \2382 , \2380 , \2381 );
xnor \U$2138 ( \2383 , \2382 , \791 );
xor \U$2139 ( \2384 , \2379 , \2383 );
and \U$2140 ( \2385 , \653 , \812 );
and \U$2141 ( \2386 , \673 , \810 );
nor \U$2142 ( \2387 , \2385 , \2386 );
xnor \U$2143 ( \2388 , \2387 , \819 );
xor \U$2144 ( \2389 , \2384 , \2388 );
xor \U$2145 ( \2390 , \2375 , \2389 );
and \U$2146 ( \2391 , \223 , \671 );
not \U$2147 ( \2392 , \2391 );
xnor \U$2148 ( \2393 , \2392 , \678 );
and \U$2149 ( \2394 , \539 , \698 );
and \U$2150 ( \2395 , \504 , \696 );
nor \U$2151 ( \2396 , \2394 , \2395 );
xnor \U$2152 ( \2397 , \2396 , \705 );
xor \U$2153 ( \2398 , \2393 , \2397 );
and \U$2154 ( \2399 , \1018 , \726 );
and \U$2155 ( \2400 , \1020 , \724 );
nor \U$2156 ( \2401 , \2399 , \2400 );
xnor \U$2157 ( \2402 , \2401 , \733 );
xor \U$2158 ( \2403 , \2398 , \2402 );
xor \U$2159 ( \2404 , \2390 , \2403 );
xor \U$2160 ( \2405 , \2371 , \2404 );
xor \U$2161 ( \2406 , \2362 , \2405 );
and \U$2162 ( \2407 , \2116 , \2137 );
and \U$2163 ( \2408 , \2137 , \2258 );
and \U$2164 ( \2409 , \2116 , \2258 );
or \U$2165 ( \2410 , \2407 , \2408 , \2409 );
nor \U$2166 ( \2411 , \2406 , \2410 );
nor \U$2167 ( \2412 , \2264 , \2411 );
and \U$2168 ( \2413 , \2366 , \2370 );
and \U$2169 ( \2414 , \2370 , \2404 );
and \U$2170 ( \2415 , \2366 , \2404 );
or \U$2171 ( \2416 , \2413 , \2414 , \2415 );
and \U$2172 ( \2417 , \2282 , \2360 );
xor \U$2173 ( \2418 , \2416 , \2417 );
and \U$2174 ( \2419 , \2286 , \2290 );
and \U$2175 ( \2420 , \2290 , \2359 );
and \U$2176 ( \2421 , \2286 , \2359 );
or \U$2177 ( \2422 , \2419 , \2420 , \2421 );
and \U$2178 ( \2423 , \2393 , \2397 );
and \U$2179 ( \2424 , \2397 , \2402 );
and \U$2180 ( \2425 , \2393 , \2402 );
or \U$2181 ( \2426 , \2423 , \2424 , \2425 );
and \U$2182 ( \2427 , \2379 , \2383 );
and \U$2183 ( \2428 , \2383 , \2388 );
and \U$2184 ( \2429 , \2379 , \2388 );
or \U$2185 ( \2430 , \2427 , \2428 , \2429 );
xor \U$2186 ( \2431 , \2426 , \2430 );
and \U$2187 ( \2432 , \2323 , \2327 );
and \U$2188 ( \2433 , \2327 , \2332 );
and \U$2189 ( \2434 , \2323 , \2332 );
or \U$2190 ( \2435 , \2432 , \2433 , \2434 );
xor \U$2191 ( \2436 , \2431 , \2435 );
not \U$2192 ( \2437 , \678 );
and \U$2193 ( \2438 , \504 , \698 );
and \U$2194 ( \2439 , \223 , \696 );
nor \U$2195 ( \2440 , \2438 , \2439 );
xnor \U$2196 ( \2441 , \2440 , \705 );
xor \U$2197 ( \2442 , \2437 , \2441 );
and \U$2198 ( \2443 , \1020 , \726 );
and \U$2199 ( \2444 , \539 , \724 );
nor \U$2200 ( \2445 , \2443 , \2444 );
xnor \U$2201 ( \2446 , \2445 , \733 );
xor \U$2202 ( \2447 , \2442 , \2446 );
and \U$2203 ( \2448 , \786 , \930 );
and \U$2204 ( \2449 , \739 , \928 );
nor \U$2205 ( \2450 , \2448 , \2449 );
xnor \U$2206 ( \2451 , \2450 , \937 );
and \U$2207 ( \2452 , \814 , \950 );
and \U$2208 ( \2453 , \766 , \948 );
nor \U$2209 ( \2454 , \2452 , \2453 );
xnor \U$2210 ( \2455 , \2454 , \957 );
xor \U$2211 ( \2456 , \2451 , \2455 );
and \U$2212 ( \2457 , \847 , \978 );
and \U$2213 ( \2458 , \794 , \961 );
nor \U$2214 ( \2459 , \2457 , \2458 );
xnor \U$2215 ( \2460 , \2459 , \568 );
xor \U$2216 ( \2461 , \2456 , \2460 );
and \U$2217 ( \2462 , \700 , \845 );
and \U$2218 ( \2463 , \653 , \843 );
nor \U$2219 ( \2464 , \2462 , \2463 );
xnor \U$2220 ( \2465 , \2464 , \852 );
and \U$2221 ( \2466 , \728 , \872 );
and \U$2222 ( \2467 , \680 , \870 );
nor \U$2223 ( \2468 , \2466 , \2467 );
xnor \U$2224 ( \2469 , \2468 , \879 );
xor \U$2225 ( \2470 , \2465 , \2469 );
and \U$2226 ( \2471 , \759 , \900 );
and \U$2227 ( \2472 , \708 , \898 );
nor \U$2228 ( \2473 , \2471 , \2472 );
xnor \U$2229 ( \2474 , \2473 , \907 );
xor \U$2230 ( \2475 , \2470 , \2474 );
xor \U$2231 ( \2476 , \2461 , \2475 );
and \U$2232 ( \2477 , \618 , \757 );
and \U$2233 ( \2478 , \1018 , \755 );
nor \U$2234 ( \2479 , \2477 , \2478 );
xnor \U$2235 ( \2480 , \2479 , \764 );
and \U$2236 ( \2481 , \643 , \784 );
and \U$2237 ( \2482 , \569 , \782 );
nor \U$2238 ( \2483 , \2481 , \2482 );
xnor \U$2239 ( \2484 , \2483 , \791 );
xor \U$2240 ( \2485 , \2480 , \2484 );
and \U$2241 ( \2486 , \673 , \812 );
and \U$2242 ( \2487 , \623 , \810 );
nor \U$2243 ( \2488 , \2486 , \2487 );
xnor \U$2244 ( \2489 , \2488 , \819 );
xor \U$2245 ( \2490 , \2485 , \2489 );
xor \U$2246 ( \2491 , \2476 , \2490 );
xor \U$2247 ( \2492 , \2447 , \2491 );
and \U$2248 ( \2493 , \2308 , \2312 );
and \U$2249 ( \2494 , \2312 , \2317 );
and \U$2250 ( \2495 , \2308 , \2317 );
or \U$2251 ( \2496 , \2493 , \2494 , \2495 );
and \U$2252 ( \2497 , \2295 , \2299 );
and \U$2253 ( \2498 , \2299 , \2303 );
and \U$2254 ( \2499 , \2295 , \2303 );
or \U$2255 ( \2500 , \2497 , \2498 , \2499 );
xor \U$2256 ( \2501 , \2496 , \2500 );
and \U$2257 ( \2502 , \874 , \1198 );
and \U$2258 ( \2503 , \827 , \1079 );
nor \U$2259 ( \2504 , \2502 , \2503 );
xnor \U$2260 ( \2505 , \2504 , \532 );
and \U$2261 ( \2506 , \902 , \497 );
and \U$2262 ( \2507 , \854 , \495 );
nor \U$2263 ( \2508 , \2506 , \2507 );
xnor \U$2264 ( \2509 , \2508 , \502 );
xor \U$2265 ( \2510 , \2505 , \2509 );
and \U$2267 ( \2511 , \882 , \505 );
nor \U$2268 ( \2512 , 1'b0 , \2511 );
not \U$2269 ( \2513 , \2512 );
xor \U$2270 ( \2514 , \2510 , \2513 );
xor \U$2271 ( \2515 , \2501 , \2514 );
xor \U$2272 ( \2516 , \2492 , \2515 );
xor \U$2273 ( \2517 , \2436 , \2516 );
and \U$2274 ( \2518 , \2348 , \2352 );
and \U$2275 ( \2519 , \2352 , \2357 );
and \U$2276 ( \2520 , \2348 , \2357 );
or \U$2277 ( \2521 , \2518 , \2519 , \2520 );
or \U$2278 ( \2522 , \2338 , \2342 );
xor \U$2279 ( \2523 , \2521 , \2522 );
and \U$2280 ( \2524 , \2304 , \2318 );
and \U$2281 ( \2525 , \2318 , \2333 );
and \U$2282 ( \2526 , \2304 , \2333 );
or \U$2283 ( \2527 , \2524 , \2525 , \2526 );
xor \U$2284 ( \2528 , \2523 , \2527 );
xor \U$2285 ( \2529 , \2517 , \2528 );
xor \U$2286 ( \2530 , \2422 , \2529 );
and \U$2287 ( \2531 , \2272 , \2276 );
and \U$2288 ( \2532 , \2276 , \2281 );
and \U$2289 ( \2533 , \2272 , \2281 );
or \U$2290 ( \2534 , \2531 , \2532 , \2533 );
and \U$2291 ( \2535 , \2375 , \2389 );
and \U$2292 ( \2536 , \2389 , \2403 );
and \U$2293 ( \2537 , \2375 , \2403 );
or \U$2294 ( \2538 , \2535 , \2536 , \2537 );
xor \U$2295 ( \2539 , \2534 , \2538 );
and \U$2296 ( \2540 , \2334 , \2343 );
and \U$2297 ( \2541 , \2343 , \2358 );
and \U$2298 ( \2542 , \2334 , \2358 );
or \U$2299 ( \2543 , \2540 , \2541 , \2542 );
xor \U$2300 ( \2544 , \2539 , \2543 );
xor \U$2301 ( \2545 , \2530 , \2544 );
xor \U$2302 ( \2546 , \2418 , \2545 );
and \U$2303 ( \2547 , \2268 , \2361 );
and \U$2304 ( \2548 , \2361 , \2405 );
and \U$2305 ( \2549 , \2268 , \2405 );
or \U$2306 ( \2550 , \2547 , \2548 , \2549 );
nor \U$2307 ( \2551 , \2546 , \2550 );
and \U$2308 ( \2552 , \2422 , \2529 );
and \U$2309 ( \2553 , \2529 , \2544 );
and \U$2310 ( \2554 , \2422 , \2544 );
or \U$2311 ( \2555 , \2552 , \2553 , \2554 );
and \U$2312 ( \2556 , \2426 , \2430 );
and \U$2313 ( \2557 , \2430 , \2435 );
and \U$2314 ( \2558 , \2426 , \2435 );
or \U$2315 ( \2559 , \2556 , \2557 , \2558 );
and \U$2316 ( \2560 , \2496 , \2500 );
and \U$2317 ( \2561 , \2500 , \2514 );
and \U$2318 ( \2562 , \2496 , \2514 );
or \U$2319 ( \2563 , \2560 , \2561 , \2562 );
xor \U$2320 ( \2564 , \2559 , \2563 );
and \U$2321 ( \2565 , \2461 , \2475 );
and \U$2322 ( \2566 , \2475 , \2490 );
and \U$2323 ( \2567 , \2461 , \2490 );
or \U$2324 ( \2568 , \2565 , \2566 , \2567 );
xor \U$2325 ( \2569 , \2564 , \2568 );
and \U$2326 ( \2570 , \2521 , \2522 );
and \U$2327 ( \2571 , \2522 , \2527 );
and \U$2328 ( \2572 , \2521 , \2527 );
or \U$2329 ( \2573 , \2570 , \2571 , \2572 );
and \U$2330 ( \2574 , \2447 , \2491 );
and \U$2331 ( \2575 , \2491 , \2515 );
and \U$2332 ( \2576 , \2447 , \2515 );
or \U$2333 ( \2577 , \2574 , \2575 , \2576 );
xor \U$2334 ( \2578 , \2573 , \2577 );
and \U$2335 ( \2579 , \2437 , \2441 );
and \U$2336 ( \2580 , \2441 , \2446 );
and \U$2337 ( \2581 , \2437 , \2446 );
or \U$2338 ( \2582 , \2579 , \2580 , \2581 );
and \U$2339 ( \2583 , \2480 , \2484 );
and \U$2340 ( \2584 , \2484 , \2489 );
and \U$2341 ( \2585 , \2480 , \2489 );
or \U$2342 ( \2586 , \2583 , \2584 , \2585 );
xor \U$2343 ( \2587 , \2582 , \2586 );
and \U$2344 ( \2588 , \2465 , \2469 );
and \U$2345 ( \2589 , \2469 , \2474 );
and \U$2346 ( \2590 , \2465 , \2474 );
or \U$2347 ( \2591 , \2588 , \2589 , \2590 );
xor \U$2348 ( \2592 , \2587 , \2591 );
xor \U$2349 ( \2593 , \2578 , \2592 );
xor \U$2350 ( \2594 , \2569 , \2593 );
xor \U$2351 ( \2595 , \2555 , \2594 );
and \U$2352 ( \2596 , \2534 , \2538 );
and \U$2353 ( \2597 , \2538 , \2543 );
and \U$2354 ( \2598 , \2534 , \2543 );
or \U$2355 ( \2599 , \2596 , \2597 , \2598 );
and \U$2356 ( \2600 , \2436 , \2516 );
and \U$2357 ( \2601 , \2516 , \2528 );
and \U$2358 ( \2602 , \2436 , \2528 );
or \U$2359 ( \2603 , \2600 , \2601 , \2602 );
xor \U$2360 ( \2604 , \2599 , \2603 );
and \U$2361 ( \2605 , \223 , \698 );
not \U$2362 ( \2606 , \2605 );
xnor \U$2363 ( \2607 , \2606 , \705 );
and \U$2364 ( \2608 , \539 , \726 );
and \U$2365 ( \2609 , \504 , \724 );
nor \U$2366 ( \2610 , \2608 , \2609 );
xnor \U$2367 ( \2611 , \2610 , \733 );
xor \U$2368 ( \2612 , \2607 , \2611 );
and \U$2369 ( \2613 , \1018 , \757 );
and \U$2370 ( \2614 , \1020 , \755 );
nor \U$2371 ( \2615 , \2613 , \2614 );
xnor \U$2372 ( \2616 , \2615 , \764 );
xor \U$2373 ( \2617 , \2612 , \2616 );
and \U$2374 ( \2618 , \766 , \950 );
and \U$2375 ( \2619 , \786 , \948 );
nor \U$2376 ( \2620 , \2618 , \2619 );
xnor \U$2377 ( \2621 , \2620 , \957 );
and \U$2378 ( \2622 , \794 , \978 );
and \U$2379 ( \2623 , \814 , \961 );
nor \U$2380 ( \2624 , \2622 , \2623 );
xnor \U$2381 ( \2625 , \2624 , \568 );
xor \U$2382 ( \2626 , \2621 , \2625 );
and \U$2383 ( \2627 , \827 , \1198 );
and \U$2384 ( \2628 , \847 , \1079 );
nor \U$2385 ( \2629 , \2627 , \2628 );
xnor \U$2386 ( \2630 , \2629 , \532 );
xor \U$2387 ( \2631 , \2626 , \2630 );
and \U$2388 ( \2632 , \680 , \872 );
and \U$2389 ( \2633 , \700 , \870 );
nor \U$2390 ( \2634 , \2632 , \2633 );
xnor \U$2391 ( \2635 , \2634 , \879 );
and \U$2392 ( \2636 , \708 , \900 );
and \U$2393 ( \2637 , \728 , \898 );
nor \U$2394 ( \2638 , \2636 , \2637 );
xnor \U$2395 ( \2639 , \2638 , \907 );
xor \U$2396 ( \2640 , \2635 , \2639 );
and \U$2397 ( \2641 , \739 , \930 );
and \U$2398 ( \2642 , \759 , \928 );
nor \U$2399 ( \2643 , \2641 , \2642 );
xnor \U$2400 ( \2644 , \2643 , \937 );
xor \U$2401 ( \2645 , \2640 , \2644 );
xor \U$2402 ( \2646 , \2631 , \2645 );
and \U$2403 ( \2647 , \569 , \784 );
and \U$2404 ( \2648 , \618 , \782 );
nor \U$2405 ( \2649 , \2647 , \2648 );
xnor \U$2406 ( \2650 , \2649 , \791 );
and \U$2407 ( \2651 , \623 , \812 );
and \U$2408 ( \2652 , \643 , \810 );
nor \U$2409 ( \2653 , \2651 , \2652 );
xnor \U$2410 ( \2654 , \2653 , \819 );
xor \U$2411 ( \2655 , \2650 , \2654 );
and \U$2412 ( \2656 , \653 , \845 );
and \U$2413 ( \2657 , \673 , \843 );
nor \U$2414 ( \2658 , \2656 , \2657 );
xnor \U$2415 ( \2659 , \2658 , \852 );
xor \U$2416 ( \2660 , \2655 , \2659 );
xor \U$2417 ( \2661 , \2646 , \2660 );
xor \U$2418 ( \2662 , \2617 , \2661 );
and \U$2419 ( \2663 , \2451 , \2455 );
and \U$2420 ( \2664 , \2455 , \2460 );
and \U$2421 ( \2665 , \2451 , \2460 );
or \U$2422 ( \2666 , \2663 , \2664 , \2665 );
and \U$2423 ( \2667 , \2505 , \2509 );
and \U$2424 ( \2668 , \2509 , \2513 );
and \U$2425 ( \2669 , \2505 , \2513 );
or \U$2426 ( \2670 , \2667 , \2668 , \2669 );
xor \U$2427 ( \2671 , \2666 , \2670 );
and \U$2428 ( \2672 , \854 , \497 );
and \U$2429 ( \2673 , \874 , \495 );
nor \U$2430 ( \2674 , \2672 , \2673 );
xnor \U$2431 ( \2675 , \2674 , \502 );
and \U$2433 ( \2676 , \902 , \505 );
nor \U$2434 ( \2677 , 1'b0 , \2676 );
not \U$2435 ( \2678 , \2677 );
xnor \U$2436 ( \2679 , \2675 , \2678 );
xor \U$2437 ( \2680 , \2671 , \2679 );
xor \U$2438 ( \2681 , \2662 , \2680 );
xor \U$2439 ( \2682 , \2604 , \2681 );
xor \U$2440 ( \2683 , \2595 , \2682 );
and \U$2441 ( \2684 , \2416 , \2417 );
and \U$2442 ( \2685 , \2417 , \2545 );
and \U$2443 ( \2686 , \2416 , \2545 );
or \U$2444 ( \2687 , \2684 , \2685 , \2686 );
nor \U$2445 ( \2688 , \2683 , \2687 );
nor \U$2446 ( \2689 , \2551 , \2688 );
nand \U$2447 ( \2690 , \2412 , \2689 );
nor \U$2448 ( \2691 , \2112 , \2690 );
and \U$2449 ( \2692 , \2599 , \2603 );
and \U$2450 ( \2693 , \2603 , \2681 );
and \U$2451 ( \2694 , \2599 , \2681 );
or \U$2452 ( \2695 , \2692 , \2693 , \2694 );
and \U$2453 ( \2696 , \2569 , \2593 );
xor \U$2454 ( \2697 , \2695 , \2696 );
and \U$2455 ( \2698 , \2573 , \2577 );
and \U$2456 ( \2699 , \2577 , \2592 );
and \U$2457 ( \2700 , \2573 , \2592 );
or \U$2458 ( \2701 , \2698 , \2699 , \2700 );
and \U$2459 ( \2702 , \2607 , \2611 );
and \U$2460 ( \2703 , \2611 , \2616 );
and \U$2461 ( \2704 , \2607 , \2616 );
or \U$2462 ( \2705 , \2702 , \2703 , \2704 );
and \U$2463 ( \2706 , \2650 , \2654 );
and \U$2464 ( \2707 , \2654 , \2659 );
and \U$2465 ( \2708 , \2650 , \2659 );
or \U$2466 ( \2709 , \2706 , \2707 , \2708 );
xor \U$2467 ( \2710 , \2705 , \2709 );
and \U$2468 ( \2711 , \2635 , \2639 );
and \U$2469 ( \2712 , \2639 , \2644 );
and \U$2470 ( \2713 , \2635 , \2644 );
or \U$2471 ( \2714 , \2711 , \2712 , \2713 );
xor \U$2472 ( \2715 , \2710 , \2714 );
and \U$2473 ( \2716 , \618 , \784 );
and \U$2474 ( \2717 , \1018 , \782 );
nor \U$2475 ( \2718 , \2716 , \2717 );
xnor \U$2476 ( \2719 , \2718 , \791 );
and \U$2477 ( \2720 , \643 , \812 );
and \U$2478 ( \2721 , \569 , \810 );
nor \U$2479 ( \2722 , \2720 , \2721 );
xnor \U$2480 ( \2723 , \2722 , \819 );
xor \U$2481 ( \2724 , \2719 , \2723 );
and \U$2482 ( \2725 , \673 , \845 );
and \U$2483 ( \2726 , \623 , \843 );
nor \U$2484 ( \2727 , \2725 , \2726 );
xnor \U$2485 ( \2728 , \2727 , \852 );
xor \U$2486 ( \2729 , \2724 , \2728 );
not \U$2487 ( \2730 , \705 );
and \U$2488 ( \2731 , \504 , \726 );
and \U$2489 ( \2732 , \223 , \724 );
nor \U$2490 ( \2733 , \2731 , \2732 );
xnor \U$2491 ( \2734 , \2733 , \733 );
xor \U$2492 ( \2735 , \2730 , \2734 );
and \U$2493 ( \2736 , \1020 , \757 );
and \U$2494 ( \2737 , \539 , \755 );
nor \U$2495 ( \2738 , \2736 , \2737 );
xnor \U$2496 ( \2739 , \2738 , \764 );
xor \U$2497 ( \2740 , \2735 , \2739 );
xor \U$2498 ( \2741 , \2729 , \2740 );
and \U$2500 ( \2742 , \854 , \505 );
nor \U$2501 ( \2743 , 1'b0 , \2742 );
not \U$2502 ( \2744 , \2743 );
and \U$2503 ( \2745 , \786 , \950 );
and \U$2504 ( \2746 , \739 , \948 );
nor \U$2505 ( \2747 , \2745 , \2746 );
xnor \U$2506 ( \2748 , \2747 , \957 );
and \U$2507 ( \2749 , \814 , \978 );
and \U$2508 ( \2750 , \766 , \961 );
nor \U$2509 ( \2751 , \2749 , \2750 );
xnor \U$2510 ( \2752 , \2751 , \568 );
xor \U$2511 ( \2753 , \2748 , \2752 );
and \U$2512 ( \2754 , \847 , \1198 );
and \U$2513 ( \2755 , \794 , \1079 );
nor \U$2514 ( \2756 , \2754 , \2755 );
xnor \U$2515 ( \2757 , \2756 , \532 );
xor \U$2516 ( \2758 , \2753 , \2757 );
xor \U$2517 ( \2759 , \2744 , \2758 );
and \U$2518 ( \2760 , \700 , \872 );
and \U$2519 ( \2761 , \653 , \870 );
nor \U$2520 ( \2762 , \2760 , \2761 );
xnor \U$2521 ( \2763 , \2762 , \879 );
and \U$2522 ( \2764 , \728 , \900 );
and \U$2523 ( \2765 , \680 , \898 );
nor \U$2524 ( \2766 , \2764 , \2765 );
xnor \U$2525 ( \2767 , \2766 , \907 );
xor \U$2526 ( \2768 , \2763 , \2767 );
and \U$2527 ( \2769 , \759 , \930 );
and \U$2528 ( \2770 , \708 , \928 );
nor \U$2529 ( \2771 , \2769 , \2770 );
xnor \U$2530 ( \2772 , \2771 , \937 );
xor \U$2531 ( \2773 , \2768 , \2772 );
xor \U$2532 ( \2774 , \2759 , \2773 );
xor \U$2533 ( \2775 , \2741 , \2774 );
xor \U$2534 ( \2776 , \2715 , \2775 );
and \U$2535 ( \2777 , \2582 , \2586 );
and \U$2536 ( \2778 , \2586 , \2591 );
and \U$2537 ( \2779 , \2582 , \2591 );
or \U$2538 ( \2780 , \2777 , \2778 , \2779 );
and \U$2539 ( \2781 , \2666 , \2670 );
and \U$2540 ( \2782 , \2670 , \2679 );
and \U$2541 ( \2783 , \2666 , \2679 );
or \U$2542 ( \2784 , \2781 , \2782 , \2783 );
xor \U$2543 ( \2785 , \2780 , \2784 );
and \U$2544 ( \2786 , \2631 , \2645 );
and \U$2545 ( \2787 , \2645 , \2660 );
and \U$2546 ( \2788 , \2631 , \2660 );
or \U$2547 ( \2789 , \2786 , \2787 , \2788 );
xor \U$2548 ( \2790 , \2785 , \2789 );
xor \U$2549 ( \2791 , \2776 , \2790 );
xor \U$2550 ( \2792 , \2701 , \2791 );
and \U$2551 ( \2793 , \2559 , \2563 );
and \U$2552 ( \2794 , \2563 , \2568 );
and \U$2553 ( \2795 , \2559 , \2568 );
or \U$2554 ( \2796 , \2793 , \2794 , \2795 );
and \U$2555 ( \2797 , \2617 , \2661 );
and \U$2556 ( \2798 , \2661 , \2680 );
and \U$2557 ( \2799 , \2617 , \2680 );
or \U$2558 ( \2800 , \2797 , \2798 , \2799 );
xor \U$2559 ( \2801 , \2796 , \2800 );
and \U$2560 ( \2802 , \2621 , \2625 );
and \U$2561 ( \2803 , \2625 , \2630 );
and \U$2562 ( \2804 , \2621 , \2630 );
or \U$2563 ( \2805 , \2802 , \2803 , \2804 );
or \U$2564 ( \2806 , \2675 , \2678 );
xor \U$2565 ( \2807 , \2805 , \2806 );
and \U$2566 ( \2808 , \874 , \497 );
and \U$2567 ( \2809 , \827 , \495 );
nor \U$2568 ( \2810 , \2808 , \2809 );
xnor \U$2569 ( \2811 , \2810 , \502 );
xor \U$2570 ( \2812 , \2807 , \2811 );
xor \U$2571 ( \2813 , \2801 , \2812 );
xor \U$2572 ( \2814 , \2792 , \2813 );
xor \U$2573 ( \2815 , \2697 , \2814 );
and \U$2574 ( \2816 , \2555 , \2594 );
and \U$2575 ( \2817 , \2594 , \2682 );
and \U$2576 ( \2818 , \2555 , \2682 );
or \U$2577 ( \2819 , \2816 , \2817 , \2818 );
nor \U$2578 ( \2820 , \2815 , \2819 );
and \U$2579 ( \2821 , \2701 , \2791 );
and \U$2580 ( \2822 , \2791 , \2813 );
and \U$2581 ( \2823 , \2701 , \2813 );
or \U$2582 ( \2824 , \2821 , \2822 , \2823 );
and \U$2583 ( \2825 , \2780 , \2784 );
and \U$2584 ( \2826 , \2784 , \2789 );
and \U$2585 ( \2827 , \2780 , \2789 );
or \U$2586 ( \2828 , \2825 , \2826 , \2827 );
and \U$2587 ( \2829 , \2729 , \2740 );
and \U$2588 ( \2830 , \2740 , \2774 );
and \U$2589 ( \2831 , \2729 , \2774 );
or \U$2590 ( \2832 , \2829 , \2830 , \2831 );
xor \U$2591 ( \2833 , \2828 , \2832 );
and \U$2592 ( \2834 , \680 , \900 );
and \U$2593 ( \2835 , \700 , \898 );
nor \U$2594 ( \2836 , \2834 , \2835 );
xnor \U$2595 ( \2837 , \2836 , \907 );
and \U$2596 ( \2838 , \708 , \930 );
and \U$2597 ( \2839 , \728 , \928 );
nor \U$2598 ( \2840 , \2838 , \2839 );
xnor \U$2599 ( \2841 , \2840 , \937 );
xor \U$2600 ( \2842 , \2837 , \2841 );
and \U$2601 ( \2843 , \739 , \950 );
and \U$2602 ( \2844 , \759 , \948 );
nor \U$2603 ( \2845 , \2843 , \2844 );
xnor \U$2604 ( \2846 , \2845 , \957 );
xor \U$2605 ( \2847 , \2842 , \2846 );
and \U$2606 ( \2848 , \569 , \812 );
and \U$2607 ( \2849 , \618 , \810 );
nor \U$2608 ( \2850 , \2848 , \2849 );
xnor \U$2609 ( \2851 , \2850 , \819 );
and \U$2610 ( \2852 , \623 , \845 );
and \U$2611 ( \2853 , \643 , \843 );
nor \U$2612 ( \2854 , \2852 , \2853 );
xnor \U$2613 ( \2855 , \2854 , \852 );
xor \U$2614 ( \2856 , \2851 , \2855 );
and \U$2615 ( \2857 , \653 , \872 );
and \U$2616 ( \2858 , \673 , \870 );
nor \U$2617 ( \2859 , \2857 , \2858 );
xnor \U$2618 ( \2860 , \2859 , \879 );
xor \U$2619 ( \2861 , \2856 , \2860 );
xor \U$2620 ( \2862 , \2847 , \2861 );
and \U$2621 ( \2863 , \223 , \726 );
not \U$2622 ( \2864 , \2863 );
xnor \U$2623 ( \2865 , \2864 , \733 );
and \U$2624 ( \2866 , \539 , \757 );
and \U$2625 ( \2867 , \504 , \755 );
nor \U$2626 ( \2868 , \2866 , \2867 );
xnor \U$2627 ( \2869 , \2868 , \764 );
xor \U$2628 ( \2870 , \2865 , \2869 );
and \U$2629 ( \2871 , \1018 , \784 );
and \U$2630 ( \2872 , \1020 , \782 );
nor \U$2631 ( \2873 , \2871 , \2872 );
xnor \U$2632 ( \2874 , \2873 , \791 );
xor \U$2633 ( \2875 , \2870 , \2874 );
xor \U$2634 ( \2876 , \2862 , \2875 );
and \U$2635 ( \2877 , \2748 , \2752 );
and \U$2636 ( \2878 , \2752 , \2757 );
and \U$2637 ( \2879 , \2748 , \2757 );
or \U$2638 ( \2880 , \2877 , \2878 , \2879 );
and \U$2640 ( \2881 , \874 , \505 );
nor \U$2641 ( \2882 , 1'b0 , \2881 );
xor \U$2642 ( \2883 , \2880 , \2882 );
and \U$2643 ( \2884 , \766 , \978 );
and \U$2644 ( \2885 , \786 , \961 );
nor \U$2645 ( \2886 , \2884 , \2885 );
xnor \U$2646 ( \2887 , \2886 , \568 );
and \U$2647 ( \2888 , \794 , \1198 );
and \U$2648 ( \2889 , \814 , \1079 );
nor \U$2649 ( \2890 , \2888 , \2889 );
xnor \U$2650 ( \2891 , \2890 , \532 );
xor \U$2651 ( \2892 , \2887 , \2891 );
and \U$2652 ( \2893 , \827 , \497 );
and \U$2653 ( \2894 , \847 , \495 );
nor \U$2654 ( \2895 , \2893 , \2894 );
xnor \U$2655 ( \2896 , \2895 , \502 );
xor \U$2656 ( \2897 , \2892 , \2896 );
xor \U$2657 ( \2898 , \2883 , \2897 );
xor \U$2658 ( \2899 , \2876 , \2898 );
and \U$2659 ( \2900 , \2730 , \2734 );
and \U$2660 ( \2901 , \2734 , \2739 );
and \U$2661 ( \2902 , \2730 , \2739 );
or \U$2662 ( \2903 , \2900 , \2901 , \2902 );
and \U$2663 ( \2904 , \2719 , \2723 );
and \U$2664 ( \2905 , \2723 , \2728 );
and \U$2665 ( \2906 , \2719 , \2728 );
or \U$2666 ( \2907 , \2904 , \2905 , \2906 );
xor \U$2667 ( \2908 , \2903 , \2907 );
and \U$2668 ( \2909 , \2763 , \2767 );
and \U$2669 ( \2910 , \2767 , \2772 );
and \U$2670 ( \2911 , \2763 , \2772 );
or \U$2671 ( \2912 , \2909 , \2910 , \2911 );
xor \U$2672 ( \2913 , \2908 , \2912 );
xor \U$2673 ( \2914 , \2899 , \2913 );
xor \U$2674 ( \2915 , \2833 , \2914 );
xor \U$2675 ( \2916 , \2824 , \2915 );
and \U$2676 ( \2917 , \2796 , \2800 );
and \U$2677 ( \2918 , \2800 , \2812 );
and \U$2678 ( \2919 , \2796 , \2812 );
or \U$2679 ( \2920 , \2917 , \2918 , \2919 );
and \U$2680 ( \2921 , \2715 , \2775 );
and \U$2681 ( \2922 , \2775 , \2790 );
and \U$2682 ( \2923 , \2715 , \2790 );
or \U$2683 ( \2924 , \2921 , \2922 , \2923 );
xor \U$2684 ( \2925 , \2920 , \2924 );
and \U$2685 ( \2926 , \2705 , \2709 );
and \U$2686 ( \2927 , \2709 , \2714 );
and \U$2687 ( \2928 , \2705 , \2714 );
or \U$2688 ( \2929 , \2926 , \2927 , \2928 );
and \U$2689 ( \2930 , \2805 , \2806 );
and \U$2690 ( \2931 , \2806 , \2811 );
and \U$2691 ( \2932 , \2805 , \2811 );
or \U$2692 ( \2933 , \2930 , \2931 , \2932 );
xor \U$2693 ( \2934 , \2929 , \2933 );
and \U$2694 ( \2935 , \2744 , \2758 );
and \U$2695 ( \2936 , \2758 , \2773 );
and \U$2696 ( \2937 , \2744 , \2773 );
or \U$2697 ( \2938 , \2935 , \2936 , \2937 );
xor \U$2698 ( \2939 , \2934 , \2938 );
xor \U$2699 ( \2940 , \2925 , \2939 );
xor \U$2700 ( \2941 , \2916 , \2940 );
and \U$2701 ( \2942 , \2695 , \2696 );
and \U$2702 ( \2943 , \2696 , \2814 );
and \U$2703 ( \2944 , \2695 , \2814 );
or \U$2704 ( \2945 , \2942 , \2943 , \2944 );
nor \U$2705 ( \2946 , \2941 , \2945 );
nor \U$2706 ( \2947 , \2820 , \2946 );
and \U$2707 ( \2948 , \2920 , \2924 );
and \U$2708 ( \2949 , \2924 , \2939 );
and \U$2709 ( \2950 , \2920 , \2939 );
or \U$2710 ( \2951 , \2948 , \2949 , \2950 );
and \U$2711 ( \2952 , \2828 , \2832 );
and \U$2712 ( \2953 , \2832 , \2914 );
and \U$2713 ( \2954 , \2828 , \2914 );
or \U$2714 ( \2955 , \2952 , \2953 , \2954 );
not \U$2715 ( \2956 , \733 );
and \U$2716 ( \2957 , \504 , \757 );
and \U$2717 ( \2958 , \223 , \755 );
nor \U$2718 ( \2959 , \2957 , \2958 );
xnor \U$2719 ( \2960 , \2959 , \764 );
xor \U$2720 ( \2961 , \2956 , \2960 );
and \U$2721 ( \2962 , \1020 , \784 );
and \U$2722 ( \2963 , \539 , \782 );
nor \U$2723 ( \2964 , \2962 , \2963 );
xnor \U$2724 ( \2965 , \2964 , \791 );
xor \U$2725 ( \2966 , \2961 , \2965 );
and \U$2726 ( \2967 , \786 , \978 );
and \U$2727 ( \2968 , \739 , \961 );
nor \U$2728 ( \2969 , \2967 , \2968 );
xnor \U$2729 ( \2970 , \2969 , \568 );
and \U$2730 ( \2971 , \814 , \1198 );
and \U$2731 ( \2972 , \766 , \1079 );
nor \U$2732 ( \2973 , \2971 , \2972 );
xnor \U$2733 ( \2974 , \2973 , \532 );
xor \U$2734 ( \2975 , \2970 , \2974 );
and \U$2735 ( \2976 , \847 , \497 );
and \U$2736 ( \2977 , \794 , \495 );
nor \U$2737 ( \2978 , \2976 , \2977 );
xnor \U$2738 ( \2979 , \2978 , \502 );
xor \U$2739 ( \2980 , \2975 , \2979 );
and \U$2740 ( \2981 , \700 , \900 );
and \U$2741 ( \2982 , \653 , \898 );
nor \U$2742 ( \2983 , \2981 , \2982 );
xnor \U$2743 ( \2984 , \2983 , \907 );
and \U$2744 ( \2985 , \728 , \930 );
and \U$2745 ( \2986 , \680 , \928 );
nor \U$2746 ( \2987 , \2985 , \2986 );
xnor \U$2747 ( \2988 , \2987 , \937 );
xor \U$2748 ( \2989 , \2984 , \2988 );
and \U$2749 ( \2990 , \759 , \950 );
and \U$2750 ( \2991 , \708 , \948 );
nor \U$2751 ( \2992 , \2990 , \2991 );
xnor \U$2752 ( \2993 , \2992 , \957 );
xor \U$2753 ( \2994 , \2989 , \2993 );
xor \U$2754 ( \2995 , \2980 , \2994 );
and \U$2755 ( \2996 , \618 , \812 );
and \U$2756 ( \2997 , \1018 , \810 );
nor \U$2757 ( \2998 , \2996 , \2997 );
xnor \U$2758 ( \2999 , \2998 , \819 );
and \U$2759 ( \3000 , \643 , \845 );
and \U$2760 ( \3001 , \569 , \843 );
nor \U$2761 ( \3002 , \3000 , \3001 );
xnor \U$2762 ( \3003 , \3002 , \852 );
xor \U$2763 ( \3004 , \2999 , \3003 );
and \U$2764 ( \3005 , \673 , \872 );
and \U$2765 ( \3006 , \623 , \870 );
nor \U$2766 ( \3007 , \3005 , \3006 );
xnor \U$2767 ( \3008 , \3007 , \879 );
xor \U$2768 ( \3009 , \3004 , \3008 );
xor \U$2769 ( \3010 , \2995 , \3009 );
xor \U$2770 ( \3011 , \2966 , \3010 );
and \U$2771 ( \3012 , \2887 , \2891 );
and \U$2772 ( \3013 , \2891 , \2896 );
and \U$2773 ( \3014 , \2887 , \2896 );
or \U$2774 ( \3015 , \3012 , \3013 , \3014 );
not \U$2775 ( \3016 , \2882 );
xor \U$2776 ( \3017 , \3015 , \3016 );
and \U$2778 ( \3018 , \827 , \505 );
nor \U$2779 ( \3019 , 1'b0 , \3018 );
not \U$2780 ( \3020 , \3019 );
xor \U$2781 ( \3021 , \3017 , \3020 );
xor \U$2782 ( \3022 , \3011 , \3021 );
and \U$2783 ( \3023 , \2903 , \2907 );
and \U$2784 ( \3024 , \2907 , \2912 );
and \U$2785 ( \3025 , \2903 , \2912 );
or \U$2786 ( \3026 , \3023 , \3024 , \3025 );
and \U$2787 ( \3027 , \2880 , \2882 );
and \U$2788 ( \3028 , \2882 , \2897 );
and \U$2789 ( \3029 , \2880 , \2897 );
or \U$2790 ( \3030 , \3027 , \3028 , \3029 );
xor \U$2791 ( \3031 , \3026 , \3030 );
and \U$2792 ( \3032 , \2847 , \2861 );
and \U$2793 ( \3033 , \2861 , \2875 );
and \U$2794 ( \3034 , \2847 , \2875 );
or \U$2795 ( \3035 , \3032 , \3033 , \3034 );
xor \U$2796 ( \3036 , \3031 , \3035 );
xor \U$2797 ( \3037 , \3022 , \3036 );
xor \U$2798 ( \3038 , \2955 , \3037 );
and \U$2799 ( \3039 , \2929 , \2933 );
and \U$2800 ( \3040 , \2933 , \2938 );
and \U$2801 ( \3041 , \2929 , \2938 );
or \U$2802 ( \3042 , \3039 , \3040 , \3041 );
and \U$2803 ( \3043 , \2876 , \2898 );
and \U$2804 ( \3044 , \2898 , \2913 );
and \U$2805 ( \3045 , \2876 , \2913 );
or \U$2806 ( \3046 , \3043 , \3044 , \3045 );
xor \U$2807 ( \3047 , \3042 , \3046 );
and \U$2808 ( \3048 , \2865 , \2869 );
and \U$2809 ( \3049 , \2869 , \2874 );
and \U$2810 ( \3050 , \2865 , \2874 );
or \U$2811 ( \3051 , \3048 , \3049 , \3050 );
and \U$2812 ( \3052 , \2851 , \2855 );
and \U$2813 ( \3053 , \2855 , \2860 );
and \U$2814 ( \3054 , \2851 , \2860 );
or \U$2815 ( \3055 , \3052 , \3053 , \3054 );
xor \U$2816 ( \3056 , \3051 , \3055 );
and \U$2817 ( \3057 , \2837 , \2841 );
and \U$2818 ( \3058 , \2841 , \2846 );
and \U$2819 ( \3059 , \2837 , \2846 );
or \U$2820 ( \3060 , \3057 , \3058 , \3059 );
xor \U$2821 ( \3061 , \3056 , \3060 );
xor \U$2822 ( \3062 , \3047 , \3061 );
xor \U$2823 ( \3063 , \3038 , \3062 );
xor \U$2824 ( \3064 , \2951 , \3063 );
and \U$2825 ( \3065 , \2824 , \2915 );
and \U$2826 ( \3066 , \2915 , \2940 );
and \U$2827 ( \3067 , \2824 , \2940 );
or \U$2828 ( \3068 , \3065 , \3066 , \3067 );
nor \U$2829 ( \3069 , \3064 , \3068 );
and \U$2830 ( \3070 , \2955 , \3037 );
and \U$2831 ( \3071 , \3037 , \3062 );
and \U$2832 ( \3072 , \2955 , \3062 );
or \U$2833 ( \3073 , \3070 , \3071 , \3072 );
and \U$2834 ( \3074 , \3026 , \3030 );
and \U$2835 ( \3075 , \3030 , \3035 );
and \U$2836 ( \3076 , \3026 , \3035 );
or \U$2837 ( \3077 , \3074 , \3075 , \3076 );
and \U$2838 ( \3078 , \2966 , \3010 );
and \U$2839 ( \3079 , \3010 , \3021 );
and \U$2840 ( \3080 , \2966 , \3021 );
or \U$2841 ( \3081 , \3078 , \3079 , \3080 );
xor \U$2842 ( \3082 , \3077 , \3081 );
and \U$2843 ( \3083 , \680 , \930 );
and \U$2844 ( \3084 , \700 , \928 );
nor \U$2845 ( \3085 , \3083 , \3084 );
xnor \U$2846 ( \3086 , \3085 , \937 );
and \U$2847 ( \3087 , \708 , \950 );
and \U$2848 ( \3088 , \728 , \948 );
nor \U$2849 ( \3089 , \3087 , \3088 );
xnor \U$2850 ( \3090 , \3089 , \957 );
xor \U$2851 ( \3091 , \3086 , \3090 );
and \U$2852 ( \3092 , \739 , \978 );
and \U$2853 ( \3093 , \759 , \961 );
nor \U$2854 ( \3094 , \3092 , \3093 );
xnor \U$2855 ( \3095 , \3094 , \568 );
xor \U$2856 ( \3096 , \3091 , \3095 );
and \U$2857 ( \3097 , \569 , \845 );
and \U$2858 ( \3098 , \618 , \843 );
nor \U$2859 ( \3099 , \3097 , \3098 );
xnor \U$2860 ( \3100 , \3099 , \852 );
and \U$2861 ( \3101 , \623 , \872 );
and \U$2862 ( \3102 , \643 , \870 );
nor \U$2863 ( \3103 , \3101 , \3102 );
xnor \U$2864 ( \3104 , \3103 , \879 );
xor \U$2865 ( \3105 , \3100 , \3104 );
and \U$2866 ( \3106 , \653 , \900 );
and \U$2867 ( \3107 , \673 , \898 );
nor \U$2868 ( \3108 , \3106 , \3107 );
xnor \U$2869 ( \3109 , \3108 , \907 );
xor \U$2870 ( \3110 , \3105 , \3109 );
xor \U$2871 ( \3111 , \3096 , \3110 );
and \U$2872 ( \3112 , \223 , \757 );
not \U$2873 ( \3113 , \3112 );
xnor \U$2874 ( \3114 , \3113 , \764 );
and \U$2875 ( \3115 , \539 , \784 );
and \U$2876 ( \3116 , \504 , \782 );
nor \U$2877 ( \3117 , \3115 , \3116 );
xnor \U$2878 ( \3118 , \3117 , \791 );
xor \U$2879 ( \3119 , \3114 , \3118 );
and \U$2880 ( \3120 , \1018 , \812 );
and \U$2881 ( \3121 , \1020 , \810 );
nor \U$2882 ( \3122 , \3120 , \3121 );
xnor \U$2883 ( \3123 , \3122 , \819 );
xor \U$2884 ( \3124 , \3119 , \3123 );
xor \U$2885 ( \3125 , \3111 , \3124 );
and \U$2886 ( \3126 , \2970 , \2974 );
and \U$2887 ( \3127 , \2974 , \2979 );
and \U$2888 ( \3128 , \2970 , \2979 );
or \U$2889 ( \3129 , \3126 , \3127 , \3128 );
and \U$2890 ( \3130 , \766 , \1198 );
and \U$2891 ( \3131 , \786 , \1079 );
nor \U$2892 ( \3132 , \3130 , \3131 );
xnor \U$2893 ( \3133 , \3132 , \532 );
and \U$2894 ( \3134 , \794 , \497 );
and \U$2895 ( \3135 , \814 , \495 );
nor \U$2896 ( \3136 , \3134 , \3135 );
xnor \U$2897 ( \3137 , \3136 , \502 );
xor \U$2898 ( \3138 , \3133 , \3137 );
and \U$2900 ( \3139 , \847 , \505 );
nor \U$2901 ( \3140 , 1'b0 , \3139 );
not \U$2902 ( \3141 , \3140 );
xor \U$2903 ( \3142 , \3138 , \3141 );
xnor \U$2904 ( \3143 , \3129 , \3142 );
xor \U$2905 ( \3144 , \3125 , \3143 );
and \U$2906 ( \3145 , \2956 , \2960 );
and \U$2907 ( \3146 , \2960 , \2965 );
and \U$2908 ( \3147 , \2956 , \2965 );
or \U$2909 ( \3148 , \3145 , \3146 , \3147 );
and \U$2910 ( \3149 , \2999 , \3003 );
and \U$2911 ( \3150 , \3003 , \3008 );
and \U$2912 ( \3151 , \2999 , \3008 );
or \U$2913 ( \3152 , \3149 , \3150 , \3151 );
xor \U$2914 ( \3153 , \3148 , \3152 );
and \U$2915 ( \3154 , \2984 , \2988 );
and \U$2916 ( \3155 , \2988 , \2993 );
and \U$2917 ( \3156 , \2984 , \2993 );
or \U$2918 ( \3157 , \3154 , \3155 , \3156 );
xor \U$2919 ( \3158 , \3153 , \3157 );
xor \U$2920 ( \3159 , \3144 , \3158 );
xor \U$2921 ( \3160 , \3082 , \3159 );
xor \U$2922 ( \3161 , \3073 , \3160 );
and \U$2923 ( \3162 , \3042 , \3046 );
and \U$2924 ( \3163 , \3046 , \3061 );
and \U$2925 ( \3164 , \3042 , \3061 );
or \U$2926 ( \3165 , \3162 , \3163 , \3164 );
and \U$2927 ( \3166 , \3022 , \3036 );
xor \U$2928 ( \3167 , \3165 , \3166 );
and \U$2929 ( \3168 , \3051 , \3055 );
and \U$2930 ( \3169 , \3055 , \3060 );
and \U$2931 ( \3170 , \3051 , \3060 );
or \U$2932 ( \3171 , \3168 , \3169 , \3170 );
and \U$2933 ( \3172 , \3015 , \3016 );
and \U$2934 ( \3173 , \3016 , \3020 );
and \U$2935 ( \3174 , \3015 , \3020 );
or \U$2936 ( \3175 , \3172 , \3173 , \3174 );
xor \U$2937 ( \3176 , \3171 , \3175 );
and \U$2938 ( \3177 , \2980 , \2994 );
and \U$2939 ( \3178 , \2994 , \3009 );
and \U$2940 ( \3179 , \2980 , \3009 );
or \U$2941 ( \3180 , \3177 , \3178 , \3179 );
xor \U$2942 ( \3181 , \3176 , \3180 );
xor \U$2943 ( \3182 , \3167 , \3181 );
xor \U$2944 ( \3183 , \3161 , \3182 );
and \U$2945 ( \3184 , \2951 , \3063 );
nor \U$2946 ( \3185 , \3183 , \3184 );
nor \U$2947 ( \3186 , \3069 , \3185 );
nand \U$2948 ( \3187 , \2947 , \3186 );
and \U$2949 ( \3188 , \3165 , \3166 );
and \U$2950 ( \3189 , \3166 , \3181 );
and \U$2951 ( \3190 , \3165 , \3181 );
or \U$2952 ( \3191 , \3188 , \3189 , \3190 );
and \U$2953 ( \3192 , \3077 , \3081 );
and \U$2954 ( \3193 , \3081 , \3159 );
and \U$2955 ( \3194 , \3077 , \3159 );
or \U$2956 ( \3195 , \3192 , \3193 , \3194 );
and \U$2957 ( \3196 , \3148 , \3152 );
and \U$2958 ( \3197 , \3152 , \3157 );
and \U$2959 ( \3198 , \3148 , \3157 );
or \U$2960 ( \3199 , \3196 , \3197 , \3198 );
or \U$2961 ( \3200 , \3129 , \3142 );
xor \U$2962 ( \3201 , \3199 , \3200 );
and \U$2963 ( \3202 , \3096 , \3110 );
and \U$2964 ( \3203 , \3110 , \3124 );
and \U$2965 ( \3204 , \3096 , \3124 );
or \U$2966 ( \3205 , \3202 , \3203 , \3204 );
xor \U$2967 ( \3206 , \3201 , \3205 );
xor \U$2968 ( \3207 , \3195 , \3206 );
and \U$2969 ( \3208 , \3171 , \3175 );
and \U$2970 ( \3209 , \3175 , \3180 );
and \U$2971 ( \3210 , \3171 , \3180 );
or \U$2972 ( \3211 , \3208 , \3209 , \3210 );
and \U$2973 ( \3212 , \3125 , \3143 );
and \U$2974 ( \3213 , \3143 , \3158 );
and \U$2975 ( \3214 , \3125 , \3158 );
or \U$2976 ( \3215 , \3212 , \3213 , \3214 );
xor \U$2977 ( \3216 , \3211 , \3215 );
and \U$2978 ( \3217 , \618 , \845 );
and \U$2979 ( \3218 , \1018 , \843 );
nor \U$2980 ( \3219 , \3217 , \3218 );
xnor \U$2981 ( \3220 , \3219 , \852 );
and \U$2982 ( \3221 , \643 , \872 );
and \U$2983 ( \3222 , \569 , \870 );
nor \U$2984 ( \3223 , \3221 , \3222 );
xnor \U$2985 ( \3224 , \3223 , \879 );
xor \U$2986 ( \3225 , \3220 , \3224 );
and \U$2987 ( \3226 , \673 , \900 );
and \U$2988 ( \3227 , \623 , \898 );
nor \U$2989 ( \3228 , \3226 , \3227 );
xnor \U$2990 ( \3229 , \3228 , \907 );
xor \U$2991 ( \3230 , \3225 , \3229 );
not \U$2992 ( \3231 , \764 );
and \U$2993 ( \3232 , \504 , \784 );
and \U$2994 ( \3233 , \223 , \782 );
nor \U$2995 ( \3234 , \3232 , \3233 );
xnor \U$2996 ( \3235 , \3234 , \791 );
xor \U$2997 ( \3236 , \3231 , \3235 );
and \U$2998 ( \3237 , \1020 , \812 );
and \U$2999 ( \3238 , \539 , \810 );
nor \U$3000 ( \3239 , \3237 , \3238 );
xnor \U$3001 ( \3240 , \3239 , \819 );
xor \U$3002 ( \3241 , \3236 , \3240 );
xor \U$3003 ( \3242 , \3230 , \3241 );
and \U$3004 ( \3243 , \3133 , \3137 );
and \U$3005 ( \3244 , \3137 , \3141 );
and \U$3006 ( \3245 , \3133 , \3141 );
or \U$3007 ( \3246 , \3243 , \3244 , \3245 );
and \U$3008 ( \3247 , \786 , \1198 );
and \U$3009 ( \3248 , \739 , \1079 );
nor \U$3010 ( \3249 , \3247 , \3248 );
xnor \U$3011 ( \3250 , \3249 , \532 );
and \U$3012 ( \3251 , \814 , \497 );
and \U$3013 ( \3252 , \766 , \495 );
nor \U$3014 ( \3253 , \3251 , \3252 );
xnor \U$3015 ( \3254 , \3253 , \502 );
xor \U$3016 ( \3255 , \3250 , \3254 );
and \U$3018 ( \3256 , \794 , \505 );
nor \U$3019 ( \3257 , 1'b0 , \3256 );
not \U$3020 ( \3258 , \3257 );
xor \U$3021 ( \3259 , \3255 , \3258 );
xor \U$3022 ( \3260 , \3246 , \3259 );
and \U$3023 ( \3261 , \700 , \930 );
and \U$3024 ( \3262 , \653 , \928 );
nor \U$3025 ( \3263 , \3261 , \3262 );
xnor \U$3026 ( \3264 , \3263 , \937 );
and \U$3027 ( \3265 , \728 , \950 );
and \U$3028 ( \3266 , \680 , \948 );
nor \U$3029 ( \3267 , \3265 , \3266 );
xnor \U$3030 ( \3268 , \3267 , \957 );
xor \U$3031 ( \3269 , \3264 , \3268 );
and \U$3032 ( \3270 , \759 , \978 );
and \U$3033 ( \3271 , \708 , \961 );
nor \U$3034 ( \3272 , \3270 , \3271 );
xnor \U$3035 ( \3273 , \3272 , \568 );
xor \U$3036 ( \3274 , \3269 , \3273 );
xor \U$3037 ( \3275 , \3260 , \3274 );
xor \U$3038 ( \3276 , \3242 , \3275 );
and \U$3039 ( \3277 , \3114 , \3118 );
and \U$3040 ( \3278 , \3118 , \3123 );
and \U$3041 ( \3279 , \3114 , \3123 );
or \U$3042 ( \3280 , \3277 , \3278 , \3279 );
and \U$3043 ( \3281 , \3100 , \3104 );
and \U$3044 ( \3282 , \3104 , \3109 );
and \U$3045 ( \3283 , \3100 , \3109 );
or \U$3046 ( \3284 , \3281 , \3282 , \3283 );
xor \U$3047 ( \3285 , \3280 , \3284 );
and \U$3048 ( \3286 , \3086 , \3090 );
and \U$3049 ( \3287 , \3090 , \3095 );
and \U$3050 ( \3288 , \3086 , \3095 );
or \U$3051 ( \3289 , \3286 , \3287 , \3288 );
xor \U$3052 ( \3290 , \3285 , \3289 );
xor \U$3053 ( \3291 , \3276 , \3290 );
xor \U$3054 ( \3292 , \3216 , \3291 );
xor \U$3055 ( \3293 , \3207 , \3292 );
xor \U$3056 ( \3294 , \3191 , \3293 );
and \U$3057 ( \3295 , \3073 , \3160 );
and \U$3058 ( \3296 , \3160 , \3182 );
and \U$3059 ( \3297 , \3073 , \3182 );
or \U$3060 ( \3298 , \3295 , \3296 , \3297 );
nor \U$3061 ( \3299 , \3294 , \3298 );
and \U$3062 ( \3300 , \3195 , \3206 );
and \U$3063 ( \3301 , \3206 , \3292 );
and \U$3064 ( \3302 , \3195 , \3292 );
or \U$3065 ( \3303 , \3300 , \3301 , \3302 );
and \U$3066 ( \3304 , \3211 , \3215 );
and \U$3067 ( \3305 , \3215 , \3291 );
and \U$3068 ( \3306 , \3211 , \3291 );
or \U$3069 ( \3307 , \3304 , \3305 , \3306 );
and \U$3070 ( \3308 , \3280 , \3284 );
and \U$3071 ( \3309 , \3284 , \3289 );
and \U$3072 ( \3310 , \3280 , \3289 );
or \U$3073 ( \3311 , \3308 , \3309 , \3310 );
and \U$3074 ( \3312 , \3246 , \3259 );
and \U$3075 ( \3313 , \3259 , \3274 );
and \U$3076 ( \3314 , \3246 , \3274 );
or \U$3077 ( \3315 , \3312 , \3313 , \3314 );
xor \U$3078 ( \3316 , \3311 , \3315 );
and \U$3079 ( \3317 , \3230 , \3241 );
xor \U$3080 ( \3318 , \3316 , \3317 );
xor \U$3081 ( \3319 , \3307 , \3318 );
and \U$3082 ( \3320 , \3199 , \3200 );
and \U$3083 ( \3321 , \3200 , \3205 );
and \U$3084 ( \3322 , \3199 , \3205 );
or \U$3085 ( \3323 , \3320 , \3321 , \3322 );
and \U$3086 ( \3324 , \3242 , \3275 );
and \U$3087 ( \3325 , \3275 , \3290 );
and \U$3088 ( \3326 , \3242 , \3290 );
or \U$3089 ( \3327 , \3324 , \3325 , \3326 );
xor \U$3090 ( \3328 , \3323 , \3327 );
and \U$3091 ( \3329 , \569 , \872 );
and \U$3092 ( \3330 , \618 , \870 );
nor \U$3093 ( \3331 , \3329 , \3330 );
xnor \U$3094 ( \3332 , \3331 , \879 );
and \U$3095 ( \3333 , \623 , \900 );
and \U$3096 ( \3334 , \643 , \898 );
nor \U$3097 ( \3335 , \3333 , \3334 );
xnor \U$3098 ( \3336 , \3335 , \907 );
xor \U$3099 ( \3337 , \3332 , \3336 );
and \U$3100 ( \3338 , \653 , \930 );
and \U$3101 ( \3339 , \673 , \928 );
nor \U$3102 ( \3340 , \3338 , \3339 );
xnor \U$3103 ( \3341 , \3340 , \937 );
xor \U$3104 ( \3342 , \3337 , \3341 );
and \U$3105 ( \3343 , \223 , \784 );
not \U$3106 ( \3344 , \3343 );
xnor \U$3107 ( \3345 , \3344 , \791 );
and \U$3108 ( \3346 , \539 , \812 );
and \U$3109 ( \3347 , \504 , \810 );
nor \U$3110 ( \3348 , \3346 , \3347 );
xnor \U$3111 ( \3349 , \3348 , \819 );
xor \U$3112 ( \3350 , \3345 , \3349 );
and \U$3113 ( \3351 , \1018 , \845 );
and \U$3114 ( \3352 , \1020 , \843 );
nor \U$3115 ( \3353 , \3351 , \3352 );
xnor \U$3116 ( \3354 , \3353 , \852 );
xor \U$3117 ( \3355 , \3350 , \3354 );
xor \U$3118 ( \3356 , \3342 , \3355 );
and \U$3119 ( \3357 , \3250 , \3254 );
and \U$3120 ( \3358 , \3254 , \3258 );
and \U$3121 ( \3359 , \3250 , \3258 );
or \U$3122 ( \3360 , \3357 , \3358 , \3359 );
and \U$3123 ( \3361 , \766 , \497 );
and \U$3124 ( \3362 , \786 , \495 );
nor \U$3125 ( \3363 , \3361 , \3362 );
xnor \U$3126 ( \3364 , \3363 , \502 );
and \U$3128 ( \3365 , \814 , \505 );
nor \U$3129 ( \3366 , 1'b0 , \3365 );
not \U$3130 ( \3367 , \3366 );
xnor \U$3131 ( \3368 , \3364 , \3367 );
xor \U$3132 ( \3369 , \3360 , \3368 );
and \U$3133 ( \3370 , \680 , \950 );
and \U$3134 ( \3371 , \700 , \948 );
nor \U$3135 ( \3372 , \3370 , \3371 );
xnor \U$3136 ( \3373 , \3372 , \957 );
and \U$3137 ( \3374 , \708 , \978 );
and \U$3138 ( \3375 , \728 , \961 );
nor \U$3139 ( \3376 , \3374 , \3375 );
xnor \U$3140 ( \3377 , \3376 , \568 );
xor \U$3141 ( \3378 , \3373 , \3377 );
and \U$3142 ( \3379 , \739 , \1198 );
and \U$3143 ( \3380 , \759 , \1079 );
nor \U$3144 ( \3381 , \3379 , \3380 );
xnor \U$3145 ( \3382 , \3381 , \532 );
xor \U$3146 ( \3383 , \3378 , \3382 );
xor \U$3147 ( \3384 , \3369 , \3383 );
xor \U$3148 ( \3385 , \3356 , \3384 );
and \U$3149 ( \3386 , \3231 , \3235 );
and \U$3150 ( \3387 , \3235 , \3240 );
and \U$3151 ( \3388 , \3231 , \3240 );
or \U$3152 ( \3389 , \3386 , \3387 , \3388 );
and \U$3153 ( \3390 , \3220 , \3224 );
and \U$3154 ( \3391 , \3224 , \3229 );
and \U$3155 ( \3392 , \3220 , \3229 );
or \U$3156 ( \3393 , \3390 , \3391 , \3392 );
xor \U$3157 ( \3394 , \3389 , \3393 );
and \U$3158 ( \3395 , \3264 , \3268 );
and \U$3159 ( \3396 , \3268 , \3273 );
and \U$3160 ( \3397 , \3264 , \3273 );
or \U$3161 ( \3398 , \3395 , \3396 , \3397 );
xor \U$3162 ( \3399 , \3394 , \3398 );
xor \U$3163 ( \3400 , \3385 , \3399 );
xor \U$3164 ( \3401 , \3328 , \3400 );
xor \U$3165 ( \3402 , \3319 , \3401 );
xor \U$3166 ( \3403 , \3303 , \3402 );
and \U$3167 ( \3404 , \3191 , \3293 );
nor \U$3168 ( \3405 , \3403 , \3404 );
nor \U$3169 ( \3406 , \3299 , \3405 );
and \U$3170 ( \3407 , \3307 , \3318 );
and \U$3171 ( \3408 , \3318 , \3401 );
and \U$3172 ( \3409 , \3307 , \3401 );
or \U$3173 ( \3410 , \3407 , \3408 , \3409 );
and \U$3174 ( \3411 , \3323 , \3327 );
and \U$3175 ( \3412 , \3327 , \3400 );
and \U$3176 ( \3413 , \3323 , \3400 );
or \U$3177 ( \3414 , \3411 , \3412 , \3413 );
and \U$3178 ( \3415 , \3389 , \3393 );
and \U$3179 ( \3416 , \3393 , \3398 );
and \U$3180 ( \3417 , \3389 , \3398 );
or \U$3181 ( \3418 , \3415 , \3416 , \3417 );
and \U$3182 ( \3419 , \3360 , \3368 );
and \U$3183 ( \3420 , \3368 , \3383 );
and \U$3184 ( \3421 , \3360 , \3383 );
or \U$3185 ( \3422 , \3419 , \3420 , \3421 );
xor \U$3186 ( \3423 , \3418 , \3422 );
and \U$3187 ( \3424 , \3342 , \3355 );
xor \U$3188 ( \3425 , \3423 , \3424 );
xor \U$3189 ( \3426 , \3414 , \3425 );
and \U$3190 ( \3427 , \3311 , \3315 );
and \U$3191 ( \3428 , \3315 , \3317 );
and \U$3192 ( \3429 , \3311 , \3317 );
or \U$3193 ( \3430 , \3427 , \3428 , \3429 );
and \U$3194 ( \3431 , \3356 , \3384 );
and \U$3195 ( \3432 , \3384 , \3399 );
and \U$3196 ( \3433 , \3356 , \3399 );
or \U$3197 ( \3434 , \3431 , \3432 , \3433 );
xor \U$3198 ( \3435 , \3430 , \3434 );
and \U$3199 ( \3436 , \700 , \950 );
and \U$3200 ( \3437 , \653 , \948 );
nor \U$3201 ( \3438 , \3436 , \3437 );
xnor \U$3202 ( \3439 , \3438 , \957 );
and \U$3203 ( \3440 , \728 , \978 );
and \U$3204 ( \3441 , \680 , \961 );
nor \U$3205 ( \3442 , \3440 , \3441 );
xnor \U$3206 ( \3443 , \3442 , \568 );
xor \U$3207 ( \3444 , \3439 , \3443 );
and \U$3208 ( \3445 , \759 , \1198 );
and \U$3209 ( \3446 , \708 , \1079 );
nor \U$3210 ( \3447 , \3445 , \3446 );
xnor \U$3211 ( \3448 , \3447 , \532 );
xor \U$3212 ( \3449 , \3444 , \3448 );
and \U$3213 ( \3450 , \618 , \872 );
and \U$3214 ( \3451 , \1018 , \870 );
nor \U$3215 ( \3452 , \3450 , \3451 );
xnor \U$3216 ( \3453 , \3452 , \879 );
and \U$3217 ( \3454 , \643 , \900 );
and \U$3218 ( \3455 , \569 , \898 );
nor \U$3219 ( \3456 , \3454 , \3455 );
xnor \U$3220 ( \3457 , \3456 , \907 );
xor \U$3221 ( \3458 , \3453 , \3457 );
and \U$3222 ( \3459 , \673 , \930 );
and \U$3223 ( \3460 , \623 , \928 );
nor \U$3224 ( \3461 , \3459 , \3460 );
xnor \U$3225 ( \3462 , \3461 , \937 );
xor \U$3226 ( \3463 , \3458 , \3462 );
xor \U$3227 ( \3464 , \3449 , \3463 );
not \U$3228 ( \3465 , \791 );
and \U$3229 ( \3466 , \504 , \812 );
and \U$3230 ( \3467 , \223 , \810 );
nor \U$3231 ( \3468 , \3466 , \3467 );
xnor \U$3232 ( \3469 , \3468 , \819 );
xor \U$3233 ( \3470 , \3465 , \3469 );
and \U$3234 ( \3471 , \1020 , \845 );
and \U$3235 ( \3472 , \539 , \843 );
nor \U$3236 ( \3473 , \3471 , \3472 );
xnor \U$3237 ( \3474 , \3473 , \852 );
xor \U$3238 ( \3475 , \3470 , \3474 );
xor \U$3239 ( \3476 , \3464 , \3475 );
or \U$3240 ( \3477 , \3364 , \3367 );
and \U$3241 ( \3478 , \786 , \497 );
and \U$3242 ( \3479 , \739 , \495 );
nor \U$3243 ( \3480 , \3478 , \3479 );
xnor \U$3244 ( \3481 , \3480 , \502 );
xor \U$3245 ( \3482 , \3477 , \3481 );
and \U$3247 ( \3483 , \766 , \505 );
nor \U$3248 ( \3484 , 1'b0 , \3483 );
not \U$3249 ( \3485 , \3484 );
xor \U$3250 ( \3486 , \3482 , \3485 );
xor \U$3251 ( \3487 , \3476 , \3486 );
and \U$3252 ( \3488 , \3345 , \3349 );
and \U$3253 ( \3489 , \3349 , \3354 );
and \U$3254 ( \3490 , \3345 , \3354 );
or \U$3255 ( \3491 , \3488 , \3489 , \3490 );
and \U$3256 ( \3492 , \3332 , \3336 );
and \U$3257 ( \3493 , \3336 , \3341 );
and \U$3258 ( \3494 , \3332 , \3341 );
or \U$3259 ( \3495 , \3492 , \3493 , \3494 );
xor \U$3260 ( \3496 , \3491 , \3495 );
and \U$3261 ( \3497 , \3373 , \3377 );
and \U$3262 ( \3498 , \3377 , \3382 );
and \U$3263 ( \3499 , \3373 , \3382 );
or \U$3264 ( \3500 , \3497 , \3498 , \3499 );
xor \U$3265 ( \3501 , \3496 , \3500 );
xor \U$3266 ( \3502 , \3487 , \3501 );
xor \U$3267 ( \3503 , \3435 , \3502 );
xor \U$3268 ( \3504 , \3426 , \3503 );
xor \U$3269 ( \3505 , \3410 , \3504 );
and \U$3270 ( \3506 , \3303 , \3402 );
nor \U$3271 ( \3507 , \3505 , \3506 );
and \U$3272 ( \3508 , \3414 , \3425 );
and \U$3273 ( \3509 , \3425 , \3503 );
and \U$3274 ( \3510 , \3414 , \3503 );
or \U$3275 ( \3511 , \3508 , \3509 , \3510 );
and \U$3276 ( \3512 , \3430 , \3434 );
and \U$3277 ( \3513 , \3434 , \3502 );
and \U$3278 ( \3514 , \3430 , \3502 );
or \U$3279 ( \3515 , \3512 , \3513 , \3514 );
and \U$3280 ( \3516 , \3491 , \3495 );
and \U$3281 ( \3517 , \3495 , \3500 );
and \U$3282 ( \3518 , \3491 , \3500 );
or \U$3283 ( \3519 , \3516 , \3517 , \3518 );
and \U$3284 ( \3520 , \3477 , \3481 );
and \U$3285 ( \3521 , \3481 , \3485 );
and \U$3286 ( \3522 , \3477 , \3485 );
or \U$3287 ( \3523 , \3520 , \3521 , \3522 );
xor \U$3288 ( \3524 , \3519 , \3523 );
and \U$3289 ( \3525 , \3449 , \3463 );
and \U$3290 ( \3526 , \3463 , \3475 );
and \U$3291 ( \3527 , \3449 , \3475 );
or \U$3292 ( \3528 , \3525 , \3526 , \3527 );
xor \U$3293 ( \3529 , \3524 , \3528 );
xor \U$3294 ( \3530 , \3515 , \3529 );
and \U$3295 ( \3531 , \3418 , \3422 );
and \U$3296 ( \3532 , \3422 , \3424 );
and \U$3297 ( \3533 , \3418 , \3424 );
or \U$3298 ( \3534 , \3531 , \3532 , \3533 );
and \U$3299 ( \3535 , \3476 , \3486 );
and \U$3300 ( \3536 , \3486 , \3501 );
and \U$3301 ( \3537 , \3476 , \3501 );
or \U$3302 ( \3538 , \3535 , \3536 , \3537 );
xor \U$3303 ( \3539 , \3534 , \3538 );
and \U$3304 ( \3540 , \569 , \900 );
and \U$3305 ( \3541 , \618 , \898 );
nor \U$3306 ( \3542 , \3540 , \3541 );
xnor \U$3307 ( \3543 , \3542 , \907 );
and \U$3308 ( \3544 , \623 , \930 );
and \U$3309 ( \3545 , \643 , \928 );
nor \U$3310 ( \3546 , \3544 , \3545 );
xnor \U$3311 ( \3547 , \3546 , \937 );
xor \U$3312 ( \3548 , \3543 , \3547 );
and \U$3313 ( \3549 , \653 , \950 );
and \U$3314 ( \3550 , \673 , \948 );
nor \U$3315 ( \3551 , \3549 , \3550 );
xnor \U$3316 ( \3552 , \3551 , \957 );
xor \U$3317 ( \3553 , \3548 , \3552 );
and \U$3318 ( \3554 , \223 , \812 );
not \U$3319 ( \3555 , \3554 );
xnor \U$3320 ( \3556 , \3555 , \819 );
and \U$3321 ( \3557 , \539 , \845 );
and \U$3322 ( \3558 , \504 , \843 );
nor \U$3323 ( \3559 , \3557 , \3558 );
xnor \U$3324 ( \3560 , \3559 , \852 );
xor \U$3325 ( \3561 , \3556 , \3560 );
and \U$3326 ( \3562 , \1018 , \872 );
and \U$3327 ( \3563 , \1020 , \870 );
nor \U$3328 ( \3564 , \3562 , \3563 );
xnor \U$3329 ( \3565 , \3564 , \879 );
xor \U$3330 ( \3566 , \3561 , \3565 );
xor \U$3331 ( \3567 , \3553 , \3566 );
and \U$3333 ( \3568 , \786 , \505 );
nor \U$3334 ( \3569 , 1'b0 , \3568 );
not \U$3335 ( \3570 , \3569 );
and \U$3336 ( \3571 , \680 , \978 );
and \U$3337 ( \3572 , \700 , \961 );
nor \U$3338 ( \3573 , \3571 , \3572 );
xnor \U$3339 ( \3574 , \3573 , \568 );
and \U$3340 ( \3575 , \708 , \1198 );
and \U$3341 ( \3576 , \728 , \1079 );
nor \U$3342 ( \3577 , \3575 , \3576 );
xnor \U$3343 ( \3578 , \3577 , \532 );
xor \U$3344 ( \3579 , \3574 , \3578 );
and \U$3345 ( \3580 , \739 , \497 );
and \U$3346 ( \3581 , \759 , \495 );
nor \U$3347 ( \3582 , \3580 , \3581 );
xnor \U$3348 ( \3583 , \3582 , \502 );
xor \U$3349 ( \3584 , \3579 , \3583 );
xnor \U$3350 ( \3585 , \3570 , \3584 );
xor \U$3351 ( \3586 , \3567 , \3585 );
and \U$3352 ( \3587 , \3465 , \3469 );
and \U$3353 ( \3588 , \3469 , \3474 );
and \U$3354 ( \3589 , \3465 , \3474 );
or \U$3355 ( \3590 , \3587 , \3588 , \3589 );
and \U$3356 ( \3591 , \3453 , \3457 );
and \U$3357 ( \3592 , \3457 , \3462 );
and \U$3358 ( \3593 , \3453 , \3462 );
or \U$3359 ( \3594 , \3591 , \3592 , \3593 );
xor \U$3360 ( \3595 , \3590 , \3594 );
and \U$3361 ( \3596 , \3439 , \3443 );
and \U$3362 ( \3597 , \3443 , \3448 );
and \U$3363 ( \3598 , \3439 , \3448 );
or \U$3364 ( \3599 , \3596 , \3597 , \3598 );
xor \U$3365 ( \3600 , \3595 , \3599 );
xor \U$3366 ( \3601 , \3586 , \3600 );
xor \U$3367 ( \3602 , \3539 , \3601 );
xor \U$3368 ( \3603 , \3530 , \3602 );
xor \U$3369 ( \3604 , \3511 , \3603 );
and \U$3370 ( \3605 , \3410 , \3504 );
nor \U$3371 ( \3606 , \3604 , \3605 );
nor \U$3372 ( \3607 , \3507 , \3606 );
nand \U$3373 ( \3608 , \3406 , \3607 );
nor \U$3374 ( \3609 , \3187 , \3608 );
nand \U$3375 ( \3610 , \2691 , \3609 );
and \U$3376 ( \3611 , \3515 , \3529 );
and \U$3377 ( \3612 , \3529 , \3602 );
and \U$3378 ( \3613 , \3515 , \3602 );
or \U$3379 ( \3614 , \3611 , \3612 , \3613 );
and \U$3380 ( \3615 , \3534 , \3538 );
and \U$3381 ( \3616 , \3538 , \3601 );
and \U$3382 ( \3617 , \3534 , \3601 );
or \U$3383 ( \3618 , \3615 , \3616 , \3617 );
and \U$3384 ( \3619 , \3590 , \3594 );
and \U$3385 ( \3620 , \3594 , \3599 );
and \U$3386 ( \3621 , \3590 , \3599 );
or \U$3387 ( \3622 , \3619 , \3620 , \3621 );
or \U$3388 ( \3623 , \3570 , \3584 );
xor \U$3389 ( \3624 , \3622 , \3623 );
and \U$3390 ( \3625 , \3553 , \3566 );
xor \U$3391 ( \3626 , \3624 , \3625 );
xor \U$3392 ( \3627 , \3618 , \3626 );
and \U$3393 ( \3628 , \3519 , \3523 );
and \U$3394 ( \3629 , \3523 , \3528 );
and \U$3395 ( \3630 , \3519 , \3528 );
or \U$3396 ( \3631 , \3628 , \3629 , \3630 );
and \U$3397 ( \3632 , \3567 , \3585 );
and \U$3398 ( \3633 , \3585 , \3600 );
and \U$3399 ( \3634 , \3567 , \3600 );
or \U$3400 ( \3635 , \3632 , \3633 , \3634 );
xor \U$3401 ( \3636 , \3631 , \3635 );
not \U$3402 ( \3637 , \819 );
and \U$3403 ( \3638 , \504 , \845 );
and \U$3404 ( \3639 , \223 , \843 );
nor \U$3405 ( \3640 , \3638 , \3639 );
xnor \U$3406 ( \3641 , \3640 , \852 );
xor \U$3407 ( \3642 , \3637 , \3641 );
and \U$3408 ( \3643 , \1020 , \872 );
and \U$3409 ( \3644 , \539 , \870 );
nor \U$3410 ( \3645 , \3643 , \3644 );
xnor \U$3411 ( \3646 , \3645 , \879 );
xor \U$3412 ( \3647 , \3642 , \3646 );
and \U$3414 ( \3648 , \739 , \505 );
nor \U$3415 ( \3649 , 1'b0 , \3648 );
not \U$3416 ( \3650 , \3649 );
and \U$3417 ( \3651 , \700 , \978 );
and \U$3418 ( \3652 , \653 , \961 );
nor \U$3419 ( \3653 , \3651 , \3652 );
xnor \U$3420 ( \3654 , \3653 , \568 );
and \U$3421 ( \3655 , \728 , \1198 );
and \U$3422 ( \3656 , \680 , \1079 );
nor \U$3423 ( \3657 , \3655 , \3656 );
xnor \U$3424 ( \3658 , \3657 , \532 );
xor \U$3425 ( \3659 , \3654 , \3658 );
and \U$3426 ( \3660 , \759 , \497 );
and \U$3427 ( \3661 , \708 , \495 );
nor \U$3428 ( \3662 , \3660 , \3661 );
xnor \U$3429 ( \3663 , \3662 , \502 );
xor \U$3430 ( \3664 , \3659 , \3663 );
xor \U$3431 ( \3665 , \3650 , \3664 );
and \U$3432 ( \3666 , \618 , \900 );
and \U$3433 ( \3667 , \1018 , \898 );
nor \U$3434 ( \3668 , \3666 , \3667 );
xnor \U$3435 ( \3669 , \3668 , \907 );
and \U$3436 ( \3670 , \643 , \930 );
and \U$3437 ( \3671 , \569 , \928 );
nor \U$3438 ( \3672 , \3670 , \3671 );
xnor \U$3439 ( \3673 , \3672 , \937 );
xor \U$3440 ( \3674 , \3669 , \3673 );
and \U$3441 ( \3675 , \673 , \950 );
and \U$3442 ( \3676 , \623 , \948 );
nor \U$3443 ( \3677 , \3675 , \3676 );
xnor \U$3444 ( \3678 , \3677 , \957 );
xor \U$3445 ( \3679 , \3674 , \3678 );
xor \U$3446 ( \3680 , \3665 , \3679 );
xor \U$3447 ( \3681 , \3647 , \3680 );
and \U$3448 ( \3682 , \3556 , \3560 );
and \U$3449 ( \3683 , \3560 , \3565 );
and \U$3450 ( \3684 , \3556 , \3565 );
or \U$3451 ( \3685 , \3682 , \3683 , \3684 );
and \U$3452 ( \3686 , \3543 , \3547 );
and \U$3453 ( \3687 , \3547 , \3552 );
and \U$3454 ( \3688 , \3543 , \3552 );
or \U$3455 ( \3689 , \3686 , \3687 , \3688 );
xor \U$3456 ( \3690 , \3685 , \3689 );
and \U$3457 ( \3691 , \3574 , \3578 );
and \U$3458 ( \3692 , \3578 , \3583 );
and \U$3459 ( \3693 , \3574 , \3583 );
or \U$3460 ( \3694 , \3691 , \3692 , \3693 );
xor \U$3461 ( \3695 , \3690 , \3694 );
xor \U$3462 ( \3696 , \3681 , \3695 );
xor \U$3463 ( \3697 , \3636 , \3696 );
xor \U$3464 ( \3698 , \3627 , \3697 );
xor \U$3465 ( \3699 , \3614 , \3698 );
and \U$3466 ( \3700 , \3511 , \3603 );
nor \U$3467 ( \3701 , \3699 , \3700 );
and \U$3468 ( \3702 , \3618 , \3626 );
and \U$3469 ( \3703 , \3626 , \3697 );
and \U$3470 ( \3704 , \3618 , \3697 );
or \U$3471 ( \3705 , \3702 , \3703 , \3704 );
and \U$3472 ( \3706 , \3631 , \3635 );
and \U$3473 ( \3707 , \3635 , \3696 );
and \U$3474 ( \3708 , \3631 , \3696 );
or \U$3475 ( \3709 , \3706 , \3707 , \3708 );
and \U$3476 ( \3710 , \3637 , \3641 );
and \U$3477 ( \3711 , \3641 , \3646 );
and \U$3478 ( \3712 , \3637 , \3646 );
or \U$3479 ( \3713 , \3710 , \3711 , \3712 );
and \U$3480 ( \3714 , \3669 , \3673 );
and \U$3481 ( \3715 , \3673 , \3678 );
and \U$3482 ( \3716 , \3669 , \3678 );
or \U$3483 ( \3717 , \3714 , \3715 , \3716 );
xor \U$3484 ( \3718 , \3713 , \3717 );
and \U$3485 ( \3719 , \3654 , \3658 );
and \U$3486 ( \3720 , \3658 , \3663 );
and \U$3487 ( \3721 , \3654 , \3663 );
or \U$3488 ( \3722 , \3719 , \3720 , \3721 );
xor \U$3489 ( \3723 , \3718 , \3722 );
and \U$3490 ( \3724 , \3685 , \3689 );
and \U$3491 ( \3725 , \3689 , \3694 );
and \U$3492 ( \3726 , \3685 , \3694 );
or \U$3493 ( \3727 , \3724 , \3725 , \3726 );
and \U$3494 ( \3728 , \3650 , \3664 );
and \U$3495 ( \3729 , \3664 , \3679 );
and \U$3496 ( \3730 , \3650 , \3679 );
or \U$3497 ( \3731 , \3728 , \3729 , \3730 );
xor \U$3498 ( \3732 , \3727 , \3731 );
and \U$3499 ( \3733 , \223 , \845 );
not \U$3500 ( \3734 , \3733 );
xnor \U$3501 ( \3735 , \3734 , \852 );
and \U$3502 ( \3736 , \539 , \872 );
and \U$3503 ( \3737 , \504 , \870 );
nor \U$3504 ( \3738 , \3736 , \3737 );
xnor \U$3505 ( \3739 , \3738 , \879 );
xor \U$3506 ( \3740 , \3735 , \3739 );
and \U$3507 ( \3741 , \1018 , \900 );
and \U$3508 ( \3742 , \1020 , \898 );
nor \U$3509 ( \3743 , \3741 , \3742 );
xnor \U$3510 ( \3744 , \3743 , \907 );
xor \U$3511 ( \3745 , \3740 , \3744 );
xor \U$3512 ( \3746 , \3732 , \3745 );
xor \U$3513 ( \3747 , \3723 , \3746 );
xor \U$3514 ( \3748 , \3709 , \3747 );
and \U$3515 ( \3749 , \3622 , \3623 );
and \U$3516 ( \3750 , \3623 , \3625 );
and \U$3517 ( \3751 , \3622 , \3625 );
or \U$3518 ( \3752 , \3749 , \3750 , \3751 );
and \U$3519 ( \3753 , \3647 , \3680 );
and \U$3520 ( \3754 , \3680 , \3695 );
and \U$3521 ( \3755 , \3647 , \3695 );
or \U$3522 ( \3756 , \3753 , \3754 , \3755 );
xor \U$3523 ( \3757 , \3752 , \3756 );
and \U$3524 ( \3758 , \680 , \1198 );
and \U$3525 ( \3759 , \700 , \1079 );
nor \U$3526 ( \3760 , \3758 , \3759 );
xnor \U$3527 ( \3761 , \3760 , \532 );
and \U$3528 ( \3762 , \708 , \497 );
and \U$3529 ( \3763 , \728 , \495 );
nor \U$3530 ( \3764 , \3762 , \3763 );
xnor \U$3531 ( \3765 , \3764 , \502 );
xor \U$3532 ( \3766 , \3761 , \3765 );
and \U$3534 ( \3767 , \759 , \505 );
nor \U$3535 ( \3768 , 1'b0 , \3767 );
not \U$3536 ( \3769 , \3768 );
xor \U$3537 ( \3770 , \3766 , \3769 );
and \U$3538 ( \3771 , \569 , \930 );
and \U$3539 ( \3772 , \618 , \928 );
nor \U$3540 ( \3773 , \3771 , \3772 );
xnor \U$3541 ( \3774 , \3773 , \937 );
and \U$3542 ( \3775 , \623 , \950 );
and \U$3543 ( \3776 , \643 , \948 );
nor \U$3544 ( \3777 , \3775 , \3776 );
xnor \U$3545 ( \3778 , \3777 , \957 );
xor \U$3546 ( \3779 , \3774 , \3778 );
and \U$3547 ( \3780 , \653 , \978 );
and \U$3548 ( \3781 , \673 , \961 );
nor \U$3549 ( \3782 , \3780 , \3781 );
xnor \U$3550 ( \3783 , \3782 , \568 );
xor \U$3551 ( \3784 , \3779 , \3783 );
xnor \U$3552 ( \3785 , \3770 , \3784 );
xor \U$3553 ( \3786 , \3757 , \3785 );
xor \U$3554 ( \3787 , \3748 , \3786 );
xor \U$3555 ( \3788 , \3705 , \3787 );
and \U$3556 ( \3789 , \3614 , \3698 );
nor \U$3557 ( \3790 , \3788 , \3789 );
nor \U$3558 ( \3791 , \3701 , \3790 );
and \U$3559 ( \3792 , \3709 , \3747 );
and \U$3560 ( \3793 , \3747 , \3786 );
and \U$3561 ( \3794 , \3709 , \3786 );
or \U$3562 ( \3795 , \3792 , \3793 , \3794 );
and \U$3563 ( \3796 , \3752 , \3756 );
and \U$3564 ( \3797 , \3756 , \3785 );
and \U$3565 ( \3798 , \3752 , \3785 );
or \U$3566 ( \3799 , \3796 , \3797 , \3798 );
and \U$3567 ( \3800 , \3723 , \3746 );
xor \U$3568 ( \3801 , \3799 , \3800 );
and \U$3569 ( \3802 , \3727 , \3731 );
and \U$3570 ( \3803 , \3731 , \3745 );
and \U$3571 ( \3804 , \3727 , \3745 );
or \U$3572 ( \3805 , \3802 , \3803 , \3804 );
and \U$3573 ( \3806 , \3735 , \3739 );
and \U$3574 ( \3807 , \3739 , \3744 );
and \U$3575 ( \3808 , \3735 , \3744 );
or \U$3576 ( \3809 , \3806 , \3807 , \3808 );
and \U$3577 ( \3810 , \3774 , \3778 );
and \U$3578 ( \3811 , \3778 , \3783 );
and \U$3579 ( \3812 , \3774 , \3783 );
or \U$3580 ( \3813 , \3810 , \3811 , \3812 );
xor \U$3581 ( \3814 , \3809 , \3813 );
and \U$3582 ( \3815 , \3761 , \3765 );
and \U$3583 ( \3816 , \3765 , \3769 );
and \U$3584 ( \3817 , \3761 , \3769 );
or \U$3585 ( \3818 , \3815 , \3816 , \3817 );
xor \U$3586 ( \3819 , \3814 , \3818 );
xor \U$3587 ( \3820 , \3805 , \3819 );
and \U$3588 ( \3821 , \3713 , \3717 );
and \U$3589 ( \3822 , \3717 , \3722 );
and \U$3590 ( \3823 , \3713 , \3722 );
or \U$3591 ( \3824 , \3821 , \3822 , \3823 );
or \U$3592 ( \3825 , \3770 , \3784 );
xor \U$3593 ( \3826 , \3824 , \3825 );
and \U$3594 ( \3827 , \700 , \1198 );
and \U$3595 ( \3828 , \653 , \1079 );
nor \U$3596 ( \3829 , \3827 , \3828 );
xnor \U$3597 ( \3830 , \3829 , \532 );
and \U$3598 ( \3831 , \728 , \497 );
and \U$3599 ( \3832 , \680 , \495 );
nor \U$3600 ( \3833 , \3831 , \3832 );
xnor \U$3601 ( \3834 , \3833 , \502 );
xor \U$3602 ( \3835 , \3830 , \3834 );
and \U$3604 ( \3836 , \708 , \505 );
nor \U$3605 ( \3837 , 1'b0 , \3836 );
not \U$3606 ( \3838 , \3837 );
xor \U$3607 ( \3839 , \3835 , \3838 );
and \U$3608 ( \3840 , \618 , \930 );
and \U$3609 ( \3841 , \1018 , \928 );
nor \U$3610 ( \3842 , \3840 , \3841 );
xnor \U$3611 ( \3843 , \3842 , \937 );
and \U$3612 ( \3844 , \643 , \950 );
and \U$3613 ( \3845 , \569 , \948 );
nor \U$3614 ( \3846 , \3844 , \3845 );
xnor \U$3615 ( \3847 , \3846 , \957 );
xor \U$3616 ( \3848 , \3843 , \3847 );
and \U$3617 ( \3849 , \673 , \978 );
and \U$3618 ( \3850 , \623 , \961 );
nor \U$3619 ( \3851 , \3849 , \3850 );
xnor \U$3620 ( \3852 , \3851 , \568 );
xor \U$3621 ( \3853 , \3848 , \3852 );
xor \U$3622 ( \3854 , \3839 , \3853 );
not \U$3623 ( \3855 , \852 );
and \U$3624 ( \3856 , \504 , \872 );
and \U$3625 ( \3857 , \223 , \870 );
nor \U$3626 ( \3858 , \3856 , \3857 );
xnor \U$3627 ( \3859 , \3858 , \879 );
xor \U$3628 ( \3860 , \3855 , \3859 );
and \U$3629 ( \3861 , \1020 , \900 );
and \U$3630 ( \3862 , \539 , \898 );
nor \U$3631 ( \3863 , \3861 , \3862 );
xnor \U$3632 ( \3864 , \3863 , \907 );
xor \U$3633 ( \3865 , \3860 , \3864 );
xor \U$3634 ( \3866 , \3854 , \3865 );
xor \U$3635 ( \3867 , \3826 , \3866 );
xor \U$3636 ( \3868 , \3820 , \3867 );
xor \U$3637 ( \3869 , \3801 , \3868 );
xor \U$3638 ( \3870 , \3795 , \3869 );
and \U$3639 ( \3871 , \3705 , \3787 );
nor \U$3640 ( \3872 , \3870 , \3871 );
and \U$3641 ( \3873 , \3799 , \3800 );
and \U$3642 ( \3874 , \3800 , \3868 );
and \U$3643 ( \3875 , \3799 , \3868 );
or \U$3644 ( \3876 , \3873 , \3874 , \3875 );
and \U$3645 ( \3877 , \3805 , \3819 );
and \U$3646 ( \3878 , \3819 , \3867 );
and \U$3647 ( \3879 , \3805 , \3867 );
or \U$3648 ( \3880 , \3877 , \3878 , \3879 );
xor \U$3649 ( \3881 , \3876 , \3880 );
and \U$3650 ( \3882 , \3824 , \3825 );
and \U$3651 ( \3883 , \3825 , \3866 );
and \U$3652 ( \3884 , \3824 , \3866 );
or \U$3653 ( \3885 , \3882 , \3883 , \3884 );
and \U$3654 ( \3886 , \3855 , \3859 );
and \U$3655 ( \3887 , \3859 , \3864 );
and \U$3656 ( \3888 , \3855 , \3864 );
or \U$3657 ( \3889 , \3886 , \3887 , \3888 );
and \U$3658 ( \3890 , \3843 , \3847 );
and \U$3659 ( \3891 , \3847 , \3852 );
and \U$3660 ( \3892 , \3843 , \3852 );
or \U$3661 ( \3893 , \3890 , \3891 , \3892 );
xor \U$3662 ( \3894 , \3889 , \3893 );
and \U$3663 ( \3895 , \3830 , \3834 );
and \U$3664 ( \3896 , \3834 , \3838 );
and \U$3665 ( \3897 , \3830 , \3838 );
or \U$3666 ( \3898 , \3895 , \3896 , \3897 );
xor \U$3667 ( \3899 , \3894 , \3898 );
xor \U$3668 ( \3900 , \3885 , \3899 );
and \U$3669 ( \3901 , \3809 , \3813 );
and \U$3670 ( \3902 , \3813 , \3818 );
and \U$3671 ( \3903 , \3809 , \3818 );
or \U$3672 ( \3904 , \3901 , \3902 , \3903 );
and \U$3673 ( \3905 , \3839 , \3853 );
and \U$3674 ( \3906 , \3853 , \3865 );
and \U$3675 ( \3907 , \3839 , \3865 );
or \U$3676 ( \3908 , \3905 , \3906 , \3907 );
xor \U$3677 ( \3909 , \3904 , \3908 );
and \U$3678 ( \3910 , \680 , \497 );
and \U$3679 ( \3911 , \700 , \495 );
nor \U$3680 ( \3912 , \3910 , \3911 );
xnor \U$3681 ( \3913 , \3912 , \502 );
and \U$3683 ( \3914 , \728 , \505 );
nor \U$3684 ( \3915 , 1'b0 , \3914 );
not \U$3685 ( \3916 , \3915 );
xnor \U$3686 ( \3917 , \3913 , \3916 );
and \U$3687 ( \3918 , \569 , \950 );
and \U$3688 ( \3919 , \618 , \948 );
nor \U$3689 ( \3920 , \3918 , \3919 );
xnor \U$3690 ( \3921 , \3920 , \957 );
and \U$3691 ( \3922 , \623 , \978 );
and \U$3692 ( \3923 , \643 , \961 );
nor \U$3693 ( \3924 , \3922 , \3923 );
xnor \U$3694 ( \3925 , \3924 , \568 );
xor \U$3695 ( \3926 , \3921 , \3925 );
and \U$3696 ( \3927 , \653 , \1198 );
and \U$3697 ( \3928 , \673 , \1079 );
nor \U$3698 ( \3929 , \3927 , \3928 );
xnor \U$3699 ( \3930 , \3929 , \532 );
xor \U$3700 ( \3931 , \3926 , \3930 );
xor \U$3701 ( \3932 , \3917 , \3931 );
and \U$3702 ( \3933 , \223 , \872 );
not \U$3703 ( \3934 , \3933 );
xnor \U$3704 ( \3935 , \3934 , \879 );
and \U$3705 ( \3936 , \539 , \900 );
and \U$3706 ( \3937 , \504 , \898 );
nor \U$3707 ( \3938 , \3936 , \3937 );
xnor \U$3708 ( \3939 , \3938 , \907 );
xor \U$3709 ( \3940 , \3935 , \3939 );
and \U$3710 ( \3941 , \1018 , \930 );
and \U$3711 ( \3942 , \1020 , \928 );
nor \U$3712 ( \3943 , \3941 , \3942 );
xnor \U$3713 ( \3944 , \3943 , \937 );
xor \U$3714 ( \3945 , \3940 , \3944 );
xor \U$3715 ( \3946 , \3932 , \3945 );
xor \U$3716 ( \3947 , \3909 , \3946 );
xor \U$3717 ( \3948 , \3900 , \3947 );
xor \U$3718 ( \3949 , \3881 , \3948 );
and \U$3719 ( \3950 , \3795 , \3869 );
nor \U$3720 ( \3951 , \3949 , \3950 );
nor \U$3721 ( \3952 , \3872 , \3951 );
nand \U$3722 ( \3953 , \3791 , \3952 );
and \U$3723 ( \3954 , \3885 , \3899 );
and \U$3724 ( \3955 , \3899 , \3947 );
and \U$3725 ( \3956 , \3885 , \3947 );
or \U$3726 ( \3957 , \3954 , \3955 , \3956 );
and \U$3727 ( \3958 , \3904 , \3908 );
and \U$3728 ( \3959 , \3908 , \3946 );
and \U$3729 ( \3960 , \3904 , \3946 );
or \U$3730 ( \3961 , \3958 , \3959 , \3960 );
and \U$3731 ( \3962 , \3935 , \3939 );
and \U$3732 ( \3963 , \3939 , \3944 );
and \U$3733 ( \3964 , \3935 , \3944 );
or \U$3734 ( \3965 , \3962 , \3963 , \3964 );
and \U$3735 ( \3966 , \3921 , \3925 );
and \U$3736 ( \3967 , \3925 , \3930 );
and \U$3737 ( \3968 , \3921 , \3930 );
or \U$3738 ( \3969 , \3966 , \3967 , \3968 );
xor \U$3739 ( \3970 , \3965 , \3969 );
or \U$3740 ( \3971 , \3913 , \3916 );
xor \U$3741 ( \3972 , \3970 , \3971 );
xor \U$3742 ( \3973 , \3961 , \3972 );
and \U$3743 ( \3974 , \3889 , \3893 );
and \U$3744 ( \3975 , \3893 , \3898 );
and \U$3745 ( \3976 , \3889 , \3898 );
or \U$3746 ( \3977 , \3974 , \3975 , \3976 );
and \U$3747 ( \3978 , \3917 , \3931 );
and \U$3748 ( \3979 , \3931 , \3945 );
and \U$3749 ( \3980 , \3917 , \3945 );
or \U$3750 ( \3981 , \3978 , \3979 , \3980 );
xor \U$3751 ( \3982 , \3977 , \3981 );
and \U$3752 ( \3983 , \700 , \497 );
and \U$3753 ( \3984 , \653 , \495 );
nor \U$3754 ( \3985 , \3983 , \3984 );
xnor \U$3755 ( \3986 , \3985 , \502 );
and \U$3757 ( \3987 , \680 , \505 );
nor \U$3758 ( \3988 , 1'b0 , \3987 );
not \U$3759 ( \3989 , \3988 );
xor \U$3760 ( \3990 , \3986 , \3989 );
and \U$3761 ( \3991 , \618 , \950 );
and \U$3762 ( \3992 , \1018 , \948 );
nor \U$3763 ( \3993 , \3991 , \3992 );
xnor \U$3764 ( \3994 , \3993 , \957 );
and \U$3765 ( \3995 , \643 , \978 );
and \U$3766 ( \3996 , \569 , \961 );
nor \U$3767 ( \3997 , \3995 , \3996 );
xnor \U$3768 ( \3998 , \3997 , \568 );
xor \U$3769 ( \3999 , \3994 , \3998 );
and \U$3770 ( \4000 , \673 , \1198 );
and \U$3771 ( \4001 , \623 , \1079 );
nor \U$3772 ( \4002 , \4000 , \4001 );
xnor \U$3773 ( \4003 , \4002 , \532 );
xor \U$3774 ( \4004 , \3999 , \4003 );
xor \U$3775 ( \4005 , \3990 , \4004 );
not \U$3776 ( \4006 , \879 );
and \U$3777 ( \4007 , \504 , \900 );
and \U$3778 ( \4008 , \223 , \898 );
nor \U$3779 ( \4009 , \4007 , \4008 );
xnor \U$3780 ( \4010 , \4009 , \907 );
xor \U$3781 ( \4011 , \4006 , \4010 );
and \U$3782 ( \4012 , \1020 , \930 );
and \U$3783 ( \4013 , \539 , \928 );
nor \U$3784 ( \4014 , \4012 , \4013 );
xnor \U$3785 ( \4015 , \4014 , \937 );
xor \U$3786 ( \4016 , \4011 , \4015 );
xor \U$3787 ( \4017 , \4005 , \4016 );
xor \U$3788 ( \4018 , \3982 , \4017 );
xor \U$3789 ( \4019 , \3973 , \4018 );
xor \U$3790 ( \4020 , \3957 , \4019 );
and \U$3791 ( \4021 , \3876 , \3880 );
and \U$3792 ( \4022 , \3880 , \3948 );
and \U$3793 ( \4023 , \3876 , \3948 );
or \U$3794 ( \4024 , \4021 , \4022 , \4023 );
nor \U$3795 ( \4025 , \4020 , \4024 );
and \U$3796 ( \4026 , \3961 , \3972 );
and \U$3797 ( \4027 , \3972 , \4018 );
and \U$3798 ( \4028 , \3961 , \4018 );
or \U$3799 ( \4029 , \4026 , \4027 , \4028 );
and \U$3800 ( \4030 , \3977 , \3981 );
and \U$3801 ( \4031 , \3981 , \4017 );
and \U$3802 ( \4032 , \3977 , \4017 );
or \U$3803 ( \4033 , \4030 , \4031 , \4032 );
and \U$3804 ( \4034 , \4006 , \4010 );
and \U$3805 ( \4035 , \4010 , \4015 );
and \U$3806 ( \4036 , \4006 , \4015 );
or \U$3807 ( \4037 , \4034 , \4035 , \4036 );
and \U$3808 ( \4038 , \3994 , \3998 );
and \U$3809 ( \4039 , \3998 , \4003 );
and \U$3810 ( \4040 , \3994 , \4003 );
or \U$3811 ( \4041 , \4038 , \4039 , \4040 );
xor \U$3812 ( \4042 , \4037 , \4041 );
and \U$3813 ( \4043 , \3986 , \3989 );
xor \U$3814 ( \4044 , \4042 , \4043 );
xor \U$3815 ( \4045 , \4033 , \4044 );
and \U$3816 ( \4046 , \3965 , \3969 );
and \U$3817 ( \4047 , \3969 , \3971 );
and \U$3818 ( \4048 , \3965 , \3971 );
or \U$3819 ( \4049 , \4046 , \4047 , \4048 );
and \U$3820 ( \4050 , \3990 , \4004 );
and \U$3821 ( \4051 , \4004 , \4016 );
and \U$3822 ( \4052 , \3990 , \4016 );
or \U$3823 ( \4053 , \4050 , \4051 , \4052 );
xor \U$3824 ( \4054 , \4049 , \4053 );
and \U$3826 ( \4055 , \700 , \505 );
nor \U$3827 ( \4056 , 1'b0 , \4055 );
and \U$3828 ( \4057 , \569 , \978 );
and \U$3829 ( \4058 , \618 , \961 );
nor \U$3830 ( \4059 , \4057 , \4058 );
xnor \U$3831 ( \4060 , \4059 , \568 );
and \U$3832 ( \4061 , \623 , \1198 );
and \U$3833 ( \4062 , \643 , \1079 );
nor \U$3834 ( \4063 , \4061 , \4062 );
xnor \U$3835 ( \4064 , \4063 , \532 );
xor \U$3836 ( \4065 , \4060 , \4064 );
and \U$3837 ( \4066 , \653 , \497 );
and \U$3838 ( \4067 , \673 , \495 );
nor \U$3839 ( \4068 , \4066 , \4067 );
xnor \U$3840 ( \4069 , \4068 , \502 );
xor \U$3841 ( \4070 , \4065 , \4069 );
xor \U$3842 ( \4071 , \4056 , \4070 );
and \U$3843 ( \4072 , \223 , \900 );
not \U$3844 ( \4073 , \4072 );
xnor \U$3845 ( \4074 , \4073 , \907 );
and \U$3846 ( \4075 , \539 , \930 );
and \U$3847 ( \4076 , \504 , \928 );
nor \U$3848 ( \4077 , \4075 , \4076 );
xnor \U$3849 ( \4078 , \4077 , \937 );
xor \U$3850 ( \4079 , \4074 , \4078 );
and \U$3851 ( \4080 , \1018 , \950 );
and \U$3852 ( \4081 , \1020 , \948 );
nor \U$3853 ( \4082 , \4080 , \4081 );
xnor \U$3854 ( \4083 , \4082 , \957 );
xor \U$3855 ( \4084 , \4079 , \4083 );
xor \U$3856 ( \4085 , \4071 , \4084 );
xor \U$3857 ( \4086 , \4054 , \4085 );
xor \U$3858 ( \4087 , \4045 , \4086 );
xor \U$3859 ( \4088 , \4029 , \4087 );
and \U$3860 ( \4089 , \3957 , \4019 );
nor \U$3861 ( \4090 , \4088 , \4089 );
nor \U$3862 ( \4091 , \4025 , \4090 );
and \U$3863 ( \4092 , \4033 , \4044 );
and \U$3864 ( \4093 , \4044 , \4086 );
and \U$3865 ( \4094 , \4033 , \4086 );
or \U$3866 ( \4095 , \4092 , \4093 , \4094 );
and \U$3867 ( \4096 , \4049 , \4053 );
and \U$3868 ( \4097 , \4053 , \4085 );
and \U$3869 ( \4098 , \4049 , \4085 );
or \U$3870 ( \4099 , \4096 , \4097 , \4098 );
and \U$3871 ( \4100 , \4074 , \4078 );
and \U$3872 ( \4101 , \4078 , \4083 );
and \U$3873 ( \4102 , \4074 , \4083 );
or \U$3874 ( \4103 , \4100 , \4101 , \4102 );
and \U$3875 ( \4104 , \4060 , \4064 );
and \U$3876 ( \4105 , \4064 , \4069 );
and \U$3877 ( \4106 , \4060 , \4069 );
or \U$3878 ( \4107 , \4104 , \4105 , \4106 );
xor \U$3879 ( \4108 , \4103 , \4107 );
not \U$3880 ( \4109 , \4056 );
xor \U$3881 ( \4110 , \4108 , \4109 );
xor \U$3882 ( \4111 , \4099 , \4110 );
and \U$3883 ( \4112 , \4037 , \4041 );
and \U$3884 ( \4113 , \4041 , \4043 );
and \U$3885 ( \4114 , \4037 , \4043 );
or \U$3886 ( \4115 , \4112 , \4113 , \4114 );
and \U$3887 ( \4116 , \4056 , \4070 );
and \U$3888 ( \4117 , \4070 , \4084 );
and \U$3889 ( \4118 , \4056 , \4084 );
or \U$3890 ( \4119 , \4116 , \4117 , \4118 );
xor \U$3891 ( \4120 , \4115 , \4119 );
and \U$3893 ( \4121 , \653 , \505 );
nor \U$3894 ( \4122 , 1'b0 , \4121 );
not \U$3895 ( \4123 , \4122 );
and \U$3896 ( \4124 , \618 , \978 );
and \U$3897 ( \4125 , \1018 , \961 );
nor \U$3898 ( \4126 , \4124 , \4125 );
xnor \U$3899 ( \4127 , \4126 , \568 );
and \U$3900 ( \4128 , \643 , \1198 );
and \U$3901 ( \4129 , \569 , \1079 );
nor \U$3902 ( \4130 , \4128 , \4129 );
xnor \U$3903 ( \4131 , \4130 , \532 );
xor \U$3904 ( \4132 , \4127 , \4131 );
and \U$3905 ( \4133 , \673 , \497 );
and \U$3906 ( \4134 , \623 , \495 );
nor \U$3907 ( \4135 , \4133 , \4134 );
xnor \U$3908 ( \4136 , \4135 , \502 );
xor \U$3909 ( \4137 , \4132 , \4136 );
xor \U$3910 ( \4138 , \4123 , \4137 );
not \U$3911 ( \4139 , \907 );
and \U$3912 ( \4140 , \504 , \930 );
and \U$3913 ( \4141 , \223 , \928 );
nor \U$3914 ( \4142 , \4140 , \4141 );
xnor \U$3915 ( \4143 , \4142 , \937 );
xor \U$3916 ( \4144 , \4139 , \4143 );
and \U$3917 ( \4145 , \1020 , \950 );
and \U$3918 ( \4146 , \539 , \948 );
nor \U$3919 ( \4147 , \4145 , \4146 );
xnor \U$3920 ( \4148 , \4147 , \957 );
xor \U$3921 ( \4149 , \4144 , \4148 );
xor \U$3922 ( \4150 , \4138 , \4149 );
xor \U$3923 ( \4151 , \4120 , \4150 );
xor \U$3924 ( \4152 , \4111 , \4151 );
xor \U$3925 ( \4153 , \4095 , \4152 );
and \U$3926 ( \4154 , \4029 , \4087 );
nor \U$3927 ( \4155 , \4153 , \4154 );
and \U$3928 ( \4156 , \4099 , \4110 );
and \U$3929 ( \4157 , \4110 , \4151 );
and \U$3930 ( \4158 , \4099 , \4151 );
or \U$3931 ( \4159 , \4156 , \4157 , \4158 );
and \U$3932 ( \4160 , \4115 , \4119 );
and \U$3933 ( \4161 , \4119 , \4150 );
and \U$3934 ( \4162 , \4115 , \4150 );
or \U$3935 ( \4163 , \4160 , \4161 , \4162 );
and \U$3936 ( \4164 , \223 , \930 );
not \U$3937 ( \4165 , \4164 );
xnor \U$3938 ( \4166 , \4165 , \937 );
and \U$3939 ( \4167 , \539 , \950 );
and \U$3940 ( \4168 , \504 , \948 );
nor \U$3941 ( \4169 , \4167 , \4168 );
xnor \U$3942 ( \4170 , \4169 , \957 );
xor \U$3943 ( \4171 , \4166 , \4170 );
and \U$3944 ( \4172 , \1018 , \978 );
and \U$3945 ( \4173 , \1020 , \961 );
nor \U$3946 ( \4174 , \4172 , \4173 );
xnor \U$3947 ( \4175 , \4174 , \568 );
xor \U$3948 ( \4176 , \4171 , \4175 );
and \U$3949 ( \4177 , \4139 , \4143 );
and \U$3950 ( \4178 , \4143 , \4148 );
and \U$3951 ( \4179 , \4139 , \4148 );
or \U$3952 ( \4180 , \4177 , \4178 , \4179 );
and \U$3953 ( \4181 , \4127 , \4131 );
and \U$3954 ( \4182 , \4131 , \4136 );
and \U$3955 ( \4183 , \4127 , \4136 );
or \U$3956 ( \4184 , \4181 , \4182 , \4183 );
xnor \U$3957 ( \4185 , \4180 , \4184 );
xor \U$3958 ( \4186 , \4176 , \4185 );
xor \U$3959 ( \4187 , \4163 , \4186 );
and \U$3960 ( \4188 , \4103 , \4107 );
and \U$3961 ( \4189 , \4107 , \4109 );
and \U$3962 ( \4190 , \4103 , \4109 );
or \U$3963 ( \4191 , \4188 , \4189 , \4190 );
and \U$3964 ( \4192 , \4123 , \4137 );
and \U$3965 ( \4193 , \4137 , \4149 );
and \U$3966 ( \4194 , \4123 , \4149 );
or \U$3967 ( \4195 , \4192 , \4193 , \4194 );
xor \U$3968 ( \4196 , \4191 , \4195 );
and \U$3969 ( \4197 , \569 , \1198 );
and \U$3970 ( \4198 , \618 , \1079 );
nor \U$3971 ( \4199 , \4197 , \4198 );
xnor \U$3972 ( \4200 , \4199 , \532 );
and \U$3973 ( \4201 , \623 , \497 );
and \U$3974 ( \4202 , \643 , \495 );
nor \U$3975 ( \4203 , \4201 , \4202 );
xnor \U$3976 ( \4204 , \4203 , \502 );
xor \U$3977 ( \4205 , \4200 , \4204 );
and \U$3979 ( \4206 , \673 , \505 );
nor \U$3980 ( \4207 , 1'b0 , \4206 );
not \U$3981 ( \4208 , \4207 );
xor \U$3982 ( \4209 , \4205 , \4208 );
xor \U$3983 ( \4210 , \4196 , \4209 );
xor \U$3984 ( \4211 , \4187 , \4210 );
xor \U$3985 ( \4212 , \4159 , \4211 );
and \U$3986 ( \4213 , \4095 , \4152 );
nor \U$3987 ( \4214 , \4212 , \4213 );
nor \U$3988 ( \4215 , \4155 , \4214 );
nand \U$3989 ( \4216 , \4091 , \4215 );
nor \U$3990 ( \4217 , \3953 , \4216 );
and \U$3991 ( \4218 , \4163 , \4186 );
and \U$3992 ( \4219 , \4186 , \4210 );
and \U$3993 ( \4220 , \4163 , \4210 );
or \U$3994 ( \4221 , \4218 , \4219 , \4220 );
and \U$3995 ( \4222 , \4191 , \4195 );
and \U$3996 ( \4223 , \4195 , \4209 );
and \U$3997 ( \4224 , \4191 , \4209 );
or \U$3998 ( \4225 , \4222 , \4223 , \4224 );
and \U$3999 ( \4226 , \4176 , \4185 );
xor \U$4000 ( \4227 , \4225 , \4226 );
or \U$4001 ( \4228 , \4180 , \4184 );
not \U$4002 ( \4229 , \937 );
and \U$4003 ( \4230 , \504 , \950 );
and \U$4004 ( \4231 , \223 , \948 );
nor \U$4005 ( \4232 , \4230 , \4231 );
xnor \U$4006 ( \4233 , \4232 , \957 );
xor \U$4007 ( \4234 , \4229 , \4233 );
and \U$4008 ( \4235 , \1020 , \978 );
and \U$4009 ( \4236 , \539 , \961 );
nor \U$4010 ( \4237 , \4235 , \4236 );
xnor \U$4011 ( \4238 , \4237 , \568 );
xor \U$4012 ( \4239 , \4234 , \4238 );
xor \U$4013 ( \4240 , \4228 , \4239 );
and \U$4014 ( \4241 , \4166 , \4170 );
and \U$4015 ( \4242 , \4170 , \4175 );
and \U$4016 ( \4243 , \4166 , \4175 );
or \U$4017 ( \4244 , \4241 , \4242 , \4243 );
and \U$4018 ( \4245 , \4200 , \4204 );
and \U$4019 ( \4246 , \4204 , \4208 );
and \U$4020 ( \4247 , \4200 , \4208 );
or \U$4021 ( \4248 , \4245 , \4246 , \4247 );
xor \U$4022 ( \4249 , \4244 , \4248 );
and \U$4023 ( \4250 , \618 , \1198 );
and \U$4024 ( \4251 , \1018 , \1079 );
nor \U$4025 ( \4252 , \4250 , \4251 );
xnor \U$4026 ( \4253 , \4252 , \532 );
and \U$4027 ( \4254 , \643 , \497 );
and \U$4028 ( \4255 , \569 , \495 );
nor \U$4029 ( \4256 , \4254 , \4255 );
xnor \U$4030 ( \4257 , \4256 , \502 );
xor \U$4031 ( \4258 , \4253 , \4257 );
and \U$4033 ( \4259 , \623 , \505 );
nor \U$4034 ( \4260 , 1'b0 , \4259 );
not \U$4035 ( \4261 , \4260 );
xor \U$4036 ( \4262 , \4258 , \4261 );
xor \U$4037 ( \4263 , \4249 , \4262 );
xor \U$4038 ( \4264 , \4240 , \4263 );
xor \U$4039 ( \4265 , \4227 , \4264 );
xor \U$4040 ( \4266 , \4221 , \4265 );
and \U$4041 ( \4267 , \4159 , \4211 );
nor \U$4042 ( \4268 , \4266 , \4267 );
and \U$4043 ( \4269 , \4225 , \4226 );
and \U$4044 ( \4270 , \4226 , \4264 );
and \U$4045 ( \4271 , \4225 , \4264 );
or \U$4046 ( \4272 , \4269 , \4270 , \4271 );
and \U$4047 ( \4273 , \4228 , \4239 );
and \U$4048 ( \4274 , \4239 , \4263 );
and \U$4049 ( \4275 , \4228 , \4263 );
or \U$4050 ( \4276 , \4273 , \4274 , \4275 );
xor \U$4051 ( \4277 , \4272 , \4276 );
and \U$4052 ( \4278 , \4244 , \4248 );
and \U$4053 ( \4279 , \4248 , \4262 );
and \U$4054 ( \4280 , \4244 , \4262 );
or \U$4055 ( \4281 , \4278 , \4279 , \4280 );
and \U$4056 ( \4282 , \223 , \950 );
not \U$4057 ( \4283 , \4282 );
xnor \U$4058 ( \4284 , \4283 , \957 );
and \U$4059 ( \4285 , \539 , \978 );
and \U$4060 ( \4286 , \504 , \961 );
nor \U$4061 ( \4287 , \4285 , \4286 );
xnor \U$4062 ( \4288 , \4287 , \568 );
xor \U$4063 ( \4289 , \4284 , \4288 );
and \U$4064 ( \4290 , \1018 , \1198 );
and \U$4065 ( \4291 , \1020 , \1079 );
nor \U$4066 ( \4292 , \4290 , \4291 );
xnor \U$4067 ( \4293 , \4292 , \532 );
xor \U$4068 ( \4294 , \4289 , \4293 );
xor \U$4069 ( \4295 , \4281 , \4294 );
and \U$4070 ( \4296 , \4229 , \4233 );
and \U$4071 ( \4297 , \4233 , \4238 );
and \U$4072 ( \4298 , \4229 , \4238 );
or \U$4073 ( \4299 , \4296 , \4297 , \4298 );
and \U$4074 ( \4300 , \4253 , \4257 );
and \U$4075 ( \4301 , \4257 , \4261 );
and \U$4076 ( \4302 , \4253 , \4261 );
or \U$4077 ( \4303 , \4300 , \4301 , \4302 );
xor \U$4078 ( \4304 , \4299 , \4303 );
and \U$4079 ( \4305 , \569 , \497 );
and \U$4080 ( \4306 , \618 , \495 );
nor \U$4081 ( \4307 , \4305 , \4306 );
xnor \U$4082 ( \4308 , \4307 , \502 );
and \U$4084 ( \4309 , \643 , \505 );
nor \U$4085 ( \4310 , 1'b0 , \4309 );
not \U$4086 ( \4311 , \4310 );
xnor \U$4087 ( \4312 , \4308 , \4311 );
xor \U$4088 ( \4313 , \4304 , \4312 );
xor \U$4089 ( \4314 , \4295 , \4313 );
xor \U$4090 ( \4315 , \4277 , \4314 );
and \U$4091 ( \4316 , \4221 , \4265 );
nor \U$4092 ( \4317 , \4315 , \4316 );
nor \U$4093 ( \4318 , \4268 , \4317 );
and \U$4094 ( \4319 , \4281 , \4294 );
and \U$4095 ( \4320 , \4294 , \4313 );
and \U$4096 ( \4321 , \4281 , \4313 );
or \U$4097 ( \4322 , \4319 , \4320 , \4321 );
and \U$4098 ( \4323 , \4299 , \4303 );
and \U$4099 ( \4324 , \4303 , \4312 );
and \U$4100 ( \4325 , \4299 , \4312 );
or \U$4101 ( \4326 , \4323 , \4324 , \4325 );
and \U$4103 ( \4327 , \569 , \505 );
nor \U$4104 ( \4328 , 1'b0 , \4327 );
not \U$4105 ( \4329 , \4328 );
not \U$4106 ( \4330 , \957 );
and \U$4107 ( \4331 , \504 , \978 );
and \U$4108 ( \4332 , \223 , \961 );
nor \U$4109 ( \4333 , \4331 , \4332 );
xnor \U$4110 ( \4334 , \4333 , \568 );
xor \U$4111 ( \4335 , \4330 , \4334 );
and \U$4112 ( \4336 , \1020 , \1198 );
and \U$4113 ( \4337 , \539 , \1079 );
nor \U$4114 ( \4338 , \4336 , \4337 );
xnor \U$4115 ( \4339 , \4338 , \532 );
xor \U$4116 ( \4340 , \4335 , \4339 );
xor \U$4117 ( \4341 , \4329 , \4340 );
xor \U$4118 ( \4342 , \4326 , \4341 );
and \U$4119 ( \4343 , \4284 , \4288 );
and \U$4120 ( \4344 , \4288 , \4293 );
and \U$4121 ( \4345 , \4284 , \4293 );
or \U$4122 ( \4346 , \4343 , \4344 , \4345 );
or \U$4123 ( \4347 , \4308 , \4311 );
xor \U$4124 ( \4348 , \4346 , \4347 );
and \U$4125 ( \4349 , \618 , \497 );
and \U$4126 ( \4350 , \1018 , \495 );
nor \U$4127 ( \4351 , \4349 , \4350 );
xnor \U$4128 ( \4352 , \4351 , \502 );
xor \U$4129 ( \4353 , \4348 , \4352 );
xor \U$4130 ( \4354 , \4342 , \4353 );
xor \U$4131 ( \4355 , \4322 , \4354 );
and \U$4132 ( \4356 , \4272 , \4276 );
and \U$4133 ( \4357 , \4276 , \4314 );
and \U$4134 ( \4358 , \4272 , \4314 );
or \U$4135 ( \4359 , \4356 , \4357 , \4358 );
nor \U$4136 ( \4360 , \4355 , \4359 );
and \U$4137 ( \4361 , \4326 , \4341 );
and \U$4138 ( \4362 , \4341 , \4353 );
and \U$4139 ( \4363 , \4326 , \4353 );
or \U$4140 ( \4364 , \4361 , \4362 , \4363 );
and \U$4141 ( \4365 , \4346 , \4347 );
and \U$4142 ( \4366 , \4347 , \4352 );
and \U$4143 ( \4367 , \4346 , \4352 );
or \U$4144 ( \4368 , \4365 , \4366 , \4367 );
and \U$4145 ( \4369 , \4329 , \4340 );
xor \U$4146 ( \4370 , \4368 , \4369 );
and \U$4147 ( \4371 , \4330 , \4334 );
and \U$4148 ( \4372 , \4334 , \4339 );
and \U$4149 ( \4373 , \4330 , \4339 );
or \U$4150 ( \4374 , \4371 , \4372 , \4373 );
and \U$4152 ( \4375 , \618 , \505 );
nor \U$4153 ( \4376 , 1'b0 , \4375 );
xor \U$4154 ( \4377 , \4374 , \4376 );
and \U$4155 ( \4378 , \223 , \978 );
not \U$4156 ( \4379 , \4378 );
xnor \U$4157 ( \4380 , \4379 , \568 );
and \U$4158 ( \4381 , \539 , \1198 );
and \U$4159 ( \4382 , \504 , \1079 );
nor \U$4160 ( \4383 , \4381 , \4382 );
xnor \U$4161 ( \4384 , \4383 , \532 );
xor \U$4162 ( \4385 , \4380 , \4384 );
and \U$4163 ( \4386 , \1018 , \497 );
and \U$4164 ( \4387 , \1020 , \495 );
nor \U$4165 ( \4388 , \4386 , \4387 );
xnor \U$4166 ( \4389 , \4388 , \502 );
xor \U$4167 ( \4390 , \4385 , \4389 );
xor \U$4168 ( \4391 , \4377 , \4390 );
xor \U$4169 ( \4392 , \4370 , \4391 );
xor \U$4170 ( \4393 , \4364 , \4392 );
and \U$4171 ( \4394 , \4322 , \4354 );
nor \U$4172 ( \4395 , \4393 , \4394 );
nor \U$4173 ( \4396 , \4360 , \4395 );
nand \U$4174 ( \4397 , \4318 , \4396 );
and \U$4175 ( \4398 , \4368 , \4369 );
and \U$4176 ( \4399 , \4369 , \4391 );
and \U$4177 ( \4400 , \4368 , \4391 );
or \U$4178 ( \4401 , \4398 , \4399 , \4400 );
and \U$4179 ( \4402 , \4374 , \4376 );
and \U$4180 ( \4403 , \4376 , \4390 );
and \U$4181 ( \4404 , \4374 , \4390 );
or \U$4182 ( \4405 , \4402 , \4403 , \4404 );
not \U$4183 ( \4406 , \568 );
and \U$4184 ( \4407 , \504 , \1198 );
and \U$4185 ( \4408 , \223 , \1079 );
nor \U$4186 ( \4409 , \4407 , \4408 );
xnor \U$4187 ( \4410 , \4409 , \532 );
xor \U$4188 ( \4411 , \4406 , \4410 );
and \U$4189 ( \4412 , \1020 , \497 );
and \U$4190 ( \4413 , \539 , \495 );
nor \U$4191 ( \4414 , \4412 , \4413 );
xnor \U$4192 ( \4415 , \4414 , \502 );
xor \U$4193 ( \4416 , \4411 , \4415 );
xor \U$4194 ( \4417 , \4405 , \4416 );
and \U$4195 ( \4418 , \4380 , \4384 );
and \U$4196 ( \4419 , \4384 , \4389 );
and \U$4197 ( \4420 , \4380 , \4389 );
or \U$4198 ( \4421 , \4418 , \4419 , \4420 );
not \U$4199 ( \4422 , \4376 );
xor \U$4200 ( \4423 , \4421 , \4422 );
and \U$4202 ( \4424 , \1018 , \505 );
nor \U$4203 ( \4425 , 1'b0 , \4424 );
not \U$4204 ( \4426 , \4425 );
xor \U$4205 ( \4427 , \4423 , \4426 );
xor \U$4206 ( \4428 , \4417 , \4427 );
xor \U$4207 ( \4429 , \4401 , \4428 );
and \U$4208 ( \4430 , \4364 , \4392 );
nor \U$4209 ( \4431 , \4429 , \4430 );
and \U$4210 ( \4432 , \4405 , \4416 );
and \U$4211 ( \4433 , \4416 , \4427 );
and \U$4212 ( \4434 , \4405 , \4427 );
or \U$4213 ( \4435 , \4432 , \4433 , \4434 );
and \U$4214 ( \4436 , \4421 , \4422 );
and \U$4215 ( \4437 , \4422 , \4426 );
and \U$4216 ( \4438 , \4421 , \4426 );
or \U$4217 ( \4439 , \4436 , \4437 , \4438 );
xor \U$4218 ( \4440 , \4435 , \4439 );
and \U$4219 ( \4441 , \4406 , \4410 );
and \U$4220 ( \4442 , \4410 , \4415 );
and \U$4221 ( \4443 , \4406 , \4415 );
or \U$4222 ( \4444 , \4441 , \4442 , \4443 );
and \U$4223 ( \4445 , \223 , \1198 );
not \U$4224 ( \4446 , \4445 );
xnor \U$4225 ( \4447 , \4446 , \532 );
and \U$4226 ( \4448 , \539 , \497 );
and \U$4227 ( \4449 , \504 , \495 );
nor \U$4228 ( \4450 , \4448 , \4449 );
xnor \U$4229 ( \4451 , \4450 , \502 );
xor \U$4230 ( \4452 , \4447 , \4451 );
and \U$4232 ( \4453 , \1020 , \505 );
nor \U$4233 ( \4454 , 1'b0 , \4453 );
not \U$4234 ( \4455 , \4454 );
xor \U$4235 ( \4456 , \4452 , \4455 );
xnor \U$4236 ( \4457 , \4444 , \4456 );
xor \U$4237 ( \4458 , \4440 , \4457 );
and \U$4238 ( \4459 , \4401 , \4428 );
nor \U$4239 ( \4460 , \4458 , \4459 );
nor \U$4240 ( \4461 , \4431 , \4460 );
or \U$4241 ( \4462 , \4444 , \4456 );
and \U$4242 ( \4463 , \4447 , \4451 );
and \U$4243 ( \4464 , \4451 , \4455 );
and \U$4244 ( \4465 , \4447 , \4455 );
or \U$4245 ( \4466 , \4463 , \4464 , \4465 );
xor \U$4246 ( \4467 , \4462 , \4466 );
xor \U$4247 ( \4468 , \533 , \537 );
xor \U$4248 ( \4469 , \4468 , \542 );
xor \U$4249 ( \4470 , \4467 , \4469 );
and \U$4250 ( \4471 , \4435 , \4439 );
and \U$4251 ( \4472 , \4439 , \4457 );
and \U$4252 ( \4473 , \4435 , \4457 );
or \U$4253 ( \4474 , \4471 , \4472 , \4473 );
nor \U$4254 ( \4475 , \4470 , \4474 );
xor \U$4255 ( \4476 , \545 , \546 );
and \U$4256 ( \4477 , \4462 , \4466 );
and \U$4257 ( \4478 , \4466 , \4469 );
and \U$4258 ( \4479 , \4462 , \4469 );
or \U$4259 ( \4480 , \4477 , \4478 , \4479 );
nor \U$4260 ( \4481 , \4476 , \4480 );
nor \U$4261 ( \4482 , \4475 , \4481 );
nand \U$4262 ( \4483 , \4461 , \4482 );
nor \U$4263 ( \4484 , \4397 , \4483 );
nand \U$4264 ( \4485 , \4217 , \4484 );
nor \U$4265 ( \4486 , \3610 , \4485 );
and \U$4266 ( \4487 , \794 , \616 );
and \U$4267 ( \4488 , \814 , \613 );
nor \U$4268 ( \4489 , \4487 , \4488 );
xnor \U$4269 ( \4490 , \4489 , \576 );
and \U$4270 ( \4491 , \791 , \4490 );
and \U$4271 ( \4492 , \827 , \641 );
and \U$4272 ( \4493 , \847 , \639 );
nor \U$4273 ( \4494 , \4492 , \4493 );
xnor \U$4274 ( \4495 , \4494 , \648 );
and \U$4275 ( \4496 , \4490 , \4495 );
and \U$4276 ( \4497 , \791 , \4495 );
or \U$4277 ( \4498 , \4491 , \4496 , \4497 );
and \U$4278 ( \4499 , \854 , \671 );
and \U$4279 ( \4500 , \874 , \669 );
nor \U$4280 ( \4501 , \4499 , \4500 );
xnor \U$4281 ( \4502 , \4501 , \678 );
and \U$4282 ( \4503 , \882 , \698 );
and \U$4283 ( \4504 , \902 , \696 );
nor \U$4284 ( \4505 , \4503 , \4504 );
xnor \U$4285 ( \4506 , \4505 , \705 );
and \U$4286 ( \4507 , \4502 , \4506 );
and \U$4287 ( \4508 , \912 , \726 );
and \U$4288 ( \4509 , \932 , \724 );
nor \U$4289 ( \4510 , \4508 , \4509 );
xnor \U$4290 ( \4511 , \4510 , \733 );
and \U$4291 ( \4512 , \4506 , \4511 );
and \U$4292 ( \4513 , \4502 , \4511 );
or \U$4293 ( \4514 , \4507 , \4512 , \4513 );
and \U$4294 ( \4515 , \4498 , \4514 );
and \U$4295 ( \4516 , \960 , \784 );
and \U$4296 ( \4517 , \939 , \782 );
nor \U$4297 ( \4518 , \4516 , \4517 );
xnor \U$4298 ( \4519 , \4518 , \791 );
and \U$4299 ( \4520 , \4514 , \4519 );
and \U$4300 ( \4521 , \4498 , \4519 );
or \U$4301 ( \4522 , \4515 , \4520 , \4521 );
and \U$4302 ( \4523 , \827 , \671 );
and \U$4303 ( \4524 , \847 , \669 );
nor \U$4304 ( \4525 , \4523 , \4524 );
xnor \U$4305 ( \4526 , \4525 , \678 );
and \U$4306 ( \4527 , \854 , \698 );
and \U$4307 ( \4528 , \874 , \696 );
nor \U$4308 ( \4529 , \4527 , \4528 );
xnor \U$4309 ( \4530 , \4529 , \705 );
xor \U$4310 ( \4531 , \4526 , \4530 );
and \U$4311 ( \4532 , \882 , \726 );
and \U$4312 ( \4533 , \902 , \724 );
nor \U$4313 ( \4534 , \4532 , \4533 );
xnor \U$4314 ( \4535 , \4534 , \733 );
xor \U$4315 ( \4536 , \4531 , \4535 );
and \U$4316 ( \4537 , \766 , \616 );
and \U$4317 ( \4538 , \786 , \613 );
nor \U$4318 ( \4539 , \4537 , \4538 );
xnor \U$4319 ( \4540 , \4539 , \576 );
xor \U$4320 ( \4541 , \819 , \4540 );
and \U$4321 ( \4542 , \794 , \641 );
and \U$4322 ( \4543 , \814 , \639 );
nor \U$4323 ( \4544 , \4542 , \4543 );
xnor \U$4324 ( \4545 , \4544 , \648 );
xor \U$4325 ( \4546 , \4541 , \4545 );
xor \U$4326 ( \4547 , \4536 , \4546 );
and \U$4327 ( \4548 , \4522 , \4547 );
and \U$4328 ( \4549 , \814 , \616 );
and \U$4329 ( \4550 , \766 , \613 );
nor \U$4330 ( \4551 , \4549 , \4550 );
xnor \U$4331 ( \4552 , \4551 , \576 );
and \U$4332 ( \4553 , \847 , \641 );
and \U$4333 ( \4554 , \794 , \639 );
nor \U$4334 ( \4555 , \4553 , \4554 );
xnor \U$4335 ( \4556 , \4555 , \648 );
and \U$4336 ( \4557 , \4552 , \4556 );
and \U$4337 ( \4558 , \874 , \671 );
and \U$4338 ( \4559 , \827 , \669 );
nor \U$4339 ( \4560 , \4558 , \4559 );
xnor \U$4340 ( \4561 , \4560 , \678 );
and \U$4341 ( \4562 , \4556 , \4561 );
and \U$4342 ( \4563 , \4552 , \4561 );
or \U$4343 ( \4564 , \4557 , \4562 , \4563 );
and \U$4344 ( \4565 , \902 , \698 );
and \U$4345 ( \4566 , \854 , \696 );
nor \U$4346 ( \4567 , \4565 , \4566 );
xnor \U$4347 ( \4568 , \4567 , \705 );
and \U$4348 ( \4569 , \932 , \726 );
and \U$4349 ( \4570 , \882 , \724 );
nor \U$4350 ( \4571 , \4569 , \4570 );
xnor \U$4351 ( \4572 , \4571 , \733 );
and \U$4352 ( \4573 , \4568 , \4572 );
and \U$4353 ( \4574 , \952 , \757 );
and \U$4354 ( \4575 , \912 , \755 );
nor \U$4355 ( \4576 , \4574 , \4575 );
xnor \U$4356 ( \4577 , \4576 , \764 );
and \U$4357 ( \4578 , \4572 , \4577 );
and \U$4358 ( \4579 , \4568 , \4577 );
or \U$4359 ( \4580 , \4573 , \4578 , \4579 );
xor \U$4360 ( \4581 , \4564 , \4580 );
and \U$4361 ( \4582 , \912 , \757 );
and \U$4362 ( \4583 , \932 , \755 );
nor \U$4363 ( \4584 , \4582 , \4583 );
xnor \U$4364 ( \4585 , \4584 , \764 );
and \U$4365 ( \4586 , \939 , \784 );
and \U$4366 ( \4587 , \952 , \782 );
nor \U$4367 ( \4588 , \4586 , \4587 );
xnor \U$4368 ( \4589 , \4588 , \791 );
xor \U$4369 ( \4590 , \4585 , \4589 );
nand \U$4370 ( \4591 , \960 , \810 );
xnor \U$4371 ( \4592 , \4591 , \819 );
xor \U$4372 ( \4593 , \4590 , \4592 );
xor \U$4373 ( \4594 , \4581 , \4593 );
and \U$4374 ( \4595 , \4547 , \4594 );
and \U$4375 ( \4596 , \4522 , \4594 );
or \U$4376 ( \4597 , \4548 , \4595 , \4596 );
and \U$4377 ( \4598 , \819 , \4540 );
and \U$4378 ( \4599 , \4540 , \4545 );
and \U$4379 ( \4600 , \819 , \4545 );
or \U$4380 ( \4601 , \4598 , \4599 , \4600 );
and \U$4381 ( \4602 , \4526 , \4530 );
and \U$4382 ( \4603 , \4530 , \4535 );
and \U$4383 ( \4604 , \4526 , \4535 );
or \U$4384 ( \4605 , \4602 , \4603 , \4604 );
xor \U$4385 ( \4606 , \4601 , \4605 );
and \U$4386 ( \4607 , \4585 , \4589 );
and \U$4387 ( \4608 , \4589 , \4592 );
and \U$4388 ( \4609 , \4585 , \4592 );
or \U$4389 ( \4610 , \4607 , \4608 , \4609 );
xor \U$4390 ( \4611 , \4606 , \4610 );
xor \U$4391 ( \4612 , \4597 , \4611 );
and \U$4392 ( \4613 , \4564 , \4580 );
and \U$4393 ( \4614 , \4580 , \4593 );
and \U$4394 ( \4615 , \4564 , \4593 );
or \U$4395 ( \4616 , \4613 , \4614 , \4615 );
and \U$4396 ( \4617 , \4536 , \4546 );
xor \U$4397 ( \4618 , \4616 , \4617 );
and \U$4398 ( \4619 , \952 , \784 );
and \U$4399 ( \4620 , \912 , \782 );
nor \U$4400 ( \4621 , \4619 , \4620 );
xnor \U$4401 ( \4622 , \4621 , \791 );
and \U$4402 ( \4623 , \960 , \812 );
and \U$4403 ( \4624 , \939 , \810 );
nor \U$4404 ( \4625 , \4623 , \4624 );
xnor \U$4405 ( \4626 , \4625 , \819 );
xor \U$4406 ( \4627 , \4622 , \4626 );
and \U$4407 ( \4628 , \874 , \698 );
and \U$4408 ( \4629 , \827 , \696 );
nor \U$4409 ( \4630 , \4628 , \4629 );
xnor \U$4410 ( \4631 , \4630 , \705 );
and \U$4411 ( \4632 , \902 , \726 );
and \U$4412 ( \4633 , \854 , \724 );
nor \U$4413 ( \4634 , \4632 , \4633 );
xnor \U$4414 ( \4635 , \4634 , \733 );
xor \U$4415 ( \4636 , \4631 , \4635 );
and \U$4416 ( \4637 , \932 , \757 );
and \U$4417 ( \4638 , \882 , \755 );
nor \U$4418 ( \4639 , \4637 , \4638 );
xnor \U$4419 ( \4640 , \4639 , \764 );
xor \U$4420 ( \4641 , \4636 , \4640 );
xor \U$4421 ( \4642 , \4627 , \4641 );
and \U$4422 ( \4643 , \786 , \616 );
and \U$4423 ( \4644 , \739 , \613 );
nor \U$4424 ( \4645 , \4643 , \4644 );
xnor \U$4425 ( \4646 , \4645 , \576 );
and \U$4426 ( \4647 , \814 , \641 );
and \U$4427 ( \4648 , \766 , \639 );
nor \U$4428 ( \4649 , \4647 , \4648 );
xnor \U$4429 ( \4650 , \4649 , \648 );
xor \U$4430 ( \4651 , \4646 , \4650 );
and \U$4431 ( \4652 , \847 , \671 );
and \U$4432 ( \4653 , \794 , \669 );
nor \U$4433 ( \4654 , \4652 , \4653 );
xnor \U$4434 ( \4655 , \4654 , \678 );
xor \U$4435 ( \4656 , \4651 , \4655 );
xor \U$4436 ( \4657 , \4642 , \4656 );
xor \U$4437 ( \4658 , \4618 , \4657 );
xor \U$4438 ( \4659 , \4612 , \4658 );
and \U$4439 ( \4660 , \847 , \616 );
and \U$4440 ( \4661 , \794 , \613 );
nor \U$4441 ( \4662 , \4660 , \4661 );
xnor \U$4442 ( \4663 , \4662 , \576 );
and \U$4443 ( \4664 , \874 , \641 );
and \U$4444 ( \4665 , \827 , \639 );
nor \U$4445 ( \4666 , \4664 , \4665 );
xnor \U$4446 ( \4667 , \4666 , \648 );
and \U$4447 ( \4668 , \4663 , \4667 );
and \U$4448 ( \4669 , \902 , \671 );
and \U$4449 ( \4670 , \854 , \669 );
nor \U$4450 ( \4671 , \4669 , \4670 );
xnor \U$4451 ( \4672 , \4671 , \678 );
and \U$4452 ( \4673 , \4667 , \4672 );
and \U$4453 ( \4674 , \4663 , \4672 );
or \U$4454 ( \4675 , \4668 , \4673 , \4674 );
and \U$4455 ( \4676 , \932 , \698 );
and \U$4456 ( \4677 , \882 , \696 );
nor \U$4457 ( \4678 , \4676 , \4677 );
xnor \U$4458 ( \4679 , \4678 , \705 );
and \U$4459 ( \4680 , \952 , \726 );
and \U$4460 ( \4681 , \912 , \724 );
nor \U$4461 ( \4682 , \4680 , \4681 );
xnor \U$4462 ( \4683 , \4682 , \733 );
and \U$4463 ( \4684 , \4679 , \4683 );
and \U$4464 ( \4685 , \960 , \757 );
and \U$4465 ( \4686 , \939 , \755 );
nor \U$4466 ( \4687 , \4685 , \4686 );
xnor \U$4467 ( \4688 , \4687 , \764 );
and \U$4468 ( \4689 , \4683 , \4688 );
and \U$4469 ( \4690 , \4679 , \4688 );
or \U$4470 ( \4691 , \4684 , \4689 , \4690 );
and \U$4471 ( \4692 , \4675 , \4691 );
and \U$4472 ( \4693 , \939 , \757 );
and \U$4473 ( \4694 , \952 , \755 );
nor \U$4474 ( \4695 , \4693 , \4694 );
xnor \U$4475 ( \4696 , \4695 , \764 );
and \U$4476 ( \4697 , \4691 , \4696 );
and \U$4477 ( \4698 , \4675 , \4696 );
or \U$4478 ( \4699 , \4692 , \4697 , \4698 );
nand \U$4479 ( \4700 , \960 , \782 );
xnor \U$4480 ( \4701 , \4700 , \791 );
xor \U$4481 ( \4702 , \4502 , \4506 );
xor \U$4482 ( \4703 , \4702 , \4511 );
and \U$4483 ( \4704 , \4701 , \4703 );
xor \U$4484 ( \4705 , \791 , \4490 );
xor \U$4485 ( \4706 , \4705 , \4495 );
and \U$4486 ( \4707 , \4703 , \4706 );
and \U$4487 ( \4708 , \4701 , \4706 );
or \U$4488 ( \4709 , \4704 , \4707 , \4708 );
and \U$4489 ( \4710 , \4699 , \4709 );
xor \U$4490 ( \4711 , \4568 , \4572 );
xor \U$4491 ( \4712 , \4711 , \4577 );
and \U$4492 ( \4713 , \4709 , \4712 );
and \U$4493 ( \4714 , \4699 , \4712 );
or \U$4494 ( \4715 , \4710 , \4713 , \4714 );
xor \U$4495 ( \4716 , \4552 , \4556 );
xor \U$4496 ( \4717 , \4716 , \4561 );
xor \U$4497 ( \4718 , \4498 , \4514 );
xor \U$4498 ( \4719 , \4718 , \4519 );
and \U$4499 ( \4720 , \4717 , \4719 );
and \U$4500 ( \4721 , \4715 , \4720 );
xor \U$4501 ( \4722 , \4522 , \4547 );
xor \U$4502 ( \4723 , \4722 , \4594 );
and \U$4503 ( \4724 , \4720 , \4723 );
and \U$4504 ( \4725 , \4715 , \4723 );
or \U$4505 ( \4726 , \4721 , \4724 , \4725 );
nor \U$4506 ( \4727 , \4659 , \4726 );
and \U$4507 ( \4728 , \4616 , \4617 );
and \U$4508 ( \4729 , \4617 , \4657 );
and \U$4509 ( \4730 , \4616 , \4657 );
or \U$4510 ( \4731 , \4728 , \4729 , \4730 );
nand \U$4511 ( \4732 , \960 , \843 );
xnor \U$4512 ( \4733 , \4732 , \852 );
and \U$4513 ( \4734 , \882 , \757 );
and \U$4514 ( \4735 , \902 , \755 );
nor \U$4515 ( \4736 , \4734 , \4735 );
xnor \U$4516 ( \4737 , \4736 , \764 );
and \U$4517 ( \4738 , \912 , \784 );
and \U$4518 ( \4739 , \932 , \782 );
nor \U$4519 ( \4740 , \4738 , \4739 );
xnor \U$4520 ( \4741 , \4740 , \791 );
xor \U$4521 ( \4742 , \4737 , \4741 );
and \U$4522 ( \4743 , \939 , \812 );
and \U$4523 ( \4744 , \952 , \810 );
nor \U$4524 ( \4745 , \4743 , \4744 );
xnor \U$4525 ( \4746 , \4745 , \819 );
xor \U$4526 ( \4747 , \4742 , \4746 );
xor \U$4527 ( \4748 , \4733 , \4747 );
and \U$4528 ( \4749 , \794 , \671 );
and \U$4529 ( \4750 , \814 , \669 );
nor \U$4530 ( \4751 , \4749 , \4750 );
xnor \U$4531 ( \4752 , \4751 , \678 );
and \U$4532 ( \4753 , \827 , \698 );
and \U$4533 ( \4754 , \847 , \696 );
nor \U$4534 ( \4755 , \4753 , \4754 );
xnor \U$4535 ( \4756 , \4755 , \705 );
xor \U$4536 ( \4757 , \4752 , \4756 );
and \U$4537 ( \4758 , \854 , \726 );
and \U$4538 ( \4759 , \874 , \724 );
nor \U$4539 ( \4760 , \4758 , \4759 );
xnor \U$4540 ( \4761 , \4760 , \733 );
xor \U$4541 ( \4762 , \4757 , \4761 );
xor \U$4542 ( \4763 , \4748 , \4762 );
and \U$4543 ( \4764 , \4646 , \4650 );
and \U$4544 ( \4765 , \4650 , \4655 );
and \U$4545 ( \4766 , \4646 , \4655 );
or \U$4546 ( \4767 , \4764 , \4765 , \4766 );
and \U$4547 ( \4768 , \4631 , \4635 );
and \U$4548 ( \4769 , \4635 , \4640 );
and \U$4549 ( \4770 , \4631 , \4640 );
or \U$4550 ( \4771 , \4768 , \4769 , \4770 );
xor \U$4551 ( \4772 , \4767 , \4771 );
and \U$4552 ( \4773 , \4622 , \4626 );
xor \U$4553 ( \4774 , \4772 , \4773 );
xor \U$4554 ( \4775 , \4763 , \4774 );
xor \U$4555 ( \4776 , \4731 , \4775 );
and \U$4556 ( \4777 , \4601 , \4605 );
and \U$4557 ( \4778 , \4605 , \4610 );
and \U$4558 ( \4779 , \4601 , \4610 );
or \U$4559 ( \4780 , \4777 , \4778 , \4779 );
and \U$4560 ( \4781 , \4627 , \4641 );
and \U$4561 ( \4782 , \4641 , \4656 );
and \U$4562 ( \4783 , \4627 , \4656 );
or \U$4563 ( \4784 , \4781 , \4782 , \4783 );
xor \U$4564 ( \4785 , \4780 , \4784 );
and \U$4565 ( \4786 , \739 , \616 );
and \U$4566 ( \4787 , \759 , \613 );
nor \U$4567 ( \4788 , \4786 , \4787 );
xnor \U$4568 ( \4789 , \4788 , \576 );
xor \U$4569 ( \4790 , \852 , \4789 );
and \U$4570 ( \4791 , \766 , \641 );
and \U$4571 ( \4792 , \786 , \639 );
nor \U$4572 ( \4793 , \4791 , \4792 );
xnor \U$4573 ( \4794 , \4793 , \648 );
xor \U$4574 ( \4795 , \4790 , \4794 );
xor \U$4575 ( \4796 , \4785 , \4795 );
xor \U$4576 ( \4797 , \4776 , \4796 );
and \U$4577 ( \4798 , \4597 , \4611 );
and \U$4578 ( \4799 , \4611 , \4658 );
and \U$4579 ( \4800 , \4597 , \4658 );
or \U$4580 ( \4801 , \4798 , \4799 , \4800 );
nor \U$4581 ( \4802 , \4797 , \4801 );
nor \U$4582 ( \4803 , \4727 , \4802 );
and \U$4583 ( \4804 , \4767 , \4771 );
and \U$4584 ( \4805 , \4771 , \4773 );
and \U$4585 ( \4806 , \4767 , \4773 );
or \U$4586 ( \4807 , \4804 , \4805 , \4806 );
and \U$4587 ( \4808 , \4733 , \4747 );
and \U$4588 ( \4809 , \4747 , \4762 );
and \U$4589 ( \4810 , \4733 , \4762 );
or \U$4590 ( \4811 , \4808 , \4809 , \4810 );
xor \U$4591 ( \4812 , \4807 , \4811 );
and \U$4592 ( \4813 , \932 , \784 );
and \U$4593 ( \4814 , \882 , \782 );
nor \U$4594 ( \4815 , \4813 , \4814 );
xnor \U$4595 ( \4816 , \4815 , \791 );
and \U$4596 ( \4817 , \952 , \812 );
and \U$4597 ( \4818 , \912 , \810 );
nor \U$4598 ( \4819 , \4817 , \4818 );
xnor \U$4599 ( \4820 , \4819 , \819 );
xor \U$4600 ( \4821 , \4816 , \4820 );
and \U$4601 ( \4822 , \960 , \845 );
and \U$4602 ( \4823 , \939 , \843 );
nor \U$4603 ( \4824 , \4822 , \4823 );
xnor \U$4604 ( \4825 , \4824 , \852 );
xor \U$4605 ( \4826 , \4821 , \4825 );
and \U$4606 ( \4827 , \847 , \698 );
and \U$4607 ( \4828 , \794 , \696 );
nor \U$4608 ( \4829 , \4827 , \4828 );
xnor \U$4609 ( \4830 , \4829 , \705 );
and \U$4610 ( \4831 , \874 , \726 );
and \U$4611 ( \4832 , \827 , \724 );
nor \U$4612 ( \4833 , \4831 , \4832 );
xnor \U$4613 ( \4834 , \4833 , \733 );
xor \U$4614 ( \4835 , \4830 , \4834 );
and \U$4615 ( \4836 , \902 , \757 );
and \U$4616 ( \4837 , \854 , \755 );
nor \U$4617 ( \4838 , \4836 , \4837 );
xnor \U$4618 ( \4839 , \4838 , \764 );
xor \U$4619 ( \4840 , \4835 , \4839 );
xor \U$4620 ( \4841 , \4826 , \4840 );
and \U$4621 ( \4842 , \759 , \616 );
and \U$4622 ( \4843 , \708 , \613 );
nor \U$4623 ( \4844 , \4842 , \4843 );
xnor \U$4624 ( \4845 , \4844 , \576 );
and \U$4625 ( \4846 , \786 , \641 );
and \U$4626 ( \4847 , \739 , \639 );
nor \U$4627 ( \4848 , \4846 , \4847 );
xnor \U$4628 ( \4849 , \4848 , \648 );
xor \U$4629 ( \4850 , \4845 , \4849 );
and \U$4630 ( \4851 , \814 , \671 );
and \U$4631 ( \4852 , \766 , \669 );
nor \U$4632 ( \4853 , \4851 , \4852 );
xnor \U$4633 ( \4854 , \4853 , \678 );
xor \U$4634 ( \4855 , \4850 , \4854 );
xor \U$4635 ( \4856 , \4841 , \4855 );
xor \U$4636 ( \4857 , \4812 , \4856 );
and \U$4637 ( \4858 , \4780 , \4784 );
and \U$4638 ( \4859 , \4784 , \4795 );
and \U$4639 ( \4860 , \4780 , \4795 );
or \U$4640 ( \4861 , \4858 , \4859 , \4860 );
and \U$4641 ( \4862 , \4763 , \4774 );
xor \U$4642 ( \4863 , \4861 , \4862 );
and \U$4643 ( \4864 , \852 , \4789 );
and \U$4644 ( \4865 , \4789 , \4794 );
and \U$4645 ( \4866 , \852 , \4794 );
or \U$4646 ( \4867 , \4864 , \4865 , \4866 );
and \U$4647 ( \4868 , \4752 , \4756 );
and \U$4648 ( \4869 , \4756 , \4761 );
and \U$4649 ( \4870 , \4752 , \4761 );
or \U$4650 ( \4871 , \4868 , \4869 , \4870 );
xor \U$4651 ( \4872 , \4867 , \4871 );
and \U$4652 ( \4873 , \4737 , \4741 );
and \U$4653 ( \4874 , \4741 , \4746 );
and \U$4654 ( \4875 , \4737 , \4746 );
or \U$4655 ( \4876 , \4873 , \4874 , \4875 );
xor \U$4656 ( \4877 , \4872 , \4876 );
xor \U$4657 ( \4878 , \4863 , \4877 );
xor \U$4658 ( \4879 , \4857 , \4878 );
and \U$4659 ( \4880 , \4731 , \4775 );
and \U$4660 ( \4881 , \4775 , \4796 );
and \U$4661 ( \4882 , \4731 , \4796 );
or \U$4662 ( \4883 , \4880 , \4881 , \4882 );
nor \U$4663 ( \4884 , \4879 , \4883 );
and \U$4664 ( \4885 , \4861 , \4862 );
and \U$4665 ( \4886 , \4862 , \4877 );
and \U$4666 ( \4887 , \4861 , \4877 );
or \U$4667 ( \4888 , \4885 , \4886 , \4887 );
and \U$4668 ( \4889 , \4807 , \4811 );
and \U$4669 ( \4890 , \4811 , \4856 );
and \U$4670 ( \4891 , \4807 , \4856 );
or \U$4671 ( \4892 , \4889 , \4890 , \4891 );
and \U$4672 ( \4893 , \708 , \616 );
and \U$4673 ( \4894 , \728 , \613 );
nor \U$4674 ( \4895 , \4893 , \4894 );
xnor \U$4675 ( \4896 , \4895 , \576 );
xor \U$4676 ( \4897 , \879 , \4896 );
and \U$4677 ( \4898 , \739 , \641 );
and \U$4678 ( \4899 , \759 , \639 );
nor \U$4679 ( \4900 , \4898 , \4899 );
xnor \U$4680 ( \4901 , \4900 , \648 );
xor \U$4681 ( \4902 , \4897 , \4901 );
and \U$4682 ( \4903 , \939 , \845 );
and \U$4683 ( \4904 , \952 , \843 );
nor \U$4684 ( \4905 , \4903 , \4904 );
xnor \U$4685 ( \4906 , \4905 , \852 );
nand \U$4686 ( \4907 , \960 , \870 );
xnor \U$4687 ( \4908 , \4907 , \879 );
xor \U$4688 ( \4909 , \4906 , \4908 );
and \U$4689 ( \4910 , \854 , \757 );
and \U$4690 ( \4911 , \874 , \755 );
nor \U$4691 ( \4912 , \4910 , \4911 );
xnor \U$4692 ( \4913 , \4912 , \764 );
and \U$4693 ( \4914 , \882 , \784 );
and \U$4694 ( \4915 , \902 , \782 );
nor \U$4695 ( \4916 , \4914 , \4915 );
xnor \U$4696 ( \4917 , \4916 , \791 );
xor \U$4697 ( \4918 , \4913 , \4917 );
and \U$4698 ( \4919 , \912 , \812 );
and \U$4699 ( \4920 , \932 , \810 );
nor \U$4700 ( \4921 , \4919 , \4920 );
xnor \U$4701 ( \4922 , \4921 , \819 );
xor \U$4702 ( \4923 , \4918 , \4922 );
xor \U$4703 ( \4924 , \4909 , \4923 );
xor \U$4704 ( \4925 , \4902 , \4924 );
and \U$4705 ( \4926 , \4845 , \4849 );
and \U$4706 ( \4927 , \4849 , \4854 );
and \U$4707 ( \4928 , \4845 , \4854 );
or \U$4708 ( \4929 , \4926 , \4927 , \4928 );
and \U$4709 ( \4930 , \4830 , \4834 );
and \U$4710 ( \4931 , \4834 , \4839 );
and \U$4711 ( \4932 , \4830 , \4839 );
or \U$4712 ( \4933 , \4930 , \4931 , \4932 );
xor \U$4713 ( \4934 , \4929 , \4933 );
and \U$4714 ( \4935 , \4816 , \4820 );
and \U$4715 ( \4936 , \4820 , \4825 );
and \U$4716 ( \4937 , \4816 , \4825 );
or \U$4717 ( \4938 , \4935 , \4936 , \4937 );
xor \U$4718 ( \4939 , \4934 , \4938 );
xor \U$4719 ( \4940 , \4925 , \4939 );
xor \U$4720 ( \4941 , \4892 , \4940 );
and \U$4721 ( \4942 , \4867 , \4871 );
and \U$4722 ( \4943 , \4871 , \4876 );
and \U$4723 ( \4944 , \4867 , \4876 );
or \U$4724 ( \4945 , \4942 , \4943 , \4944 );
and \U$4725 ( \4946 , \4826 , \4840 );
and \U$4726 ( \4947 , \4840 , \4855 );
and \U$4727 ( \4948 , \4826 , \4855 );
or \U$4728 ( \4949 , \4946 , \4947 , \4948 );
xor \U$4729 ( \4950 , \4945 , \4949 );
and \U$4730 ( \4951 , \766 , \671 );
and \U$4731 ( \4952 , \786 , \669 );
nor \U$4732 ( \4953 , \4951 , \4952 );
xnor \U$4733 ( \4954 , \4953 , \678 );
and \U$4734 ( \4955 , \794 , \698 );
and \U$4735 ( \4956 , \814 , \696 );
nor \U$4736 ( \4957 , \4955 , \4956 );
xnor \U$4737 ( \4958 , \4957 , \705 );
xor \U$4738 ( \4959 , \4954 , \4958 );
and \U$4739 ( \4960 , \827 , \726 );
and \U$4740 ( \4961 , \847 , \724 );
nor \U$4741 ( \4962 , \4960 , \4961 );
xnor \U$4742 ( \4963 , \4962 , \733 );
xor \U$4743 ( \4964 , \4959 , \4963 );
xor \U$4744 ( \4965 , \4950 , \4964 );
xor \U$4745 ( \4966 , \4941 , \4965 );
xor \U$4746 ( \4967 , \4888 , \4966 );
and \U$4747 ( \4968 , \4857 , \4878 );
nor \U$4748 ( \4969 , \4967 , \4968 );
nor \U$4749 ( \4970 , \4884 , \4969 );
nand \U$4750 ( \4971 , \4803 , \4970 );
and \U$4751 ( \4972 , \4892 , \4940 );
and \U$4752 ( \4973 , \4940 , \4965 );
and \U$4753 ( \4974 , \4892 , \4965 );
or \U$4754 ( \4975 , \4972 , \4973 , \4974 );
and \U$4755 ( \4976 , \879 , \4896 );
and \U$4756 ( \4977 , \4896 , \4901 );
and \U$4757 ( \4978 , \879 , \4901 );
or \U$4758 ( \4979 , \4976 , \4977 , \4978 );
and \U$4759 ( \4980 , \4954 , \4958 );
and \U$4760 ( \4981 , \4958 , \4963 );
and \U$4761 ( \4982 , \4954 , \4963 );
or \U$4762 ( \4983 , \4980 , \4981 , \4982 );
xor \U$4763 ( \4984 , \4979 , \4983 );
and \U$4764 ( \4985 , \4913 , \4917 );
and \U$4765 ( \4986 , \4917 , \4922 );
and \U$4766 ( \4987 , \4913 , \4922 );
or \U$4767 ( \4988 , \4985 , \4986 , \4987 );
xor \U$4768 ( \4989 , \4984 , \4988 );
and \U$4769 ( \4990 , \4929 , \4933 );
and \U$4770 ( \4991 , \4933 , \4938 );
and \U$4771 ( \4992 , \4929 , \4938 );
or \U$4772 ( \4993 , \4990 , \4991 , \4992 );
and \U$4773 ( \4994 , \4906 , \4908 );
and \U$4774 ( \4995 , \4908 , \4923 );
and \U$4775 ( \4996 , \4906 , \4923 );
or \U$4776 ( \4997 , \4994 , \4995 , \4996 );
xor \U$4777 ( \4998 , \4993 , \4997 );
and \U$4778 ( \4999 , \728 , \616 );
and \U$4779 ( \5000 , \680 , \613 );
nor \U$4780 ( \5001 , \4999 , \5000 );
xnor \U$4781 ( \5002 , \5001 , \576 );
and \U$4782 ( \5003 , \759 , \641 );
and \U$4783 ( \5004 , \708 , \639 );
nor \U$4784 ( \5005 , \5003 , \5004 );
xnor \U$4785 ( \5006 , \5005 , \648 );
xor \U$4786 ( \5007 , \5002 , \5006 );
and \U$4787 ( \5008 , \786 , \671 );
and \U$4788 ( \5009 , \739 , \669 );
nor \U$4789 ( \5010 , \5008 , \5009 );
xnor \U$4790 ( \5011 , \5010 , \678 );
xor \U$4791 ( \5012 , \5007 , \5011 );
xor \U$4792 ( \5013 , \4998 , \5012 );
xor \U$4793 ( \5014 , \4989 , \5013 );
xor \U$4794 ( \5015 , \4975 , \5014 );
and \U$4795 ( \5016 , \4945 , \4949 );
and \U$4796 ( \5017 , \4949 , \4964 );
and \U$4797 ( \5018 , \4945 , \4964 );
or \U$4798 ( \5019 , \5016 , \5017 , \5018 );
and \U$4799 ( \5020 , \4902 , \4924 );
and \U$4800 ( \5021 , \4924 , \4939 );
and \U$4801 ( \5022 , \4902 , \4939 );
or \U$4802 ( \5023 , \5020 , \5021 , \5022 );
xor \U$4803 ( \5024 , \5019 , \5023 );
and \U$4804 ( \5025 , \960 , \872 );
and \U$4805 ( \5026 , \939 , \870 );
nor \U$4806 ( \5027 , \5025 , \5026 );
xnor \U$4807 ( \5028 , \5027 , \879 );
and \U$4808 ( \5029 , \902 , \784 );
and \U$4809 ( \5030 , \854 , \782 );
nor \U$4810 ( \5031 , \5029 , \5030 );
xnor \U$4811 ( \5032 , \5031 , \791 );
and \U$4812 ( \5033 , \932 , \812 );
and \U$4813 ( \5034 , \882 , \810 );
nor \U$4814 ( \5035 , \5033 , \5034 );
xnor \U$4815 ( \5036 , \5035 , \819 );
xor \U$4816 ( \5037 , \5032 , \5036 );
and \U$4817 ( \5038 , \952 , \845 );
and \U$4818 ( \5039 , \912 , \843 );
nor \U$4819 ( \5040 , \5038 , \5039 );
xnor \U$4820 ( \5041 , \5040 , \852 );
xor \U$4821 ( \5042 , \5037 , \5041 );
xor \U$4822 ( \5043 , \5028 , \5042 );
and \U$4823 ( \5044 , \814 , \698 );
and \U$4824 ( \5045 , \766 , \696 );
nor \U$4825 ( \5046 , \5044 , \5045 );
xnor \U$4826 ( \5047 , \5046 , \705 );
and \U$4827 ( \5048 , \847 , \726 );
and \U$4828 ( \5049 , \794 , \724 );
nor \U$4829 ( \5050 , \5048 , \5049 );
xnor \U$4830 ( \5051 , \5050 , \733 );
xor \U$4831 ( \5052 , \5047 , \5051 );
and \U$4832 ( \5053 , \874 , \757 );
and \U$4833 ( \5054 , \827 , \755 );
nor \U$4834 ( \5055 , \5053 , \5054 );
xnor \U$4835 ( \5056 , \5055 , \764 );
xor \U$4836 ( \5057 , \5052 , \5056 );
xor \U$4837 ( \5058 , \5043 , \5057 );
xor \U$4838 ( \5059 , \5024 , \5058 );
xor \U$4839 ( \5060 , \5015 , \5059 );
and \U$4840 ( \5061 , \4888 , \4966 );
nor \U$4841 ( \5062 , \5060 , \5061 );
and \U$4842 ( \5063 , \5019 , \5023 );
and \U$4843 ( \5064 , \5023 , \5058 );
and \U$4844 ( \5065 , \5019 , \5058 );
or \U$4845 ( \5066 , \5063 , \5064 , \5065 );
and \U$4846 ( \5067 , \4989 , \5013 );
xor \U$4847 ( \5068 , \5066 , \5067 );
and \U$4848 ( \5069 , \4993 , \4997 );
and \U$4849 ( \5070 , \4997 , \5012 );
and \U$4850 ( \5071 , \4993 , \5012 );
or \U$4851 ( \5072 , \5069 , \5070 , \5071 );
and \U$4852 ( \5073 , \912 , \845 );
and \U$4853 ( \5074 , \932 , \843 );
nor \U$4854 ( \5075 , \5073 , \5074 );
xnor \U$4855 ( \5076 , \5075 , \852 );
and \U$4856 ( \5077 , \939 , \872 );
and \U$4857 ( \5078 , \952 , \870 );
nor \U$4858 ( \5079 , \5077 , \5078 );
xnor \U$4859 ( \5080 , \5079 , \879 );
xor \U$4860 ( \5081 , \5076 , \5080 );
nand \U$4861 ( \5082 , \960 , \898 );
xnor \U$4862 ( \5083 , \5082 , \907 );
xor \U$4863 ( \5084 , \5081 , \5083 );
and \U$4864 ( \5085 , \827 , \757 );
and \U$4865 ( \5086 , \847 , \755 );
nor \U$4866 ( \5087 , \5085 , \5086 );
xnor \U$4867 ( \5088 , \5087 , \764 );
and \U$4868 ( \5089 , \854 , \784 );
and \U$4869 ( \5090 , \874 , \782 );
nor \U$4870 ( \5091 , \5089 , \5090 );
xnor \U$4871 ( \5092 , \5091 , \791 );
xor \U$4872 ( \5093 , \5088 , \5092 );
and \U$4873 ( \5094 , \882 , \812 );
and \U$4874 ( \5095 , \902 , \810 );
nor \U$4875 ( \5096 , \5094 , \5095 );
xnor \U$4876 ( \5097 , \5096 , \819 );
xor \U$4877 ( \5098 , \5093 , \5097 );
xor \U$4878 ( \5099 , \5084 , \5098 );
and \U$4879 ( \5100 , \739 , \671 );
and \U$4880 ( \5101 , \759 , \669 );
nor \U$4881 ( \5102 , \5100 , \5101 );
xnor \U$4882 ( \5103 , \5102 , \678 );
and \U$4883 ( \5104 , \766 , \698 );
and \U$4884 ( \5105 , \786 , \696 );
nor \U$4885 ( \5106 , \5104 , \5105 );
xnor \U$4886 ( \5107 , \5106 , \705 );
xor \U$4887 ( \5108 , \5103 , \5107 );
and \U$4888 ( \5109 , \794 , \726 );
and \U$4889 ( \5110 , \814 , \724 );
nor \U$4890 ( \5111 , \5109 , \5110 );
xnor \U$4891 ( \5112 , \5111 , \733 );
xor \U$4892 ( \5113 , \5108 , \5112 );
xor \U$4893 ( \5114 , \5099 , \5113 );
and \U$4894 ( \5115 , \5002 , \5006 );
and \U$4895 ( \5116 , \5006 , \5011 );
and \U$4896 ( \5117 , \5002 , \5011 );
or \U$4897 ( \5118 , \5115 , \5116 , \5117 );
and \U$4898 ( \5119 , \5047 , \5051 );
and \U$4899 ( \5120 , \5051 , \5056 );
and \U$4900 ( \5121 , \5047 , \5056 );
or \U$4901 ( \5122 , \5119 , \5120 , \5121 );
xor \U$4902 ( \5123 , \5118 , \5122 );
and \U$4903 ( \5124 , \5032 , \5036 );
and \U$4904 ( \5125 , \5036 , \5041 );
and \U$4905 ( \5126 , \5032 , \5041 );
or \U$4906 ( \5127 , \5124 , \5125 , \5126 );
xor \U$4907 ( \5128 , \5123 , \5127 );
xor \U$4908 ( \5129 , \5114 , \5128 );
xor \U$4909 ( \5130 , \5072 , \5129 );
and \U$4910 ( \5131 , \4979 , \4983 );
and \U$4911 ( \5132 , \4983 , \4988 );
and \U$4912 ( \5133 , \4979 , \4988 );
or \U$4913 ( \5134 , \5131 , \5132 , \5133 );
and \U$4914 ( \5135 , \5028 , \5042 );
and \U$4915 ( \5136 , \5042 , \5057 );
and \U$4916 ( \5137 , \5028 , \5057 );
or \U$4917 ( \5138 , \5135 , \5136 , \5137 );
xor \U$4918 ( \5139 , \5134 , \5138 );
and \U$4919 ( \5140 , \680 , \616 );
and \U$4920 ( \5141 , \700 , \613 );
nor \U$4921 ( \5142 , \5140 , \5141 );
xnor \U$4922 ( \5143 , \5142 , \576 );
xor \U$4923 ( \5144 , \907 , \5143 );
and \U$4924 ( \5145 , \708 , \641 );
and \U$4925 ( \5146 , \728 , \639 );
nor \U$4926 ( \5147 , \5145 , \5146 );
xnor \U$4927 ( \5148 , \5147 , \648 );
xor \U$4928 ( \5149 , \5144 , \5148 );
xor \U$4929 ( \5150 , \5139 , \5149 );
xor \U$4930 ( \5151 , \5130 , \5150 );
xor \U$4931 ( \5152 , \5068 , \5151 );
and \U$4932 ( \5153 , \4975 , \5014 );
and \U$4933 ( \5154 , \5014 , \5059 );
and \U$4934 ( \5155 , \4975 , \5059 );
or \U$4935 ( \5156 , \5153 , \5154 , \5155 );
nor \U$4936 ( \5157 , \5152 , \5156 );
nor \U$4937 ( \5158 , \5062 , \5157 );
and \U$4938 ( \5159 , \5072 , \5129 );
and \U$4939 ( \5160 , \5129 , \5150 );
and \U$4940 ( \5161 , \5072 , \5150 );
or \U$4941 ( \5162 , \5159 , \5160 , \5161 );
and \U$4942 ( \5163 , \907 , \5143 );
and \U$4943 ( \5164 , \5143 , \5148 );
and \U$4944 ( \5165 , \907 , \5148 );
or \U$4945 ( \5166 , \5163 , \5164 , \5165 );
and \U$4946 ( \5167 , \5103 , \5107 );
and \U$4947 ( \5168 , \5107 , \5112 );
and \U$4948 ( \5169 , \5103 , \5112 );
or \U$4949 ( \5170 , \5167 , \5168 , \5169 );
xor \U$4950 ( \5171 , \5166 , \5170 );
and \U$4951 ( \5172 , \5088 , \5092 );
and \U$4952 ( \5173 , \5092 , \5097 );
and \U$4953 ( \5174 , \5088 , \5097 );
or \U$4954 ( \5175 , \5172 , \5173 , \5174 );
xor \U$4955 ( \5176 , \5171 , \5175 );
and \U$4956 ( \5177 , \5118 , \5122 );
and \U$4957 ( \5178 , \5122 , \5127 );
and \U$4958 ( \5179 , \5118 , \5127 );
or \U$4959 ( \5180 , \5177 , \5178 , \5179 );
and \U$4960 ( \5181 , \5084 , \5098 );
and \U$4961 ( \5182 , \5098 , \5113 );
and \U$4962 ( \5183 , \5084 , \5113 );
or \U$4963 ( \5184 , \5181 , \5182 , \5183 );
xor \U$4964 ( \5185 , \5180 , \5184 );
and \U$4965 ( \5186 , \874 , \784 );
and \U$4966 ( \5187 , \827 , \782 );
nor \U$4967 ( \5188 , \5186 , \5187 );
xnor \U$4968 ( \5189 , \5188 , \791 );
and \U$4969 ( \5190 , \902 , \812 );
and \U$4970 ( \5191 , \854 , \810 );
nor \U$4971 ( \5192 , \5190 , \5191 );
xnor \U$4972 ( \5193 , \5192 , \819 );
xor \U$4973 ( \5194 , \5189 , \5193 );
and \U$4974 ( \5195 , \932 , \845 );
and \U$4975 ( \5196 , \882 , \843 );
nor \U$4976 ( \5197 , \5195 , \5196 );
xnor \U$4977 ( \5198 , \5197 , \852 );
xor \U$4978 ( \5199 , \5194 , \5198 );
and \U$4979 ( \5200 , \786 , \698 );
and \U$4980 ( \5201 , \739 , \696 );
nor \U$4981 ( \5202 , \5200 , \5201 );
xnor \U$4982 ( \5203 , \5202 , \705 );
and \U$4983 ( \5204 , \814 , \726 );
and \U$4984 ( \5205 , \766 , \724 );
nor \U$4985 ( \5206 , \5204 , \5205 );
xnor \U$4986 ( \5207 , \5206 , \733 );
xor \U$4987 ( \5208 , \5203 , \5207 );
and \U$4988 ( \5209 , \847 , \757 );
and \U$4989 ( \5210 , \794 , \755 );
nor \U$4990 ( \5211 , \5209 , \5210 );
xnor \U$4991 ( \5212 , \5211 , \764 );
xor \U$4992 ( \5213 , \5208 , \5212 );
xor \U$4993 ( \5214 , \5199 , \5213 );
and \U$4994 ( \5215 , \700 , \616 );
and \U$4995 ( \5216 , \653 , \613 );
nor \U$4996 ( \5217 , \5215 , \5216 );
xnor \U$4997 ( \5218 , \5217 , \576 );
and \U$4998 ( \5219 , \728 , \641 );
and \U$4999 ( \5220 , \680 , \639 );
nor \U$5000 ( \5221 , \5219 , \5220 );
xnor \U$5001 ( \5222 , \5221 , \648 );
xor \U$5002 ( \5223 , \5218 , \5222 );
and \U$5003 ( \5224 , \759 , \671 );
and \U$5004 ( \5225 , \708 , \669 );
nor \U$5005 ( \5226 , \5224 , \5225 );
xnor \U$5006 ( \5227 , \5226 , \678 );
xor \U$5007 ( \5228 , \5223 , \5227 );
xor \U$5008 ( \5229 , \5214 , \5228 );
xor \U$5009 ( \5230 , \5185 , \5229 );
xor \U$5010 ( \5231 , \5176 , \5230 );
xor \U$5011 ( \5232 , \5162 , \5231 );
and \U$5012 ( \5233 , \5134 , \5138 );
and \U$5013 ( \5234 , \5138 , \5149 );
and \U$5014 ( \5235 , \5134 , \5149 );
or \U$5015 ( \5236 , \5233 , \5234 , \5235 );
and \U$5016 ( \5237 , \5114 , \5128 );
xor \U$5017 ( \5238 , \5236 , \5237 );
and \U$5018 ( \5239 , \5076 , \5080 );
and \U$5019 ( \5240 , \5080 , \5083 );
and \U$5020 ( \5241 , \5076 , \5083 );
or \U$5021 ( \5242 , \5239 , \5240 , \5241 );
and \U$5022 ( \5243 , \952 , \872 );
and \U$5023 ( \5244 , \912 , \870 );
nor \U$5024 ( \5245 , \5243 , \5244 );
xnor \U$5025 ( \5246 , \5245 , \879 );
xor \U$5026 ( \5247 , \5242 , \5246 );
and \U$5027 ( \5248 , \960 , \900 );
and \U$5028 ( \5249 , \939 , \898 );
nor \U$5029 ( \5250 , \5248 , \5249 );
xnor \U$5030 ( \5251 , \5250 , \907 );
xor \U$5031 ( \5252 , \5247 , \5251 );
xor \U$5032 ( \5253 , \5238 , \5252 );
xor \U$5033 ( \5254 , \5232 , \5253 );
and \U$5034 ( \5255 , \5066 , \5067 );
and \U$5035 ( \5256 , \5067 , \5151 );
and \U$5036 ( \5257 , \5066 , \5151 );
or \U$5037 ( \5258 , \5255 , \5256 , \5257 );
nor \U$5038 ( \5259 , \5254 , \5258 );
and \U$5039 ( \5260 , \5236 , \5237 );
and \U$5040 ( \5261 , \5237 , \5252 );
and \U$5041 ( \5262 , \5236 , \5252 );
or \U$5042 ( \5263 , \5260 , \5261 , \5262 );
and \U$5043 ( \5264 , \5176 , \5230 );
xor \U$5044 ( \5265 , \5263 , \5264 );
and \U$5045 ( \5266 , \5180 , \5184 );
and \U$5046 ( \5267 , \5184 , \5229 );
and \U$5047 ( \5268 , \5180 , \5229 );
or \U$5048 ( \5269 , \5266 , \5267 , \5268 );
and \U$5049 ( \5270 , \708 , \671 );
and \U$5050 ( \5271 , \728 , \669 );
nor \U$5051 ( \5272 , \5270 , \5271 );
xnor \U$5052 ( \5273 , \5272 , \678 );
and \U$5053 ( \5274 , \739 , \698 );
and \U$5054 ( \5275 , \759 , \696 );
nor \U$5055 ( \5276 , \5274 , \5275 );
xnor \U$5056 ( \5277 , \5276 , \705 );
xor \U$5057 ( \5278 , \5273 , \5277 );
and \U$5058 ( \5279 , \766 , \726 );
and \U$5059 ( \5280 , \786 , \724 );
nor \U$5060 ( \5281 , \5279 , \5280 );
xnor \U$5061 ( \5282 , \5281 , \733 );
xor \U$5062 ( \5283 , \5278 , \5282 );
and \U$5063 ( \5284 , \653 , \616 );
and \U$5064 ( \5285 , \673 , \613 );
nor \U$5065 ( \5286 , \5284 , \5285 );
xnor \U$5066 ( \5287 , \5286 , \576 );
xor \U$5067 ( \5288 , \937 , \5287 );
and \U$5068 ( \5289 , \680 , \641 );
and \U$5069 ( \5290 , \700 , \639 );
nor \U$5070 ( \5291 , \5289 , \5290 );
xnor \U$5071 ( \5292 , \5291 , \648 );
xor \U$5072 ( \5293 , \5288 , \5292 );
xor \U$5073 ( \5294 , \5283 , \5293 );
nand \U$5074 ( \5295 , \960 , \928 );
xnor \U$5075 ( \5296 , \5295 , \937 );
and \U$5076 ( \5297 , \882 , \845 );
and \U$5077 ( \5298 , \902 , \843 );
nor \U$5078 ( \5299 , \5297 , \5298 );
xnor \U$5079 ( \5300 , \5299 , \852 );
and \U$5080 ( \5301 , \912 , \872 );
and \U$5081 ( \5302 , \932 , \870 );
nor \U$5082 ( \5303 , \5301 , \5302 );
xnor \U$5083 ( \5304 , \5303 , \879 );
xor \U$5084 ( \5305 , \5300 , \5304 );
and \U$5085 ( \5306 , \939 , \900 );
and \U$5086 ( \5307 , \952 , \898 );
nor \U$5087 ( \5308 , \5306 , \5307 );
xnor \U$5088 ( \5309 , \5308 , \907 );
xor \U$5089 ( \5310 , \5305 , \5309 );
xor \U$5090 ( \5311 , \5296 , \5310 );
and \U$5091 ( \5312 , \794 , \757 );
and \U$5092 ( \5313 , \814 , \755 );
nor \U$5093 ( \5314 , \5312 , \5313 );
xnor \U$5094 ( \5315 , \5314 , \764 );
and \U$5095 ( \5316 , \827 , \784 );
and \U$5096 ( \5317 , \847 , \782 );
nor \U$5097 ( \5318 , \5316 , \5317 );
xnor \U$5098 ( \5319 , \5318 , \791 );
xor \U$5099 ( \5320 , \5315 , \5319 );
and \U$5100 ( \5321 , \854 , \812 );
and \U$5101 ( \5322 , \874 , \810 );
nor \U$5102 ( \5323 , \5321 , \5322 );
xnor \U$5103 ( \5324 , \5323 , \819 );
xor \U$5104 ( \5325 , \5320 , \5324 );
xor \U$5105 ( \5326 , \5311 , \5325 );
xor \U$5106 ( \5327 , \5294 , \5326 );
and \U$5107 ( \5328 , \5218 , \5222 );
and \U$5108 ( \5329 , \5222 , \5227 );
and \U$5109 ( \5330 , \5218 , \5227 );
or \U$5110 ( \5331 , \5328 , \5329 , \5330 );
and \U$5111 ( \5332 , \5203 , \5207 );
and \U$5112 ( \5333 , \5207 , \5212 );
and \U$5113 ( \5334 , \5203 , \5212 );
or \U$5114 ( \5335 , \5332 , \5333 , \5334 );
xor \U$5115 ( \5336 , \5331 , \5335 );
and \U$5116 ( \5337 , \5189 , \5193 );
and \U$5117 ( \5338 , \5193 , \5198 );
and \U$5118 ( \5339 , \5189 , \5198 );
or \U$5119 ( \5340 , \5337 , \5338 , \5339 );
xor \U$5120 ( \5341 , \5336 , \5340 );
xor \U$5121 ( \5342 , \5327 , \5341 );
xor \U$5122 ( \5343 , \5269 , \5342 );
and \U$5123 ( \5344 , \5166 , \5170 );
and \U$5124 ( \5345 , \5170 , \5175 );
and \U$5125 ( \5346 , \5166 , \5175 );
or \U$5126 ( \5347 , \5344 , \5345 , \5346 );
and \U$5127 ( \5348 , \5242 , \5246 );
and \U$5128 ( \5349 , \5246 , \5251 );
and \U$5129 ( \5350 , \5242 , \5251 );
or \U$5130 ( \5351 , \5348 , \5349 , \5350 );
xor \U$5131 ( \5352 , \5347 , \5351 );
and \U$5132 ( \5353 , \5199 , \5213 );
and \U$5133 ( \5354 , \5213 , \5228 );
and \U$5134 ( \5355 , \5199 , \5228 );
or \U$5135 ( \5356 , \5353 , \5354 , \5355 );
xor \U$5136 ( \5357 , \5352 , \5356 );
xor \U$5137 ( \5358 , \5343 , \5357 );
xor \U$5138 ( \5359 , \5265 , \5358 );
and \U$5139 ( \5360 , \5162 , \5231 );
and \U$5140 ( \5361 , \5231 , \5253 );
and \U$5141 ( \5362 , \5162 , \5253 );
or \U$5142 ( \5363 , \5360 , \5361 , \5362 );
nor \U$5143 ( \5364 , \5359 , \5363 );
nor \U$5144 ( \5365 , \5259 , \5364 );
nand \U$5145 ( \5366 , \5158 , \5365 );
nor \U$5146 ( \5367 , \4971 , \5366 );
and \U$5147 ( \5368 , \5269 , \5342 );
and \U$5148 ( \5369 , \5342 , \5357 );
and \U$5149 ( \5370 , \5269 , \5357 );
or \U$5150 ( \5371 , \5368 , \5369 , \5370 );
and \U$5151 ( \5372 , \5331 , \5335 );
and \U$5152 ( \5373 , \5335 , \5340 );
and \U$5153 ( \5374 , \5331 , \5340 );
or \U$5154 ( \5375 , \5372 , \5373 , \5374 );
and \U$5155 ( \5376 , \5296 , \5310 );
and \U$5156 ( \5377 , \5310 , \5325 );
and \U$5157 ( \5378 , \5296 , \5325 );
or \U$5158 ( \5379 , \5376 , \5377 , \5378 );
xor \U$5159 ( \5380 , \5375 , \5379 );
and \U$5160 ( \5381 , \5283 , \5293 );
xor \U$5161 ( \5382 , \5380 , \5381 );
xor \U$5162 ( \5383 , \5371 , \5382 );
and \U$5163 ( \5384 , \5347 , \5351 );
and \U$5164 ( \5385 , \5351 , \5356 );
and \U$5165 ( \5386 , \5347 , \5356 );
or \U$5166 ( \5387 , \5384 , \5385 , \5386 );
and \U$5167 ( \5388 , \5294 , \5326 );
and \U$5168 ( \5389 , \5326 , \5341 );
and \U$5169 ( \5390 , \5294 , \5341 );
or \U$5170 ( \5391 , \5388 , \5389 , \5390 );
xor \U$5171 ( \5392 , \5387 , \5391 );
and \U$5172 ( \5393 , \759 , \698 );
and \U$5173 ( \5394 , \708 , \696 );
nor \U$5174 ( \5395 , \5393 , \5394 );
xnor \U$5175 ( \5396 , \5395 , \705 );
and \U$5176 ( \5397 , \786 , \726 );
and \U$5177 ( \5398 , \739 , \724 );
nor \U$5178 ( \5399 , \5397 , \5398 );
xnor \U$5179 ( \5400 , \5399 , \733 );
xor \U$5180 ( \5401 , \5396 , \5400 );
and \U$5181 ( \5402 , \814 , \757 );
and \U$5182 ( \5403 , \766 , \755 );
nor \U$5183 ( \5404 , \5402 , \5403 );
xnor \U$5184 ( \5405 , \5404 , \764 );
xor \U$5185 ( \5406 , \5401 , \5405 );
and \U$5186 ( \5407 , \673 , \616 );
and \U$5187 ( \5408 , \623 , \613 );
nor \U$5188 ( \5409 , \5407 , \5408 );
xnor \U$5189 ( \5410 , \5409 , \576 );
and \U$5190 ( \5411 , \700 , \641 );
and \U$5191 ( \5412 , \653 , \639 );
nor \U$5192 ( \5413 , \5411 , \5412 );
xnor \U$5193 ( \5414 , \5413 , \648 );
xor \U$5194 ( \5415 , \5410 , \5414 );
and \U$5195 ( \5416 , \728 , \671 );
and \U$5196 ( \5417 , \680 , \669 );
nor \U$5197 ( \5418 , \5416 , \5417 );
xnor \U$5198 ( \5419 , \5418 , \678 );
xor \U$5199 ( \5420 , \5415 , \5419 );
xor \U$5200 ( \5421 , \5406 , \5420 );
and \U$5201 ( \5422 , \5300 , \5304 );
and \U$5202 ( \5423 , \5304 , \5309 );
and \U$5203 ( \5424 , \5300 , \5309 );
or \U$5204 ( \5425 , \5422 , \5423 , \5424 );
and \U$5205 ( \5426 , \932 , \872 );
and \U$5206 ( \5427 , \882 , \870 );
nor \U$5207 ( \5428 , \5426 , \5427 );
xnor \U$5208 ( \5429 , \5428 , \879 );
and \U$5209 ( \5430 , \952 , \900 );
and \U$5210 ( \5431 , \912 , \898 );
nor \U$5211 ( \5432 , \5430 , \5431 );
xnor \U$5212 ( \5433 , \5432 , \907 );
xor \U$5213 ( \5434 , \5429 , \5433 );
and \U$5214 ( \5435 , \960 , \930 );
and \U$5215 ( \5436 , \939 , \928 );
nor \U$5216 ( \5437 , \5435 , \5436 );
xnor \U$5217 ( \5438 , \5437 , \937 );
xor \U$5218 ( \5439 , \5434 , \5438 );
xor \U$5219 ( \5440 , \5425 , \5439 );
and \U$5220 ( \5441 , \847 , \784 );
and \U$5221 ( \5442 , \794 , \782 );
nor \U$5222 ( \5443 , \5441 , \5442 );
xnor \U$5223 ( \5444 , \5443 , \791 );
and \U$5224 ( \5445 , \874 , \812 );
and \U$5225 ( \5446 , \827 , \810 );
nor \U$5226 ( \5447 , \5445 , \5446 );
xnor \U$5227 ( \5448 , \5447 , \819 );
xor \U$5228 ( \5449 , \5444 , \5448 );
and \U$5229 ( \5450 , \902 , \845 );
and \U$5230 ( \5451 , \854 , \843 );
nor \U$5231 ( \5452 , \5450 , \5451 );
xnor \U$5232 ( \5453 , \5452 , \852 );
xor \U$5233 ( \5454 , \5449 , \5453 );
xor \U$5234 ( \5455 , \5440 , \5454 );
xor \U$5235 ( \5456 , \5421 , \5455 );
and \U$5236 ( \5457 , \937 , \5287 );
and \U$5237 ( \5458 , \5287 , \5292 );
and \U$5238 ( \5459 , \937 , \5292 );
or \U$5239 ( \5460 , \5457 , \5458 , \5459 );
and \U$5240 ( \5461 , \5273 , \5277 );
and \U$5241 ( \5462 , \5277 , \5282 );
and \U$5242 ( \5463 , \5273 , \5282 );
or \U$5243 ( \5464 , \5461 , \5462 , \5463 );
xor \U$5244 ( \5465 , \5460 , \5464 );
and \U$5245 ( \5466 , \5315 , \5319 );
and \U$5246 ( \5467 , \5319 , \5324 );
and \U$5247 ( \5468 , \5315 , \5324 );
or \U$5248 ( \5469 , \5466 , \5467 , \5468 );
xor \U$5249 ( \5470 , \5465 , \5469 );
xor \U$5250 ( \5471 , \5456 , \5470 );
xor \U$5251 ( \5472 , \5392 , \5471 );
xor \U$5252 ( \5473 , \5383 , \5472 );
and \U$5253 ( \5474 , \5263 , \5264 );
and \U$5254 ( \5475 , \5264 , \5358 );
and \U$5255 ( \5476 , \5263 , \5358 );
or \U$5256 ( \5477 , \5474 , \5475 , \5476 );
nor \U$5257 ( \5478 , \5473 , \5477 );
and \U$5258 ( \5479 , \5387 , \5391 );
and \U$5259 ( \5480 , \5391 , \5471 );
and \U$5260 ( \5481 , \5387 , \5471 );
or \U$5261 ( \5482 , \5479 , \5480 , \5481 );
and \U$5262 ( \5483 , \5460 , \5464 );
and \U$5263 ( \5484 , \5464 , \5469 );
and \U$5264 ( \5485 , \5460 , \5469 );
or \U$5265 ( \5486 , \5483 , \5484 , \5485 );
and \U$5266 ( \5487 , \5425 , \5439 );
and \U$5267 ( \5488 , \5439 , \5454 );
and \U$5268 ( \5489 , \5425 , \5454 );
or \U$5269 ( \5490 , \5487 , \5488 , \5489 );
xor \U$5270 ( \5491 , \5486 , \5490 );
and \U$5271 ( \5492 , \5406 , \5420 );
xor \U$5272 ( \5493 , \5491 , \5492 );
xor \U$5273 ( \5494 , \5482 , \5493 );
and \U$5274 ( \5495 , \5375 , \5379 );
and \U$5275 ( \5496 , \5379 , \5381 );
and \U$5276 ( \5497 , \5375 , \5381 );
or \U$5277 ( \5498 , \5495 , \5496 , \5497 );
and \U$5278 ( \5499 , \5421 , \5455 );
and \U$5279 ( \5500 , \5455 , \5470 );
and \U$5280 ( \5501 , \5421 , \5470 );
or \U$5281 ( \5502 , \5499 , \5500 , \5501 );
xor \U$5282 ( \5503 , \5498 , \5502 );
and \U$5283 ( \5504 , \766 , \757 );
and \U$5284 ( \5505 , \786 , \755 );
nor \U$5285 ( \5506 , \5504 , \5505 );
xnor \U$5286 ( \5507 , \5506 , \764 );
and \U$5287 ( \5508 , \794 , \784 );
and \U$5288 ( \5509 , \814 , \782 );
nor \U$5289 ( \5510 , \5508 , \5509 );
xnor \U$5290 ( \5511 , \5510 , \791 );
xor \U$5291 ( \5512 , \5507 , \5511 );
and \U$5292 ( \5513 , \827 , \812 );
and \U$5293 ( \5514 , \847 , \810 );
nor \U$5294 ( \5515 , \5513 , \5514 );
xnor \U$5295 ( \5516 , \5515 , \819 );
xor \U$5296 ( \5517 , \5512 , \5516 );
and \U$5297 ( \5518 , \680 , \671 );
and \U$5298 ( \5519 , \700 , \669 );
nor \U$5299 ( \5520 , \5518 , \5519 );
xnor \U$5300 ( \5521 , \5520 , \678 );
and \U$5301 ( \5522 , \708 , \698 );
and \U$5302 ( \5523 , \728 , \696 );
nor \U$5303 ( \5524 , \5522 , \5523 );
xnor \U$5304 ( \5525 , \5524 , \705 );
xor \U$5305 ( \5526 , \5521 , \5525 );
and \U$5306 ( \5527 , \739 , \726 );
and \U$5307 ( \5528 , \759 , \724 );
nor \U$5308 ( \5529 , \5527 , \5528 );
xnor \U$5309 ( \5530 , \5529 , \733 );
xor \U$5310 ( \5531 , \5526 , \5530 );
xor \U$5311 ( \5532 , \5517 , \5531 );
and \U$5312 ( \5533 , \623 , \616 );
and \U$5313 ( \5534 , \643 , \613 );
nor \U$5314 ( \5535 , \5533 , \5534 );
xnor \U$5315 ( \5536 , \5535 , \576 );
xor \U$5316 ( \5537 , \957 , \5536 );
and \U$5317 ( \5538 , \653 , \641 );
and \U$5318 ( \5539 , \673 , \639 );
nor \U$5319 ( \5540 , \5538 , \5539 );
xnor \U$5320 ( \5541 , \5540 , \648 );
xor \U$5321 ( \5542 , \5537 , \5541 );
xor \U$5322 ( \5543 , \5532 , \5542 );
and \U$5323 ( \5544 , \5429 , \5433 );
and \U$5324 ( \5545 , \5433 , \5438 );
and \U$5325 ( \5546 , \5429 , \5438 );
or \U$5326 ( \5547 , \5544 , \5545 , \5546 );
and \U$5327 ( \5548 , \939 , \930 );
and \U$5328 ( \5549 , \952 , \928 );
nor \U$5329 ( \5550 , \5548 , \5549 );
xnor \U$5330 ( \5551 , \5550 , \937 );
nand \U$5331 ( \5552 , \960 , \948 );
xnor \U$5332 ( \5553 , \5552 , \957 );
xor \U$5333 ( \5554 , \5551 , \5553 );
xor \U$5334 ( \5555 , \5547 , \5554 );
and \U$5335 ( \5556 , \854 , \845 );
and \U$5336 ( \5557 , \874 , \843 );
nor \U$5337 ( \5558 , \5556 , \5557 );
xnor \U$5338 ( \5559 , \5558 , \852 );
and \U$5339 ( \5560 , \882 , \872 );
and \U$5340 ( \5561 , \902 , \870 );
nor \U$5341 ( \5562 , \5560 , \5561 );
xnor \U$5342 ( \5563 , \5562 , \879 );
xor \U$5343 ( \5564 , \5559 , \5563 );
and \U$5344 ( \5565 , \912 , \900 );
and \U$5345 ( \5566 , \932 , \898 );
nor \U$5346 ( \5567 , \5565 , \5566 );
xnor \U$5347 ( \5568 , \5567 , \907 );
xor \U$5348 ( \5569 , \5564 , \5568 );
xor \U$5349 ( \5570 , \5555 , \5569 );
xor \U$5350 ( \5571 , \5543 , \5570 );
and \U$5351 ( \5572 , \5410 , \5414 );
and \U$5352 ( \5573 , \5414 , \5419 );
and \U$5353 ( \5574 , \5410 , \5419 );
or \U$5354 ( \5575 , \5572 , \5573 , \5574 );
and \U$5355 ( \5576 , \5396 , \5400 );
and \U$5356 ( \5577 , \5400 , \5405 );
and \U$5357 ( \5578 , \5396 , \5405 );
or \U$5358 ( \5579 , \5576 , \5577 , \5578 );
xor \U$5359 ( \5580 , \5575 , \5579 );
and \U$5360 ( \5581 , \5444 , \5448 );
and \U$5361 ( \5582 , \5448 , \5453 );
and \U$5362 ( \5583 , \5444 , \5453 );
or \U$5363 ( \5584 , \5581 , \5582 , \5583 );
xor \U$5364 ( \5585 , \5580 , \5584 );
xor \U$5365 ( \5586 , \5571 , \5585 );
xor \U$5366 ( \5587 , \5503 , \5586 );
xor \U$5367 ( \5588 , \5494 , \5587 );
and \U$5368 ( \5589 , \5371 , \5382 );
and \U$5369 ( \5590 , \5382 , \5472 );
and \U$5370 ( \5591 , \5371 , \5472 );
or \U$5371 ( \5592 , \5589 , \5590 , \5591 );
nor \U$5372 ( \5593 , \5588 , \5592 );
nor \U$5373 ( \5594 , \5478 , \5593 );
and \U$5374 ( \5595 , \5498 , \5502 );
and \U$5375 ( \5596 , \5502 , \5586 );
and \U$5376 ( \5597 , \5498 , \5586 );
or \U$5377 ( \5598 , \5595 , \5596 , \5597 );
xor \U$5378 ( \5599 , \1532 , \1536 );
xor \U$5379 ( \5600 , \5599 , \1541 );
xor \U$5380 ( \5601 , \1584 , \1588 );
xor \U$5381 ( \5602 , \5601 , \1593 );
xor \U$5382 ( \5603 , \1565 , \1569 );
xor \U$5383 ( \5604 , \5603 , \1574 );
xor \U$5384 ( \5605 , \5602 , \5604 );
xor \U$5385 ( \5606 , \1548 , \1552 );
xor \U$5386 ( \5607 , \5606 , \1557 );
xor \U$5387 ( \5608 , \5605 , \5607 );
xor \U$5388 ( \5609 , \5600 , \5608 );
and \U$5389 ( \5610 , \5559 , \5563 );
and \U$5390 ( \5611 , \5563 , \5568 );
and \U$5391 ( \5612 , \5559 , \5568 );
or \U$5392 ( \5613 , \5610 , \5611 , \5612 );
and \U$5393 ( \5614 , \5551 , \5553 );
xor \U$5394 ( \5615 , \5613 , \5614 );
and \U$5395 ( \5616 , \960 , \950 );
and \U$5396 ( \5617 , \939 , \948 );
nor \U$5397 ( \5618 , \5616 , \5617 );
xnor \U$5398 ( \5619 , \5618 , \957 );
xor \U$5399 ( \5620 , \5615 , \5619 );
xor \U$5400 ( \5621 , \5609 , \5620 );
and \U$5401 ( \5622 , \5575 , \5579 );
and \U$5402 ( \5623 , \5579 , \5584 );
and \U$5403 ( \5624 , \5575 , \5584 );
or \U$5404 ( \5625 , \5622 , \5623 , \5624 );
and \U$5405 ( \5626 , \5547 , \5554 );
and \U$5406 ( \5627 , \5554 , \5569 );
and \U$5407 ( \5628 , \5547 , \5569 );
or \U$5408 ( \5629 , \5626 , \5627 , \5628 );
xor \U$5409 ( \5630 , \5625 , \5629 );
and \U$5410 ( \5631 , \5517 , \5531 );
and \U$5411 ( \5632 , \5531 , \5542 );
and \U$5412 ( \5633 , \5517 , \5542 );
or \U$5413 ( \5634 , \5631 , \5632 , \5633 );
xor \U$5414 ( \5635 , \5630 , \5634 );
xor \U$5415 ( \5636 , \5621 , \5635 );
xor \U$5416 ( \5637 , \5598 , \5636 );
and \U$5417 ( \5638 , \5486 , \5490 );
and \U$5418 ( \5639 , \5490 , \5492 );
and \U$5419 ( \5640 , \5486 , \5492 );
or \U$5420 ( \5641 , \5638 , \5639 , \5640 );
and \U$5421 ( \5642 , \5543 , \5570 );
and \U$5422 ( \5643 , \5570 , \5585 );
and \U$5423 ( \5644 , \5543 , \5585 );
or \U$5424 ( \5645 , \5642 , \5643 , \5644 );
xor \U$5425 ( \5646 , \5641 , \5645 );
and \U$5426 ( \5647 , \957 , \5536 );
and \U$5427 ( \5648 , \5536 , \5541 );
and \U$5428 ( \5649 , \957 , \5541 );
or \U$5429 ( \5650 , \5647 , \5648 , \5649 );
and \U$5430 ( \5651 , \5521 , \5525 );
and \U$5431 ( \5652 , \5525 , \5530 );
and \U$5432 ( \5653 , \5521 , \5530 );
or \U$5433 ( \5654 , \5651 , \5652 , \5653 );
xor \U$5434 ( \5655 , \5650 , \5654 );
and \U$5435 ( \5656 , \5507 , \5511 );
and \U$5436 ( \5657 , \5511 , \5516 );
and \U$5437 ( \5658 , \5507 , \5516 );
or \U$5438 ( \5659 , \5656 , \5657 , \5658 );
xor \U$5439 ( \5660 , \5655 , \5659 );
xor \U$5440 ( \5661 , \5646 , \5660 );
xor \U$5441 ( \5662 , \5637 , \5661 );
and \U$5442 ( \5663 , \5482 , \5493 );
and \U$5443 ( \5664 , \5493 , \5587 );
and \U$5444 ( \5665 , \5482 , \5587 );
or \U$5445 ( \5666 , \5663 , \5664 , \5665 );
nor \U$5446 ( \5667 , \5662 , \5666 );
and \U$5447 ( \5668 , \5625 , \5629 );
and \U$5448 ( \5669 , \5629 , \5634 );
and \U$5449 ( \5670 , \5625 , \5634 );
or \U$5450 ( \5671 , \5668 , \5669 , \5670 );
and \U$5451 ( \5672 , \5600 , \5608 );
and \U$5452 ( \5673 , \5608 , \5620 );
and \U$5453 ( \5674 , \5600 , \5620 );
or \U$5454 ( \5675 , \5672 , \5673 , \5674 );
xor \U$5455 ( \5676 , \5671 , \5675 );
xor \U$5456 ( \5677 , \1607 , \1609 );
xor \U$5457 ( \5678 , \5677 , \1612 );
xor \U$5458 ( \5679 , \1596 , \1598 );
xor \U$5459 ( \5680 , \5679 , \1601 );
xor \U$5460 ( \5681 , \5678 , \5680 );
xor \U$5461 ( \5682 , \1544 , \1560 );
xor \U$5462 ( \5683 , \5682 , \1577 );
xor \U$5463 ( \5684 , \5681 , \5683 );
xor \U$5464 ( \5685 , \5676 , \5684 );
and \U$5465 ( \5686 , \5641 , \5645 );
and \U$5466 ( \5687 , \5645 , \5660 );
and \U$5467 ( \5688 , \5641 , \5660 );
or \U$5468 ( \5689 , \5686 , \5687 , \5688 );
and \U$5469 ( \5690 , \5621 , \5635 );
xor \U$5470 ( \5691 , \5689 , \5690 );
and \U$5471 ( \5692 , \5650 , \5654 );
and \U$5472 ( \5693 , \5654 , \5659 );
and \U$5473 ( \5694 , \5650 , \5659 );
or \U$5474 ( \5695 , \5692 , \5693 , \5694 );
and \U$5475 ( \5696 , \5613 , \5614 );
and \U$5476 ( \5697 , \5614 , \5619 );
and \U$5477 ( \5698 , \5613 , \5619 );
or \U$5478 ( \5699 , \5696 , \5697 , \5698 );
xor \U$5479 ( \5700 , \5695 , \5699 );
and \U$5480 ( \5701 , \5602 , \5604 );
and \U$5481 ( \5702 , \5604 , \5607 );
and \U$5482 ( \5703 , \5602 , \5607 );
or \U$5483 ( \5704 , \5701 , \5702 , \5703 );
xor \U$5484 ( \5705 , \5700 , \5704 );
xor \U$5485 ( \5706 , \5691 , \5705 );
xor \U$5486 ( \5707 , \5685 , \5706 );
and \U$5487 ( \5708 , \5598 , \5636 );
and \U$5488 ( \5709 , \5636 , \5661 );
and \U$5489 ( \5710 , \5598 , \5661 );
or \U$5490 ( \5711 , \5708 , \5709 , \5710 );
nor \U$5491 ( \5712 , \5707 , \5711 );
nor \U$5492 ( \5713 , \5667 , \5712 );
nand \U$5493 ( \5714 , \5594 , \5713 );
and \U$5494 ( \5715 , \5689 , \5690 );
and \U$5495 ( \5716 , \5690 , \5705 );
and \U$5496 ( \5717 , \5689 , \5705 );
or \U$5497 ( \5718 , \5715 , \5716 , \5717 );
and \U$5498 ( \5719 , \5671 , \5675 );
and \U$5499 ( \5720 , \5675 , \5684 );
and \U$5500 ( \5721 , \5671 , \5684 );
or \U$5501 ( \5722 , \5719 , \5720 , \5721 );
xor \U$5502 ( \5723 , \652 , \737 );
xor \U$5503 ( \5724 , \5723 , \823 );
xor \U$5504 ( \5725 , \1620 , \1622 );
xor \U$5505 ( \5726 , \5725 , \1625 );
xor \U$5506 ( \5727 , \5724 , \5726 );
xor \U$5507 ( \5728 , \1580 , \1604 );
xor \U$5508 ( \5729 , \5728 , \1615 );
xor \U$5509 ( \5730 , \5727 , \5729 );
xor \U$5510 ( \5731 , \5722 , \5730 );
and \U$5511 ( \5732 , \5695 , \5699 );
and \U$5512 ( \5733 , \5699 , \5704 );
and \U$5513 ( \5734 , \5695 , \5704 );
or \U$5514 ( \5735 , \5732 , \5733 , \5734 );
and \U$5515 ( \5736 , \5678 , \5680 );
and \U$5516 ( \5737 , \5680 , \5683 );
and \U$5517 ( \5738 , \5678 , \5683 );
or \U$5518 ( \5739 , \5736 , \5737 , \5738 );
xor \U$5519 ( \5740 , \5735 , \5739 );
xor \U$5520 ( \5741 , \911 , \966 );
xor \U$5521 ( \5742 , \5741 , \971 );
xor \U$5522 ( \5743 , \5740 , \5742 );
xor \U$5523 ( \5744 , \5731 , \5743 );
xor \U$5524 ( \5745 , \5718 , \5744 );
and \U$5525 ( \5746 , \5685 , \5706 );
nor \U$5526 ( \5747 , \5745 , \5746 );
and \U$5527 ( \5748 , \5722 , \5730 );
and \U$5528 ( \5749 , \5730 , \5743 );
and \U$5529 ( \5750 , \5722 , \5743 );
or \U$5530 ( \5751 , \5748 , \5749 , \5750 );
xor \U$5531 ( \5752 , \826 , \974 );
xor \U$5532 ( \5753 , \5752 , \1014 );
xor \U$5533 ( \5754 , \1618 , \1628 );
xor \U$5534 ( \5755 , \5754 , \1631 );
xor \U$5535 ( \5756 , \5753 , \5755 );
xor \U$5536 ( \5757 , \5751 , \5756 );
and \U$5537 ( \5758 , \5735 , \5739 );
and \U$5538 ( \5759 , \5739 , \5742 );
and \U$5539 ( \5760 , \5735 , \5742 );
or \U$5540 ( \5761 , \5758 , \5759 , \5760 );
and \U$5541 ( \5762 , \5724 , \5726 );
and \U$5542 ( \5763 , \5726 , \5729 );
and \U$5543 ( \5764 , \5724 , \5729 );
or \U$5544 ( \5765 , \5762 , \5763 , \5764 );
xor \U$5545 ( \5766 , \5761 , \5765 );
xor \U$5546 ( \5767 , \1029 , \1073 );
xor \U$5547 ( \5768 , \5767 , \1097 );
xor \U$5548 ( \5769 , \5766 , \5768 );
xor \U$5549 ( \5770 , \5757 , \5769 );
and \U$5550 ( \5771 , \5718 , \5744 );
nor \U$5551 ( \5772 , \5770 , \5771 );
nor \U$5552 ( \5773 , \5747 , \5772 );
and \U$5553 ( \5774 , \5761 , \5765 );
and \U$5554 ( \5775 , \5765 , \5768 );
and \U$5555 ( \5776 , \5761 , \5768 );
or \U$5556 ( \5777 , \5774 , \5775 , \5776 );
and \U$5557 ( \5778 , \5753 , \5755 );
xor \U$5558 ( \5779 , \5777 , \5778 );
xor \U$5559 ( \5780 , \1634 , \1635 );
xor \U$5560 ( \5781 , \5780 , \1638 );
xor \U$5561 ( \5782 , \5779 , \5781 );
and \U$5562 ( \5783 , \5751 , \5756 );
and \U$5563 ( \5784 , \5756 , \5769 );
and \U$5564 ( \5785 , \5751 , \5769 );
or \U$5565 ( \5786 , \5783 , \5784 , \5785 );
nor \U$5566 ( \5787 , \5782 , \5786 );
xor \U$5567 ( \5788 , \1641 , \1642 );
xor \U$5568 ( \5789 , \5788 , \1645 );
and \U$5569 ( \5790 , \5777 , \5778 );
and \U$5570 ( \5791 , \5778 , \5781 );
and \U$5571 ( \5792 , \5777 , \5781 );
or \U$5572 ( \5793 , \5790 , \5791 , \5792 );
nor \U$5573 ( \5794 , \5789 , \5793 );
nor \U$5574 ( \5795 , \5787 , \5794 );
nand \U$5575 ( \5796 , \5773 , \5795 );
nor \U$5576 ( \5797 , \5714 , \5796 );
nand \U$5577 ( \5798 , \5367 , \5797 );
and \U$5578 ( \5799 , \902 , \616 );
and \U$5579 ( \5800 , \854 , \613 );
nor \U$5580 ( \5801 , \5799 , \5800 );
xnor \U$5581 ( \5802 , \5801 , \576 );
and \U$5582 ( \5803 , \932 , \641 );
and \U$5583 ( \5804 , \882 , \639 );
nor \U$5584 ( \5805 , \5803 , \5804 );
xnor \U$5585 ( \5806 , \5805 , \648 );
xor \U$5586 ( \5807 , \5802 , \5806 );
and \U$5587 ( \5808 , \952 , \671 );
and \U$5588 ( \5809 , \912 , \669 );
nor \U$5589 ( \5810 , \5808 , \5809 );
xnor \U$5590 ( \5811 , \5810 , \678 );
xor \U$5591 ( \5812 , \5807 , \5811 );
and \U$5592 ( \5813 , \882 , \616 );
and \U$5593 ( \5814 , \902 , \613 );
nor \U$5594 ( \5815 , \5813 , \5814 );
xnor \U$5595 ( \5816 , \5815 , \576 );
and \U$5596 ( \5817 , \705 , \5816 );
and \U$5597 ( \5818 , \912 , \641 );
and \U$5598 ( \5819 , \932 , \639 );
nor \U$5599 ( \5820 , \5818 , \5819 );
xnor \U$5600 ( \5821 , \5820 , \648 );
and \U$5601 ( \5822 , \5816 , \5821 );
and \U$5602 ( \5823 , \705 , \5821 );
or \U$5603 ( \5824 , \5817 , \5822 , \5823 );
and \U$5604 ( \5825 , \939 , \671 );
and \U$5605 ( \5826 , \952 , \669 );
nor \U$5606 ( \5827 , \5825 , \5826 );
xnor \U$5607 ( \5828 , \5827 , \678 );
nand \U$5608 ( \5829 , \960 , \696 );
xnor \U$5609 ( \5830 , \5829 , \705 );
and \U$5610 ( \5831 , \5828 , \5830 );
xor \U$5611 ( \5832 , \5824 , \5831 );
and \U$5612 ( \5833 , \960 , \698 );
and \U$5613 ( \5834 , \939 , \696 );
nor \U$5614 ( \5835 , \5833 , \5834 );
xnor \U$5615 ( \5836 , \5835 , \705 );
xor \U$5616 ( \5837 , \5832 , \5836 );
xor \U$5617 ( \5838 , \5812 , \5837 );
and \U$5618 ( \5839 , \932 , \616 );
and \U$5619 ( \5840 , \882 , \613 );
nor \U$5620 ( \5841 , \5839 , \5840 );
xnor \U$5621 ( \5842 , \5841 , \576 );
and \U$5622 ( \5843 , \952 , \641 );
and \U$5623 ( \5844 , \912 , \639 );
nor \U$5624 ( \5845 , \5843 , \5844 );
xnor \U$5625 ( \5846 , \5845 , \648 );
and \U$5626 ( \5847 , \5842 , \5846 );
and \U$5627 ( \5848 , \960 , \671 );
and \U$5628 ( \5849 , \939 , \669 );
nor \U$5629 ( \5850 , \5848 , \5849 );
xnor \U$5630 ( \5851 , \5850 , \678 );
and \U$5631 ( \5852 , \5846 , \5851 );
and \U$5632 ( \5853 , \5842 , \5851 );
or \U$5633 ( \5854 , \5847 , \5852 , \5853 );
xor \U$5634 ( \5855 , \5828 , \5830 );
and \U$5635 ( \5856 , \5854 , \5855 );
xor \U$5636 ( \5857 , \705 , \5816 );
xor \U$5637 ( \5858 , \5857 , \5821 );
and \U$5638 ( \5859 , \5855 , \5858 );
and \U$5639 ( \5860 , \5854 , \5858 );
or \U$5640 ( \5861 , \5856 , \5859 , \5860 );
nor \U$5641 ( \5862 , \5838 , \5861 );
and \U$5642 ( \5863 , \5824 , \5831 );
and \U$5643 ( \5864 , \5831 , \5836 );
and \U$5644 ( \5865 , \5824 , \5836 );
or \U$5645 ( \5866 , \5863 , \5864 , \5865 );
and \U$5646 ( \5867 , \5802 , \5806 );
and \U$5647 ( \5868 , \5806 , \5811 );
and \U$5648 ( \5869 , \5802 , \5811 );
or \U$5649 ( \5870 , \5867 , \5868 , \5869 );
and \U$5650 ( \5871 , \912 , \671 );
and \U$5651 ( \5872 , \932 , \669 );
nor \U$5652 ( \5873 , \5871 , \5872 );
xnor \U$5653 ( \5874 , \5873 , \678 );
and \U$5654 ( \5875 , \939 , \698 );
and \U$5655 ( \5876 , \952 , \696 );
nor \U$5656 ( \5877 , \5875 , \5876 );
xnor \U$5657 ( \5878 , \5877 , \705 );
xor \U$5658 ( \5879 , \5874 , \5878 );
nand \U$5659 ( \5880 , \960 , \724 );
xnor \U$5660 ( \5881 , \5880 , \733 );
xor \U$5661 ( \5882 , \5879 , \5881 );
xor \U$5662 ( \5883 , \5870 , \5882 );
and \U$5663 ( \5884 , \854 , \616 );
and \U$5664 ( \5885 , \874 , \613 );
nor \U$5665 ( \5886 , \5884 , \5885 );
xnor \U$5666 ( \5887 , \5886 , \576 );
xor \U$5667 ( \5888 , \733 , \5887 );
and \U$5668 ( \5889 , \882 , \641 );
and \U$5669 ( \5890 , \902 , \639 );
nor \U$5670 ( \5891 , \5889 , \5890 );
xnor \U$5671 ( \5892 , \5891 , \648 );
xor \U$5672 ( \5893 , \5888 , \5892 );
xor \U$5673 ( \5894 , \5883 , \5893 );
xor \U$5674 ( \5895 , \5866 , \5894 );
and \U$5675 ( \5896 , \5812 , \5837 );
nor \U$5676 ( \5897 , \5895 , \5896 );
nor \U$5677 ( \5898 , \5862 , \5897 );
and \U$5678 ( \5899 , \5870 , \5882 );
and \U$5679 ( \5900 , \5882 , \5893 );
and \U$5680 ( \5901 , \5870 , \5893 );
or \U$5681 ( \5902 , \5899 , \5900 , \5901 );
and \U$5682 ( \5903 , \960 , \726 );
and \U$5683 ( \5904 , \939 , \724 );
nor \U$5684 ( \5905 , \5903 , \5904 );
xnor \U$5685 ( \5906 , \5905 , \733 );
and \U$5686 ( \5907 , \874 , \616 );
and \U$5687 ( \5908 , \827 , \613 );
nor \U$5688 ( \5909 , \5907 , \5908 );
xnor \U$5689 ( \5910 , \5909 , \576 );
and \U$5690 ( \5911 , \902 , \641 );
and \U$5691 ( \5912 , \854 , \639 );
nor \U$5692 ( \5913 , \5911 , \5912 );
xnor \U$5693 ( \5914 , \5913 , \648 );
xor \U$5694 ( \5915 , \5910 , \5914 );
and \U$5695 ( \5916 , \932 , \671 );
and \U$5696 ( \5917 , \882 , \669 );
nor \U$5697 ( \5918 , \5916 , \5917 );
xnor \U$5698 ( \5919 , \5918 , \678 );
xor \U$5699 ( \5920 , \5915 , \5919 );
xor \U$5700 ( \5921 , \5906 , \5920 );
xor \U$5701 ( \5922 , \5902 , \5921 );
and \U$5702 ( \5923 , \733 , \5887 );
and \U$5703 ( \5924 , \5887 , \5892 );
and \U$5704 ( \5925 , \733 , \5892 );
or \U$5705 ( \5926 , \5923 , \5924 , \5925 );
and \U$5706 ( \5927 , \5874 , \5878 );
and \U$5707 ( \5928 , \5878 , \5881 );
and \U$5708 ( \5929 , \5874 , \5881 );
or \U$5709 ( \5930 , \5927 , \5928 , \5929 );
xor \U$5710 ( \5931 , \5926 , \5930 );
and \U$5711 ( \5932 , \952 , \698 );
and \U$5712 ( \5933 , \912 , \696 );
nor \U$5713 ( \5934 , \5932 , \5933 );
xnor \U$5714 ( \5935 , \5934 , \705 );
xor \U$5715 ( \5936 , \5931 , \5935 );
xor \U$5716 ( \5937 , \5922 , \5936 );
and \U$5717 ( \5938 , \5866 , \5894 );
nor \U$5718 ( \5939 , \5937 , \5938 );
and \U$5719 ( \5940 , \5910 , \5914 );
and \U$5720 ( \5941 , \5914 , \5919 );
and \U$5721 ( \5942 , \5910 , \5919 );
or \U$5722 ( \5943 , \5940 , \5941 , \5942 );
nand \U$5723 ( \5944 , \960 , \755 );
xnor \U$5724 ( \5945 , \5944 , \764 );
xor \U$5725 ( \5946 , \5943 , \5945 );
and \U$5726 ( \5947 , \882 , \671 );
and \U$5727 ( \5948 , \902 , \669 );
nor \U$5728 ( \5949 , \5947 , \5948 );
xnor \U$5729 ( \5950 , \5949 , \678 );
and \U$5730 ( \5951 , \912 , \698 );
and \U$5731 ( \5952 , \932 , \696 );
nor \U$5732 ( \5953 , \5951 , \5952 );
xnor \U$5733 ( \5954 , \5953 , \705 );
xor \U$5734 ( \5955 , \5950 , \5954 );
and \U$5735 ( \5956 , \939 , \726 );
and \U$5736 ( \5957 , \952 , \724 );
nor \U$5737 ( \5958 , \5956 , \5957 );
xnor \U$5738 ( \5959 , \5958 , \733 );
xor \U$5739 ( \5960 , \5955 , \5959 );
xor \U$5740 ( \5961 , \5946 , \5960 );
and \U$5741 ( \5962 , \5926 , \5930 );
and \U$5742 ( \5963 , \5930 , \5935 );
and \U$5743 ( \5964 , \5926 , \5935 );
or \U$5744 ( \5965 , \5962 , \5963 , \5964 );
and \U$5745 ( \5966 , \5906 , \5920 );
xor \U$5746 ( \5967 , \5965 , \5966 );
and \U$5747 ( \5968 , \827 , \616 );
and \U$5748 ( \5969 , \847 , \613 );
nor \U$5749 ( \5970 , \5968 , \5969 );
xnor \U$5750 ( \5971 , \5970 , \576 );
xor \U$5751 ( \5972 , \764 , \5971 );
and \U$5752 ( \5973 , \854 , \641 );
and \U$5753 ( \5974 , \874 , \639 );
nor \U$5754 ( \5975 , \5973 , \5974 );
xnor \U$5755 ( \5976 , \5975 , \648 );
xor \U$5756 ( \5977 , \5972 , \5976 );
xor \U$5757 ( \5978 , \5967 , \5977 );
xor \U$5758 ( \5979 , \5961 , \5978 );
and \U$5759 ( \5980 , \5902 , \5921 );
and \U$5760 ( \5981 , \5921 , \5936 );
and \U$5761 ( \5982 , \5902 , \5936 );
or \U$5762 ( \5983 , \5980 , \5981 , \5982 );
nor \U$5763 ( \5984 , \5979 , \5983 );
nor \U$5764 ( \5985 , \5939 , \5984 );
nand \U$5765 ( \5986 , \5898 , \5985 );
and \U$5766 ( \5987 , \5965 , \5966 );
and \U$5767 ( \5988 , \5966 , \5977 );
and \U$5768 ( \5989 , \5965 , \5977 );
or \U$5769 ( \5990 , \5987 , \5988 , \5989 );
and \U$5770 ( \5991 , \5943 , \5945 );
and \U$5771 ( \5992 , \5945 , \5960 );
and \U$5772 ( \5993 , \5943 , \5960 );
or \U$5773 ( \5994 , \5991 , \5992 , \5993 );
xor \U$5774 ( \5995 , \4663 , \4667 );
xor \U$5775 ( \5996 , \5995 , \4672 );
xor \U$5776 ( \5997 , \5994 , \5996 );
and \U$5777 ( \5998 , \764 , \5971 );
and \U$5778 ( \5999 , \5971 , \5976 );
and \U$5779 ( \6000 , \764 , \5976 );
or \U$5780 ( \6001 , \5998 , \5999 , \6000 );
and \U$5781 ( \6002 , \5950 , \5954 );
and \U$5782 ( \6003 , \5954 , \5959 );
and \U$5783 ( \6004 , \5950 , \5959 );
or \U$5784 ( \6005 , \6002 , \6003 , \6004 );
xor \U$5785 ( \6006 , \6001 , \6005 );
xor \U$5786 ( \6007 , \4679 , \4683 );
xor \U$5787 ( \6008 , \6007 , \4688 );
xor \U$5788 ( \6009 , \6006 , \6008 );
xor \U$5789 ( \6010 , \5997 , \6009 );
xor \U$5790 ( \6011 , \5990 , \6010 );
and \U$5791 ( \6012 , \5961 , \5978 );
nor \U$5792 ( \6013 , \6011 , \6012 );
and \U$5793 ( \6014 , \5994 , \5996 );
and \U$5794 ( \6015 , \5996 , \6009 );
and \U$5795 ( \6016 , \5994 , \6009 );
or \U$5796 ( \6017 , \6014 , \6015 , \6016 );
and \U$5797 ( \6018 , \6001 , \6005 );
and \U$5798 ( \6019 , \6005 , \6008 );
and \U$5799 ( \6020 , \6001 , \6008 );
or \U$5800 ( \6021 , \6018 , \6019 , \6020 );
xor \U$5801 ( \6022 , \4701 , \4703 );
xor \U$5802 ( \6023 , \6022 , \4706 );
xor \U$5803 ( \6024 , \6021 , \6023 );
xor \U$5804 ( \6025 , \4675 , \4691 );
xor \U$5805 ( \6026 , \6025 , \4696 );
xor \U$5806 ( \6027 , \6024 , \6026 );
xor \U$5807 ( \6028 , \6017 , \6027 );
and \U$5808 ( \6029 , \5990 , \6010 );
nor \U$5809 ( \6030 , \6028 , \6029 );
nor \U$5810 ( \6031 , \6013 , \6030 );
and \U$5811 ( \6032 , \6021 , \6023 );
and \U$5812 ( \6033 , \6023 , \6026 );
and \U$5813 ( \6034 , \6021 , \6026 );
or \U$5814 ( \6035 , \6032 , \6033 , \6034 );
xor \U$5815 ( \6036 , \4717 , \4719 );
xor \U$5816 ( \6037 , \6035 , \6036 );
xor \U$5817 ( \6038 , \4699 , \4709 );
xor \U$5818 ( \6039 , \6038 , \4712 );
xor \U$5819 ( \6040 , \6037 , \6039 );
and \U$5820 ( \6041 , \6017 , \6027 );
nor \U$5821 ( \6042 , \6040 , \6041 );
xor \U$5822 ( \6043 , \4715 , \4720 );
xor \U$5823 ( \6044 , \6043 , \4723 );
and \U$5824 ( \6045 , \6035 , \6036 );
and \U$5825 ( \6046 , \6036 , \6039 );
and \U$5826 ( \6047 , \6035 , \6039 );
or \U$5827 ( \6048 , \6045 , \6046 , \6047 );
nor \U$5828 ( \6049 , \6044 , \6048 );
nor \U$5829 ( \6050 , \6042 , \6049 );
nand \U$5830 ( \6051 , \6031 , \6050 );
nor \U$5831 ( \6052 , \5986 , \6051 );
and \U$5832 ( \6053 , \952 , \616 );
and \U$5833 ( \6054 , \912 , \613 );
nor \U$5834 ( \6055 , \6053 , \6054 );
xnor \U$5835 ( \6056 , \6055 , \576 );
and \U$5836 ( \6057 , \960 , \641 );
and \U$5837 ( \6058 , \939 , \639 );
nor \U$5838 ( \6059 , \6057 , \6058 );
xnor \U$5839 ( \6060 , \6059 , \648 );
xor \U$5840 ( \6061 , \6056 , \6060 );
and \U$5841 ( \6062 , \939 , \616 );
and \U$5842 ( \6063 , \952 , \613 );
nor \U$5843 ( \6064 , \6062 , \6063 );
xnor \U$5844 ( \6065 , \6064 , \576 );
and \U$5845 ( \6066 , \6065 , \648 );
nor \U$5846 ( \6067 , \6061 , \6066 );
nand \U$5847 ( \6068 , \960 , \669 );
xnor \U$5848 ( \6069 , \6068 , \678 );
and \U$5849 ( \6070 , \912 , \616 );
and \U$5850 ( \6071 , \932 , \613 );
nor \U$5851 ( \6072 , \6070 , \6071 );
xnor \U$5852 ( \6073 , \6072 , \576 );
xor \U$5853 ( \6074 , \678 , \6073 );
and \U$5854 ( \6075 , \939 , \641 );
and \U$5855 ( \6076 , \952 , \639 );
nor \U$5856 ( \6077 , \6075 , \6076 );
xnor \U$5857 ( \6078 , \6077 , \648 );
xor \U$5858 ( \6079 , \6074 , \6078 );
xor \U$5859 ( \6080 , \6069 , \6079 );
and \U$5860 ( \6081 , \6056 , \6060 );
nor \U$5861 ( \6082 , \6080 , \6081 );
nor \U$5862 ( \6083 , \6067 , \6082 );
and \U$5863 ( \6084 , \678 , \6073 );
and \U$5864 ( \6085 , \6073 , \6078 );
and \U$5865 ( \6086 , \678 , \6078 );
or \U$5866 ( \6087 , \6084 , \6085 , \6086 );
xor \U$5867 ( \6088 , \5842 , \5846 );
xor \U$5868 ( \6089 , \6088 , \5851 );
xor \U$5869 ( \6090 , \6087 , \6089 );
and \U$5870 ( \6091 , \6069 , \6079 );
nor \U$5871 ( \6092 , \6090 , \6091 );
xor \U$5872 ( \6093 , \5854 , \5855 );
xor \U$5873 ( \6094 , \6093 , \5858 );
and \U$5874 ( \6095 , \6087 , \6089 );
nor \U$5875 ( \6096 , \6094 , \6095 );
nor \U$5876 ( \6097 , \6092 , \6096 );
nand \U$5877 ( \6098 , \6083 , \6097 );
xor \U$5878 ( \6099 , \6065 , \648 );
nand \U$5879 ( \6100 , \960 , \639 );
xnor \U$5880 ( \6101 , \6100 , \648 );
nor \U$5881 ( \6102 , \6099 , \6101 );
and \U$5882 ( \6103 , \960 , \616 );
and \U$5883 ( \6104 , \939 , \613 );
nor \U$5884 ( \6105 , \6103 , \6104 );
xnor \U$5885 ( \6106 , \6105 , \576 );
nand \U$5886 ( \6107 , \960 , \613 );
xnor \U$5887 ( \6108 , \6107 , \576 );
and \U$5888 ( \6109 , \6108 , \576 );
nand \U$5889 ( \6110 , \6106 , \6109 );
or \U$5890 ( \6111 , \6102 , \6110 );
nand \U$5891 ( \6112 , \6099 , \6101 );
nand \U$5892 ( \6113 , \6111 , \6112 );
not \U$5893 ( \6114 , \6113 );
or \U$5894 ( \6115 , \6098 , \6114 );
nand \U$5895 ( \6116 , \6061 , \6066 );
or \U$5896 ( \6117 , \6082 , \6116 );
nand \U$5897 ( \6118 , \6080 , \6081 );
nand \U$5898 ( \6119 , \6117 , \6118 );
and \U$5899 ( \6120 , \6097 , \6119 );
nand \U$5900 ( \6121 , \6090 , \6091 );
or \U$5901 ( \6122 , \6096 , \6121 );
nand \U$5902 ( \6123 , \6094 , \6095 );
nand \U$5903 ( \6124 , \6122 , \6123 );
nor \U$5904 ( \6125 , \6120 , \6124 );
nand \U$5905 ( \6126 , \6115 , \6125 );
and \U$5906 ( \6127 , \6052 , \6126 );
nand \U$5907 ( \6128 , \5838 , \5861 );
or \U$5908 ( \6129 , \5897 , \6128 );
nand \U$5909 ( \6130 , \5895 , \5896 );
nand \U$5910 ( \6131 , \6129 , \6130 );
and \U$5911 ( \6132 , \5985 , \6131 );
nand \U$5912 ( \6133 , \5937 , \5938 );
or \U$5913 ( \6134 , \5984 , \6133 );
nand \U$5914 ( \6135 , \5979 , \5983 );
nand \U$5915 ( \6136 , \6134 , \6135 );
nor \U$5916 ( \6137 , \6132 , \6136 );
or \U$5917 ( \6138 , \6051 , \6137 );
nand \U$5918 ( \6139 , \6011 , \6012 );
or \U$5919 ( \6140 , \6030 , \6139 );
nand \U$5920 ( \6141 , \6028 , \6029 );
nand \U$5921 ( \6142 , \6140 , \6141 );
and \U$5922 ( \6143 , \6050 , \6142 );
nand \U$5923 ( \6144 , \6040 , \6041 );
or \U$5924 ( \6145 , \6049 , \6144 );
nand \U$5925 ( \6146 , \6044 , \6048 );
nand \U$5926 ( \6147 , \6145 , \6146 );
nor \U$5927 ( \6148 , \6143 , \6147 );
nand \U$5928 ( \6149 , \6138 , \6148 );
nor \U$5929 ( \6150 , \6127 , \6149 );
or \U$5930 ( \6151 , \5798 , \6150 );
nand \U$5931 ( \6152 , \4659 , \4726 );
or \U$5932 ( \6153 , \4802 , \6152 );
nand \U$5933 ( \6154 , \4797 , \4801 );
nand \U$5934 ( \6155 , \6153 , \6154 );
and \U$5935 ( \6156 , \4970 , \6155 );
nand \U$5936 ( \6157 , \4879 , \4883 );
or \U$5937 ( \6158 , \4969 , \6157 );
nand \U$5938 ( \6159 , \4967 , \4968 );
nand \U$5939 ( \6160 , \6158 , \6159 );
nor \U$5940 ( \6161 , \6156 , \6160 );
or \U$5941 ( \6162 , \5366 , \6161 );
nand \U$5942 ( \6163 , \5060 , \5061 );
or \U$5943 ( \6164 , \5157 , \6163 );
nand \U$5944 ( \6165 , \5152 , \5156 );
nand \U$5945 ( \6166 , \6164 , \6165 );
and \U$5946 ( \6167 , \5365 , \6166 );
nand \U$5947 ( \6168 , \5254 , \5258 );
or \U$5948 ( \6169 , \5364 , \6168 );
nand \U$5949 ( \6170 , \5359 , \5363 );
nand \U$5950 ( \6171 , \6169 , \6170 );
nor \U$5951 ( \6172 , \6167 , \6171 );
nand \U$5952 ( \6173 , \6162 , \6172 );
and \U$5953 ( \6174 , \5797 , \6173 );
nand \U$5954 ( \6175 , \5473 , \5477 );
or \U$5955 ( \6176 , \5593 , \6175 );
nand \U$5956 ( \6177 , \5588 , \5592 );
nand \U$5957 ( \6178 , \6176 , \6177 );
and \U$5958 ( \6179 , \5713 , \6178 );
nand \U$5959 ( \6180 , \5662 , \5666 );
or \U$5960 ( \6181 , \5712 , \6180 );
nand \U$5961 ( \6182 , \5707 , \5711 );
nand \U$5962 ( \6183 , \6181 , \6182 );
nor \U$5963 ( \6184 , \6179 , \6183 );
or \U$5964 ( \6185 , \5796 , \6184 );
nand \U$5965 ( \6186 , \5745 , \5746 );
or \U$5966 ( \6187 , \5772 , \6186 );
nand \U$5967 ( \6188 , \5770 , \5771 );
nand \U$5968 ( \6189 , \6187 , \6188 );
and \U$5969 ( \6190 , \5795 , \6189 );
nand \U$5970 ( \6191 , \5782 , \5786 );
or \U$5971 ( \6192 , \5794 , \6191 );
nand \U$5972 ( \6193 , \5789 , \5793 );
nand \U$5973 ( \6194 , \6192 , \6193 );
nor \U$5974 ( \6195 , \6190 , \6194 );
nand \U$5975 ( \6196 , \6185 , \6195 );
nor \U$5976 ( \6197 , \6174 , \6196 );
nand \U$5977 ( \6198 , \6151 , \6197 );
and \U$5978 ( \6199 , \4486 , \6198 );
nand \U$5979 ( \6200 , \1528 , \1648 );
or \U$5980 ( \6201 , \1802 , \6200 );
nand \U$5981 ( \6202 , \1797 , \1801 );
nand \U$5982 ( \6203 , \6201 , \6202 );
and \U$5983 ( \6204 , \2111 , \6203 );
nand \U$5984 ( \6205 , \1952 , \1956 );
or \U$5985 ( \6206 , \2110 , \6205 );
nand \U$5986 ( \6207 , \2105 , \2109 );
nand \U$5987 ( \6208 , \6206 , \6207 );
nor \U$5988 ( \6209 , \6204 , \6208 );
or \U$5989 ( \6210 , \2690 , \6209 );
nand \U$5990 ( \6211 , \2259 , \2263 );
or \U$5991 ( \6212 , \2411 , \6211 );
nand \U$5992 ( \6213 , \2406 , \2410 );
nand \U$5993 ( \6214 , \6212 , \6213 );
and \U$5994 ( \6215 , \2689 , \6214 );
nand \U$5995 ( \6216 , \2546 , \2550 );
or \U$5996 ( \6217 , \2688 , \6216 );
nand \U$5997 ( \6218 , \2683 , \2687 );
nand \U$5998 ( \6219 , \6217 , \6218 );
nor \U$5999 ( \6220 , \6215 , \6219 );
nand \U$6000 ( \6221 , \6210 , \6220 );
and \U$6001 ( \6222 , \3609 , \6221 );
nand \U$6002 ( \6223 , \2815 , \2819 );
or \U$6003 ( \6224 , \2946 , \6223 );
nand \U$6004 ( \6225 , \2941 , \2945 );
nand \U$6005 ( \6226 , \6224 , \6225 );
and \U$6006 ( \6227 , \3186 , \6226 );
nand \U$6007 ( \6228 , \3064 , \3068 );
or \U$6008 ( \6229 , \3185 , \6228 );
nand \U$6009 ( \6230 , \3183 , \3184 );
nand \U$6010 ( \6231 , \6229 , \6230 );
nor \U$6011 ( \6232 , \6227 , \6231 );
or \U$6012 ( \6233 , \3608 , \6232 );
nand \U$6013 ( \6234 , \3294 , \3298 );
or \U$6014 ( \6235 , \3405 , \6234 );
nand \U$6015 ( \6236 , \3403 , \3404 );
nand \U$6016 ( \6237 , \6235 , \6236 );
and \U$6017 ( \6238 , \3607 , \6237 );
nand \U$6018 ( \6239 , \3505 , \3506 );
or \U$6019 ( \6240 , \3606 , \6239 );
nand \U$6020 ( \6241 , \3604 , \3605 );
nand \U$6021 ( \6242 , \6240 , \6241 );
nor \U$6022 ( \6243 , \6238 , \6242 );
nand \U$6023 ( \6244 , \6233 , \6243 );
nor \U$6024 ( \6245 , \6222 , \6244 );
or \U$6025 ( \6246 , \4485 , \6245 );
nand \U$6026 ( \6247 , \3699 , \3700 );
or \U$6027 ( \6248 , \3790 , \6247 );
nand \U$6028 ( \6249 , \3788 , \3789 );
nand \U$6029 ( \6250 , \6248 , \6249 );
and \U$6030 ( \6251 , \3952 , \6250 );
nand \U$6031 ( \6252 , \3870 , \3871 );
or \U$6032 ( \6253 , \3951 , \6252 );
nand \U$6033 ( \6254 , \3949 , \3950 );
nand \U$6034 ( \6255 , \6253 , \6254 );
nor \U$6035 ( \6256 , \6251 , \6255 );
or \U$6036 ( \6257 , \4216 , \6256 );
nand \U$6037 ( \6258 , \4020 , \4024 );
or \U$6038 ( \6259 , \4090 , \6258 );
nand \U$6039 ( \6260 , \4088 , \4089 );
nand \U$6040 ( \6261 , \6259 , \6260 );
and \U$6041 ( \6262 , \4215 , \6261 );
nand \U$6042 ( \6263 , \4153 , \4154 );
or \U$6043 ( \6264 , \4214 , \6263 );
nand \U$6044 ( \6265 , \4212 , \4213 );
nand \U$6045 ( \6266 , \6264 , \6265 );
nor \U$6046 ( \6267 , \6262 , \6266 );
nand \U$6047 ( \6268 , \6257 , \6267 );
and \U$6048 ( \6269 , \4484 , \6268 );
nand \U$6049 ( \6270 , \4266 , \4267 );
or \U$6050 ( \6271 , \4317 , \6270 );
nand \U$6051 ( \6272 , \4315 , \4316 );
nand \U$6052 ( \6273 , \6271 , \6272 );
and \U$6053 ( \6274 , \4396 , \6273 );
nand \U$6054 ( \6275 , \4355 , \4359 );
or \U$6055 ( \6276 , \4395 , \6275 );
nand \U$6056 ( \6277 , \4393 , \4394 );
nand \U$6057 ( \6278 , \6276 , \6277 );
nor \U$6058 ( \6279 , \6274 , \6278 );
or \U$6059 ( \6280 , \4483 , \6279 );
nand \U$6060 ( \6281 , \4429 , \4430 );
or \U$6061 ( \6282 , \4460 , \6281 );
nand \U$6062 ( \6283 , \4458 , \4459 );
nand \U$6063 ( \6284 , \6282 , \6283 );
and \U$6064 ( \6285 , \4482 , \6284 );
nand \U$6065 ( \6286 , \4470 , \4474 );
or \U$6066 ( \6287 , \4481 , \6286 );
nand \U$6067 ( \6288 , \4476 , \4480 );
nand \U$6068 ( \6289 , \6287 , \6288 );
nor \U$6069 ( \6290 , \6285 , \6289 );
nand \U$6070 ( \6291 , \6280 , \6290 );
nor \U$6071 ( \6292 , \6269 , \6291 );
nand \U$6072 ( \6293 , \6246 , \6292 );
nor \U$6073 ( \6294 , \6199 , \6293 );
not \U$6074 ( \6295 , \6294 );
xnor \U$6075 ( \6296 , \551 , \6295 );
buf \U$6076 ( \6297 , \6296 );
buf \U$6077 ( \6298 , \6297 );
not \U$6078 ( \6299 , \4481 );
nand \U$6079 ( \6300 , \6288 , \6299 );
nor \U$6080 ( \6301 , \5794 , \1649 );
nor \U$6081 ( \6302 , \1802 , \1957 );
nand \U$6082 ( \6303 , \6301 , \6302 );
nor \U$6083 ( \6304 , \2110 , \2264 );
nor \U$6084 ( \6305 , \2411 , \2551 );
nand \U$6085 ( \6306 , \6304 , \6305 );
nor \U$6086 ( \6307 , \6303 , \6306 );
nor \U$6087 ( \6308 , \2688 , \2820 );
nor \U$6088 ( \6309 , \2946 , \3069 );
nand \U$6089 ( \6310 , \6308 , \6309 );
nor \U$6090 ( \6311 , \3185 , \3299 );
nor \U$6091 ( \6312 , \3405 , \3507 );
nand \U$6092 ( \6313 , \6311 , \6312 );
nor \U$6093 ( \6314 , \6310 , \6313 );
nand \U$6094 ( \6315 , \6307 , \6314 );
nor \U$6095 ( \6316 , \3606 , \3701 );
nor \U$6096 ( \6317 , \3790 , \3872 );
nand \U$6097 ( \6318 , \6316 , \6317 );
nor \U$6098 ( \6319 , \3951 , \4025 );
nor \U$6099 ( \6320 , \4090 , \4155 );
nand \U$6100 ( \6321 , \6319 , \6320 );
nor \U$6101 ( \6322 , \6318 , \6321 );
nor \U$6102 ( \6323 , \4214 , \4268 );
nor \U$6103 ( \6324 , \4317 , \4360 );
nand \U$6104 ( \6325 , \6323 , \6324 );
nor \U$6105 ( \6326 , \4395 , \4431 );
nor \U$6106 ( \6327 , \4460 , \4475 );
nand \U$6107 ( \6328 , \6326 , \6327 );
nor \U$6108 ( \6329 , \6325 , \6328 );
nand \U$6109 ( \6330 , \6322 , \6329 );
nor \U$6110 ( \6331 , \6315 , \6330 );
nor \U$6111 ( \6332 , \6049 , \4727 );
nor \U$6112 ( \6333 , \4802 , \4884 );
nand \U$6113 ( \6334 , \6332 , \6333 );
nor \U$6114 ( \6335 , \4969 , \5062 );
nor \U$6115 ( \6336 , \5157 , \5259 );
nand \U$6116 ( \6337 , \6335 , \6336 );
nor \U$6117 ( \6338 , \6334 , \6337 );
nor \U$6118 ( \6339 , \5364 , \5478 );
nor \U$6119 ( \6340 , \5593 , \5667 );
nand \U$6120 ( \6341 , \6339 , \6340 );
nor \U$6121 ( \6342 , \5712 , \5747 );
nor \U$6122 ( \6343 , \5772 , \5787 );
nand \U$6123 ( \6344 , \6342 , \6343 );
nor \U$6124 ( \6345 , \6341 , \6344 );
nand \U$6125 ( \6346 , \6338 , \6345 );
nor \U$6126 ( \6347 , \6096 , \5862 );
nor \U$6127 ( \6348 , \5897 , \5939 );
nand \U$6128 ( \6349 , \6347 , \6348 );
nor \U$6129 ( \6350 , \5984 , \6013 );
nor \U$6130 ( \6351 , \6030 , \6042 );
nand \U$6131 ( \6352 , \6350 , \6351 );
nor \U$6132 ( \6353 , \6349 , \6352 );
nor \U$6133 ( \6354 , \6102 , \6067 );
nor \U$6134 ( \6355 , \6082 , \6092 );
nand \U$6135 ( \6356 , \6354 , \6355 );
or \U$6136 ( \6357 , \6356 , \6110 );
or \U$6137 ( \6358 , \6067 , \6112 );
nand \U$6138 ( \6359 , \6358 , \6116 );
and \U$6139 ( \6360 , \6355 , \6359 );
or \U$6140 ( \6361 , \6092 , \6118 );
nand \U$6141 ( \6362 , \6361 , \6121 );
nor \U$6142 ( \6363 , \6360 , \6362 );
nand \U$6143 ( \6364 , \6357 , \6363 );
and \U$6144 ( \6365 , \6353 , \6364 );
or \U$6145 ( \6366 , \5862 , \6123 );
nand \U$6146 ( \6367 , \6366 , \6128 );
and \U$6147 ( \6368 , \6348 , \6367 );
or \U$6148 ( \6369 , \5939 , \6130 );
nand \U$6149 ( \6370 , \6369 , \6133 );
nor \U$6150 ( \6371 , \6368 , \6370 );
or \U$6151 ( \6372 , \6352 , \6371 );
or \U$6152 ( \6373 , \6013 , \6135 );
nand \U$6153 ( \6374 , \6373 , \6139 );
and \U$6154 ( \6375 , \6351 , \6374 );
or \U$6155 ( \6376 , \6042 , \6141 );
nand \U$6156 ( \6377 , \6376 , \6144 );
nor \U$6157 ( \6378 , \6375 , \6377 );
nand \U$6158 ( \6379 , \6372 , \6378 );
nor \U$6159 ( \6380 , \6365 , \6379 );
or \U$6160 ( \6381 , \6346 , \6380 );
or \U$6161 ( \6382 , \4727 , \6146 );
nand \U$6162 ( \6383 , \6382 , \6152 );
and \U$6163 ( \6384 , \6333 , \6383 );
or \U$6164 ( \6385 , \4884 , \6154 );
nand \U$6165 ( \6386 , \6385 , \6157 );
nor \U$6166 ( \6387 , \6384 , \6386 );
or \U$6167 ( \6388 , \6337 , \6387 );
or \U$6168 ( \6389 , \5062 , \6159 );
nand \U$6169 ( \6390 , \6389 , \6163 );
and \U$6170 ( \6391 , \6336 , \6390 );
or \U$6171 ( \6392 , \5259 , \6165 );
nand \U$6172 ( \6393 , \6392 , \6168 );
nor \U$6173 ( \6394 , \6391 , \6393 );
nand \U$6174 ( \6395 , \6388 , \6394 );
and \U$6175 ( \6396 , \6345 , \6395 );
or \U$6176 ( \6397 , \5478 , \6170 );
nand \U$6177 ( \6398 , \6397 , \6175 );
and \U$6178 ( \6399 , \6340 , \6398 );
or \U$6179 ( \6400 , \5667 , \6177 );
nand \U$6180 ( \6401 , \6400 , \6180 );
nor \U$6181 ( \6402 , \6399 , \6401 );
or \U$6182 ( \6403 , \6344 , \6402 );
or \U$6183 ( \6404 , \5747 , \6182 );
nand \U$6184 ( \6405 , \6404 , \6186 );
and \U$6185 ( \6406 , \6343 , \6405 );
or \U$6186 ( \6407 , \5787 , \6188 );
nand \U$6187 ( \6408 , \6407 , \6191 );
nor \U$6188 ( \6409 , \6406 , \6408 );
nand \U$6189 ( \6410 , \6403 , \6409 );
nor \U$6190 ( \6411 , \6396 , \6410 );
nand \U$6191 ( \6412 , \6381 , \6411 );
and \U$6192 ( \6413 , \6331 , \6412 );
or \U$6193 ( \6414 , \1649 , \6193 );
nand \U$6194 ( \6415 , \6414 , \6200 );
and \U$6195 ( \6416 , \6302 , \6415 );
or \U$6196 ( \6417 , \1957 , \6202 );
nand \U$6197 ( \6418 , \6417 , \6205 );
nor \U$6198 ( \6419 , \6416 , \6418 );
or \U$6199 ( \6420 , \6306 , \6419 );
or \U$6200 ( \6421 , \2264 , \6207 );
nand \U$6201 ( \6422 , \6421 , \6211 );
and \U$6202 ( \6423 , \6305 , \6422 );
or \U$6203 ( \6424 , \2551 , \6213 );
nand \U$6204 ( \6425 , \6424 , \6216 );
nor \U$6205 ( \6426 , \6423 , \6425 );
nand \U$6206 ( \6427 , \6420 , \6426 );
and \U$6207 ( \6428 , \6314 , \6427 );
or \U$6208 ( \6429 , \2820 , \6218 );
nand \U$6209 ( \6430 , \6429 , \6223 );
and \U$6210 ( \6431 , \6309 , \6430 );
or \U$6211 ( \6432 , \3069 , \6225 );
nand \U$6212 ( \6433 , \6432 , \6228 );
nor \U$6213 ( \6434 , \6431 , \6433 );
or \U$6214 ( \6435 , \6313 , \6434 );
or \U$6215 ( \6436 , \3299 , \6230 );
nand \U$6216 ( \6437 , \6436 , \6234 );
and \U$6217 ( \6438 , \6312 , \6437 );
or \U$6218 ( \6439 , \3507 , \6236 );
nand \U$6219 ( \6440 , \6439 , \6239 );
nor \U$6220 ( \6441 , \6438 , \6440 );
nand \U$6221 ( \6442 , \6435 , \6441 );
nor \U$6222 ( \6443 , \6428 , \6442 );
or \U$6223 ( \6444 , \6330 , \6443 );
or \U$6224 ( \6445 , \3701 , \6241 );
nand \U$6225 ( \6446 , \6445 , \6247 );
and \U$6226 ( \6447 , \6317 , \6446 );
or \U$6227 ( \6448 , \3872 , \6249 );
nand \U$6228 ( \6449 , \6448 , \6252 );
nor \U$6229 ( \6450 , \6447 , \6449 );
or \U$6230 ( \6451 , \6321 , \6450 );
or \U$6231 ( \6452 , \4025 , \6254 );
nand \U$6232 ( \6453 , \6452 , \6258 );
and \U$6233 ( \6454 , \6320 , \6453 );
or \U$6234 ( \6455 , \4155 , \6260 );
nand \U$6235 ( \6456 , \6455 , \6263 );
nor \U$6236 ( \6457 , \6454 , \6456 );
nand \U$6237 ( \6458 , \6451 , \6457 );
and \U$6238 ( \6459 , \6329 , \6458 );
or \U$6239 ( \6460 , \4268 , \6265 );
nand \U$6240 ( \6461 , \6460 , \6270 );
and \U$6241 ( \6462 , \6324 , \6461 );
or \U$6242 ( \6463 , \4360 , \6272 );
nand \U$6243 ( \6464 , \6463 , \6275 );
nor \U$6244 ( \6465 , \6462 , \6464 );
or \U$6245 ( \6466 , \6328 , \6465 );
or \U$6246 ( \6467 , \4431 , \6277 );
nand \U$6247 ( \6468 , \6467 , \6281 );
and \U$6248 ( \6469 , \6327 , \6468 );
or \U$6249 ( \6470 , \4475 , \6283 );
nand \U$6250 ( \6471 , \6470 , \6286 );
nor \U$6251 ( \6472 , \6469 , \6471 );
nand \U$6252 ( \6473 , \6466 , \6472 );
nor \U$6253 ( \6474 , \6459 , \6473 );
nand \U$6254 ( \6475 , \6444 , \6474 );
nor \U$6255 ( \6476 , \6413 , \6475 );
not \U$6256 ( \6477 , \6476 );
xnor \U$6257 ( \6478 , \6300 , \6477 );
buf \U$6258 ( \6479 , \6478 );
buf \U$6259 ( \6480 , \6479 );
not \U$6260 ( \6481 , \4475 );
nand \U$6261 ( \6482 , \6286 , \6481 );
nand \U$6262 ( \6483 , \5795 , \1803 );
nand \U$6263 ( \6484 , \2111 , \2412 );
nor \U$6264 ( \6485 , \6483 , \6484 );
nand \U$6265 ( \6486 , \2689 , \2947 );
nand \U$6266 ( \6487 , \3186 , \3406 );
nor \U$6267 ( \6488 , \6486 , \6487 );
nand \U$6268 ( \6489 , \6485 , \6488 );
nand \U$6269 ( \6490 , \3607 , \3791 );
nand \U$6270 ( \6491 , \3952 , \4091 );
nor \U$6271 ( \6492 , \6490 , \6491 );
nand \U$6272 ( \6493 , \4215 , \4318 );
nand \U$6273 ( \6494 , \4396 , \4461 );
nor \U$6274 ( \6495 , \6493 , \6494 );
nand \U$6275 ( \6496 , \6492 , \6495 );
nor \U$6276 ( \6497 , \6489 , \6496 );
nand \U$6277 ( \6498 , \6050 , \4803 );
nand \U$6278 ( \6499 , \4970 , \5158 );
nor \U$6279 ( \6500 , \6498 , \6499 );
nand \U$6280 ( \6501 , \5365 , \5594 );
nand \U$6281 ( \6502 , \5713 , \5773 );
nor \U$6282 ( \6503 , \6501 , \6502 );
nand \U$6283 ( \6504 , \6500 , \6503 );
nand \U$6284 ( \6505 , \6097 , \5898 );
nand \U$6285 ( \6506 , \5985 , \6031 );
nor \U$6286 ( \6507 , \6505 , \6506 );
and \U$6287 ( \6508 , \6083 , \6113 );
nor \U$6288 ( \6509 , \6508 , \6119 );
not \U$6289 ( \6510 , \6509 );
and \U$6290 ( \6511 , \6507 , \6510 );
and \U$6291 ( \6512 , \5898 , \6124 );
nor \U$6292 ( \6513 , \6512 , \6131 );
or \U$6293 ( \6514 , \6506 , \6513 );
and \U$6294 ( \6515 , \6031 , \6136 );
nor \U$6295 ( \6516 , \6515 , \6142 );
nand \U$6296 ( \6517 , \6514 , \6516 );
nor \U$6297 ( \6518 , \6511 , \6517 );
or \U$6298 ( \6519 , \6504 , \6518 );
and \U$6299 ( \6520 , \4803 , \6147 );
nor \U$6300 ( \6521 , \6520 , \6155 );
or \U$6301 ( \6522 , \6499 , \6521 );
and \U$6302 ( \6523 , \5158 , \6160 );
nor \U$6303 ( \6524 , \6523 , \6166 );
nand \U$6304 ( \6525 , \6522 , \6524 );
and \U$6305 ( \6526 , \6503 , \6525 );
and \U$6306 ( \6527 , \5594 , \6171 );
nor \U$6307 ( \6528 , \6527 , \6178 );
or \U$6308 ( \6529 , \6502 , \6528 );
and \U$6309 ( \6530 , \5773 , \6183 );
nor \U$6310 ( \6531 , \6530 , \6189 );
nand \U$6311 ( \6532 , \6529 , \6531 );
nor \U$6312 ( \6533 , \6526 , \6532 );
nand \U$6313 ( \6534 , \6519 , \6533 );
and \U$6314 ( \6535 , \6497 , \6534 );
and \U$6315 ( \6536 , \1803 , \6194 );
nor \U$6316 ( \6537 , \6536 , \6203 );
or \U$6317 ( \6538 , \6484 , \6537 );
and \U$6318 ( \6539 , \2412 , \6208 );
nor \U$6319 ( \6540 , \6539 , \6214 );
nand \U$6320 ( \6541 , \6538 , \6540 );
and \U$6321 ( \6542 , \6488 , \6541 );
and \U$6322 ( \6543 , \2947 , \6219 );
nor \U$6323 ( \6544 , \6543 , \6226 );
or \U$6324 ( \6545 , \6487 , \6544 );
and \U$6325 ( \6546 , \3406 , \6231 );
nor \U$6326 ( \6547 , \6546 , \6237 );
nand \U$6327 ( \6548 , \6545 , \6547 );
nor \U$6328 ( \6549 , \6542 , \6548 );
or \U$6329 ( \6550 , \6496 , \6549 );
and \U$6330 ( \6551 , \3791 , \6242 );
nor \U$6331 ( \6552 , \6551 , \6250 );
or \U$6332 ( \6553 , \6491 , \6552 );
and \U$6333 ( \6554 , \4091 , \6255 );
nor \U$6334 ( \6555 , \6554 , \6261 );
nand \U$6335 ( \6556 , \6553 , \6555 );
and \U$6336 ( \6557 , \6495 , \6556 );
and \U$6337 ( \6558 , \4318 , \6266 );
nor \U$6338 ( \6559 , \6558 , \6273 );
or \U$6339 ( \6560 , \6494 , \6559 );
and \U$6340 ( \6561 , \4461 , \6278 );
nor \U$6341 ( \6562 , \6561 , \6284 );
nand \U$6342 ( \6563 , \6560 , \6562 );
nor \U$6343 ( \6564 , \6557 , \6563 );
nand \U$6344 ( \6565 , \6550 , \6564 );
nor \U$6345 ( \6566 , \6535 , \6565 );
not \U$6346 ( \6567 , \6566 );
xnor \U$6347 ( \6568 , \6482 , \6567 );
buf \U$6348 ( \6569 , \6568 );
buf \U$6349 ( \6570 , \6569 );
not \U$6350 ( \6571 , \4460 );
nand \U$6351 ( \6572 , \6283 , \6571 );
nand \U$6352 ( \6573 , \6343 , \6301 );
nand \U$6353 ( \6574 , \6302 , \6304 );
nor \U$6354 ( \6575 , \6573 , \6574 );
nand \U$6355 ( \6576 , \6305 , \6308 );
nand \U$6356 ( \6577 , \6309 , \6311 );
nor \U$6357 ( \6578 , \6576 , \6577 );
nand \U$6358 ( \6579 , \6575 , \6578 );
nand \U$6359 ( \6580 , \6312 , \6316 );
nand \U$6360 ( \6581 , \6317 , \6319 );
nor \U$6361 ( \6582 , \6580 , \6581 );
nand \U$6362 ( \6583 , \6320 , \6323 );
nand \U$6363 ( \6584 , \6324 , \6326 );
nor \U$6364 ( \6585 , \6583 , \6584 );
nand \U$6365 ( \6586 , \6582 , \6585 );
nor \U$6366 ( \6587 , \6579 , \6586 );
nand \U$6367 ( \6588 , \6351 , \6332 );
nand \U$6368 ( \6589 , \6333 , \6335 );
nor \U$6369 ( \6590 , \6588 , \6589 );
nand \U$6370 ( \6591 , \6336 , \6339 );
nand \U$6371 ( \6592 , \6340 , \6342 );
nor \U$6372 ( \6593 , \6591 , \6592 );
nand \U$6373 ( \6594 , \6590 , \6593 );
nand \U$6374 ( \6595 , \6355 , \6347 );
nand \U$6375 ( \6596 , \6348 , \6350 );
nor \U$6376 ( \6597 , \6595 , \6596 );
not \U$6377 ( \6598 , \6110 );
and \U$6378 ( \6599 , \6354 , \6598 );
nor \U$6379 ( \6600 , \6599 , \6359 );
not \U$6380 ( \6601 , \6600 );
and \U$6381 ( \6602 , \6597 , \6601 );
and \U$6382 ( \6603 , \6347 , \6362 );
nor \U$6383 ( \6604 , \6603 , \6367 );
or \U$6384 ( \6605 , \6596 , \6604 );
and \U$6385 ( \6606 , \6350 , \6370 );
nor \U$6386 ( \6607 , \6606 , \6374 );
nand \U$6387 ( \6608 , \6605 , \6607 );
nor \U$6388 ( \6609 , \6602 , \6608 );
or \U$6389 ( \6610 , \6594 , \6609 );
and \U$6390 ( \6611 , \6332 , \6377 );
nor \U$6391 ( \6612 , \6611 , \6383 );
or \U$6392 ( \6613 , \6589 , \6612 );
and \U$6393 ( \6614 , \6335 , \6386 );
nor \U$6394 ( \6615 , \6614 , \6390 );
nand \U$6395 ( \6616 , \6613 , \6615 );
and \U$6396 ( \6617 , \6593 , \6616 );
and \U$6397 ( \6618 , \6339 , \6393 );
nor \U$6398 ( \6619 , \6618 , \6398 );
or \U$6399 ( \6620 , \6592 , \6619 );
and \U$6400 ( \6621 , \6342 , \6401 );
nor \U$6401 ( \6622 , \6621 , \6405 );
nand \U$6402 ( \6623 , \6620 , \6622 );
nor \U$6403 ( \6624 , \6617 , \6623 );
nand \U$6404 ( \6625 , \6610 , \6624 );
and \U$6405 ( \6626 , \6587 , \6625 );
and \U$6406 ( \6627 , \6301 , \6408 );
nor \U$6407 ( \6628 , \6627 , \6415 );
or \U$6408 ( \6629 , \6574 , \6628 );
and \U$6409 ( \6630 , \6304 , \6418 );
nor \U$6410 ( \6631 , \6630 , \6422 );
nand \U$6411 ( \6632 , \6629 , \6631 );
and \U$6412 ( \6633 , \6578 , \6632 );
and \U$6413 ( \6634 , \6308 , \6425 );
nor \U$6414 ( \6635 , \6634 , \6430 );
or \U$6415 ( \6636 , \6577 , \6635 );
and \U$6416 ( \6637 , \6311 , \6433 );
nor \U$6417 ( \6638 , \6637 , \6437 );
nand \U$6418 ( \6639 , \6636 , \6638 );
nor \U$6419 ( \6640 , \6633 , \6639 );
or \U$6420 ( \6641 , \6586 , \6640 );
and \U$6421 ( \6642 , \6316 , \6440 );
nor \U$6422 ( \6643 , \6642 , \6446 );
or \U$6423 ( \6644 , \6581 , \6643 );
and \U$6424 ( \6645 , \6319 , \6449 );
nor \U$6425 ( \6646 , \6645 , \6453 );
nand \U$6426 ( \6647 , \6644 , \6646 );
and \U$6427 ( \6648 , \6585 , \6647 );
and \U$6428 ( \6649 , \6323 , \6456 );
nor \U$6429 ( \6650 , \6649 , \6461 );
or \U$6430 ( \6651 , \6584 , \6650 );
and \U$6431 ( \6652 , \6326 , \6464 );
nor \U$6432 ( \6653 , \6652 , \6468 );
nand \U$6433 ( \6654 , \6651 , \6653 );
nor \U$6434 ( \6655 , \6648 , \6654 );
nand \U$6435 ( \6656 , \6641 , \6655 );
nor \U$6436 ( \6657 , \6626 , \6656 );
not \U$6437 ( \6658 , \6657 );
xnor \U$6438 ( \6659 , \6572 , \6658 );
buf \U$6439 ( \6660 , \6659 );
buf \U$6440 ( \6661 , \6660 );
not \U$6441 ( \6662 , \4431 );
nand \U$6442 ( \6663 , \6281 , \6662 );
nor \U$6443 ( \6664 , \5796 , \2112 );
nor \U$6444 ( \6665 , \2690 , \3187 );
nand \U$6445 ( \6666 , \6664 , \6665 );
nor \U$6446 ( \6667 , \3608 , \3953 );
nor \U$6447 ( \6668 , \4216 , \4397 );
nand \U$6448 ( \6669 , \6667 , \6668 );
nor \U$6449 ( \6670 , \6666 , \6669 );
nor \U$6450 ( \6671 , \6051 , \4971 );
nor \U$6451 ( \6672 , \5366 , \5714 );
nand \U$6452 ( \6673 , \6671 , \6672 );
nor \U$6453 ( \6674 , \6098 , \5986 );
and \U$6454 ( \6675 , \6674 , \6113 );
or \U$6455 ( \6676 , \5986 , \6125 );
nand \U$6456 ( \6677 , \6676 , \6137 );
nor \U$6457 ( \6678 , \6675 , \6677 );
or \U$6458 ( \6679 , \6673 , \6678 );
or \U$6459 ( \6680 , \4971 , \6148 );
nand \U$6460 ( \6681 , \6680 , \6161 );
and \U$6461 ( \6682 , \6672 , \6681 );
or \U$6462 ( \6683 , \5714 , \6172 );
nand \U$6463 ( \6684 , \6683 , \6184 );
nor \U$6464 ( \6685 , \6682 , \6684 );
nand \U$6465 ( \6686 , \6679 , \6685 );
and \U$6466 ( \6687 , \6670 , \6686 );
or \U$6467 ( \6688 , \2112 , \6195 );
nand \U$6468 ( \6689 , \6688 , \6209 );
and \U$6469 ( \6690 , \6665 , \6689 );
or \U$6470 ( \6691 , \3187 , \6220 );
nand \U$6471 ( \6692 , \6691 , \6232 );
nor \U$6472 ( \6693 , \6690 , \6692 );
or \U$6473 ( \6694 , \6669 , \6693 );
or \U$6474 ( \6695 , \3953 , \6243 );
nand \U$6475 ( \6696 , \6695 , \6256 );
and \U$6476 ( \6697 , \6668 , \6696 );
or \U$6477 ( \6698 , \4397 , \6267 );
nand \U$6478 ( \6699 , \6698 , \6279 );
nor \U$6479 ( \6700 , \6697 , \6699 );
nand \U$6480 ( \6701 , \6694 , \6700 );
nor \U$6481 ( \6702 , \6687 , \6701 );
not \U$6482 ( \6703 , \6702 );
xnor \U$6483 ( \6704 , \6663 , \6703 );
buf \U$6484 ( \6705 , \6704 );
buf \U$6485 ( \6706 , \6705 );
not \U$6486 ( \6707 , \4395 );
nand \U$6487 ( \6708 , \6277 , \6707 );
nor \U$6488 ( \6709 , \6344 , \6303 );
nor \U$6489 ( \6710 , \6306 , \6310 );
nand \U$6490 ( \6711 , \6709 , \6710 );
nor \U$6491 ( \6712 , \6313 , \6318 );
nor \U$6492 ( \6713 , \6321 , \6325 );
nand \U$6493 ( \6714 , \6712 , \6713 );
nor \U$6494 ( \6715 , \6711 , \6714 );
nor \U$6495 ( \6716 , \6352 , \6334 );
nor \U$6496 ( \6717 , \6337 , \6341 );
nand \U$6497 ( \6718 , \6716 , \6717 );
nor \U$6498 ( \6719 , \6356 , \6349 );
and \U$6499 ( \6720 , \6719 , \6598 );
or \U$6500 ( \6721 , \6349 , \6363 );
nand \U$6501 ( \6722 , \6721 , \6371 );
nor \U$6502 ( \6723 , \6720 , \6722 );
or \U$6503 ( \6724 , \6718 , \6723 );
or \U$6504 ( \6725 , \6334 , \6378 );
nand \U$6505 ( \6726 , \6725 , \6387 );
and \U$6506 ( \6727 , \6717 , \6726 );
or \U$6507 ( \6728 , \6341 , \6394 );
nand \U$6508 ( \6729 , \6728 , \6402 );
nor \U$6509 ( \6730 , \6727 , \6729 );
nand \U$6510 ( \6731 , \6724 , \6730 );
and \U$6511 ( \6732 , \6715 , \6731 );
or \U$6512 ( \6733 , \6303 , \6409 );
nand \U$6513 ( \6734 , \6733 , \6419 );
and \U$6514 ( \6735 , \6710 , \6734 );
or \U$6515 ( \6736 , \6310 , \6426 );
nand \U$6516 ( \6737 , \6736 , \6434 );
nor \U$6517 ( \6738 , \6735 , \6737 );
or \U$6518 ( \6739 , \6714 , \6738 );
or \U$6519 ( \6740 , \6318 , \6441 );
nand \U$6520 ( \6741 , \6740 , \6450 );
and \U$6521 ( \6742 , \6713 , \6741 );
or \U$6522 ( \6743 , \6325 , \6457 );
nand \U$6523 ( \6744 , \6743 , \6465 );
nor \U$6524 ( \6745 , \6742 , \6744 );
nand \U$6525 ( \6746 , \6739 , \6745 );
nor \U$6526 ( \6747 , \6732 , \6746 );
not \U$6527 ( \6748 , \6747 );
xnor \U$6528 ( \6749 , \6708 , \6748 );
buf \U$6529 ( \6750 , \6749 );
buf \U$6530 ( \6751 , \6750 );
not \U$6531 ( \6752 , \4360 );
nand \U$6532 ( \6753 , \6275 , \6752 );
nor \U$6533 ( \6754 , \6502 , \6483 );
nor \U$6534 ( \6755 , \6484 , \6486 );
nand \U$6535 ( \6756 , \6754 , \6755 );
nor \U$6536 ( \6757 , \6487 , \6490 );
nor \U$6537 ( \6758 , \6491 , \6493 );
nand \U$6538 ( \6759 , \6757 , \6758 );
nor \U$6539 ( \6760 , \6756 , \6759 );
nor \U$6540 ( \6761 , \6506 , \6498 );
nor \U$6541 ( \6762 , \6499 , \6501 );
nand \U$6542 ( \6763 , \6761 , \6762 );
or \U$6543 ( \6764 , \6505 , \6509 );
nand \U$6544 ( \6765 , \6764 , \6513 );
not \U$6545 ( \6766 , \6765 );
or \U$6546 ( \6767 , \6763 , \6766 );
or \U$6547 ( \6768 , \6498 , \6516 );
nand \U$6548 ( \6769 , \6768 , \6521 );
and \U$6549 ( \6770 , \6762 , \6769 );
or \U$6550 ( \6771 , \6501 , \6524 );
nand \U$6551 ( \6772 , \6771 , \6528 );
nor \U$6552 ( \6773 , \6770 , \6772 );
nand \U$6553 ( \6774 , \6767 , \6773 );
and \U$6554 ( \6775 , \6760 , \6774 );
or \U$6555 ( \6776 , \6483 , \6531 );
nand \U$6556 ( \6777 , \6776 , \6537 );
and \U$6557 ( \6778 , \6755 , \6777 );
or \U$6558 ( \6779 , \6486 , \6540 );
nand \U$6559 ( \6780 , \6779 , \6544 );
nor \U$6560 ( \6781 , \6778 , \6780 );
or \U$6561 ( \6782 , \6759 , \6781 );
or \U$6562 ( \6783 , \6490 , \6547 );
nand \U$6563 ( \6784 , \6783 , \6552 );
and \U$6564 ( \6785 , \6758 , \6784 );
or \U$6565 ( \6786 , \6493 , \6555 );
nand \U$6566 ( \6787 , \6786 , \6559 );
nor \U$6567 ( \6788 , \6785 , \6787 );
nand \U$6568 ( \6789 , \6782 , \6788 );
nor \U$6569 ( \6790 , \6775 , \6789 );
not \U$6570 ( \6791 , \6790 );
xnor \U$6571 ( \6792 , \6753 , \6791 );
buf \U$6572 ( \6793 , \6792 );
buf \U$6573 ( \6794 , \6793 );
not \U$6574 ( \6795 , \4317 );
nand \U$6575 ( \6796 , \6272 , \6795 );
nor \U$6576 ( \6797 , \6592 , \6573 );
nor \U$6577 ( \6798 , \6574 , \6576 );
nand \U$6578 ( \6799 , \6797 , \6798 );
nor \U$6579 ( \6800 , \6577 , \6580 );
nor \U$6580 ( \6801 , \6581 , \6583 );
nand \U$6581 ( \6802 , \6800 , \6801 );
nor \U$6582 ( \6803 , \6799 , \6802 );
nor \U$6583 ( \6804 , \6596 , \6588 );
nor \U$6584 ( \6805 , \6589 , \6591 );
nand \U$6585 ( \6806 , \6804 , \6805 );
or \U$6586 ( \6807 , \6595 , \6600 );
nand \U$6587 ( \6808 , \6807 , \6604 );
not \U$6588 ( \6809 , \6808 );
or \U$6589 ( \6810 , \6806 , \6809 );
or \U$6590 ( \6811 , \6588 , \6607 );
nand \U$6591 ( \6812 , \6811 , \6612 );
and \U$6592 ( \6813 , \6805 , \6812 );
or \U$6593 ( \6814 , \6591 , \6615 );
nand \U$6594 ( \6815 , \6814 , \6619 );
nor \U$6595 ( \6816 , \6813 , \6815 );
nand \U$6596 ( \6817 , \6810 , \6816 );
and \U$6597 ( \6818 , \6803 , \6817 );
or \U$6598 ( \6819 , \6573 , \6622 );
nand \U$6599 ( \6820 , \6819 , \6628 );
and \U$6600 ( \6821 , \6798 , \6820 );
or \U$6601 ( \6822 , \6576 , \6631 );
nand \U$6602 ( \6823 , \6822 , \6635 );
nor \U$6603 ( \6824 , \6821 , \6823 );
or \U$6604 ( \6825 , \6802 , \6824 );
or \U$6605 ( \6826 , \6580 , \6638 );
nand \U$6606 ( \6827 , \6826 , \6643 );
and \U$6607 ( \6828 , \6801 , \6827 );
or \U$6608 ( \6829 , \6583 , \6646 );
nand \U$6609 ( \6830 , \6829 , \6650 );
nor \U$6610 ( \6831 , \6828 , \6830 );
nand \U$6611 ( \6832 , \6825 , \6831 );
nor \U$6612 ( \6833 , \6818 , \6832 );
not \U$6613 ( \6834 , \6833 );
xnor \U$6614 ( \6835 , \6796 , \6834 );
buf \U$6615 ( \6836 , \6835 );
buf \U$6616 ( \6837 , \6836 );
not \U$6617 ( \6838 , \4268 );
nand \U$6618 ( \6839 , \6270 , \6838 );
nand \U$6619 ( \6840 , \5797 , \2691 );
nand \U$6620 ( \6841 , \3609 , \4217 );
nor \U$6621 ( \6842 , \6840 , \6841 );
nand \U$6622 ( \6843 , \6052 , \5367 );
not \U$6623 ( \6844 , \6126 );
or \U$6624 ( \6845 , \6843 , \6844 );
and \U$6625 ( \6846 , \5367 , \6149 );
nor \U$6626 ( \6847 , \6846 , \6173 );
nand \U$6627 ( \6848 , \6845 , \6847 );
and \U$6628 ( \6849 , \6842 , \6848 );
and \U$6629 ( \6850 , \2691 , \6196 );
nor \U$6630 ( \6851 , \6850 , \6221 );
or \U$6631 ( \6852 , \6841 , \6851 );
and \U$6632 ( \6853 , \4217 , \6244 );
nor \U$6633 ( \6854 , \6853 , \6268 );
nand \U$6634 ( \6855 , \6852 , \6854 );
nor \U$6635 ( \6856 , \6849 , \6855 );
not \U$6636 ( \6857 , \6856 );
xnor \U$6637 ( \6858 , \6839 , \6857 );
buf \U$6638 ( \6859 , \6858 );
buf \U$6639 ( \6860 , \6859 );
not \U$6640 ( \6861 , \4214 );
nand \U$6641 ( \6862 , \6265 , \6861 );
nand \U$6642 ( \6863 , \6345 , \6307 );
nand \U$6643 ( \6864 , \6314 , \6322 );
nor \U$6644 ( \6865 , \6863 , \6864 );
nand \U$6645 ( \6866 , \6353 , \6338 );
not \U$6646 ( \6867 , \6364 );
or \U$6647 ( \6868 , \6866 , \6867 );
and \U$6648 ( \6869 , \6338 , \6379 );
nor \U$6649 ( \6870 , \6869 , \6395 );
nand \U$6650 ( \6871 , \6868 , \6870 );
and \U$6651 ( \6872 , \6865 , \6871 );
and \U$6652 ( \6873 , \6307 , \6410 );
nor \U$6653 ( \6874 , \6873 , \6427 );
or \U$6654 ( \6875 , \6864 , \6874 );
and \U$6655 ( \6876 , \6322 , \6442 );
nor \U$6656 ( \6877 , \6876 , \6458 );
nand \U$6657 ( \6878 , \6875 , \6877 );
nor \U$6658 ( \6879 , \6872 , \6878 );
not \U$6659 ( \6880 , \6879 );
xnor \U$6660 ( \6881 , \6862 , \6880 );
buf \U$6661 ( \6882 , \6881 );
buf \U$6662 ( \6883 , \6882 );
not \U$6663 ( \6884 , \4155 );
nand \U$6664 ( \6885 , \6263 , \6884 );
nand \U$6665 ( \6886 , \6503 , \6485 );
nand \U$6666 ( \6887 , \6488 , \6492 );
nor \U$6667 ( \6888 , \6886 , \6887 );
nand \U$6668 ( \6889 , \6507 , \6500 );
or \U$6669 ( \6890 , \6889 , \6509 );
and \U$6670 ( \6891 , \6500 , \6517 );
nor \U$6671 ( \6892 , \6891 , \6525 );
nand \U$6672 ( \6893 , \6890 , \6892 );
and \U$6673 ( \6894 , \6888 , \6893 );
and \U$6674 ( \6895 , \6485 , \6532 );
nor \U$6675 ( \6896 , \6895 , \6541 );
or \U$6676 ( \6897 , \6887 , \6896 );
and \U$6677 ( \6898 , \6492 , \6548 );
nor \U$6678 ( \6899 , \6898 , \6556 );
nand \U$6679 ( \6900 , \6897 , \6899 );
nor \U$6680 ( \6901 , \6894 , \6900 );
not \U$6681 ( \6902 , \6901 );
xnor \U$6682 ( \6903 , \6885 , \6902 );
buf \U$6683 ( \6904 , \6903 );
buf \U$6684 ( \6905 , \6904 );
not \U$6685 ( \6906 , \4090 );
nand \U$6686 ( \6907 , \6260 , \6906 );
nand \U$6687 ( \6908 , \6593 , \6575 );
nand \U$6688 ( \6909 , \6578 , \6582 );
nor \U$6689 ( \6910 , \6908 , \6909 );
nand \U$6690 ( \6911 , \6597 , \6590 );
or \U$6691 ( \6912 , \6911 , \6600 );
and \U$6692 ( \6913 , \6590 , \6608 );
nor \U$6693 ( \6914 , \6913 , \6616 );
nand \U$6694 ( \6915 , \6912 , \6914 );
and \U$6695 ( \6916 , \6910 , \6915 );
and \U$6696 ( \6917 , \6575 , \6623 );
nor \U$6697 ( \6918 , \6917 , \6632 );
or \U$6698 ( \6919 , \6909 , \6918 );
and \U$6699 ( \6920 , \6582 , \6639 );
nor \U$6700 ( \6921 , \6920 , \6647 );
nand \U$6701 ( \6922 , \6919 , \6921 );
nor \U$6702 ( \6923 , \6916 , \6922 );
not \U$6703 ( \6924 , \6923 );
xnor \U$6704 ( \6925 , \6907 , \6924 );
buf \U$6705 ( \6926 , \6925 );
buf \U$6706 ( \6927 , \6926 );
not \U$6707 ( \6928 , \4025 );
nand \U$6708 ( \6929 , \6258 , \6928 );
nand \U$6709 ( \6930 , \6672 , \6664 );
nand \U$6710 ( \6931 , \6665 , \6667 );
nor \U$6711 ( \6932 , \6930 , \6931 );
nand \U$6712 ( \6933 , \6674 , \6671 );
or \U$6713 ( \6934 , \6933 , \6114 );
and \U$6714 ( \6935 , \6671 , \6677 );
nor \U$6715 ( \6936 , \6935 , \6681 );
nand \U$6716 ( \6937 , \6934 , \6936 );
and \U$6717 ( \6938 , \6932 , \6937 );
and \U$6718 ( \6939 , \6664 , \6684 );
nor \U$6719 ( \6940 , \6939 , \6689 );
or \U$6720 ( \6941 , \6931 , \6940 );
and \U$6721 ( \6942 , \6667 , \6692 );
nor \U$6722 ( \6943 , \6942 , \6696 );
nand \U$6723 ( \6944 , \6941 , \6943 );
nor \U$6724 ( \6945 , \6938 , \6944 );
not \U$6725 ( \6946 , \6945 );
xnor \U$6726 ( \6947 , \6929 , \6946 );
buf \U$6727 ( \6948 , \6947 );
buf \U$6728 ( \6949 , \6948 );
not \U$6729 ( \6950 , \3951 );
nand \U$6730 ( \6951 , \6254 , \6950 );
nand \U$6731 ( \6952 , \6717 , \6709 );
nand \U$6732 ( \6953 , \6710 , \6712 );
nor \U$6733 ( \6954 , \6952 , \6953 );
nand \U$6734 ( \6955 , \6719 , \6716 );
or \U$6735 ( \6956 , \6955 , \6110 );
and \U$6736 ( \6957 , \6716 , \6722 );
nor \U$6737 ( \6958 , \6957 , \6726 );
nand \U$6738 ( \6959 , \6956 , \6958 );
and \U$6739 ( \6960 , \6954 , \6959 );
and \U$6740 ( \6961 , \6709 , \6729 );
nor \U$6741 ( \6962 , \6961 , \6734 );
or \U$6742 ( \6963 , \6953 , \6962 );
and \U$6743 ( \6964 , \6712 , \6737 );
nor \U$6744 ( \6965 , \6964 , \6741 );
nand \U$6745 ( \6966 , \6963 , \6965 );
nor \U$6746 ( \6967 , \6960 , \6966 );
not \U$6747 ( \6968 , \6967 );
xnor \U$6748 ( \6969 , \6951 , \6968 );
buf \U$6749 ( \6970 , \6969 );
buf \U$6750 ( \6971 , \6970 );
not \U$6751 ( \6972 , \3872 );
nand \U$6752 ( \6973 , \6252 , \6972 );
nand \U$6753 ( \6974 , \6762 , \6754 );
nand \U$6754 ( \6975 , \6755 , \6757 );
nor \U$6755 ( \6976 , \6974 , \6975 );
and \U$6756 ( \6977 , \6761 , \6765 );
nor \U$6757 ( \6978 , \6977 , \6769 );
not \U$6758 ( \6979 , \6978 );
and \U$6759 ( \6980 , \6976 , \6979 );
and \U$6760 ( \6981 , \6754 , \6772 );
nor \U$6761 ( \6982 , \6981 , \6777 );
or \U$6762 ( \6983 , \6975 , \6982 );
and \U$6763 ( \6984 , \6757 , \6780 );
nor \U$6764 ( \6985 , \6984 , \6784 );
nand \U$6765 ( \6986 , \6983 , \6985 );
nor \U$6766 ( \6987 , \6980 , \6986 );
not \U$6767 ( \6988 , \6987 );
xnor \U$6768 ( \6989 , \6973 , \6988 );
buf \U$6769 ( \6990 , \6989 );
buf \U$6770 ( \6991 , \6990 );
not \U$6771 ( \6992 , \3790 );
nand \U$6772 ( \6993 , \6249 , \6992 );
nand \U$6773 ( \6994 , \6805 , \6797 );
nand \U$6774 ( \6995 , \6798 , \6800 );
nor \U$6775 ( \6996 , \6994 , \6995 );
and \U$6776 ( \6997 , \6804 , \6808 );
nor \U$6777 ( \6998 , \6997 , \6812 );
not \U$6778 ( \6999 , \6998 );
and \U$6779 ( \7000 , \6996 , \6999 );
and \U$6780 ( \7001 , \6797 , \6815 );
nor \U$6781 ( \7002 , \7001 , \6820 );
or \U$6782 ( \7003 , \6995 , \7002 );
and \U$6783 ( \7004 , \6800 , \6823 );
nor \U$6784 ( \7005 , \7004 , \6827 );
nand \U$6785 ( \7006 , \7003 , \7005 );
nor \U$6786 ( \7007 , \7000 , \7006 );
not \U$6787 ( \7008 , \7007 );
xnor \U$6788 ( \7009 , \6993 , \7008 );
buf \U$6789 ( \7010 , \7009 );
buf \U$6790 ( \7011 , \7010 );
not \U$6791 ( \7012 , \3701 );
nand \U$6792 ( \7013 , \6247 , \7012 );
nor \U$6793 ( \7014 , \5798 , \3610 );
not \U$6794 ( \7015 , \6150 );
and \U$6795 ( \7016 , \7014 , \7015 );
or \U$6796 ( \7017 , \3610 , \6197 );
nand \U$6797 ( \7018 , \7017 , \6245 );
nor \U$6798 ( \7019 , \7016 , \7018 );
not \U$6799 ( \7020 , \7019 );
xnor \U$6800 ( \7021 , \7013 , \7020 );
buf \U$6801 ( \7022 , \7021 );
buf \U$6802 ( \7023 , \7022 );
not \U$6803 ( \7024 , \3606 );
nand \U$6804 ( \7025 , \6241 , \7024 );
nor \U$6805 ( \7026 , \6346 , \6315 );
not \U$6806 ( \7027 , \6380 );
and \U$6807 ( \7028 , \7026 , \7027 );
or \U$6808 ( \7029 , \6315 , \6411 );
nand \U$6809 ( \7030 , \7029 , \6443 );
nor \U$6810 ( \7031 , \7028 , \7030 );
not \U$6811 ( \7032 , \7031 );
xnor \U$6812 ( \7033 , \7025 , \7032 );
buf \U$6813 ( \7034 , \7033 );
buf \U$6814 ( \7035 , \7034 );
not \U$6815 ( \7036 , \3507 );
nand \U$6816 ( \7037 , \6239 , \7036 );
nor \U$6817 ( \7038 , \6504 , \6489 );
not \U$6818 ( \7039 , \6518 );
and \U$6819 ( \7040 , \7038 , \7039 );
or \U$6820 ( \7041 , \6489 , \6533 );
nand \U$6821 ( \7042 , \7041 , \6549 );
nor \U$6822 ( \7043 , \7040 , \7042 );
not \U$6823 ( \7044 , \7043 );
xnor \U$6824 ( \7045 , \7037 , \7044 );
buf \U$6825 ( \7046 , \7045 );
buf \U$6826 ( \7047 , \7046 );
not \U$6827 ( \7048 , \3405 );
nand \U$6828 ( \7049 , \6236 , \7048 );
nor \U$6829 ( \7050 , \6594 , \6579 );
not \U$6830 ( \7051 , \6609 );
and \U$6831 ( \7052 , \7050 , \7051 );
or \U$6832 ( \7053 , \6579 , \6624 );
nand \U$6833 ( \7054 , \7053 , \6640 );
nor \U$6834 ( \7055 , \7052 , \7054 );
not \U$6835 ( \7056 , \7055 );
xnor \U$6836 ( \7057 , \7049 , \7056 );
buf \U$6837 ( \7058 , \7057 );
buf \U$6838 ( \7059 , \7058 );
not \U$6839 ( \7060 , \3299 );
nand \U$6840 ( \7061 , \6234 , \7060 );
nor \U$6841 ( \7062 , \6673 , \6666 );
not \U$6842 ( \7063 , \6678 );
and \U$6843 ( \7064 , \7062 , \7063 );
or \U$6844 ( \7065 , \6666 , \6685 );
nand \U$6845 ( \7066 , \7065 , \6693 );
nor \U$6846 ( \7067 , \7064 , \7066 );
not \U$6847 ( \7068 , \7067 );
xnor \U$6848 ( \7069 , \7061 , \7068 );
buf \U$6849 ( \7070 , \7069 );
buf \U$6850 ( \7071 , \7070 );
not \U$6851 ( \7072 , \3185 );
nand \U$6852 ( \7073 , \6230 , \7072 );
nor \U$6853 ( \7074 , \6718 , \6711 );
not \U$6854 ( \7075 , \6723 );
and \U$6855 ( \7076 , \7074 , \7075 );
or \U$6856 ( \7077 , \6711 , \6730 );
nand \U$6857 ( \7078 , \7077 , \6738 );
nor \U$6858 ( \7079 , \7076 , \7078 );
not \U$6859 ( \7080 , \7079 );
xnor \U$6860 ( \7081 , \7073 , \7080 );
buf \U$6861 ( \7082 , \7081 );
buf \U$6862 ( \7083 , \7082 );
not \U$6863 ( \7084 , \3069 );
nand \U$6864 ( \7085 , \6228 , \7084 );
nor \U$6865 ( \7086 , \6763 , \6756 );
and \U$6866 ( \7087 , \7086 , \6765 );
or \U$6867 ( \7088 , \6756 , \6773 );
nand \U$6868 ( \7089 , \7088 , \6781 );
nor \U$6869 ( \7090 , \7087 , \7089 );
not \U$6870 ( \7091 , \7090 );
xnor \U$6871 ( \7092 , \7085 , \7091 );
buf \U$6872 ( \7093 , \7092 );
buf \U$6873 ( \7094 , \7093 );
not \U$6874 ( \7095 , \2946 );
nand \U$6875 ( \7096 , \6225 , \7095 );
nor \U$6876 ( \7097 , \6806 , \6799 );
and \U$6877 ( \7098 , \7097 , \6808 );
or \U$6878 ( \7099 , \6799 , \6816 );
nand \U$6879 ( \7100 , \7099 , \6824 );
nor \U$6880 ( \7101 , \7098 , \7100 );
not \U$6881 ( \7102 , \7101 );
xnor \U$6882 ( \7103 , \7096 , \7102 );
buf \U$6883 ( \7104 , \7103 );
buf \U$6884 ( \7105 , \7104 );
not \U$6885 ( \7106 , \2820 );
nand \U$6886 ( \7107 , \6223 , \7106 );
nor \U$6887 ( \7108 , \6843 , \6840 );
and \U$6888 ( \7109 , \7108 , \6126 );
or \U$6889 ( \7110 , \6840 , \6847 );
nand \U$6890 ( \7111 , \7110 , \6851 );
nor \U$6891 ( \7112 , \7109 , \7111 );
not \U$6892 ( \7113 , \7112 );
xnor \U$6893 ( \7114 , \7107 , \7113 );
buf \U$6894 ( \7115 , \7114 );
buf \U$6895 ( \7116 , \7115 );
not \U$6896 ( \7117 , \2688 );
nand \U$6897 ( \7118 , \6218 , \7117 );
nor \U$6898 ( \7119 , \6866 , \6863 );
and \U$6899 ( \7120 , \7119 , \6364 );
or \U$6900 ( \7121 , \6863 , \6870 );
nand \U$6901 ( \7122 , \7121 , \6874 );
nor \U$6902 ( \7123 , \7120 , \7122 );
not \U$6903 ( \7124 , \7123 );
xnor \U$6904 ( \7125 , \7118 , \7124 );
buf \U$6905 ( \7126 , \7125 );
buf \U$6906 ( \7127 , \7126 );
not \U$6907 ( \7128 , \2551 );
nand \U$6908 ( \7129 , \6216 , \7128 );
nor \U$6909 ( \7130 , \6889 , \6886 );
and \U$6910 ( \7131 , \7130 , \6510 );
or \U$6911 ( \7132 , \6886 , \6892 );
nand \U$6912 ( \7133 , \7132 , \6896 );
nor \U$6913 ( \7134 , \7131 , \7133 );
not \U$6914 ( \7135 , \7134 );
xnor \U$6915 ( \7136 , \7129 , \7135 );
buf \U$6916 ( \7137 , \7136 );
buf \U$6917 ( \7138 , \7137 );
not \U$6918 ( \7139 , \2411 );
nand \U$6919 ( \7140 , \6213 , \7139 );
nor \U$6920 ( \7141 , \6911 , \6908 );
and \U$6921 ( \7142 , \7141 , \6601 );
or \U$6922 ( \7143 , \6908 , \6914 );
nand \U$6923 ( \7144 , \7143 , \6918 );
nor \U$6924 ( \7145 , \7142 , \7144 );
not \U$6925 ( \7146 , \7145 );
xnor \U$6926 ( \7147 , \7140 , \7146 );
buf \U$6927 ( \7148 , \7147 );
buf \U$6928 ( \7149 , \7148 );
not \U$6929 ( \7150 , \2264 );
nand \U$6930 ( \7151 , \6211 , \7150 );
nor \U$6931 ( \7152 , \6933 , \6930 );
and \U$6932 ( \7153 , \7152 , \6113 );
or \U$6933 ( \7154 , \6930 , \6936 );
nand \U$6934 ( \7155 , \7154 , \6940 );
nor \U$6935 ( \7156 , \7153 , \7155 );
not \U$6936 ( \7157 , \7156 );
xnor \U$6937 ( \7158 , \7151 , \7157 );
buf \U$6938 ( \7159 , \7158 );
buf \U$6939 ( \7160 , \7159 );
not \U$6940 ( \7161 , \2110 );
nand \U$6941 ( \7162 , \6207 , \7161 );
nor \U$6942 ( \7163 , \6955 , \6952 );
and \U$6943 ( \7164 , \7163 , \6598 );
or \U$6944 ( \7165 , \6952 , \6958 );
nand \U$6945 ( \7166 , \7165 , \6962 );
nor \U$6946 ( \7167 , \7164 , \7166 );
not \U$6947 ( \7168 , \7167 );
xnor \U$6948 ( \7169 , \7162 , \7168 );
buf \U$6949 ( \7170 , \7169 );
buf \U$6950 ( \7171 , \7170 );
not \U$6951 ( \7172 , \1957 );
nand \U$6952 ( \7173 , \6205 , \7172 );
or \U$6953 ( \7174 , \6974 , \6978 );
nand \U$6954 ( \7175 , \7174 , \6982 );
xnor \U$6955 ( \7176 , \7173 , \7175 );
buf \U$6956 ( \7177 , \7176 );
buf \U$6957 ( \7178 , \7177 );
not \U$6958 ( \7179 , \1802 );
nand \U$6959 ( \7180 , \6202 , \7179 );
or \U$6960 ( \7181 , \6994 , \6998 );
nand \U$6961 ( \7182 , \7181 , \7002 );
xnor \U$6962 ( \7183 , \7180 , \7182 );
buf \U$6963 ( \7184 , \7183 );
buf \U$6964 ( \7185 , \7184 );
not \U$6965 ( \7186 , \1649 );
nand \U$6966 ( \7187 , \6200 , \7186 );
xnor \U$6967 ( \7188 , \7187 , \6198 );
buf \U$6968 ( \7189 , \7188 );
buf \U$6969 ( \7190 , \7189 );
not \U$6970 ( \7191 , \5794 );
nand \U$6971 ( \7192 , \6193 , \7191 );
xnor \U$6972 ( \7193 , \7192 , \6412 );
buf \U$6973 ( \7194 , \7193 );
buf \U$6974 ( \7195 , \7194 );
not \U$6975 ( \7196 , \5787 );
nand \U$6976 ( \7197 , \6191 , \7196 );
xnor \U$6977 ( \7198 , \7197 , \6534 );
buf \U$6978 ( \7199 , \7198 );
buf \U$6979 ( \7200 , \7199 );
not \U$6980 ( \7201 , \5772 );
nand \U$6981 ( \7202 , \6188 , \7201 );
xnor \U$6982 ( \7203 , \7202 , \6625 );
buf \U$6983 ( \7204 , \7203 );
buf \U$6984 ( \7205 , \7204 );
not \U$6985 ( \7206 , \5747 );
nand \U$6986 ( \7207 , \6186 , \7206 );
xnor \U$6987 ( \7208 , \7207 , \6686 );
buf \U$6988 ( \7209 , \7208 );
buf \U$6989 ( \7210 , \7209 );
not \U$6990 ( \7211 , \5712 );
nand \U$6991 ( \7212 , \6182 , \7211 );
xnor \U$6992 ( \7213 , \7212 , \6731 );
buf \U$6993 ( \7214 , \7213 );
buf \U$6994 ( \7215 , \7214 );
not \U$6995 ( \7216 , \5667 );
nand \U$6996 ( \7217 , \6180 , \7216 );
xnor \U$6997 ( \7218 , \7217 , \6774 );
buf \U$6998 ( \7219 , \7218 );
buf \U$6999 ( \7220 , \7219 );
not \U$7000 ( \7221 , \5593 );
nand \U$7001 ( \7222 , \6177 , \7221 );
xnor \U$7002 ( \7223 , \7222 , \6817 );
buf \U$7003 ( \7224 , \7223 );
buf \U$7004 ( \7225 , \7224 );
not \U$7005 ( \7226 , \5478 );
nand \U$7006 ( \7227 , \6175 , \7226 );
xnor \U$7007 ( \7228 , \7227 , \6848 );
buf \U$7008 ( \7229 , \7228 );
buf \U$7009 ( \7230 , \7229 );
not \U$7010 ( \7231 , \5364 );
nand \U$7011 ( \7232 , \6170 , \7231 );
xnor \U$7012 ( \7233 , \7232 , \6871 );
buf \U$7013 ( \7234 , \7233 );
buf \U$7014 ( \7235 , \7234 );
not \U$7015 ( \7236 , \5259 );
nand \U$7016 ( \7237 , \6168 , \7236 );
xnor \U$7017 ( \7238 , \7237 , \6893 );
buf \U$7018 ( \7239 , \7238 );
buf \U$7019 ( \7240 , \7239 );
not \U$7020 ( \7241 , \5157 );
nand \U$7021 ( \7242 , \6165 , \7241 );
xnor \U$7022 ( \7243 , \7242 , \6915 );
buf \U$7023 ( \7244 , \7243 );
buf \U$7024 ( \7245 , \7244 );
not \U$7025 ( \7246 , \5062 );
nand \U$7026 ( \7247 , \6163 , \7246 );
xnor \U$7027 ( \7248 , \7247 , \6937 );
buf \U$7028 ( \7249 , \7248 );
buf \U$7029 ( \7250 , \7249 );
not \U$7030 ( \7251 , \4969 );
nand \U$7031 ( \7252 , \6159 , \7251 );
xnor \U$7032 ( \7253 , \7252 , \6959 );
buf \U$7033 ( \7254 , \7253 );
buf \U$7034 ( \7255 , \7254 );
not \U$7035 ( \7256 , \4884 );
nand \U$7036 ( \7257 , \6157 , \7256 );
xnor \U$7037 ( \7258 , \7257 , \6979 );
buf \U$7038 ( \7259 , \7258 );
buf \U$7039 ( \7260 , \7259 );
not \U$7040 ( \7261 , \4802 );
nand \U$7041 ( \7262 , \6154 , \7261 );
xnor \U$7042 ( \7263 , \7262 , \6999 );
buf \U$7043 ( \7264 , \7263 );
buf \U$7044 ( \7265 , \7264 );
not \U$7045 ( \7266 , \4727 );
nand \U$7046 ( \7267 , \6152 , \7266 );
xnor \U$7047 ( \7268 , \7267 , \7015 );
buf \U$7048 ( \7269 , \7268 );
buf \U$7049 ( \7270 , \7269 );
not \U$7050 ( \7271 , \6049 );
nand \U$7051 ( \7272 , \6146 , \7271 );
xnor \U$7052 ( \7273 , \7272 , \7027 );
buf \U$7053 ( \7274 , \7273 );
buf \U$7054 ( \7275 , \7274 );
not \U$7055 ( \7276 , \6042 );
nand \U$7056 ( \7277 , \6144 , \7276 );
xnor \U$7057 ( \7278 , \7277 , \7039 );
buf \U$7058 ( \7279 , \7278 );
buf \U$7059 ( \7280 , \7279 );
not \U$7060 ( \7281 , \6030 );
nand \U$7061 ( \7282 , \6141 , \7281 );
xnor \U$7062 ( \7283 , \7282 , \7051 );
buf \U$7063 ( \7284 , \7283 );
buf \U$7064 ( \7285 , \7284 );
not \U$7065 ( \7286 , \6013 );
nand \U$7066 ( \7287 , \6139 , \7286 );
xnor \U$7067 ( \7288 , \7287 , \7063 );
buf \U$7068 ( \7289 , \7288 );
buf \U$7069 ( \7290 , \7289 );
not \U$7070 ( \7291 , \5984 );
nand \U$7071 ( \7292 , \6135 , \7291 );
xnor \U$7072 ( \7293 , \7292 , \7075 );
buf \U$7073 ( \7294 , \7293 );
buf \U$7074 ( \7295 , \7294 );
not \U$7075 ( \7296 , \5939 );
nand \U$7076 ( \7297 , \6133 , \7296 );
xnor \U$7077 ( \7298 , \7297 , \6765 );
buf \U$7078 ( \7299 , \7298 );
buf \U$7079 ( \7300 , \7299 );
not \U$7080 ( \7301 , \5897 );
nand \U$7081 ( \7302 , \6130 , \7301 );
xnor \U$7082 ( \7303 , \7302 , \6808 );
buf \U$7083 ( \7304 , \7303 );
buf \U$7084 ( \7305 , \7304 );
not \U$7085 ( \7306 , \5862 );
nand \U$7086 ( \7307 , \6128 , \7306 );
xnor \U$7087 ( \7308 , \7307 , \6126 );
buf \U$7088 ( \7309 , \7308 );
buf \U$7089 ( \7310 , \7309 );
not \U$7090 ( \7311 , \6096 );
nand \U$7091 ( \7312 , \6123 , \7311 );
xnor \U$7092 ( \7313 , \7312 , \6364 );
buf \U$7093 ( \7314 , \7313 );
buf \U$7094 ( \7315 , \7314 );
not \U$7095 ( \7316 , \6092 );
nand \U$7096 ( \7317 , \6121 , \7316 );
xnor \U$7097 ( \7318 , \7317 , \6510 );
buf \U$7098 ( \7319 , \7318 );
buf \U$7099 ( \7320 , \7319 );
endmodule

