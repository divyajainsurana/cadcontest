//
// Conformal-LEC Version 19.20-d255 (16-Apr-2020)
//
module top(\s[31] ,\s[30] ,\s[29] ,\s[28] ,\s[27] ,\s[26] ,\s[25] ,\s[24] ,\s[23] ,
        \s[22] ,\s[21] ,\s[20] ,\s[19] ,\s[18] ,\s[17] ,\s[16] ,\s[15] ,\s[14] ,\s[13] ,
        \s[12] ,\s[11] ,\s[10] ,\s[9] ,\s[8] ,\s[7] ,\s[6] ,\s[5] ,\s[4] ,\s[3] ,
        \s[2] ,\s[1] ,\s[0] ,\a[31] ,\a[30] ,\a[29] ,\a[28] ,\a[27] ,\a[26] ,\a[25] ,
        \a[24] ,\a[23] ,\a[22] ,\a[21] ,\a[20] ,\a[19] ,\a[18] ,\a[17] ,\a[16] ,\a[15] ,
        \a[14] ,\a[13] ,\a[12] ,\a[11] ,\a[10] ,\a[9] ,\a[8] ,\a[7] ,\a[6] ,\a[5] ,
        \a[4] ,\a[3] ,\a[2] ,\a[1] ,\a[0] ,\b[31] ,\b[30] ,\b[29] ,\b[28] ,\b[27] ,
        \b[26] ,\b[25] ,\b[24] ,\b[23] ,\b[22] ,\b[21] ,\b[20] ,\b[19] ,\b[18] ,\b[17] ,
        \b[16] ,\b[15] ,\b[14] ,\b[13] ,\b[12] ,\b[11] ,\b[10] ,\b[9] ,\b[8] ,\b[7] ,
        \b[6] ,\b[5] ,\b[4] ,\b[3] ,\b[2] ,\b[1] ,\b[0] ,\c[31] ,\c[30] ,\c[29] ,
        \c[28] ,\c[27] ,\c[26] ,\c[25] ,\c[24] ,\c[23] ,\c[22] ,\c[21] ,\c[20] ,\c[19] ,
        \c[18] ,\c[17] ,\c[16] ,\c[15] ,\c[14] ,\c[13] ,\c[12] ,\c[11] ,\c[10] ,\c[9] ,
        \c[8] ,\c[7] ,\c[6] ,\c[5] ,\c[4] ,\c[3] ,\c[2] ,\c[1] ,\c[0] ,\d[31] ,
        \d[30] ,\d[29] ,\d[28] ,\d[27] ,\d[26] ,\d[25] ,\d[24] ,\d[23] ,\d[22] ,\d[21] ,
        \d[20] ,\d[19] ,\d[18] ,\d[17] ,\d[16] ,\d[15] ,\d[14] ,\d[13] ,\d[12] ,\d[11] ,
        \d[10] ,\d[9] ,\d[8] ,\d[7] ,\d[6] ,\d[5] ,\d[4] ,\d[3] ,\d[2] ,\d[1] ,
        \d[0] ,\o[31] ,\o[30] ,\o[29] ,\o[28] ,\o[27] ,\o[26] ,\o[25] ,\o[24] ,\o[23] ,
        \o[22] ,\o[21] ,\o[20] ,\o[19] ,\o[18] ,\o[17] ,\o[16] ,\o[15] ,\o[14] ,\o[13] ,
        \o[12] ,\o[11] ,\o[10] ,\o[9] ,\o[8] ,\o[7] ,\o[6] ,\o[5] ,\o[4] ,\o[3] ,
        \o[2] ,\o[1] ,\o[0] );
input \s[31] ,\s[30] ,\s[29] ,\s[28] ,\s[27] ,\s[26] ,\s[25] ,\s[24] ,\s[23] ,
        \s[22] ,\s[21] ,\s[20] ,\s[19] ,\s[18] ,\s[17] ,\s[16] ,\s[15] ,\s[14] ,\s[13] ,
        \s[12] ,\s[11] ,\s[10] ,\s[9] ,\s[8] ,\s[7] ,\s[6] ,\s[5] ,\s[4] ,\s[3] ,
        \s[2] ,\s[1] ,\s[0] ,\a[31] ,\a[30] ,\a[29] ,\a[28] ,\a[27] ,\a[26] ,\a[25] ,
        \a[24] ,\a[23] ,\a[22] ,\a[21] ,\a[20] ,\a[19] ,\a[18] ,\a[17] ,\a[16] ,\a[15] ,
        \a[14] ,\a[13] ,\a[12] ,\a[11] ,\a[10] ,\a[9] ,\a[8] ,\a[7] ,\a[6] ,\a[5] ,
        \a[4] ,\a[3] ,\a[2] ,\a[1] ,\a[0] ,\b[31] ,\b[30] ,\b[29] ,\b[28] ,\b[27] ,
        \b[26] ,\b[25] ,\b[24] ,\b[23] ,\b[22] ,\b[21] ,\b[20] ,\b[19] ,\b[18] ,\b[17] ,
        \b[16] ,\b[15] ,\b[14] ,\b[13] ,\b[12] ,\b[11] ,\b[10] ,\b[9] ,\b[8] ,\b[7] ,
        \b[6] ,\b[5] ,\b[4] ,\b[3] ,\b[2] ,\b[1] ,\b[0] ,\c[31] ,\c[30] ,\c[29] ,
        \c[28] ,\c[27] ,\c[26] ,\c[25] ,\c[24] ,\c[23] ,\c[22] ,\c[21] ,\c[20] ,\c[19] ,
        \c[18] ,\c[17] ,\c[16] ,\c[15] ,\c[14] ,\c[13] ,\c[12] ,\c[11] ,\c[10] ,\c[9] ,
        \c[8] ,\c[7] ,\c[6] ,\c[5] ,\c[4] ,\c[3] ,\c[2] ,\c[1] ,\c[0] ,\d[31] ,
        \d[30] ,\d[29] ,\d[28] ,\d[27] ,\d[26] ,\d[25] ,\d[24] ,\d[23] ,\d[22] ,\d[21] ,
        \d[20] ,\d[19] ,\d[18] ,\d[17] ,\d[16] ,\d[15] ,\d[14] ,\d[13] ,\d[12] ,\d[11] ,
        \d[10] ,\d[9] ,\d[8] ,\d[7] ,\d[6] ,\d[5] ,\d[4] ,\d[3] ,\d[2] ,\d[1] ,
        \d[0] ;
output \o[31] ,\o[30] ,\o[29] ,\o[28] ,\o[27] ,\o[26] ,\o[25] ,\o[24] ,\o[23] ,
        \o[22] ,\o[21] ,\o[20] ,\o[19] ,\o[18] ,\o[17] ,\o[16] ,\o[15] ,\o[14] ,\o[13] ,
        \o[12] ,\o[11] ,\o[10] ,\o[9] ,\o[8] ,\o[7] ,\o[6] ,\o[5] ,\o[4] ,\o[3] ,
        \o[2] ,\o[1] ,\o[0] ;

wire \193_ZERO , \194_ONE , \195 , \196 , \197 , \198 , \199 , \200 , \201 ,
         \202 , \203 , \204 , \205 , \206 , \207 , \208 , \209 , \210 , \211 ,
         \212 , \213 , \214 , \215 , \216 , \217 , \218 , \219 , \220 , \221 ,
         \222 , \223 , \224 , \225 , \226 , \227 , \228 , \229 , \230 , \231 ,
         \232 , \233 , \234 , \235 , \236 , \237 , \238 , \239 , \240 , \241 ,
         \242 , \243 , \244 , \245 , \246 , \247 , \248 , \249 , \250 , \251 ,
         \252 , \253 , \254 , \255 , \256 , \257 , \258 , \259 , \260 , \261 ,
         \262 , \263 , \264 , \265 , \266 , \267 , \268 , \269 , \270 , \271 ,
         \272 , \273 , \274 , \275 , \276 , \277 , \278 , \279 , \280 , \281 ,
         \282 , \283 , \284 , \285 , \286 , \287 , \288 , \289 , \290 , \291 ,
         \292 , \293 , \294 , \295 , \296 , \297 , \298 , \299 , \300 , \301 ,
         \302 , \303 , \304 , \305 , \306 , \307 , \308 , \309 , \310 , \311 ,
         \312 , \313 , \314 , \315 , \316 , \317 , \318 , \319 , \320 , \321 ,
         \322 , \323 , \324 , \325 , \326 , \327 , \328 , \329 , \330 , \331 ,
         \332 , \333 , \334 , \335 , \336 , \337 , \338 , \339 , \340 , \341 ,
         \342 , \343 , \344 , \345 , \346 , \347 , \348 , \349 , \350 , \351 ,
         \352 , \353 , \354 , \355 , \356 , \357 , \358 , \359 , \360 , \361 ,
         \362 , \363 , \364 , \365 , \366 , \367 , \368 , \369 , \370 , \371 ,
         \372 , \373 , \374 , \375 , \376 , \377 , \378 , \379 , \380 , \381 ,
         \382 , \383 , \384 , \385 , \386 , \387 , \388 , \389 , \390 , \391 ,
         \392 , \393 , \394 , \395 , \396 , \397 , \398 , \399 , \400 , \401 ,
         \402 , \403 , \404 , \405 , \406 , \407 , \408 , \409 , \410 , \411 ,
         \412 , \413 , \414 , \415 , \416 , \417 , \418 , \419 , \420 , \421 ,
         \422 , \423 , \424 , \425 , \426 , \427 , \428 , \429 , \430 , \431 ,
         \432 , \433 , \434 , \435 , \436 , \437 , \438 , \439 , \440 , \441 ,
         \442 , \443 , \444 , \445 , \446 , \447 , \448 , \449 , \450 , \451 ,
         \452 , \453 , \454 , \455 , \456 , \457 , \458 , \459 , \460 , \461 ,
         \462 , \463 , \464 , \465 , \466 , \467 , \468 , \469 , \470 , \471 ,
         \472 , \473 , \474 , \475 , \476 , \477 , \478 , \479 , \480 , \481 ,
         \482 , \483 , \484 , \485 , \486 , \487 , \488 , \489 , \490 , \491 ,
         \492 , \493 , \494 , \495 , \496 , \497 , \498 , \499 , \500 , \501 ,
         \502 , \503 , \504 , \505 , \506 , \507 , \508 , \509 , \510 , \511 ,
         \512 , \513 , \514 , \515 , \516 , \517 , \518 , \519 , \520 , \521 ,
         \522 , \523 , \524 , \525 , \526 , \527 , \528 , \529 , \530 , \531 ,
         \532 , \533 , \534 , \535 , \536 , \537 , \538 , \539 , \540 , \541 ,
         \542 , \543 , \544 , \545 , \546 , \547 , \548 , \549 , \550 , \551 ,
         \552 , \553 , \554 , \555 , \556 , \557 , \558 , \559 , \560 , \561 ,
         \562 , \563 , \564 , \565 , \566 , \567 , \568 , \569 , \570 , \571 ,
         \572 , \573 , \574 , \575 , \576 , \577 , \578 , \579 , \580 , \581 ,
         \582 , \583 , \584 , \585 , \586 , \587 , \588 , \589 , \590 , \591 ,
         \592 , \593 , \594 , \595 , \596 , \597 , \598 , \599 , \600 , \601 ,
         \602 , \603 , \604 , \605 , \606 , \607 , \608 , \609 , \610 , \611 ,
         \612 , \613 , \614 , \615 , \616 , \617 , \618 , \619 , \620 , \621 ,
         \622 , \623 , \624 , \625 , \626 , \627 , \628 , \629 , \630 , \631 ,
         \632 , \633 , \634 , \635 , \636 , \637 , \638 , \639 , \640 , \641 ,
         \642 , \643 , \644 , \645 , \646 , \647 , \648 , \649 , \650 , \651 ,
         \652 , \653 , \654 , \655 , \656 , \657 , \658 , \659 , \660 , \661 ,
         \662 , \663 , \664 , \665 , \666 , \667 , \668 , \669 , \670 , \671 ,
         \672 , \673 , \674 , \675 , \676 , \677 , \678 , \679 , \680 , \681 ,
         \682 , \683 , \684 , \685 , \686 , \687 , \688 , \689 , \690 , \691 ,
         \692 , \693 , \694 , \695 , \696 , \697 , \698 , \699 , \700 , \701 ,
         \702 , \703 , \704 , \705 , \706 , \707 , \708 , \709 , \710 , \711 ,
         \712 , \713 , \714 , \715 , \716 , \717 , \718 , \719 , \720 , \721 ,
         \722 , \723 , \724 , \725 , \726 , \727 , \728 , \729 , \730 , \731 ,
         \732 , \733 , \734 , \735 , \736 , \737 , \738 , \739 , \740 , \741 ,
         \742 , \743 , \744 , \745 , \746 , \747 , \748 , \749 , \750 , \751 ,
         \752 , \753 , \754 , \755 , \756 , \757 , \758 , \759 , \760 , \761 ,
         \762 , \763 , \764 , \765 , \766 , \767 , \768 , \769 , \770 , \771 ,
         \772 , \773 , \774 , \775 , \776 , \777 , \778 , \779 , \780 , \781 ,
         \782 , \783 , \784 , \785 , \786 , \787 , \788 , \789 , \790 , \791 ,
         \792 , \793 , \794 , \795 , \796 , \797 , \798 , \799 , \800 , \801 ,
         \802 , \803 , \804 , \805 , \806 , \807 , \808 , \809 , \810 , \811 ,
         \812 , \813 , \814 , \815 , \816 , \817 , \818 , \819 , \820 , \821 ,
         \822 , \823 , \824 , \825 , \826 , \827 , \828 , \829 , \830 , \831 ,
         \832 , \833 , \834 , \835 , \836 , \837 , \838 , \839 , \840 , \841 ,
         \842 , \843 , \844 , \845 , \846 , \847 , \848 , \849 , \850 , \851 ,
         \852 , \853 , \854 , \855 , \856 , \857 , \858 , \859 , \860 , \861 ,
         \862 , \863 , \864 , \865 , \866 , \867 , \868 , \869 , \870 , \871 ,
         \872 , \873 , \874 , \875 , \876 , \877 , \878 , \879 , \880 , \881 ,
         \882 , \883 , \884 , \885 , \886 , \887 , \888 , \889 , \890 , \891 ,
         \892 , \893 , \894 , \895 , \896 , \897 , \898 , \899 , \900 , \901 ,
         \902 , \903 , \904 , \905 , \906 , \907 , \908 , \909 , \910 , \911 ,
         \912 , \913 , \914 , \915 , \916 , \917 , \918 , \919 , \920 , \921 ,
         \922 , \923 , \924 , \925 , \926 , \927 , \928 , \929 , \930 , \931 ,
         \932 , \933 , \934 , \935 , \936 , \937 , \938 , \939 , \940 , \941 ,
         \942 , \943 , \944 , \945 , \946 , \947 , \948 , \949 , \950 , \951 ,
         \952 , \953 , \954 , \955 , \956 , \957 , \958 , \959 , \960 , \961 ,
         \962 , \963 , \964 , \965 , \966 , \967 , \968 , \969 , \970 , \971 ,
         \972 , \973 , \974 , \975 , \976 , \977 , \978 , \979 , \980 , \981 ,
         \982 , \983 , \984 , \985 , \986 , \987 , \988 , \989 , \990 , \991 ,
         \992 , \993 , \994 , \995 , \996 , \997 , \998 , \999 , \1000 , \1001 ,
         \1002 , \1003 , \1004 , \1005 , \1006 , \1007 , \1008 , \1009 , \1010 , \1011 ,
         \1012 , \1013 , \1014 , \1015 , \1016 , \1017 , \1018 , \1019 , \1020 , \1021 ,
         \1022 , \1023 , \1024 , \1025 , \1026 , \1027 , \1028 , \1029 , \1030 , \1031 ,
         \1032 , \1033 , \1034 , \1035 , \1036 , \1037 , \1038 , \1039 , \1040 , \1041 ,
         \1042 , \1043 , \1044 , \1045 , \1046 , \1047 , \1048 , \1049 , \1050 , \1051 ,
         \1052 , \1053 , \1054 , \1055 , \1056 , \1057 , \1058 , \1059 , \1060 , \1061 ,
         \1062 , \1063 , \1064 , \1065 , \1066 , \1067 , \1068 , \1069 , \1070 , \1071 ,
         \1072 , \1073 , \1074 , \1075 , \1076 , \1077 , \1078 , \1079 , \1080 , \1081 ,
         \1082 , \1083 , \1084 , \1085 , \1086 , \1087 , \1088 , \1089 , \1090 , \1091 ,
         \1092 , \1093 , \1094 , \1095 , \1096 , \1097 , \1098 , \1099 , \1100 , \1101 ,
         \1102 , \1103 , \1104 , \1105 , \1106 , \1107 , \1108 , \1109 , \1110 , \1111 ,
         \1112 , \1113 , \1114 , \1115 , \1116 , \1117 , \1118 , \1119 , \1120 , \1121 ,
         \1122 , \1123 , \1124 , \1125 , \1126 , \1127 , \1128 , \1129 , \1130 , \1131 ,
         \1132 , \1133 , \1134 , \1135 , \1136 , \1137 , \1138 , \1139 , \1140 , \1141 ,
         \1142 , \1143 , \1144 , \1145 , \1146 , \1147 , \1148 , \1149 , \1150 , \1151 ,
         \1152 , \1153 , \1154 , \1155 , \1156 , \1157 , \1158 , \1159 , \1160 , \1161 ,
         \1162 , \1163 , \1164 , \1165 , \1166 , \1167 , \1168 , \1169 , \1170 , \1171 ,
         \1172 , \1173 , \1174 , \1175 , \1176 , \1177 , \1178 , \1179 , \1180 , \1181 ,
         \1182 , \1183 , \1184 , \1185 , \1186 , \1187 , \1188 , \1189 , \1190 , \1191 ,
         \1192 , \1193 , \1194 , \1195 , \1196 , \1197 , \1198 , \1199 , \1200 , \1201 ,
         \1202 , \1203 , \1204 , \1205 , \1206 , \1207 , \1208 , \1209 , \1210 , \1211 ,
         \1212 , \1213 , \1214 , \1215 , \1216 , \1217 , \1218 , \1219 , \1220 , \1221 ,
         \1222 , \1223 , \1224 , \1225 , \1226 , \1227 , \1228 , \1229 , \1230 , \1231 ,
         \1232 , \1233 , \1234 , \1235 , \1236 , \1237 , \1238 , \1239 , \1240 , \1241 ,
         \1242 , \1243 , \1244 , \1245 , \1246 , \1247 , \1248 , \1249 , \1250 , \1251 ,
         \1252 , \1253 , \1254 , \1255 , \1256 , \1257 , \1258 , \1259 , \1260 , \1261 ,
         \1262 , \1263 , \1264 , \1265 , \1266 , \1267 , \1268 , \1269 , \1270 , \1271 ,
         \1272 , \1273 , \1274 , \1275 , \1276 , \1277 , \1278 , \1279 , \1280 , \1281 ,
         \1282 , \1283 , \1284 , \1285 , \1286 , \1287 , \1288 , \1289 , \1290 , \1291 ,
         \1292 , \1293 , \1294 , \1295 , \1296 , \1297 , \1298 , \1299 , \1300 , \1301 ,
         \1302 , \1303 , \1304 , \1305 , \1306 , \1307 , \1308 , \1309 , \1310 , \1311 ,
         \1312 , \1313 , \1314 , \1315 , \1316 , \1317 , \1318 , \1319 , \1320 , \1321 ,
         \1322 , \1323 , \1324 , \1325 , \1326 , \1327 , \1328 , \1329 , \1330 , \1331 ,
         \1332 , \1333 , \1334 , \1335 , \1336 , \1337 , \1338 , \1339 , \1340 , \1341 ,
         \1342 , \1343 , \1344 , \1345 , \1346 , \1347 , \1348 , \1349 , \1350 , \1351 ,
         \1352 , \1353 , \1354 , \1355 , \1356 , \1357 , \1358 , \1359 , \1360 , \1361 ,
         \1362 , \1363 , \1364 , \1365 , \1366 , \1367 , \1368 , \1369 , \1370 , \1371 ,
         \1372 , \1373 , \1374 , \1375 , \1376 , \1377 , \1378 , \1379 , \1380 , \1381 ,
         \1382 , \1383 , \1384 , \1385 , \1386 , \1387 , \1388 , \1389 , \1390 , \1391 ,
         \1392 , \1393 , \1394 , \1395 , \1396 , \1397 , \1398 , \1399 , \1400 , \1401 ,
         \1402 , \1403 , \1404 , \1405 , \1406 , \1407 , \1408 , \1409 , \1410 , \1411 ,
         \1412 , \1413 , \1414 , \1415 , \1416 , \1417 , \1418 , \1419 , \1420 , \1421 ,
         \1422 , \1423 , \1424 , \1425 , \1426 , \1427 , \1428 , \1429 , \1430 , \1431 ,
         \1432 , \1433 , \1434 , \1435 , \1436 , \1437 , \1438 , \1439 , \1440 , \1441 ,
         \1442 , \1443 , \1444 , \1445 , \1446 , \1447 , \1448 , \1449 , \1450 , \1451 ,
         \1452 , \1453 , \1454 , \1455 , \1456 , \1457 , \1458 , \1459 , \1460 , \1461 ,
         \1462 , \1463 , \1464 , \1465 , \1466 , \1467 , \1468 , \1469 , \1470 , \1471 ,
         \1472 , \1473 , \1474 , \1475 , \1476 , \1477 , \1478 , \1479 , \1480 , \1481 ,
         \1482 , \1483 , \1484 , \1485 , \1486 , \1487 , \1488 , \1489 , \1490 , \1491 ,
         \1492 , \1493 , \1494 , \1495 , \1496 , \1497 , \1498 , \1499 , \1500 , \1501 ,
         \1502 , \1503 , \1504 , \1505 , \1506 , \1507 , \1508 , \1509 , \1510 , \1511 ,
         \1512 , \1513 , \1514 , \1515 , \1516 , \1517 , \1518 , \1519 , \1520 , \1521 ,
         \1522 , \1523 , \1524 , \1525 , \1526 , \1527 , \1528 , \1529 , \1530 , \1531 ,
         \1532 , \1533 , \1534 , \1535 , \1536 , \1537 , \1538 , \1539 , \1540 , \1541 ,
         \1542 , \1543 , \1544 , \1545 , \1546 , \1547 , \1548 , \1549 , \1550 , \1551 ,
         \1552 , \1553 , \1554 , \1555 , \1556 , \1557 , \1558 , \1559 , \1560 , \1561 ,
         \1562 , \1563 , \1564 , \1565 , \1566 , \1567 , \1568 , \1569 , \1570 , \1571 ,
         \1572 , \1573 , \1574 , \1575 , \1576 , \1577 , \1578 , \1579 , \1580 , \1581 ,
         \1582 , \1583 , \1584 , \1585 , \1586 , \1587 , \1588 , \1589 , \1590 , \1591 ,
         \1592 , \1593 , \1594 , \1595 , \1596 , \1597 , \1598 , \1599 , \1600 , \1601 ,
         \1602 , \1603 , \1604 , \1605 , \1606 , \1607 , \1608 , \1609 , \1610 , \1611 ,
         \1612 , \1613 , \1614 , \1615 , \1616 , \1617 , \1618 , \1619 , \1620 , \1621 ,
         \1622 , \1623 , \1624 , \1625 , \1626 , \1627 , \1628 , \1629 , \1630 , \1631 ,
         \1632 , \1633 , \1634 , \1635 , \1636 , \1637 , \1638 , \1639 , \1640 , \1641 ,
         \1642 , \1643 , \1644 , \1645 , \1646 , \1647 , \1648 , \1649 , \1650 , \1651 ,
         \1652 , \1653 , \1654 , \1655 , \1656 , \1657 , \1658 , \1659 , \1660 , \1661 ,
         \1662 , \1663 , \1664 , \1665 , \1666 , \1667 , \1668 , \1669 , \1670 , \1671 ,
         \1672 , \1673 , \1674 , \1675 , \1676 , \1677 , \1678 , \1679 , \1680 , \1681 ,
         \1682 , \1683 , \1684 , \1685 , \1686 , \1687 , \1688 , \1689 , \1690 , \1691 ,
         \1692 , \1693 , \1694 , \1695 , \1696 , \1697 , \1698 , \1699 , \1700 , \1701 ,
         \1702 , \1703 , \1704 , \1705 , \1706 , \1707 , \1708 , \1709 , \1710 , \1711 ,
         \1712 , \1713 , \1714 , \1715 , \1716 , \1717 , \1718 , \1719 , \1720 , \1721 ,
         \1722 , \1723 , \1724 , \1725 , \1726 , \1727 , \1728 , \1729 , \1730 , \1731 ,
         \1732 , \1733 , \1734 , \1735 , \1736 , \1737 , \1738 , \1739 , \1740 , \1741 ,
         \1742 , \1743 , \1744 , \1745 , \1746 , \1747 , \1748 , \1749 , \1750 , \1751 ,
         \1752 , \1753 , \1754 , \1755 , \1756 , \1757 , \1758 , \1759 , \1760 , \1761 ,
         \1762 , \1763 , \1764 , \1765 , \1766 , \1767 , \1768 , \1769 , \1770 , \1771 ,
         \1772 , \1773 , \1774 , \1775 , \1776 , \1777 , \1778 , \1779 , \1780 , \1781 ,
         \1782 , \1783 , \1784 , \1785 , \1786 , \1787 , \1788 , \1789 , \1790 , \1791 ,
         \1792 , \1793 , \1794 , \1795 , \1796 , \1797 , \1798 , \1799 , \1800 , \1801 ,
         \1802 , \1803 , \1804 , \1805 , \1806 , \1807 , \1808 , \1809 , \1810 , \1811 ,
         \1812 , \1813 , \1814 , \1815 , \1816 , \1817 , \1818 , \1819 , \1820 , \1821 ,
         \1822 , \1823 , \1824 , \1825 , \1826 , \1827 , \1828 , \1829 , \1830 , \1831 ,
         \1832 , \1833 , \1834 , \1835 , \1836 , \1837 , \1838 , \1839 , \1840 , \1841 ,
         \1842 , \1843 , \1844 , \1845 , \1846 , \1847 , \1848 , \1849 , \1850 , \1851 ,
         \1852 , \1853 , \1854 , \1855 , \1856 , \1857 , \1858 , \1859 , \1860 , \1861 ,
         \1862 , \1863 , \1864 , \1865 , \1866 , \1867 , \1868 , \1869 , \1870 , \1871 ,
         \1872 , \1873 , \1874 , \1875 , \1876 , \1877 , \1878 , \1879 , \1880 , \1881 ,
         \1882 , \1883 , \1884 , \1885 , \1886 , \1887 , \1888 , \1889 , \1890 , \1891 ,
         \1892 , \1893 , \1894 , \1895 , \1896 , \1897 , \1898 , \1899 , \1900 , \1901 ,
         \1902 , \1903 , \1904 , \1905 , \1906 , \1907 , \1908 , \1909 , \1910 , \1911 ,
         \1912 , \1913 , \1914 , \1915 , \1916 , \1917 , \1918 , \1919 , \1920 , \1921 ,
         \1922 , \1923 , \1924 , \1925 , \1926 , \1927 , \1928 , \1929 , \1930 , \1931 ,
         \1932 , \1933 , \1934 , \1935 , \1936 , \1937 , \1938 , \1939 , \1940 , \1941 ,
         \1942 , \1943 , \1944 , \1945 , \1946 , \1947 , \1948 , \1949 , \1950 , \1951 ,
         \1952 , \1953 , \1954 , \1955 , \1956 , \1957 , \1958 , \1959 , \1960 , \1961 ,
         \1962 , \1963 , \1964 , \1965 , \1966 , \1967 , \1968 , \1969 , \1970 , \1971 ,
         \1972 , \1973 , \1974 , \1975 , \1976 , \1977 , \1978 , \1979 , \1980 , \1981 ,
         \1982 , \1983 , \1984 , \1985 , \1986 , \1987 , \1988 , \1989 , \1990 , \1991 ,
         \1992 , \1993 , \1994 , \1995 , \1996 , \1997 , \1998 , \1999 , \2000 , \2001 ,
         \2002 , \2003 , \2004 , \2005 , \2006 , \2007 , \2008 , \2009 , \2010 , \2011 ,
         \2012 , \2013 , \2014 , \2015 , \2016 , \2017 , \2018 , \2019 , \2020 , \2021 ,
         \2022 , \2023 , \2024 , \2025 , \2026 , \2027 , \2028 , \2029 , \2030 , \2031 ,
         \2032 , \2033 , \2034 , \2035 , \2036 , \2037 , \2038 , \2039 , \2040 , \2041 ,
         \2042 , \2043 , \2044 , \2045 , \2046 , \2047 , \2048 , \2049 , \2050 , \2051 ,
         \2052 , \2053 , \2054 , \2055 , \2056 , \2057 , \2058 , \2059 , \2060 , \2061 ,
         \2062 , \2063 , \2064 , \2065 , \2066 , \2067 , \2068 , \2069 , \2070 , \2071 ,
         \2072 , \2073 , \2074 , \2075 , \2076 , \2077 , \2078 , \2079 , \2080 , \2081 ,
         \2082 , \2083 , \2084 , \2085 , \2086 , \2087 , \2088 , \2089 , \2090 , \2091 ,
         \2092 , \2093 , \2094 , \2095 , \2096 , \2097 , \2098 , \2099 , \2100 , \2101 ,
         \2102 , \2103 , \2104 , \2105 , \2106 , \2107 , \2108 , \2109 , \2110 , \2111 ,
         \2112 , \2113 , \2114 , \2115 , \2116 , \2117 , \2118 , \2119 , \2120 , \2121 ,
         \2122 , \2123 , \2124 , \2125 , \2126 , \2127 , \2128 , \2129 , \2130 , \2131 ,
         \2132 , \2133 , \2134 , \2135 , \2136 , \2137 , \2138 , \2139 , \2140 , \2141 ,
         \2142 , \2143 , \2144 , \2145 , \2146 , \2147 , \2148 , \2149 , \2150 , \2151 ,
         \2152 , \2153 , \2154 , \2155 , \2156 , \2157 , \2158 , \2159 , \2160 , \2161 ,
         \2162 , \2163 , \2164 , \2165 , \2166 , \2167 , \2168 , \2169 , \2170 , \2171 ,
         \2172 , \2173 , \2174 , \2175 , \2176 , \2177 , \2178 , \2179 , \2180 , \2181 ,
         \2182 , \2183 , \2184 , \2185 , \2186 , \2187 , \2188 , \2189 , \2190 , \2191 ,
         \2192 , \2193 , \2194 , \2195 , \2196 , \2197 , \2198 , \2199 , \2200 , \2201 ,
         \2202 , \2203 , \2204 , \2205 , \2206 , \2207 , \2208 , \2209 , \2210 , \2211 ,
         \2212 , \2213 , \2214 , \2215 , \2216 , \2217 , \2218 , \2219 , \2220 , \2221 ,
         \2222 , \2223 , \2224 , \2225 , \2226 , \2227 , \2228 , \2229 , \2230 , \2231 ,
         \2232 , \2233 , \2234 , \2235 , \2236 , \2237 , \2238 , \2239 , \2240 , \2241 ,
         \2242 , \2243 , \2244 , \2245 , \2246 , \2247 , \2248 , \2249 , \2250 , \2251 ,
         \2252 , \2253 , \2254 , \2255 , \2256 , \2257 , \2258 , \2259 , \2260 , \2261 ,
         \2262 , \2263 , \2264 , \2265 , \2266 , \2267 , \2268 , \2269 , \2270 , \2271 ,
         \2272 , \2273 , \2274 , \2275 , \2276 , \2277 , \2278 , \2279 , \2280 , \2281 ,
         \2282 , \2283 , \2284 , \2285 , \2286 , \2287 , \2288 , \2289 , \2290 , \2291 ,
         \2292 , \2293 , \2294 , \2295 , \2296 , \2297 , \2298 , \2299 , \2300 , \2301 ,
         \2302 , \2303 , \2304 , \2305 , \2306 , \2307 , \2308 , \2309 , \2310 , \2311 ,
         \2312 , \2313 , \2314 , \2315 , \2316 , \2317 , \2318 , \2319 , \2320 , \2321 ,
         \2322 , \2323 , \2324 , \2325 , \2326 , \2327 , \2328 , \2329 , \2330 , \2331 ,
         \2332 , \2333 , \2334 , \2335 , \2336 , \2337 , \2338 , \2339 , \2340 , \2341 ,
         \2342 , \2343 , \2344 , \2345 , \2346 , \2347 , \2348 , \2349 , \2350 , \2351 ,
         \2352 , \2353 , \2354 , \2355 , \2356 , \2357 , \2358 , \2359 , \2360 , \2361 ,
         \2362 , \2363 , \2364 , \2365 , \2366 , \2367 , \2368 , \2369 , \2370 , \2371 ,
         \2372 , \2373 , \2374 , \2375 , \2376 , \2377 , \2378 , \2379 , \2380 , \2381 ,
         \2382 , \2383 , \2384 , \2385 , \2386 , \2387 , \2388 , \2389 , \2390 , \2391 ,
         \2392 , \2393 , \2394 , \2395 , \2396 , \2397 , \2398 , \2399 , \2400 , \2401 ,
         \2402 , \2403 , \2404 , \2405 , \2406 , \2407 , \2408 , \2409 , \2410 , \2411 ,
         \2412 , \2413 , \2414 , \2415 , \2416 , \2417 , \2418 , \2419 , \2420 , \2421 ,
         \2422 , \2423 , \2424 , \2425 , \2426 , \2427 , \2428 , \2429 , \2430 , \2431 ,
         \2432 , \2433 , \2434 , \2435 , \2436 , \2437 , \2438 , \2439 , \2440 , \2441 ,
         \2442 , \2443 , \2444 , \2445 , \2446 , \2447 , \2448 , \2449 , \2450 , \2451 ,
         \2452 , \2453 , \2454 , \2455 , \2456 , \2457 , \2458 , \2459 , \2460 , \2461 ,
         \2462 , \2463 , \2464 , \2465 , \2466 , \2467 , \2468 , \2469 , \2470 , \2471 ,
         \2472 , \2473 , \2474 , \2475 , \2476 , \2477 , \2478 , \2479 , \2480 , \2481 ,
         \2482 , \2483 , \2484 , \2485 , \2486 , \2487 , \2488 , \2489 , \2490 , \2491 ,
         \2492 , \2493 , \2494 , \2495 , \2496 , \2497 , \2498 , \2499 , \2500 , \2501 ,
         \2502 , \2503 , \2504 , \2505 , \2506 , \2507 , \2508 , \2509 , \2510 , \2511 ,
         \2512 , \2513 , \2514 , \2515 , \2516 , \2517 , \2518 , \2519 , \2520 , \2521 ,
         \2522 , \2523 , \2524 , \2525 , \2526 , \2527 , \2528 , \2529 , \2530 , \2531 ,
         \2532 , \2533 , \2534 , \2535 , \2536 , \2537 , \2538 , \2539 , \2540 , \2541 ,
         \2542 , \2543 , \2544 , \2545 , \2546 , \2547 , \2548 , \2549 , \2550 , \2551 ,
         \2552 , \2553 , \2554 , \2555 , \2556 , \2557 , \2558 , \2559 , \2560 , \2561 ,
         \2562 , \2563 , \2564 , \2565 , \2566 , \2567 , \2568 , \2569 , \2570 , \2571 ,
         \2572 , \2573 , \2574 , \2575 , \2576 , \2577 , \2578 , \2579 , \2580 , \2581 ,
         \2582 , \2583 , \2584 , \2585 , \2586 , \2587 , \2588 , \2589 , \2590 , \2591 ,
         \2592 , \2593 , \2594 , \2595 , \2596 , \2597 , \2598 , \2599 , \2600 , \2601 ,
         \2602 , \2603 , \2604 , \2605 , \2606 , \2607 , \2608 , \2609 , \2610 , \2611 ,
         \2612 , \2613 , \2614 , \2615 , \2616 , \2617 , \2618 , \2619 , \2620 , \2621 ,
         \2622 , \2623 , \2624 , \2625 , \2626 , \2627 , \2628 , \2629 , \2630 , \2631 ,
         \2632 , \2633 , \2634 , \2635 , \2636 , \2637 , \2638 , \2639 , \2640 , \2641 ,
         \2642 , \2643 , \2644 , \2645 , \2646 , \2647 , \2648 , \2649 , \2650 , \2651 ,
         \2652 , \2653 , \2654 , \2655 , \2656 , \2657 , \2658 , \2659 , \2660 , \2661 ,
         \2662 , \2663 , \2664 , \2665 , \2666 , \2667 , \2668 , \2669 , \2670 , \2671 ,
         \2672 , \2673 , \2674 , \2675 , \2676 , \2677 , \2678 , \2679 , \2680 , \2681 ,
         \2682 , \2683 , \2684 , \2685 , \2686 , \2687 , \2688 , \2689 , \2690 , \2691 ,
         \2692 , \2693 , \2694 , \2695 , \2696 , \2697 , \2698 , \2699 , \2700 , \2701 ,
         \2702 , \2703 , \2704 , \2705 , \2706 , \2707 , \2708 , \2709 , \2710 , \2711 ,
         \2712 , \2713 , \2714 , \2715 , \2716 , \2717 , \2718 , \2719 , \2720 , \2721 ,
         \2722 , \2723 , \2724 , \2725 , \2726 , \2727 , \2728 , \2729 , \2730 , \2731 ,
         \2732 , \2733 , \2734 , \2735 , \2736 , \2737 , \2738 , \2739 , \2740 , \2741 ,
         \2742 , \2743 , \2744 , \2745 , \2746 , \2747 , \2748 , \2749 , \2750 , \2751 ,
         \2752 , \2753 , \2754 , \2755 , \2756 , \2757 , \2758 , \2759 , \2760 , \2761 ,
         \2762 , \2763 , \2764 , \2765 , \2766 , \2767 , \2768 , \2769 , \2770 , \2771 ,
         \2772 , \2773 , \2774 , \2775 , \2776 , \2777 , \2778 , \2779 , \2780 , \2781 ,
         \2782 , \2783 , \2784 , \2785 , \2786 , \2787 , \2788 , \2789 , \2790 , \2791 ,
         \2792 , \2793 , \2794 , \2795 , \2796 , \2797 , \2798 , \2799 , \2800 , \2801 ,
         \2802 , \2803 , \2804 , \2805 , \2806 , \2807 , \2808 , \2809 , \2810 , \2811 ,
         \2812 , \2813 , \2814 , \2815 , \2816 , \2817 , \2818 , \2819 , \2820 , \2821 ,
         \2822 , \2823 , \2824 , \2825 , \2826 , \2827 , \2828 , \2829 , \2830 , \2831 ,
         \2832 , \2833 , \2834 , \2835 , \2836 , \2837 , \2838 , \2839 , \2840 , \2841 ,
         \2842 , \2843 , \2844 , \2845 , \2846 , \2847 , \2848 , \2849 , \2850 , \2851 ,
         \2852 , \2853 , \2854 , \2855 , \2856 , \2857 , \2858 , \2859 , \2860 , \2861 ,
         \2862 , \2863 , \2864 , \2865 , \2866 , \2867 , \2868 , \2869 , \2870 , \2871 ,
         \2872 , \2873 , \2874 , \2875 , \2876 , \2877 , \2878 , \2879 , \2880 , \2881 ,
         \2882 , \2883 , \2884 , \2885 , \2886 , \2887 , \2888 , \2889 , \2890 , \2891 ,
         \2892 , \2893 , \2894 , \2895 , \2896 , \2897 , \2898 , \2899 , \2900 , \2901 ,
         \2902 , \2903 , \2904 , \2905 , \2906 , \2907 , \2908 , \2909 , \2910 , \2911 ,
         \2912 , \2913 , \2914 , \2915 , \2916 , \2917 , \2918 , \2919 , \2920 , \2921 ,
         \2922 , \2923 , \2924 , \2925 , \2926 , \2927 , \2928 , \2929 , \2930 , \2931 ,
         \2932 , \2933 , \2934 , \2935 , \2936 , \2937 , \2938 , \2939 , \2940 , \2941 ,
         \2942 , \2943 , \2944 , \2945 , \2946 , \2947 , \2948 , \2949 , \2950 , \2951 ,
         \2952 , \2953 , \2954 , \2955 , \2956 , \2957 , \2958 , \2959 , \2960 , \2961 ,
         \2962 , \2963 , \2964 , \2965 , \2966 , \2967 , \2968 , \2969 , \2970 , \2971 ,
         \2972 , \2973 , \2974 , \2975 , \2976 , \2977 , \2978 , \2979 , \2980 , \2981 ,
         \2982 , \2983 , \2984 , \2985 , \2986 , \2987 , \2988 , \2989 , \2990 , \2991 ,
         \2992 , \2993 , \2994 , \2995 , \2996 , \2997 , \2998 , \2999 , \3000 , \3001 ,
         \3002 , \3003 , \3004 , \3005 , \3006 , \3007 , \3008 , \3009 , \3010 , \3011 ,
         \3012 , \3013 , \3014 , \3015 , \3016 , \3017 , \3018 , \3019 , \3020 , \3021 ,
         \3022 , \3023 , \3024 , \3025 , \3026 , \3027 , \3028 , \3029 , \3030 , \3031 ,
         \3032 , \3033 , \3034 , \3035 , \3036 , \3037 , \3038 , \3039 , \3040 , \3041 ,
         \3042 , \3043 , \3044 , \3045 , \3046 , \3047 , \3048 , \3049 , \3050 , \3051 ,
         \3052 , \3053 , \3054 , \3055 , \3056 , \3057 , \3058 , \3059 , \3060 , \3061 ,
         \3062 , \3063 , \3064 , \3065 , \3066 , \3067 , \3068 , \3069 , \3070 , \3071 ,
         \3072 , \3073 , \3074 , \3075 , \3076 , \3077 , \3078 , \3079 , \3080 , \3081 ,
         \3082 , \3083 , \3084 , \3085 , \3086 , \3087 , \3088 , \3089 , \3090 , \3091 ,
         \3092 , \3093 , \3094 , \3095 , \3096 , \3097 , \3098 , \3099 , \3100 , \3101 ,
         \3102 , \3103 , \3104 , \3105 , \3106 , \3107 , \3108 , \3109 , \3110 , \3111 ,
         \3112 , \3113 , \3114 , \3115 , \3116 , \3117 , \3118 , \3119 , \3120 , \3121 ,
         \3122 , \3123 , \3124 , \3125 , \3126 , \3127 , \3128 , \3129 , \3130 , \3131 ,
         \3132 , \3133 , \3134 , \3135 , \3136 , \3137 , \3138 , \3139 , \3140 , \3141 ,
         \3142 , \3143 , \3144 , \3145 , \3146 , \3147 , \3148 , \3149 , \3150 , \3151 ,
         \3152 , \3153 , \3154 , \3155 , \3156 , \3157 , \3158 , \3159 , \3160 , \3161 ,
         \3162 , \3163 , \3164 , \3165 , \3166 , \3167 , \3168 , \3169 , \3170 , \3171 ,
         \3172 , \3173 , \3174 , \3175 , \3176 , \3177 , \3178 , \3179 , \3180 , \3181 ,
         \3182 , \3183 , \3184 , \3185 , \3186 , \3187 , \3188 , \3189 , \3190 , \3191 ,
         \3192 , \3193 , \3194 , \3195 , \3196 , \3197 , \3198 , \3199 , \3200 , \3201 ,
         \3202 , \3203 , \3204 , \3205 , \3206 , \3207 , \3208 , \3209 , \3210 , \3211 ,
         \3212 , \3213 , \3214 , \3215 , \3216 , \3217 , \3218 , \3219 , \3220 , \3221 ,
         \3222 , \3223 , \3224 , \3225 , \3226 , \3227 , \3228 , \3229 , \3230 , \3231 ,
         \3232 , \3233 , \3234 , \3235 , \3236 , \3237 , \3238 , \3239 , \3240 , \3241 ,
         \3242 , \3243 , \3244 , \3245 , \3246 , \3247 , \3248 , \3249 , \3250 , \3251 ,
         \3252 , \3253 , \3254 , \3255 , \3256 , \3257 , \3258 , \3259 , \3260 , \3261 ,
         \3262 , \3263 , \3264 , \3265 , \3266 , \3267 , \3268 , \3269 , \3270 , \3271 ,
         \3272 , \3273 , \3274 , \3275 , \3276 , \3277 , \3278 , \3279 , \3280 , \3281 ,
         \3282 , \3283 , \3284 , \3285 , \3286 , \3287 , \3288 , \3289 , \3290 , \3291 ,
         \3292 , \3293 , \3294 , \3295 , \3296 , \3297 , \3298 , \3299 , \3300 , \3301 ,
         \3302 , \3303 , \3304 , \3305 , \3306 , \3307 , \3308 , \3309 , \3310 , \3311 ,
         \3312 , \3313 , \3314 , \3315 , \3316 , \3317 , \3318 , \3319 , \3320 , \3321 ,
         \3322 , \3323 , \3324 , \3325 , \3326 , \3327 , \3328 , \3329 , \3330 , \3331 ,
         \3332 , \3333 , \3334 , \3335 , \3336 , \3337 , \3338 , \3339 , \3340 , \3341 ,
         \3342 , \3343 , \3344 , \3345 , \3346 , \3347 , \3348 , \3349 , \3350 , \3351 ,
         \3352 , \3353 , \3354 , \3355 , \3356 , \3357 , \3358 , \3359 , \3360 , \3361 ,
         \3362 , \3363 , \3364 , \3365 , \3366 , \3367 , \3368 , \3369 , \3370 , \3371 ,
         \3372 , \3373 , \3374 , \3375 , \3376 , \3377 , \3378 , \3379 , \3380 , \3381 ,
         \3382 , \3383 , \3384 , \3385 , \3386 , \3387 , \3388 , \3389 , \3390 , \3391 ,
         \3392 , \3393 , \3394 , \3395 , \3396 , \3397 , \3398 , \3399 , \3400 , \3401 ,
         \3402 , \3403 , \3404 , \3405 , \3406 , \3407 , \3408 , \3409 , \3410 , \3411 ,
         \3412 , \3413 , \3414 , \3415 , \3416 , \3417 , \3418 , \3419 , \3420 , \3421 ,
         \3422 , \3423 , \3424 , \3425 , \3426 , \3427 , \3428 , \3429 , \3430 , \3431 ,
         \3432 , \3433 , \3434 , \3435 , \3436 , \3437 , \3438 , \3439 , \3440 , \3441 ,
         \3442 , \3443 , \3444 , \3445 , \3446 , \3447 , \3448 , \3449 , \3450 , \3451 ,
         \3452 , \3453 , \3454 , \3455 , \3456 , \3457 , \3458 , \3459 , \3460 , \3461 ,
         \3462 , \3463 , \3464 , \3465 , \3466 , \3467 , \3468 , \3469 , \3470 , \3471 ,
         \3472 , \3473 , \3474 , \3475 , \3476 , \3477 , \3478 , \3479 , \3480 , \3481 ,
         \3482 , \3483 , \3484 , \3485 , \3486 , \3487 , \3488 , \3489 , \3490 , \3491 ,
         \3492 , \3493 , \3494 , \3495 , \3496 , \3497 , \3498 , \3499 , \3500 , \3501 ,
         \3502 , \3503 , \3504 , \3505 , \3506 , \3507 , \3508 , \3509 , \3510 , \3511 ,
         \3512 , \3513 , \3514 , \3515 , \3516 , \3517 , \3518 , \3519 , \3520 , \3521 ,
         \3522 , \3523 , \3524 , \3525 , \3526 , \3527 , \3528 , \3529 , \3530 , \3531 ,
         \3532 , \3533 , \3534 , \3535 , \3536 , \3537 , \3538 , \3539 , \3540 , \3541 ,
         \3542 , \3543 , \3544 , \3545 , \3546 , \3547 , \3548 , \3549 , \3550 , \3551 ,
         \3552 , \3553 , \3554 , \3555 , \3556 , \3557 , \3558 , \3559 , \3560 , \3561 ,
         \3562 , \3563 , \3564 , \3565 , \3566 , \3567 , \3568 , \3569 , \3570 , \3571 ,
         \3572 , \3573 , \3574 , \3575 , \3576 , \3577 , \3578 , \3579 , \3580 , \3581 ,
         \3582 , \3583 , \3584 , \3585 , \3586 , \3587 , \3588 , \3589 , \3590 , \3591 ,
         \3592 , \3593 , \3594 , \3595 , \3596 , \3597 , \3598 , \3599 , \3600 , \3601 ,
         \3602 , \3603 , \3604 , \3605 , \3606 , \3607 , \3608 , \3609 , \3610 , \3611 ,
         \3612 , \3613 , \3614 , \3615 , \3616 , \3617 , \3618 , \3619 , \3620 , \3621 ,
         \3622 , \3623 , \3624 , \3625 , \3626 , \3627 , \3628 , \3629 , \3630 , \3631 ,
         \3632 , \3633 , \3634 , \3635 , \3636 , \3637 , \3638 , \3639 , \3640 , \3641 ,
         \3642 , \3643 , \3644 , \3645 , \3646 , \3647 , \3648 , \3649 , \3650 , \3651 ,
         \3652 , \3653 , \3654 , \3655 , \3656 , \3657 , \3658 , \3659 , \3660 , \3661 ,
         \3662 , \3663 , \3664 , \3665 , \3666 , \3667 , \3668 , \3669 , \3670 , \3671 ,
         \3672 , \3673 , \3674 , \3675 , \3676 , \3677 , \3678 , \3679 , \3680 , \3681 ,
         \3682 , \3683 , \3684 , \3685 , \3686 , \3687 , \3688 , \3689 , \3690 , \3691 ,
         \3692 , \3693 , \3694 , \3695 , \3696 , \3697 , \3698 , \3699 , \3700 , \3701 ,
         \3702 , \3703 , \3704 , \3705 , \3706 , \3707 , \3708 , \3709 , \3710 , \3711 ,
         \3712 , \3713 , \3714 , \3715 , \3716 , \3717 , \3718 , \3719 , \3720 , \3721 ,
         \3722 , \3723 , \3724 , \3725 , \3726 , \3727 , \3728 , \3729 , \3730 , \3731 ,
         \3732 , \3733 , \3734 , \3735 , \3736 , \3737 , \3738 , \3739 , \3740 , \3741 ,
         \3742 , \3743 , \3744 , \3745 , \3746 , \3747 , \3748 , \3749 , \3750 , \3751 ,
         \3752 , \3753 , \3754 , \3755 , \3756 , \3757 , \3758 , \3759 , \3760 , \3761 ,
         \3762 , \3763 , \3764 , \3765 , \3766 , \3767 , \3768 , \3769 , \3770 , \3771 ,
         \3772 , \3773 , \3774 , \3775 , \3776 , \3777 , \3778 , \3779 , \3780 , \3781 ,
         \3782 , \3783 , \3784 , \3785 , \3786 , \3787 , \3788 , \3789 , \3790 , \3791 ,
         \3792 , \3793 , \3794 , \3795 , \3796 , \3797 , \3798 , \3799 , \3800 , \3801 ,
         \3802 , \3803 , \3804 , \3805 , \3806 , \3807 , \3808 , \3809 , \3810 , \3811 ,
         \3812 , \3813 , \3814 , \3815 , \3816 , \3817 , \3818 , \3819 , \3820 , \3821 ,
         \3822 , \3823 , \3824 , \3825 , \3826 , \3827 , \3828 , \3829 , \3830 , \3831 ,
         \3832 , \3833 , \3834 , \3835 , \3836 , \3837 , \3838 , \3839 , \3840 , \3841 ,
         \3842 , \3843 , \3844 , \3845 , \3846 , \3847 , \3848 , \3849 , \3850 , \3851 ,
         \3852 , \3853 , \3854 , \3855 , \3856 , \3857 , \3858 , \3859 , \3860 , \3861 ,
         \3862 , \3863 , \3864 , \3865 , \3866 , \3867 , \3868 , \3869 , \3870 , \3871 ,
         \3872 , \3873 , \3874 , \3875 , \3876 , \3877 , \3878 , \3879 , \3880 , \3881 ,
         \3882 , \3883 , \3884 , \3885 , \3886 , \3887 , \3888 , \3889 , \3890 , \3891 ,
         \3892 , \3893 , \3894 , \3895 , \3896 , \3897 , \3898 , \3899 , \3900 , \3901 ,
         \3902 , \3903 , \3904 , \3905 , \3906 , \3907 , \3908 , \3909 , \3910 , \3911 ,
         \3912 , \3913 , \3914 , \3915 , \3916 , \3917 , \3918 , \3919 , \3920 , \3921 ,
         \3922 , \3923 , \3924 , \3925 , \3926 , \3927 , \3928 , \3929 , \3930 , \3931 ,
         \3932 , \3933 , \3934 , \3935 , \3936 , \3937 , \3938 , \3939 , \3940 , \3941 ,
         \3942 , \3943 , \3944 , \3945 , \3946 , \3947 , \3948 , \3949 , \3950 , \3951 ,
         \3952 , \3953 , \3954 , \3955 , \3956 , \3957 , \3958 , \3959 , \3960 , \3961 ,
         \3962 , \3963 , \3964 , \3965 , \3966 , \3967 , \3968 , \3969 , \3970 , \3971 ,
         \3972 , \3973 , \3974 , \3975 , \3976 , \3977 , \3978 , \3979 , \3980 , \3981 ,
         \3982 , \3983 , \3984 , \3985 , \3986 , \3987 , \3988 , \3989 , \3990 , \3991 ,
         \3992 , \3993 , \3994 , \3995 , \3996 , \3997 , \3998 , \3999 , \4000 , \4001 ,
         \4002 , \4003 , \4004 , \4005 , \4006 , \4007 , \4008 , \4009 , \4010 , \4011 ,
         \4012 , \4013 , \4014 , \4015 , \4016 , \4017 , \4018 , \4019 , \4020 , \4021 ,
         \4022 , \4023 , \4024 , \4025 , \4026 , \4027 , \4028 , \4029 , \4030 , \4031 ,
         \4032 , \4033 , \4034 , \4035 , \4036 , \4037 , \4038 , \4039 , \4040 , \4041 ,
         \4042 , \4043 , \4044 , \4045 , \4046 , \4047 , \4048 , \4049 , \4050 , \4051 ,
         \4052 , \4053 , \4054 , \4055 , \4056 , \4057 , \4058 , \4059 , \4060 , \4061 ,
         \4062 , \4063 , \4064 , \4065 , \4066 , \4067 , \4068 , \4069 , \4070 , \4071 ,
         \4072 , \4073 , \4074 , \4075 , \4076 , \4077 , \4078 , \4079 , \4080 , \4081 ,
         \4082 , \4083 , \4084 , \4085 , \4086 , \4087 , \4088 , \4089 , \4090 , \4091 ,
         \4092 , \4093 , \4094 , \4095 , \4096 , \4097 , \4098 , \4099 , \4100 , \4101 ,
         \4102 , \4103 , \4104 , \4105 , \4106 , \4107 , \4108 , \4109 , \4110 , \4111 ,
         \4112 , \4113 , \4114 , \4115 , \4116 , \4117 , \4118 , \4119 , \4120 , \4121 ,
         \4122 , \4123 , \4124 , \4125 , \4126 , \4127 , \4128 , \4129 , \4130 , \4131 ,
         \4132 , \4133 , \4134 , \4135 , \4136 , \4137 , \4138 , \4139 , \4140 , \4141 ,
         \4142 , \4143 , \4144 , \4145 , \4146 , \4147 , \4148 , \4149 , \4150 , \4151 ,
         \4152 , \4153 , \4154 , \4155 , \4156 , \4157 , \4158 , \4159 , \4160 , \4161 ,
         \4162 , \4163 , \4164 , \4165 , \4166 , \4167 , \4168 , \4169 , \4170 , \4171 ,
         \4172 , \4173 , \4174 , \4175 , \4176 , \4177 , \4178 , \4179 , \4180 , \4181 ,
         \4182 , \4183 , \4184 , \4185 , \4186 , \4187 , \4188 , \4189 , \4190 , \4191 ,
         \4192 , \4193 , \4194 , \4195 , \4196 , \4197 , \4198 , \4199 , \4200 , \4201 ,
         \4202 , \4203 , \4204 , \4205 , \4206 , \4207 , \4208 , \4209 , \4210 , \4211 ,
         \4212 , \4213 , \4214 , \4215 , \4216 , \4217 , \4218 , \4219 , \4220 , \4221 ,
         \4222 , \4223 , \4224 , \4225 , \4226 , \4227 , \4228 , \4229 , \4230 , \4231 ,
         \4232 , \4233 , \4234 , \4235 , \4236 , \4237 , \4238 , \4239 , \4240 , \4241 ,
         \4242 , \4243 , \4244 , \4245 , \4246 , \4247 , \4248 , \4249 , \4250 , \4251 ,
         \4252 , \4253 , \4254 , \4255 , \4256 , \4257 , \4258 , \4259 , \4260 , \4261 ,
         \4262 , \4263 , \4264 , \4265 , \4266 , \4267 , \4268 , \4269 , \4270 , \4271 ,
         \4272 , \4273 , \4274 , \4275 , \4276 , \4277 , \4278 , \4279 , \4280 , \4281 ,
         \4282 , \4283 , \4284 , \4285 , \4286 , \4287 , \4288 , \4289 , \4290 , \4291 ,
         \4292 , \4293 , \4294 , \4295 , \4296 , \4297 , \4298 , \4299 , \4300 , \4301 ,
         \4302 , \4303 , \4304 , \4305 , \4306 , \4307 , \4308 , \4309 , \4310 , \4311 ,
         \4312 , \4313 , \4314 , \4315 , \4316 , \4317 , \4318 , \4319 , \4320 , \4321 ,
         \4322 , \4323 , \4324 , \4325 , \4326 , \4327 , \4328 , \4329 , \4330 , \4331 ,
         \4332 , \4333 , \4334 , \4335 , \4336 , \4337 , \4338 , \4339 , \4340 , \4341 ,
         \4342 , \4343 , \4344 , \4345 , \4346 , \4347 , \4348 , \4349 , \4350 , \4351 ,
         \4352 , \4353 , \4354 , \4355 , \4356 , \4357 , \4358 , \4359 , \4360 , \4361 ,
         \4362 , \4363 , \4364 , \4365 , \4366 , \4367 , \4368 , \4369 , \4370 , \4371 ,
         \4372 , \4373 , \4374 , \4375 , \4376 , \4377 , \4378 , \4379 , \4380 , \4381 ,
         \4382 , \4383 , \4384 , \4385 , \4386 , \4387 , \4388 , \4389 , \4390 , \4391 ,
         \4392 , \4393 , \4394 , \4395 , \4396 , \4397 , \4398 , \4399 , \4400 , \4401 ,
         \4402 , \4403 , \4404 , \4405 , \4406 , \4407 , \4408 , \4409 , \4410 , \4411 ,
         \4412 , \4413 , \4414 , \4415 , \4416 , \4417 , \4418 , \4419 , \4420 , \4421 ,
         \4422 , \4423 , \4424 , \4425 , \4426 , \4427 , \4428 , \4429 , \4430 , \4431 ,
         \4432 , \4433 , \4434 , \4435 , \4436 , \4437 , \4438 , \4439 , \4440 , \4441 ,
         \4442 , \4443 , \4444 , \4445 , \4446 , \4447 , \4448 , \4449 , \4450 , \4451 ,
         \4452 , \4453 , \4454 , \4455 , \4456 , \4457 , \4458 , \4459 , \4460 , \4461 ,
         \4462 , \4463 , \4464 , \4465 , \4466 , \4467 , \4468 , \4469 , \4470 , \4471 ,
         \4472 , \4473 , \4474 , \4475 , \4476 , \4477 , \4478 , \4479 , \4480 , \4481 ,
         \4482 , \4483 , \4484 , \4485 , \4486 , \4487 , \4488 , \4489 , \4490 , \4491 ,
         \4492 , \4493 , \4494 , \4495 , \4496 , \4497 , \4498 , \4499 , \4500 , \4501 ,
         \4502 , \4503 , \4504 , \4505 , \4506 , \4507 , \4508 , \4509 , \4510 , \4511 ,
         \4512 , \4513 , \4514 , \4515 , \4516 , \4517 , \4518 , \4519 , \4520 , \4521 ,
         \4522 , \4523 , \4524 , \4525 , \4526 , \4527 , \4528 , \4529 , \4530 , \4531 ,
         \4532 , \4533 , \4534 , \4535 , \4536 , \4537 , \4538 , \4539 , \4540 , \4541 ,
         \4542 , \4543 , \4544 , \4545 , \4546 , \4547 , \4548 , \4549 , \4550 , \4551 ,
         \4552 , \4553 , \4554 , \4555 , \4556 , \4557 , \4558 , \4559 , \4560 , \4561 ,
         \4562 , \4563 , \4564 , \4565 , \4566 , \4567 , \4568 , \4569 , \4570 , \4571 ,
         \4572 , \4573 , \4574 , \4575 , \4576 , \4577 , \4578 , \4579 , \4580 , \4581 ,
         \4582 , \4583 , \4584 , \4585 , \4586 , \4587 , \4588 , \4589 , \4590 , \4591 ,
         \4592 , \4593 , \4594 , \4595 , \4596 , \4597 , \4598 , \4599 , \4600 , \4601 ,
         \4602 , \4603 , \4604 , \4605 , \4606 , \4607 , \4608 , \4609 , \4610 , \4611 ,
         \4612 , \4613 , \4614 , \4615 , \4616 , \4617 , \4618 , \4619 , \4620 , \4621 ,
         \4622 , \4623 , \4624 , \4625 , \4626 , \4627 , \4628 , \4629 , \4630 , \4631 ,
         \4632 , \4633 , \4634 , \4635 , \4636 , \4637 , \4638 , \4639 , \4640 , \4641 ,
         \4642 , \4643 , \4644 , \4645 , \4646 , \4647 , \4648 , \4649 , \4650 , \4651 ,
         \4652 , \4653 , \4654 , \4655 , \4656 , \4657 , \4658 , \4659 , \4660 , \4661 ,
         \4662 , \4663 , \4664 , \4665 , \4666 , \4667 , \4668 , \4669 , \4670 , \4671 ,
         \4672 , \4673 , \4674 , \4675 , \4676 , \4677 , \4678 , \4679 , \4680 , \4681 ,
         \4682 , \4683 , \4684 , \4685 , \4686 , \4687 , \4688 , \4689 , \4690 , \4691 ,
         \4692 , \4693 , \4694 , \4695 , \4696 , \4697 , \4698 , \4699 , \4700 , \4701 ,
         \4702 , \4703 , \4704 , \4705 , \4706 , \4707 , \4708 , \4709 , \4710 , \4711 ,
         \4712 , \4713 , \4714 , \4715 , \4716 , \4717 , \4718 , \4719 , \4720 , \4721 ,
         \4722 , \4723 , \4724 , \4725 , \4726 , \4727 , \4728 , \4729 , \4730 , \4731 ,
         \4732 , \4733 , \4734 , \4735 , \4736 , \4737 , \4738 , \4739 , \4740 , \4741 ,
         \4742 , \4743 , \4744 , \4745 , \4746 , \4747 , \4748 , \4749 , \4750 , \4751 ,
         \4752 , \4753 , \4754 , \4755 , \4756 , \4757 , \4758 , \4759 , \4760 , \4761 ,
         \4762 , \4763 , \4764 , \4765 , \4766 , \4767 , \4768 , \4769 , \4770 , \4771 ,
         \4772 , \4773 , \4774 , \4775 , \4776 , \4777 , \4778 , \4779 , \4780 , \4781 ,
         \4782 , \4783 , \4784 , \4785 , \4786 , \4787 , \4788 , \4789 , \4790 , \4791 ,
         \4792 , \4793 , \4794 , \4795 , \4796 , \4797 , \4798 , \4799 , \4800 , \4801 ,
         \4802 , \4803 , \4804 , \4805 , \4806 , \4807 , \4808 , \4809 , \4810 , \4811 ,
         \4812 , \4813 , \4814 , \4815 , \4816 , \4817 , \4818 , \4819 , \4820 , \4821 ,
         \4822 , \4823 , \4824 , \4825 , \4826 , \4827 , \4828 , \4829 , \4830 , \4831 ,
         \4832 , \4833 , \4834 , \4835 , \4836 , \4837 , \4838 , \4839 , \4840 , \4841 ,
         \4842 , \4843 , \4844 , \4845 , \4846 , \4847 , \4848 , \4849 , \4850 , \4851 ,
         \4852 , \4853 , \4854 , \4855 , \4856 , \4857 , \4858 , \4859 , \4860 , \4861 ,
         \4862 , \4863 , \4864 , \4865 , \4866 , \4867 , \4868 , \4869 , \4870 , \4871 ,
         \4872 , \4873 , \4874 , \4875 , \4876 , \4877 , \4878 , \4879 , \4880 , \4881 ,
         \4882 , \4883 , \4884 , \4885 , \4886 , \4887 , \4888 , \4889 , \4890 , \4891 ,
         \4892 , \4893 , \4894 , \4895 , \4896 , \4897 , \4898 , \4899 , \4900 , \4901 ,
         \4902 , \4903 , \4904 , \4905 , \4906 , \4907 , \4908 , \4909 , \4910 , \4911 ,
         \4912 , \4913 , \4914 , \4915 , \4916 , \4917 , \4918 , \4919 , \4920 , \4921 ,
         \4922 , \4923 , \4924 , \4925 , \4926 , \4927 , \4928 , \4929 , \4930 , \4931 ,
         \4932 , \4933 , \4934 , \4935 , \4936 , \4937 , \4938 , \4939 , \4940 , \4941 ,
         \4942 , \4943 , \4944 , \4945 , \4946 , \4947 , \4948 , \4949 , \4950 , \4951 ,
         \4952 , \4953 , \4954 , \4955 , \4956 , \4957 , \4958 , \4959 , \4960 , \4961 ,
         \4962 , \4963 , \4964 , \4965 , \4966 , \4967 , \4968 , \4969 , \4970 , \4971 ,
         \4972 , \4973 , \4974 , \4975 , \4976 , \4977 , \4978 , \4979 , \4980 , \4981 ,
         \4982 , \4983 , \4984 , \4985 , \4986 , \4987 , \4988 , \4989 , \4990 , \4991 ,
         \4992 , \4993 , \4994 , \4995 , \4996 , \4997 , \4998 , \4999 , \5000 , \5001 ,
         \5002 , \5003 , \5004 , \5005 , \5006 , \5007 , \5008 , \5009 , \5010 , \5011 ,
         \5012 , \5013 , \5014 , \5015 , \5016 , \5017 , \5018 , \5019 , \5020 , \5021 ,
         \5022 , \5023 , \5024 , \5025 , \5026 , \5027 , \5028 , \5029 , \5030 , \5031 ,
         \5032 , \5033 , \5034 , \5035 , \5036 , \5037 , \5038 , \5039 , \5040 , \5041 ,
         \5042 , \5043 , \5044 , \5045 , \5046 , \5047 , \5048 , \5049 , \5050 , \5051 ,
         \5052 , \5053 , \5054 , \5055 , \5056 , \5057 , \5058 , \5059 , \5060 , \5061 ,
         \5062 , \5063 , \5064 , \5065 , \5066 , \5067 , \5068 , \5069 , \5070 , \5071 ,
         \5072 , \5073 , \5074 , \5075 , \5076 , \5077 , \5078 , \5079 , \5080 , \5081 ,
         \5082 , \5083 , \5084 , \5085 , \5086 , \5087 , \5088 , \5089 , \5090 , \5091 ,
         \5092 , \5093 , \5094 , \5095 , \5096 , \5097 , \5098 , \5099 , \5100 , \5101 ,
         \5102 , \5103 , \5104 , \5105 , \5106 , \5107 , \5108 , \5109 , \5110 , \5111 ,
         \5112 , \5113 , \5114 , \5115 , \5116 , \5117 , \5118 , \5119 , \5120 , \5121 ,
         \5122 , \5123 , \5124 , \5125 , \5126 , \5127 , \5128 , \5129 , \5130 , \5131 ,
         \5132 , \5133 , \5134 , \5135 , \5136 , \5137 , \5138 , \5139 , \5140 , \5141 ,
         \5142 , \5143 , \5144 , \5145 , \5146 , \5147 , \5148 , \5149 , \5150 , \5151 ,
         \5152 , \5153 , \5154 , \5155 , \5156 , \5157 , \5158 , \5159 , \5160 , \5161 ,
         \5162 , \5163 , \5164 , \5165 , \5166 , \5167 , \5168 , \5169 , \5170 , \5171 ,
         \5172 , \5173 , \5174 , \5175 , \5176 , \5177 , \5178 , \5179 , \5180 , \5181 ,
         \5182 , \5183 , \5184 , \5185 , \5186 , \5187 , \5188 , \5189 , \5190 , \5191 ,
         \5192 , \5193 , \5194 , \5195 , \5196 , \5197 , \5198 , \5199 , \5200 , \5201 ,
         \5202 , \5203 , \5204 , \5205 , \5206 , \5207 , \5208 , \5209 , \5210 , \5211 ,
         \5212 , \5213 , \5214 , \5215 , \5216 , \5217 , \5218 , \5219 , \5220 , \5221 ,
         \5222 , \5223 , \5224 , \5225 , \5226 , \5227 , \5228 , \5229 , \5230 , \5231 ,
         \5232 , \5233 , \5234 , \5235 , \5236 , \5237 , \5238 , \5239 , \5240 , \5241 ,
         \5242 , \5243 , \5244 , \5245 , \5246 , \5247 , \5248 , \5249 , \5250 , \5251 ,
         \5252 , \5253 , \5254 , \5255 , \5256 , \5257 , \5258 , \5259 , \5260 , \5261 ,
         \5262 , \5263 , \5264 , \5265 , \5266 , \5267 , \5268 , \5269 , \5270 , \5271 ,
         \5272 , \5273 , \5274 , \5275 , \5276 , \5277 , \5278 , \5279 , \5280 , \5281 ,
         \5282 , \5283 , \5284 , \5285 , \5286 , \5287 , \5288 , \5289 , \5290 , \5291 ,
         \5292 , \5293 , \5294 , \5295 , \5296 , \5297 , \5298 , \5299 , \5300 , \5301 ,
         \5302 , \5303 , \5304 , \5305 , \5306 , \5307 , \5308 , \5309 , \5310 , \5311 ,
         \5312 , \5313 , \5314 , \5315 , \5316 , \5317 , \5318 , \5319 , \5320 , \5321 ,
         \5322 , \5323 , \5324 , \5325 , \5326 , \5327 , \5328 , \5329 , \5330 , \5331 ,
         \5332 , \5333 , \5334 , \5335 , \5336 , \5337 , \5338 , \5339 , \5340 , \5341 ,
         \5342 , \5343 , \5344 , \5345 , \5346 , \5347 , \5348 , \5349 , \5350 , \5351 ,
         \5352 , \5353 , \5354 , \5355 , \5356 , \5357 , \5358 , \5359 , \5360 , \5361 ,
         \5362 , \5363 , \5364 , \5365 , \5366 , \5367 , \5368 , \5369 , \5370 , \5371 ,
         \5372 , \5373 , \5374 , \5375 , \5376 , \5377 , \5378 , \5379 , \5380 , \5381 ,
         \5382 , \5383 , \5384 , \5385 , \5386 , \5387 , \5388 , \5389 , \5390 , \5391 ,
         \5392 , \5393 , \5394 , \5395 , \5396 , \5397 , \5398 , \5399 , \5400 , \5401 ,
         \5402 , \5403 , \5404 , \5405 , \5406 , \5407 , \5408 , \5409 , \5410 , \5411 ,
         \5412 , \5413 , \5414 , \5415 , \5416 , \5417 , \5418 , \5419 , \5420 , \5421 ,
         \5422 , \5423 , \5424 , \5425 , \5426 , \5427 , \5428 , \5429 , \5430 , \5431 ,
         \5432 , \5433 , \5434 , \5435 , \5436 , \5437 , \5438 , \5439 , \5440 , \5441 ,
         \5442 , \5443 , \5444 , \5445 , \5446 , \5447 , \5448 , \5449 , \5450 , \5451 ,
         \5452 , \5453 , \5454 , \5455 , \5456 , \5457 , \5458 , \5459 , \5460 , \5461 ,
         \5462 , \5463 , \5464 , \5465 , \5466 , \5467 , \5468 , \5469 , \5470 , \5471 ,
         \5472 , \5473 , \5474 , \5475 , \5476 , \5477 , \5478 , \5479 , \5480 , \5481 ,
         \5482 , \5483 , \5484 , \5485 , \5486 , \5487 , \5488 , \5489 , \5490 , \5491 ,
         \5492 , \5493 , \5494 , \5495 , \5496 , \5497 , \5498 , \5499 , \5500 , \5501 ,
         \5502 , \5503 , \5504 , \5505 , \5506 , \5507 , \5508 , \5509 , \5510 , \5511 ,
         \5512 , \5513 , \5514 , \5515 , \5516 , \5517 , \5518 , \5519 , \5520 , \5521 ,
         \5522 , \5523 , \5524 , \5525 , \5526 , \5527 , \5528 , \5529 , \5530 , \5531 ,
         \5532 , \5533 , \5534 , \5535 , \5536 , \5537 , \5538 , \5539 , \5540 , \5541 ,
         \5542 , \5543 , \5544 , \5545 , \5546 , \5547 , \5548 , \5549 , \5550 , \5551 ,
         \5552 , \5553 , \5554 , \5555 , \5556 , \5557 , \5558 , \5559 , \5560 , \5561 ,
         \5562 , \5563 , \5564 , \5565 , \5566 , \5567 , \5568 , \5569 , \5570 , \5571 ,
         \5572 , \5573 , \5574 , \5575 , \5576 , \5577 , \5578 , \5579 , \5580 , \5581 ,
         \5582 , \5583 , \5584 , \5585 , \5586 , \5587 , \5588 , \5589 , \5590 , \5591 ,
         \5592 , \5593 , \5594 , \5595 , \5596 , \5597 , \5598 , \5599 , \5600 , \5601 ,
         \5602 , \5603 , \5604 , \5605 , \5606 , \5607 , \5608 , \5609 , \5610 , \5611 ,
         \5612 , \5613 , \5614 , \5615 , \5616 , \5617 , \5618 , \5619 , \5620 , \5621 ,
         \5622 , \5623 , \5624 , \5625 , \5626 , \5627 , \5628 , \5629 , \5630 , \5631 ,
         \5632 , \5633 , \5634 , \5635 , \5636 , \5637 , \5638 , \5639 , \5640 , \5641 ,
         \5642 , \5643 , \5644 , \5645 , \5646 , \5647 , \5648 , \5649 , \5650 , \5651 ,
         \5652 , \5653 , \5654 , \5655 , \5656 , \5657 , \5658 , \5659 , \5660 , \5661 ,
         \5662 , \5663 , \5664 , \5665 , \5666 , \5667 , \5668 , \5669 , \5670 , \5671 ,
         \5672 , \5673 , \5674 , \5675 , \5676 , \5677 , \5678 , \5679 , \5680 , \5681 ,
         \5682 , \5683 , \5684 , \5685 , \5686 , \5687 , \5688 , \5689 , \5690 , \5691 ,
         \5692 , \5693 , \5694 , \5695 , \5696 , \5697 , \5698 , \5699 , \5700 , \5701 ,
         \5702 , \5703 , \5704 , \5705 , \5706 , \5707 , \5708 , \5709 , \5710 , \5711 ,
         \5712 , \5713 , \5714 , \5715 , \5716 , \5717 , \5718 , \5719 , \5720 , \5721 ,
         \5722 , \5723 , \5724 , \5725 , \5726 , \5727 , \5728 , \5729 , \5730 , \5731 ,
         \5732 , \5733 , \5734 , \5735 , \5736 , \5737 , \5738 , \5739 , \5740 , \5741 ,
         \5742 , \5743 , \5744 , \5745 , \5746 , \5747 , \5748 , \5749 , \5750 , \5751 ,
         \5752 , \5753 , \5754 , \5755 , \5756 , \5757 , \5758 , \5759 , \5760 , \5761 ,
         \5762 , \5763 , \5764 , \5765 , \5766 , \5767 , \5768 , \5769 , \5770 , \5771 ,
         \5772 , \5773 , \5774 , \5775 , \5776 , \5777 , \5778 , \5779 , \5780 , \5781 ,
         \5782 , \5783 , \5784 , \5785 , \5786 , \5787 , \5788 , \5789 , \5790 , \5791 ,
         \5792 , \5793 , \5794 , \5795 , \5796 , \5797 , \5798 , \5799 , \5800 , \5801 ,
         \5802 , \5803 , \5804 , \5805 , \5806 , \5807 , \5808 , \5809 , \5810 , \5811 ,
         \5812 , \5813 , \5814 , \5815 , \5816 , \5817 , \5818 , \5819 , \5820 , \5821 ,
         \5822 , \5823 , \5824 , \5825 , \5826 , \5827 , \5828 , \5829 , \5830 , \5831 ,
         \5832 , \5833 , \5834 , \5835 , \5836 , \5837 , \5838 , \5839 , \5840 , \5841 ,
         \5842 , \5843 , \5844 , \5845 , \5846 , \5847 , \5848 , \5849 , \5850 , \5851 ,
         \5852 , \5853 , \5854 , \5855 , \5856 , \5857 , \5858 , \5859 , \5860 , \5861 ,
         \5862 , \5863 , \5864 , \5865 , \5866 , \5867 , \5868 , \5869 , \5870 , \5871 ,
         \5872 , \5873 , \5874 , \5875 , \5876 , \5877 , \5878 , \5879 , \5880 , \5881 ,
         \5882 , \5883 , \5884 , \5885 , \5886 , \5887 , \5888 , \5889 , \5890 , \5891 ,
         \5892 , \5893 , \5894 , \5895 , \5896 , \5897 , \5898 , \5899 , \5900 , \5901 ,
         \5902 , \5903 , \5904 , \5905 , \5906 , \5907 , \5908 , \5909 , \5910 , \5911 ,
         \5912 , \5913 , \5914 , \5915 , \5916 , \5917 , \5918 , \5919 , \5920 , \5921 ,
         \5922 , \5923 , \5924 , \5925 , \5926 , \5927 , \5928 , \5929 , \5930 , \5931 ,
         \5932 , \5933 , \5934 , \5935 , \5936 , \5937 , \5938 , \5939 , \5940 , \5941 ,
         \5942 , \5943 , \5944 , \5945 , \5946 , \5947 , \5948 , \5949 , \5950 , \5951 ,
         \5952 , \5953 , \5954 , \5955 , \5956 , \5957 , \5958 , \5959 , \5960 , \5961 ,
         \5962 , \5963 , \5964 , \5965 , \5966 , \5967 , \5968 , \5969 , \5970 , \5971 ,
         \5972 , \5973 , \5974 , \5975 , \5976 , \5977 , \5978 , \5979 , \5980 , \5981 ,
         \5982 , \5983 , \5984 , \5985 , \5986 , \5987 , \5988 , \5989 , \5990 , \5991 ,
         \5992 , \5993 , \5994 , \5995 , \5996 , \5997 , \5998 , \5999 , \6000 , \6001 ,
         \6002 , \6003 , \6004 , \6005 , \6006 , \6007 , \6008 , \6009 , \6010 , \6011 ,
         \6012 , \6013 , \6014 , \6015 , \6016 , \6017 , \6018 , \6019 , \6020 , \6021 ,
         \6022 , \6023 , \6024 , \6025 , \6026 , \6027 , \6028 , \6029 , \6030 , \6031 ,
         \6032 , \6033 , \6034 , \6035 , \6036 , \6037 , \6038 , \6039 , \6040 , \6041 ,
         \6042 , \6043 , \6044 , \6045 , \6046 , \6047 , \6048 , \6049 , \6050 , \6051 ,
         \6052 , \6053 , \6054 , \6055 , \6056 , \6057 , \6058 , \6059 , \6060 , \6061 ,
         \6062 , \6063 , \6064 , \6065 , \6066 , \6067 , \6068 , \6069 , \6070 , \6071 ,
         \6072 , \6073 , \6074 , \6075 , \6076 , \6077 , \6078 , \6079 , \6080 , \6081 ,
         \6082 , \6083 , \6084 , \6085 , \6086 , \6087 , \6088 , \6089 , \6090 , \6091 ,
         \6092 , \6093 , \6094 , \6095 , \6096 , \6097 , \6098 , \6099 , \6100 , \6101 ,
         \6102 , \6103 , \6104 , \6105 , \6106 , \6107 , \6108 , \6109 , \6110 , \6111 ,
         \6112 , \6113 , \6114 , \6115 , \6116 , \6117 , \6118 , \6119 , \6120 , \6121 ,
         \6122 , \6123 , \6124 , \6125 , \6126 , \6127 , \6128 , \6129 , \6130 , \6131 ,
         \6132 , \6133 , \6134 , \6135 , \6136 , \6137 , \6138 , \6139 , \6140 , \6141 ,
         \6142 , \6143 , \6144 , \6145 , \6146 , \6147 , \6148 , \6149 , \6150 , \6151 ,
         \6152 , \6153 , \6154 , \6155 , \6156 , \6157 , \6158 , \6159 , \6160 , \6161 ,
         \6162 , \6163 , \6164 , \6165 , \6166 , \6167 , \6168 , \6169 , \6170 , \6171 ,
         \6172 , \6173 , \6174 , \6175 , \6176 , \6177 , \6178 , \6179 , \6180 , \6181 ,
         \6182 , \6183 , \6184 , \6185 , \6186 , \6187 , \6188 , \6189 , \6190 , \6191 ,
         \6192 , \6193 , \6194 , \6195 , \6196 , \6197 , \6198 , \6199 , \6200 , \6201 ,
         \6202 , \6203 , \6204 , \6205 , \6206 , \6207 , \6208 , \6209 , \6210 , \6211 ,
         \6212 , \6213 , \6214 , \6215 , \6216 , \6217 , \6218 , \6219 , \6220 , \6221 ,
         \6222 , \6223 , \6224 , \6225 , \6226 , \6227 , \6228 , \6229 , \6230 , \6231 ,
         \6232 , \6233 , \6234 , \6235 , \6236 , \6237 , \6238 , \6239 , \6240 , \6241 ,
         \6242 , \6243 , \6244 , \6245 , \6246 , \6247 , \6248 , \6249 , \6250 , \6251 ,
         \6252 , \6253 , \6254 , \6255 , \6256 , \6257 , \6258 , \6259 , \6260 , \6261 ,
         \6262 , \6263 , \6264 , \6265 , \6266 , \6267 , \6268 , \6269 , \6270 , \6271 ,
         \6272 , \6273 , \6274 , \6275 , \6276 , \6277 , \6278 , \6279 , \6280 , \6281 ,
         \6282 , \6283 , \6284 , \6285 , \6286 , \6287 , \6288 , \6289 , \6290 , \6291 ,
         \6292 , \6293 , \6294 , \6295 , \6296 , \6297 , \6298 , \6299 , \6300 , \6301 ,
         \6302 , \6303 , \6304 , \6305 , \6306 , \6307 , \6308 , \6309 , \6310 , \6311 ,
         \6312 , \6313 , \6314 , \6315 , \6316 , \6317 , \6318 , \6319 , \6320 , \6321 ,
         \6322 , \6323 , \6324 , \6325 , \6326 , \6327 , \6328 , \6329 , \6330 , \6331 ,
         \6332 , \6333 , \6334 , \6335 , \6336 , \6337 , \6338 , \6339 , \6340 , \6341 ,
         \6342 , \6343 , \6344 , \6345 , \6346 , \6347 , \6348 , \6349 , \6350 , \6351 ,
         \6352 , \6353 , \6354 , \6355 , \6356 , \6357 , \6358 , \6359 , \6360 , \6361 ,
         \6362 , \6363 , \6364 , \6365 , \6366 , \6367 , \6368 , \6369 , \6370 , \6371 ,
         \6372 , \6373 , \6374 , \6375 , \6376 , \6377 , \6378 , \6379 , \6380 , \6381 ,
         \6382 , \6383 , \6384 , \6385 , \6386 , \6387 , \6388 , \6389 , \6390 , \6391 ,
         \6392 , \6393 , \6394 , \6395 , \6396 , \6397 , \6398 , \6399 , \6400 , \6401 ,
         \6402 , \6403 , \6404 , \6405 , \6406 , \6407 , \6408 , \6409 , \6410 , \6411 ,
         \6412 , \6413 , \6414 , \6415 , \6416 , \6417 , \6418 , \6419 , \6420 , \6421 ,
         \6422 , \6423 , \6424 , \6425 , \6426 , \6427 , \6428 , \6429 , \6430 , \6431 ,
         \6432 , \6433 , \6434 , \6435 , \6436 , \6437 , \6438 , \6439 , \6440 , \6441 ,
         \6442 , \6443 , \6444 , \6445 , \6446 , \6447 , \6448 , \6449 , \6450 , \6451 ,
         \6452 , \6453 , \6454 , \6455 , \6456 , \6457 , \6458 , \6459 , \6460 , \6461 ,
         \6462 , \6463 , \6464 , \6465 , \6466 , \6467 , \6468 , \6469 , \6470 , \6471 ,
         \6472 , \6473 , \6474 , \6475 , \6476 , \6477 , \6478 , \6479 , \6480 , \6481 ,
         \6482 , \6483 , \6484 , \6485 , \6486 , \6487 , \6488 , \6489 , \6490 , \6491 ,
         \6492 , \6493 , \6494 , \6495 , \6496 , \6497 , \6498 , \6499 , \6500 , \6501 ,
         \6502 , \6503 , \6504 , \6505 , \6506 , \6507 , \6508 , \6509 , \6510 , \6511 ,
         \6512 , \6513 , \6514 , \6515 , \6516 , \6517 , \6518 , \6519 , \6520 , \6521 ,
         \6522 , \6523 , \6524 , \6525 , \6526 , \6527 , \6528 , \6529 , \6530 , \6531 ,
         \6532 , \6533 , \6534 , \6535 , \6536 , \6537 , \6538 , \6539 , \6540 , \6541 ,
         \6542 , \6543 , \6544 , \6545 , \6546 , \6547 , \6548 , \6549 , \6550 , \6551 ,
         \6552 , \6553 , \6554 , \6555 , \6556 , \6557 , \6558 , \6559 , \6560 , \6561 ,
         \6562 , \6563 , \6564 , \6565 , \6566 , \6567 , \6568 , \6569 , \6570 , \6571 ,
         \6572 , \6573 , \6574 , \6575 , \6576 , \6577 , \6578 , \6579 , \6580 , \6581 ,
         \6582 , \6583 , \6584 , \6585 , \6586 , \6587 , \6588 , \6589 , \6590 , \6591 ,
         \6592 , \6593 , \6594 , \6595 , \6596 , \6597 , \6598 , \6599 , \6600 , \6601 ,
         \6602 , \6603 , \6604 , \6605 , \6606 , \6607 , \6608 , \6609 , \6610 , \6611 ,
         \6612 , \6613 , \6614 , \6615 , \6616 , \6617 , \6618 , \6619 , \6620 , \6621 ,
         \6622 , \6623 , \6624 , \6625 , \6626 , \6627 , \6628 , \6629 , \6630 , \6631 ,
         \6632 , \6633 , \6634 , \6635 , \6636 , \6637 , \6638 , \6639 , \6640 , \6641 ,
         \6642 , \6643 , \6644 , \6645 , \6646 , \6647 , \6648 , \6649 , \6650 , \6651 ,
         \6652 , \6653 , \6654 , \6655 , \6656 , \6657 , \6658 , \6659 , \6660 , \6661 ,
         \6662 , \6663 , \6664 , \6665 , \6666 , \6667 , \6668 , \6669 , \6670 , \6671 ,
         \6672 , \6673 , \6674 , \6675 , \6676 , \6677 , \6678 , \6679 , \6680 , \6681 ,
         \6682 , \6683 , \6684 , \6685 , \6686 , \6687 , \6688 , \6689 , \6690 , \6691 ,
         \6692 , \6693 , \6694 , \6695 , \6696 , \6697 , \6698 , \6699 , \6700 , \6701 ,
         \6702 , \6703 , \6704 , \6705 , \6706 , \6707 , \6708 , \6709 , \6710 , \6711 ,
         \6712 , \6713 , \6714 , \6715 , \6716 , \6717 , \6718 , \6719 , \6720 , \6721 ,
         \6722 , \6723 , \6724 , \6725 , \6726 , \6727 , \6728 , \6729 , \6730 , \6731 ,
         \6732 , \6733 , \6734 , \6735 , \6736 , \6737 , \6738 , \6739 , \6740 , \6741 ,
         \6742 , \6743 , \6744 , \6745 , \6746 , \6747 , \6748 , \6749 , \6750 , \6751 ,
         \6752 , \6753 , \6754 , \6755 , \6756 , \6757 , \6758 , \6759 , \6760 , \6761 ,
         \6762 , \6763 , \6764 , \6765 , \6766 , \6767 , \6768 , \6769 , \6770 , \6771 ,
         \6772 , \6773 , \6774 , \6775 , \6776 , \6777 , \6778 , \6779 , \6780 , \6781 ,
         \6782 , \6783 , \6784 , \6785 , \6786 , \6787 , \6788 , \6789 , \6790 , \6791 ,
         \6792 , \6793 , \6794 , \6795 , \6796 , \6797 , \6798 , \6799 , \6800 , \6801 ,
         \6802 , \6803 , \6804 , \6805 , \6806 , \6807 , \6808 , \6809 , \6810 , \6811 ,
         \6812 , \6813 , \6814 , \6815 , \6816 , \6817 , \6818 , \6819 , \6820 , \6821 ,
         \6822 , \6823 , \6824 , \6825 , \6826 , \6827 , \6828 , \6829 , \6830 , \6831 ,
         \6832 , \6833 , \6834 , \6835 , \6836 , \6837 , \6838 , \6839 , \6840 , \6841 ,
         \6842 , \6843 , \6844 , \6845 , \6846 , \6847 , \6848 , \6849 , \6850 , \6851 ,
         \6852 , \6853 , \6854 , \6855 , \6856 , \6857 , \6858 , \6859 , \6860 , \6861 ,
         \6862 , \6863 , \6864 , \6865 , \6866 , \6867 , \6868 , \6869 , \6870 , \6871 ,
         \6872 , \6873 , \6874 , \6875 , \6876 , \6877 , \6878 , \6879 , \6880 , \6881 ,
         \6882 , \6883 , \6884 , \6885 , \6886 , \6887 , \6888 , \6889 , \6890 , \6891 ,
         \6892 , \6893 , \6894 , \6895 , \6896 , \6897 , \6898 , \6899 , \6900 , \6901 ,
         \6902 , \6903 , \6904 , \6905 , \6906 , \6907 , \6908 , \6909 , \6910 , \6911 ,
         \6912 , \6913 , \6914 , \6915 , \6916 , \6917 , \6918 , \6919 , \6920 , \6921 ,
         \6922 , \6923 , \6924 , \6925 , \6926 , \6927 , \6928 , \6929 , \6930 , \6931 ,
         \6932 , \6933 , \6934 , \6935 , \6936 , \6937 , \6938 , \6939 , \6940 , \6941 ,
         \6942 , \6943 , \6944 , \6945 , \6946 , \6947 , \6948 , \6949 , \6950 , \6951 ,
         \6952 , \6953 , \6954 , \6955 , \6956 , \6957 , \6958 , \6959 , \6960 , \6961 ,
         \6962 , \6963 , \6964 , \6965 , \6966 , \6967 , \6968 , \6969 , \6970 , \6971 ,
         \6972 , \6973 , \6974 , \6975 , \6976 , \6977 , \6978 , \6979 , \6980 , \6981 ,
         \6982 , \6983 , \6984 , \6985 , \6986 , \6987 , \6988 , \6989 , \6990 , \6991 ,
         \6992 , \6993 , \6994 , \6995 , \6996 , \6997 , \6998 , \6999 , \7000 , \7001 ,
         \7002 , \7003 , \7004 , \7005 , \7006 , \7007 , \7008 , \7009 , \7010 , \7011 ,
         \7012 , \7013 , \7014 , \7015 , \7016 , \7017 , \7018 , \7019 , \7020 , \7021 ,
         \7022 , \7023 , \7024 , \7025 , \7026 , \7027 , \7028 , \7029 , \7030 , \7031 ,
         \7032 , \7033 , \7034 , \7035 , \7036 , \7037 , \7038 , \7039 , \7040 , \7041 ,
         \7042 , \7043 , \7044 , \7045 , \7046 , \7047 , \7048 , \7049 , \7050 , \7051 ,
         \7052 , \7053 , \7054 , \7055 , \7056 , \7057 , \7058 , \7059 , \7060 , \7061 ,
         \7062 , \7063 , \7064 , \7065 , \7066 , \7067 , \7068 , \7069 , \7070 , \7071 ,
         \7072 , \7073 , \7074 , \7075 , \7076 , \7077 , \7078 , \7079 , \7080 , \7081 ,
         \7082 , \7083 , \7084 , \7085 , \7086 , \7087 , \7088 , \7089 , \7090 , \7091 ,
         \7092 , \7093 , \7094 , \7095 , \7096 , \7097 , \7098 , \7099 , \7100 , \7101 ,
         \7102 , \7103 , \7104 , \7105 , \7106 , \7107 , \7108 , \7109 , \7110 , \7111 ,
         \7112 , \7113 , \7114 , \7115 , \7116 , \7117 , \7118 , \7119 , \7120 , \7121 ,
         \7122 , \7123 , \7124 , \7125 , \7126 , \7127 , \7128 , \7129 , \7130 , \7131 ,
         \7132 , \7133 , \7134 , \7135 , \7136 , \7137 , \7138 , \7139 , \7140 , \7141 ,
         \7142 , \7143 , \7144 , \7145 , \7146 , \7147 , \7148 , \7149 , \7150 , \7151 ,
         \7152 , \7153 , \7154 , \7155 , \7156 , \7157 , \7158 , \7159 , \7160 , \7161 ,
         \7162 , \7163 , \7164 , \7165 , \7166 , \7167 , \7168 , \7169 , \7170 , \7171 ,
         \7172 , \7173 , \7174 , \7175 , \7176 , \7177 , \7178 , \7179 , \7180 , \7181 ,
         \7182 , \7183 , \7184 , \7185 , \7186 , \7187 , \7188 , \7189 , \7190 , \7191 ,
         \7192 , \7193 , \7194 , \7195 , \7196 , \7197 , \7198 , \7199 , \7200 , \7201 ,
         \7202 , \7203 , \7204 , \7205 , \7206 , \7207 , \7208 , \7209 , \7210 , \7211 ,
         \7212 , \7213 , \7214 , \7215 , \7216 , \7217 , \7218 , \7219 , \7220 , \7221 ,
         \7222 , \7223 , \7224 , \7225 , \7226 , \7227 , \7228 , \7229 , \7230 , \7231 ,
         \7232 , \7233 , \7234 , \7235 , \7236 , \7237 , \7238 , \7239 , \7240 , \7241 ,
         \7242 , \7243 , \7244 , \7245 , \7246 , \7247 , \7248 , \7249 , \7250 , \7251 ,
         \7252 , \7253 , \7254 , \7255 , \7256 , \7257 , \7258 , \7259 , \7260 , \7261 ,
         \7262 , \7263 , \7264 , \7265 , \7266 , \7267 , \7268 , \7269 , \7270 , \7271 ,
         \7272 , \7273 , \7274 , \7275 , \7276 , \7277 , \7278 , \7279 , \7280 , \7281 ,
         \7282 , \7283 , \7284 , \7285 , \7286 , \7287 , \7288 , \7289 , \7290 , \7291 ,
         \7292 , \7293 , \7294 , \7295 , \7296 , \7297 , \7298 , \7299 , \7300 , \7301 ,
         \7302 , \7303 , \7304 , \7305 , \7306 , \7307 , \7308 , \7309 , \7310 , \7311 ,
         \7312 , \7313 , \7314 , \7315 , \7316 , \7317 , \7318 , \7319 , \7320 , \7321 ,
         \7322 , \7323 , \7324 , \7325 , \7326 , \7327 , \7328 , \7329 , \7330 , \7331 ,
         \7332 , \7333 , \7334 , \7335 , \7336 , \7337 , \7338 , \7339 , \7340 , \7341 ,
         \7342 , \7343 , \7344 , \7345 , \7346 , \7347 , \7348 , \7349 , \7350 , \7351 ,
         \7352 , \7353 , \7354 , \7355 , \7356 , \7357 , \7358 , \7359 , \7360 , \7361 ,
         \7362 , \7363 , \7364 , \7365 , \7366 , \7367 , \7368 , \7369 , \7370 , \7371 ,
         \7372 , \7373 , \7374 , \7375 , \7376 , \7377 , \7378 , \7379 , \7380 , \7381 ,
         \7382 , \7383 , \7384 , \7385 , \7386 , \7387 , \7388 , \7389 , \7390 , \7391 ,
         \7392 , \7393 , \7394 , \7395 , \7396 , \7397 , \7398 , \7399 , \7400 , \7401 ,
         \7402 , \7403 , \7404 , \7405 , \7406 , \7407 , \7408 , \7409 , \7410 , \7411 ,
         \7412 , \7413 , \7414 , \7415 , \7416 , \7417 , \7418 , \7419 , \7420 , \7421 ,
         \7422 , \7423 , \7424 , \7425 , \7426 , \7427 , \7428 , \7429 , \7430 , \7431 ,
         \7432 , \7433 , \7434 , \7435 , \7436 , \7437 , \7438 , \7439 , \7440 , \7441 ,
         \7442 , \7443 , \7444 , \7445 , \7446 , \7447 , \7448 , \7449 , \7450 , \7451 ,
         \7452 , \7453 , \7454 , \7455 , \7456 , \7457 , \7458 , \7459 , \7460 , \7461 ,
         \7462 , \7463 , \7464 , \7465 , \7466 , \7467 , \7468 , \7469 , \7470 , \7471 ,
         \7472 , \7473 , \7474 , \7475 , \7476 , \7477 , \7478 , \7479 , \7480 , \7481 ,
         \7482 , \7483 , \7484 , \7485 , \7486 , \7487 , \7488 , \7489 , \7490 , \7491 ,
         \7492 , \7493 , \7494 , \7495 , \7496 , \7497 , \7498 , \7499 , \7500 , \7501 ,
         \7502 , \7503 , \7504 , \7505 , \7506 , \7507 , \7508 , \7509 , \7510 , \7511 ,
         \7512 , \7513 , \7514 , \7515 , \7516 , \7517 , \7518 , \7519 , \7520 , \7521 ,
         \7522 , \7523 , \7524 , \7525 , \7526 , \7527 , \7528 , \7529 , \7530 , \7531 ,
         \7532 , \7533 , \7534 , \7535 , \7536 , \7537 , \7538 ;
buf \U$labaj781 ( \o[31] , \7297 );
buf \U$labaj782 ( \o[30] , \7310 );
buf \U$labaj783 ( \o[29] , \7323 );
buf \U$labaj784 ( \o[28] , \7330 );
buf \U$labaj785 ( \o[27] , \7340 );
buf \U$labaj786 ( \o[26] , \7352 );
buf \U$labaj787 ( \o[25] , \7364 );
buf \U$labaj788 ( \o[24] , \7371 );
buf \U$labaj789 ( \o[23] , \7393 );
buf \U$labaj790 ( \o[22] , \7400 );
buf \U$labaj791 ( \o[21] , \7411 );
buf \U$labaj792 ( \o[20] , \7435 );
buf \U$labaj793 ( \o[19] , \7429 );
buf \U$labaj794 ( \o[18] , \7441 );
buf \U$labaj795 ( \o[17] , \7452 );
buf \U$labaj796 ( \o[16] , \7471 );
buf \U$labaj797 ( \o[15] , \7465 );
buf \U$labaj798 ( \o[14] , \7477 );
buf \U$labaj799 ( \o[13] , \7490 );
buf \U$labaj800 ( \o[12] , \7496 );
buf \U$labaj801 ( \o[11] , \7509 );
buf \U$labaj802 ( \o[10] , \7538 );
buf \U$labaj803 ( \o[9] , \7530 );
buf \U$labaj804 ( \o[8] , \7529 );
buf \U$labaj805 ( \o[7] , \7514 );
buf \U$labaj806 ( \o[6] , \7531 );
buf \U$labaj807 ( \o[5] , \7533 );
buf \U$labaj808 ( \o[4] , \7534 );
buf \U$labaj809 ( \o[3] , \7535 );
buf \U$labaj810 ( \o[2] , \7536 );
buf \U$labaj811 ( \o[1] , \7525 );
buf \U$labaj812 ( \o[0] , \7526 );
xor \g45314/U$1 ( \195 , \s[22] , \s[4] );
and \g3018/U$2 ( \196 , \s[12] , \s[6] );
not \g3018/U$4 ( \197 , \s[12] );
not \g3044/U$1 ( \198 , \s[6] );
and \g3018/U$3 ( \199 , \197 , \198 );
nor \g3018/U$1 ( \200 , \196 , \199 );
xor \g2987/U$1 ( \201 , \195 , \200 );
not \g2975/U$3 ( \202 , \201 );
xnor \g3084/U$1 ( \203 , \s[20] , \s[19] );
not \g2995/U$3 ( \204 , \203 );
and \g3026/U$2 ( \205 , \s[26] , \s[16] );
not \g3026/U$4 ( \206 , \s[26] );
not \g3052/U$1 ( \207 , \s[16] );
and \g3026/U$3 ( \208 , \206 , \207 );
nor \g3026/U$1 ( \209 , \205 , \208 );
not \g2995/U$4 ( \210 , \209 );
and \g2995/U$2 ( \211 , \204 , \210 );
and \g2995/U$5 ( \212 , \203 , \209 );
nor \g2995/U$1 ( \213 , \211 , \212 );
not \g2975/U$4 ( \214 , \213 );
or \g2975/U$2 ( \215 , \202 , \214 );
or \g2975/U$5 ( \216 , \213 , \201 );
nand \g2975/U$1 ( \217 , \215 , \216 );
not \g2974/U$1 ( \218 , \217 );
not \g45820/U$3 ( \219 , \218 );
xor \g45317/U$1 ( \220 , \s[31] , \s[0] );
and \g3001/U$2 ( \221 , \s[14] , \s[13] );
not \g3001/U$4 ( \222 , \s[14] );
not \g3046/U$1 ( \223 , \s[13] );
and \g3001/U$3 ( \224 , \222 , \223 );
nor \g3001/U$1 ( \225 , \221 , \224 );
xor \g2986/U$1 ( \226 , \220 , \225 );
not \g2981/U$3 ( \227 , \226 );
xor \g45833/U$1 ( \228 , \s[30] , \s[1] );
and \g3031/U$2 ( \229 , \s[10] , \s[2] );
not \g3031/U$4 ( \230 , \s[10] );
not \g3059/U$1 ( \231 , \s[2] );
and \g3031/U$3 ( \232 , \230 , \231 );
nor \g3031/U$1 ( \233 , \229 , \232 );
xnor \g2992/U$1 ( \234 , \228 , \233 );
not \g2981/U$4 ( \235 , \234 );
and \g2981/U$2 ( \236 , \227 , \235 );
and \g2981/U$5 ( \237 , \234 , \226 );
nor \g2981/U$1 ( \238 , \236 , \237 );
not \g2980/U$1 ( \239 , \238 );
not \g45820/U$4 ( \240 , \239 );
or \g45820/U$2 ( \241 , \219 , \240 );
nand \g2969/U$1 ( \242 , \238 , \217 );
nand \g45820/U$1 ( \243 , \241 , \242 );
and \g3006/U$2 ( \244 , \s[29] , \s[3] );
not \g3006/U$4 ( \245 , \s[29] );
not \g3056/U$1 ( \246 , \s[3] );
and \g3006/U$3 ( \247 , \245 , \246 );
nor \g3006/U$1 ( \248 , \244 , \247 );
xor \g45664/U$1 ( \249 , \s[27] , \s[15] );
xor \g45562/U$1 ( \250 , \248 , \249 );
not \g2973/U$3 ( \251 , \250 );
and \g3017/U$2 ( \252 , \s[24] , \s[17] );
not \g3017/U$4 ( \253 , \s[24] );
not \g3051/U$1 ( \254 , \s[17] );
and \g3017/U$3 ( \255 , \253 , \254 );
nor \g3017/U$1 ( \256 , \252 , \255 );
not \g3016/U$1 ( \257 , \256 );
not \g2988/U$3 ( \258 , \257 );
and \g3013/U$2 ( \259 , \s[11] , \s[5] );
not \g3013/U$4 ( \260 , \s[11] );
not \g3050/U$1 ( \261 , \s[5] );
and \g3013/U$3 ( \262 , \260 , \261 );
nor \g3013/U$1 ( \263 , \259 , \262 );
not \g2988/U$4 ( \264 , \263 );
and \g2988/U$2 ( \265 , \258 , \264 );
and \g2988/U$5 ( \266 , \257 , \263 );
nor \g2988/U$1 ( \267 , \265 , \266 );
not \g2973/U$4 ( \268 , \267 );
or \g2973/U$2 ( \269 , \251 , \268 );
or \g2973/U$5 ( \270 , \250 , \267 );
nand \g2973/U$1 ( \271 , \269 , \270 );
and \g3033/U$2 ( \272 , \s[21] , \s[9] );
not \g3033/U$4 ( \273 , \s[21] );
not \g3045/U$1 ( \274 , \s[9] );
and \g3033/U$3 ( \275 , \273 , \274 );
nor \g3033/U$1 ( \276 , \272 , \275 );
xor \g3096/U$1 ( \277 , \s[23] , \s[18] );
xor \g3/U$1 ( \278 , \276 , \277 );
and \g3024/U$2 ( \279 , \s[28] , \s[7] );
not \g3024/U$4 ( \280 , \s[28] );
not \g3064/U$1 ( \281 , \s[7] );
and \g3024/U$3 ( \282 , \280 , \281 );
nor \g3024/U$1 ( \283 , \279 , \282 );
and \g3028/U$2 ( \284 , \s[25] , \s[8] );
not \g3028/U$4 ( \285 , \s[25] );
not \g3058/U$1 ( \286 , \s[8] );
and \g3028/U$3 ( \287 , \285 , \286 );
nor \g3028/U$1 ( \288 , \284 , \287 );
xor \g2994/U$1 ( \289 , \283 , \288 );
xnor \g3/U$1_r1 ( \290 , \278 , \289 );
xor \g45547/U$1 ( \291 , \271 , \290 );
xor \g45311/U$1 ( \292 , \243 , \291 );
buf \g2939/U$1 ( \293 , \292 );
not \g2932/U$1 ( \294 , \293 );
buf \g2920/U$1 ( \295 , \294 );
buf \g2929/U$1 ( \296 , \295 );
buf \g2928/U$1 ( \297 , \296 );
not \g2924/U$1 ( \298 , \297 );
xor \g45767/U$1 ( \299 , \c[31] , \d[31] );
not \sub_5_33_g9561/U$2 ( \300 , \c[19] );
nand \sub_5_33_g9561/U$1 ( \301 , \300 , \d[19] );
not \sub_5_33_g9581/U$2 ( \302 , \c[18] );
nand \sub_5_33_g9581/U$1 ( \303 , \302 , \d[18] );
and \sub_5_33_g9332/U$1 ( \304 , \301 , \303 );
not \sub_5_33_g9547/U$2 ( \305 , \304 );
not \sub_5_33_g9557/U$2 ( \306 , \c[17] );
nand \sub_5_33_g9557/U$1 ( \307 , \306 , \d[17] );
not \sub_5_33_g9563/U$2 ( \308 , \c[16] );
nand \sub_5_33_g9563/U$1 ( \309 , \308 , \d[16] );
nand \sub_5_33_g9351/U$1 ( \310 , \307 , \309 );
nor \sub_5_33_g9547/U$1 ( \311 , \305 , \310 );
not \sub_5_33_g9309/U$3 ( \312 , \d[21] );
not \sub_5_33_g9500/U$1 ( \313 , \c[21] );
not \sub_5_33_g9309/U$4 ( \314 , \313 );
or \sub_5_33_g9309/U$2 ( \315 , \312 , \314 );
not \sub_5_33_g9580/U$2 ( \316 , \c[20] );
nand \sub_5_33_g9580/U$1 ( \317 , \316 , \d[20] );
nand \sub_5_33_g9309/U$1 ( \318 , \315 , \317 );
not \sub_5_33_g9585/U$2 ( \319 , \c[23] );
nand \sub_5_33_g9585/U$1 ( \320 , \319 , \d[23] );
not \sub_5_33_g9571/U$2 ( \321 , \c[22] );
nand \sub_5_33_g9571/U$1 ( \322 , \321 , \d[22] );
nand \sub_5_33_g9334/U$1 ( \323 , \320 , \322 );
nor \sub_5_33_g9227/U$1 ( \324 , \318 , \323 );
nand \sub_5_33_g9207/U$1 ( \325 , \311 , \324 );
not \sub_5_33_g9206/U$1 ( \326 , \325 );
not \sub_5_33_g9503/U$1 ( \327 , \d[28] );
or \sub_5_33_g9449/U$1 ( \328 , \327 , \c[28] );
not \sub_5_33_g9446/U$2 ( \329 , \c[29] );
nand \sub_5_33_g9446/U$1 ( \330 , \329 , \d[29] );
nand \sub_5_33_g9354/U$1 ( \331 , \328 , \330 );
not \sub_5_33_g9222/U$2 ( \332 , \331 );
not \sub_5_33_g9361/U$2 ( \333 , \c[30] );
nand \sub_5_33_g9361/U$1 ( \334 , \333 , \d[30] );
nand \sub_5_33_g9222/U$1 ( \335 , \332 , \334 );
not \sub_5_33_g9568/U$2 ( \336 , \c[27] );
nand \sub_5_33_g9568/U$1 ( \337 , \336 , \d[27] );
not \sub_5_33_g9579/U$2 ( \338 , \c[26] );
nand \sub_5_33_g9579/U$1 ( \339 , \338 , \d[26] );
and \sub_5_33_g9314/U$1 ( \340 , \337 , \339 );
not \sub_5_33_g9545/U$2 ( \341 , \340 );
not \sub_5_33_g9564/U$2 ( \342 , \c[25] );
nand \sub_5_33_g9564/U$1 ( \343 , \342 , \d[25] );
not \sub_5_33_g9573/U$2 ( \344 , \c[24] );
nand \sub_5_33_g9573/U$1 ( \345 , \344 , \d[24] );
nand \sub_5_33_g9284/U$1 ( \346 , \343 , \345 );
nor \sub_5_33_g9545/U$1 ( \347 , \341 , \346 );
not \sub_5_33_g9225/U$1 ( \348 , \347 );
nor \sub_5_33_g9208/U$1 ( \349 , \335 , \348 );
and \sub_5_33_g9175/U$1 ( \350 , \326 , \349 );
not \sub_5_33_g9089/U$3 ( \351 , \350 );
not \sub_5_33_g9588/U$2 ( \352 , \c[15] );
nand \sub_5_33_g9588/U$1 ( \353 , \352 , \d[15] );
not \g45697/U$2 ( \354 , \c[14] );
nand \g45697/U$1 ( \355 , \354 , \d[14] );
and \sub_5_33_g9531/U$1 ( \356 , \353 , \355 );
not \sub_5_33_g9198/U$3 ( \357 , \356 );
not \sub_5_33_g9592/U$2 ( \358 , \c[13] );
nand \sub_5_33_g9592/U$1 ( \359 , \358 , \d[13] );
not \sub_5_33_g9266/U$3 ( \360 , \359 );
not \sub_5_33_g45808/U$2 ( \361 , \c[12] );
nor \sub_5_33_g45808/U$1 ( \362 , \361 , \d[12] );
not \sub_5_33_g9266/U$4 ( \363 , \362 );
or \sub_5_33_g9266/U$2 ( \364 , \360 , \363 );
not \sub_5_33_g9582/U$2 ( \365 , \d[13] );
nand \sub_5_33_g9582/U$1 ( \366 , \365 , \c[13] );
nand \sub_5_33_g9266/U$1 ( \367 , \364 , \366 );
not \sub_5_33_g9198/U$4 ( \368 , \367 );
or \sub_5_33_g9198/U$2 ( \369 , \357 , \368 );
not \sub_5_33_g9396/U$2 ( \370 , \c[14] );
nor \sub_5_33_g9396/U$1 ( \371 , \370 , \d[14] );
and \sub_5_33_g9264/U$2 ( \372 , \371 , \353 );
not \sub_5_33_g9587/U$2 ( \373 , \c[15] );
nor \sub_5_33_g9587/U$1 ( \374 , \373 , \d[15] );
nor \sub_5_33_g9264/U$1 ( \375 , \372 , \374 );
nand \sub_5_33_g9198/U$1 ( \376 , \369 , \375 );
not \sub_5_33_g9197/U$1 ( \377 , \376 );
not \sub_5_33_g9562/U$2 ( \378 , \c[7] );
nand \sub_5_33_g9562/U$1 ( \379 , \378 , \d[7] );
not \sub_5_33_g9558/U$2 ( \380 , \c[11] );
nand \sub_5_33_g9558/U$1 ( \381 , \380 , \d[11] );
and \sub_5_33_g9529/U$1 ( \382 , \379 , \359 , \353 , \381 );
not \sub_5_33_g9578/U$2 ( \383 , \c[9] );
nand \sub_5_33_g9578/U$1 ( \384 , \383 , \d[9] );
not \sub_5_33_g9565/U$2 ( \385 , \c[8] );
nand \sub_5_33_g9565/U$1 ( \386 , \385 , \d[8] );
and \sub_5_33_g9289/U$1 ( \387 , \384 , \386 );
not \sub_5_33_g45650/U$2 ( \388 , \c[5] );
nand \sub_5_33_g45650/U$1 ( \389 , \388 , \d[5] );
not \g45699/U$2 ( \390 , \c[4] );
nand \g45699/U$1 ( \391 , \390 , \d[4] );
nand \sub_5_33_g9300/U$1 ( \392 , \389 , \391 );
not \sub_5_33_g9299/U$1 ( \393 , \392 );
not \sub_5_33_g9455/U$2 ( \394 , \c[12] );
nand \sub_5_33_g9455/U$1 ( \395 , \394 , \d[12] );
not \sub_5_33_g9567/U$2 ( \396 , \c[6] );
nand \sub_5_33_g9567/U$1 ( \397 , \396 , \d[6] );
nand \sub_5_33_g9323/U$1 ( \398 , \395 , \397 );
not \sub_5_33_g9434/U$2 ( \399 , \c[14] );
nand \sub_5_33_g9434/U$1 ( \400 , \399 , \d[14] );
not \g45698/U$2 ( \401 , \c[10] );
nand \g45698/U$1 ( \402 , \401 , \d[10] );
nand \sub_5_33_g9316/U$1 ( \403 , \400 , \402 );
nor \sub_5_33_g9277/U$1 ( \404 , \398 , \403 );
and \sub_5_33_g9189/U$1 ( \405 , \382 , \387 , \393 , \404 );
not \sub_5_33_g9377/U$2 ( \406 , \c[0] );
nand \sub_5_33_g9377/U$1 ( \407 , \406 , \d[0] );
not \sub_5_33_g9187/U$3 ( \408 , \407 );
not \sub_5_33_g9368/U$2 ( \409 , \c[1] );
nand \sub_5_33_g9368/U$1 ( \410 , \409 , \d[1] );
not \sub_5_33_g9187/U$4 ( \411 , \410 );
or \sub_5_33_g9187/U$2 ( \412 , \408 , \411 );
not \sub_5_33_g9575/U$2 ( \413 , \d[1] );
nand \sub_5_33_g9575/U$1 ( \414 , \413 , \c[1] );
nand \sub_5_33_g9187/U$1 ( \415 , \412 , \414 );
not \sub_5_33_g9521/U$3 ( \416 , \415 );
not \sub_5_33_g9472/U$2 ( \417 , \c[3] );
nand \sub_5_33_g9472/U$1 ( \418 , \417 , \d[3] );
not \sub_5_33_g9589/U$2 ( \419 , \c[2] );
nand \sub_5_33_g9589/U$1 ( \420 , \419 , \d[2] );
and \sub_5_33_g9355/U$1 ( \421 , \418 , \420 );
not \sub_5_33_g9521/U$4 ( \422 , \421 );
or \sub_5_33_g9521/U$2 ( \423 , \416 , \422 );
not \sub_5_33_g9474/U$2 ( \424 , \c[2] );
nor \sub_5_33_g9474/U$1 ( \425 , \424 , \d[2] );
not \sub_5_33_g9268/U$3 ( \426 , \425 );
not \sub_5_33_g9268/U$4 ( \427 , \418 );
or \sub_5_33_g9268/U$2 ( \428 , \426 , \427 );
not \sub_5_33_g9577/U$2 ( \429 , \d[3] );
nand \sub_5_33_g9577/U$1 ( \430 , \429 , \c[3] );
nand \sub_5_33_g9268/U$1 ( \431 , \428 , \430 );
not \sub_5_33_g9267/U$1 ( \432 , \431 );
nand \sub_5_33_g9521/U$1 ( \433 , \423 , \432 );
nand \sub_5_33_g9125/U$1 ( \434 , \405 , \433 );
not \sub_5_33_g9569/U$2 ( \435 , \c[12] );
nand \sub_5_33_g9569/U$1 ( \436 , \435 , \d[12] );
nand \sub_5_33_g9348/U$1 ( \437 , \359 , \436 );
not \sub_5_33_g9347/U$1 ( \438 , \437 );
nand \sub_5_33_g9232/U$1 ( \439 , \356 , \438 );
not \sub_5_33_g9534/U$2 ( \440 , \439 );
and \sub_5_33_g9530/U$1 ( \441 , \381 , \402 );
not \sub_5_33_g9196/U$3 ( \442 , \441 );
not \sub_5_33_g9404/U$2 ( \443 , \c[8] );
nor \sub_5_33_g9404/U$1 ( \444 , \443 , \d[8] );
not \sub_5_33_g9260/U$3 ( \445 , \444 );
not \sub_5_33_g9260/U$4 ( \446 , \384 );
or \sub_5_33_g9260/U$2 ( \447 , \445 , \446 );
not \sub_5_33_g9591/U$2 ( \448 , \d[9] );
nand \sub_5_33_g9591/U$1 ( \449 , \448 , \c[9] );
nand \sub_5_33_g9260/U$1 ( \450 , \447 , \449 );
not \sub_5_33_g9196/U$4 ( \451 , \450 );
or \sub_5_33_g9196/U$2 ( \452 , \442 , \451 );
not \sub_5_33_g9255/U$3 ( \453 , \381 );
not \sub_5_33_g9429/U$2 ( \454 , \c[10] );
nor \sub_5_33_g9429/U$1 ( \455 , \454 , \d[10] );
not \sub_5_33_g9255/U$4 ( \456 , \455 );
or \sub_5_33_g9255/U$2 ( \457 , \453 , \456 );
not \sub_5_33_g9590/U$2 ( \458 , \d[11] );
nand \sub_5_33_g9590/U$1 ( \459 , \458 , \c[11] );
nand \sub_5_33_g9255/U$1 ( \460 , \457 , \459 );
not \sub_5_33_g9254/U$1 ( \461 , \460 );
nand \sub_5_33_g9196/U$1 ( \462 , \452 , \461 );
nand \sub_5_33_g9534/U$1 ( \463 , \440 , \462 );
nand \sub_5_33_g9237/U$1 ( \464 , \387 , \441 );
nor \sub_5_33_g9216/U$1 ( \465 , \464 , \439 );
not \sub_5_33_g9249/U$3 ( \466 , \389 );
not \sub_5_33_g9379/U$2 ( \467 , \c[4] );
nor \sub_5_33_g9379/U$1 ( \468 , \467 , \d[4] );
not \sub_5_33_g9249/U$4 ( \469 , \468 );
or \sub_5_33_g9249/U$2 ( \470 , \466 , \469 );
not \sub_5_33_g9593/U$2 ( \471 , \d[5] );
nand \sub_5_33_g9593/U$1 ( \472 , \471 , \c[5] );
nand \sub_5_33_g9249/U$1 ( \473 , \470 , \472 );
not \sub_5_33_g9200/U$3 ( \474 , \473 );
and \sub_5_33_g9282/U$1 ( \475 , \379 , \397 );
not \sub_5_33_g9200/U$4 ( \476 , \475 );
or \sub_5_33_g9200/U$2 ( \477 , \474 , \476 );
not \sub_5_33_g9394/U$2 ( \478 , \c[6] );
nor \sub_5_33_g9394/U$1 ( \479 , \478 , \d[6] );
not \sub_5_33_g9257/U$3 ( \480 , \479 );
not \sub_5_33_g9257/U$4 ( \481 , \379 );
or \sub_5_33_g9257/U$2 ( \482 , \480 , \481 );
not \sub_5_33_g9566/U$2 ( \483 , \d[7] );
nand \sub_5_33_g9566/U$1 ( \484 , \483 , \c[7] );
nand \sub_5_33_g9257/U$1 ( \485 , \482 , \484 );
not \sub_5_33_g9256/U$1 ( \486 , \485 );
nand \sub_5_33_g9200/U$1 ( \487 , \477 , \486 );
nand \sub_5_33_g9168/U$1 ( \488 , \465 , \487 );
nand \sub_5_33_g9119/U$1 ( \489 , \377 , \434 , \463 , \488 );
buf \fopt45582/U$1 ( \490 , \489 );
not \sub_5_33_g9089/U$4 ( \491 , \490 );
or \sub_5_33_g9089/U$2 ( \492 , \351 , \491 );
not \sub_5_33_g9155/U$3 ( \493 , \324 );
not \sub_5_33_g9263/U$3 ( \494 , \307 );
not \sub_5_33_g9360/U$2 ( \495 , \c[16] );
nor \sub_5_33_g9360/U$1 ( \496 , \495 , \d[16] );
not \sub_5_33_g9263/U$4 ( \497 , \496 );
or \sub_5_33_g9263/U$2 ( \498 , \494 , \497 );
not \sub_5_33_g9559/U$2 ( \499 , \d[17] );
nand \sub_5_33_g9559/U$1 ( \500 , \499 , \c[17] );
nand \sub_5_33_g9263/U$1 ( \501 , \498 , \500 );
not \sub_5_33_g9191/U$3 ( \502 , \501 );
not \sub_5_33_g9191/U$4 ( \503 , \304 );
or \sub_5_33_g9191/U$2 ( \504 , \502 , \503 );
not \sub_5_33_g9458/U$2 ( \505 , \c[18] );
nor \sub_5_33_g9458/U$1 ( \506 , \505 , \d[18] );
not \sub_5_33_g9253/U$3 ( \507 , \506 );
not \sub_5_33_g9253/U$4 ( \508 , \301 );
or \sub_5_33_g9253/U$2 ( \509 , \507 , \508 );
not \sub_5_33_g9576/U$2 ( \510 , \d[19] );
nand \sub_5_33_g9576/U$1 ( \511 , \510 , \c[19] );
nand \sub_5_33_g9253/U$1 ( \512 , \509 , \511 );
not \sub_5_33_g9252/U$1 ( \513 , \512 );
nand \sub_5_33_g9191/U$1 ( \514 , \504 , \513 );
not \sub_5_33_g9155/U$4 ( \515 , \514 );
or \sub_5_33_g9155/U$2 ( \516 , \493 , \515 );
not \sub_5_33_g9333/U$1 ( \517 , \323 );
not \sub_5_33_g9202/U$3 ( \518 , \517 );
not \sub_5_33_g9476/U$2 ( \519 , \c[20] );
nor \sub_5_33_g9476/U$1 ( \520 , \519 , \d[20] );
not \sub_5_33_g9246/U$3 ( \521 , \520 );
nand \sub_5_33_g9437/U$1 ( \522 , \313 , \d[21] );
not \sub_5_33_g9246/U$4 ( \523 , \522 );
or \sub_5_33_g9246/U$2 ( \524 , \521 , \523 );
not \sub_5_33_g9584/U$2 ( \525 , \d[21] );
nand \sub_5_33_g9584/U$1 ( \526 , \525 , \c[21] );
nand \sub_5_33_g9246/U$1 ( \527 , \524 , \526 );
not \sub_5_33_g9202/U$4 ( \528 , \527 );
or \sub_5_33_g9202/U$2 ( \529 , \518 , \528 );
not \sub_5_33_g9270/U$3 ( \530 , \320 );
not \sub_5_33_g9468/U$2 ( \531 , \c[22] );
nor \sub_5_33_g9468/U$1 ( \532 , \531 , \d[22] );
not \sub_5_33_g9270/U$4 ( \533 , \532 );
or \sub_5_33_g9270/U$2 ( \534 , \530 , \533 );
not \sub_5_33_g9570/U$2 ( \535 , \d[23] );
nand \sub_5_33_g9570/U$1 ( \536 , \535 , \c[23] );
nand \sub_5_33_g9270/U$1 ( \537 , \534 , \536 );
not \sub_5_33_g9269/U$1 ( \538 , \537 );
nand \sub_5_33_g9202/U$1 ( \539 , \529 , \538 );
not \sub_5_33_g9201/U$1 ( \540 , \539 );
nand \sub_5_33_g9155/U$1 ( \541 , \516 , \540 );
and \sub_5_33_g9130/U$2 ( \542 , \541 , \349 );
not \sub_5_33_g9251/U$3 ( \543 , \343 );
not \sub_5_33_g9451/U$2 ( \544 , \c[24] );
nor \sub_5_33_g9451/U$1 ( \545 , \544 , \d[24] );
not \sub_5_33_g9251/U$4 ( \546 , \545 );
or \sub_5_33_g9251/U$2 ( \547 , \543 , \546 );
not \sub_5_33_g9560/U$2 ( \548 , \d[25] );
nand \sub_5_33_g9560/U$1 ( \549 , \548 , \c[25] );
nand \sub_5_33_g9251/U$1 ( \550 , \547 , \549 );
not \sub_5_33_g9193/U$3 ( \551 , \550 );
not \sub_5_33_g9193/U$4 ( \552 , \340 );
or \sub_5_33_g9193/U$2 ( \553 , \551 , \552 );
not \sub_5_33_g9444/U$2 ( \554 , \c[26] );
nor \sub_5_33_g9444/U$1 ( \555 , \554 , \d[26] );
not \sub_5_33_g9272/U$3 ( \556 , \555 );
not \sub_5_33_g9272/U$4 ( \557 , \337 );
or \sub_5_33_g9272/U$2 ( \558 , \556 , \557 );
not \sub_5_33_g9583/U$2 ( \559 , \d[27] );
nand \sub_5_33_g9583/U$1 ( \560 , \559 , \c[27] );
nand \sub_5_33_g9272/U$1 ( \561 , \558 , \560 );
not \sub_5_33_g9271/U$1 ( \562 , \561 );
nand \sub_5_33_g9193/U$1 ( \563 , \553 , \562 );
not \sub_5_33_g9192/U$1 ( \564 , \563 );
or \sub_5_33_g9161/U$2 ( \565 , \564 , \335 );
not \sub_5_33_g9445/U$1 ( \566 , \330 );
nand \sub_5_33_g9443/U$1 ( \567 , \327 , \c[28] );
or \sub_5_33_g9243/U$2 ( \568 , \566 , \567 );
not \sub_5_33_g9400/U$2 ( \569 , \d[29] );
nand \sub_5_33_g9400/U$1 ( \570 , \569 , \c[29] );
nand \sub_5_33_g9243/U$1 ( \571 , \568 , \570 );
and \sub_5_33_g9182/U$2 ( \572 , \571 , \334 );
not \sub_5_33_g9366/U$2 ( \573 , \c[30] );
nor \sub_5_33_g9366/U$1 ( \574 , \573 , \d[30] );
nor \sub_5_33_g9182/U$1 ( \575 , \572 , \574 );
nand \sub_5_33_g9161/U$1 ( \576 , \565 , \575 );
nor \sub_5_33_g9130/U$1 ( \577 , \542 , \576 );
nand \sub_5_33_g9089/U$1 ( \578 , \492 , \577 );
xnor \g45767/U$1_r1 ( \579 , \299 , \578 );
and \g2878/U$2 ( \580 , \298 , \579 );
not \g2878/U$4 ( \581 , \298 );
nor \add_5_20_g13942/U$1 ( \582 , \c[19] , \d[19] );
nor \add_5_20_g13970/U$1 ( \583 , \c[18] , \d[18] );
nor \add_5_20_g13837/U$1 ( \584 , \582 , \583 );
nor \add_5_20_g13975/U$1 ( \585 , \c[17] , \d[17] );
nor \add_5_20_g13899/U$1 ( \586 , \c[16] , \d[16] );
nor \add_5_20_g13815/U$1 ( \587 , \585 , \586 );
and \add_5_20_g13747/U$1 ( \588 , \584 , \587 );
nor \add_5_20_g13912/U$1 ( \589 , \c[21] , \d[21] );
nor \add_5_20_g13885/U$1 ( \590 , \c[20] , \d[20] );
nor \add_5_20_g13825/U$1 ( \591 , \589 , \590 );
nor \add_5_20_g13991/U$1 ( \592 , \c[22] , \d[22] );
nor \add_5_20_g13877/U$1 ( \593 , \c[23] , \d[23] );
nor \add_5_20_g13799/U$1 ( \594 , \592 , \593 );
and \add_5_20_g2/U$1 ( \595 , \591 , \594 );
nand \add_5_20_g13727/U$1 ( \596 , \588 , \595 );
not \add_5_20_g13725/U$1 ( \597 , \596 );
nor \add_5_20_g13869/U$1 ( \598 , \c[30] , \d[30] );
not \add_5_20_g13755/U$2 ( \599 , \598 );
nor \add_5_20_g13895/U$1 ( \600 , \c[29] , \d[29] );
nor \add_5_20_g13928/U$1 ( \601 , \c[28] , \d[28] );
nor \add_5_20_g13855/U$1 ( \602 , \600 , \601 );
nand \add_5_20_g13755/U$1 ( \603 , \599 , \602 );
nor \add_5_20_g13958/U$1 ( \604 , \c[27] , \d[27] );
nor \add_5_20_g13930/U$1 ( \605 , \c[26] , \d[26] );
nor \add_5_20_g13836/U$1 ( \606 , \604 , \605 );
nor \add_5_20_g13995/U$1 ( \607 , \c[25] , \d[25] );
nor \add_5_20_g13873/U$1 ( \608 , \c[24] , \d[24] );
nor \add_5_20_g13811/U$1 ( \609 , \607 , \608 );
and \add_5_20_g13752/U$1 ( \610 , \606 , \609 );
not \add_5_20_g13751/U$1 ( \611 , \610 );
nor \add_5_20_g13735/U$1 ( \612 , \603 , \611 );
and \add_5_20_g13691/U$1 ( \613 , \597 , \612 );
not \add_5_20_g13616/U$3 ( \614 , \613 );
nor \add_5_20_g14006/U$1 ( \615 , \c[3] , \d[3] );
nor \add_5_20_g13946/U$1 ( \616 , \c[2] , \d[2] );
nor \add_5_20_g13856/U$1 ( \617 , \615 , \616 );
not \add_5_20_g13664/U$3 ( \618 , \617 );
nor \add_5_20_g13879/U$1 ( \619 , \c[1] , \d[1] );
nand \g45804/U$2 ( \620 , \c[0] , \d[0] );
or \add_5_20_g13695/U$2 ( \621 , \619 , \620 );
nand \add_5_20_g13926/U$1 ( \622 , \c[1] , \d[1] );
nand \add_5_20_g13695/U$1 ( \623 , \621 , \622 );
not \add_5_20_g13664/U$4 ( \624 , \623 );
or \add_5_20_g13664/U$2 ( \625 , \618 , \624 );
not \add_5_20_g13768/U$3 ( \626 , \615 );
nand \add_5_20_g14007/U$1 ( \627 , \c[2] , \d[2] );
not \add_5_20_g13768/U$4 ( \628 , \627 );
and \add_5_20_g13768/U$2 ( \629 , \626 , \628 );
nand \add_5_20_g13966/U$1 ( \630 , \c[3] , \d[3] );
not \add_5_20_g13965/U$1 ( \631 , \630 );
nor \add_5_20_g13768/U$1 ( \632 , \629 , \631 );
nand \add_5_20_g13664/U$1 ( \633 , \625 , \632 );
nor \add_5_20_g13998/U$1 ( \634 , \c[7] , \d[7] );
not \add_5_20_g13997/U$1 ( \635 , \634 );
nor \add_5_20_g14008/U$1 ( \636 , \c[11] , \d[11] );
not \add_5_20_g13923/U$1 ( \637 , \636 );
or \g45657/U$1 ( \638 , \c[13] , \d[13] );
or \add_5_20_g14037/U$1 ( \639 , \d[15] , \c[15] );
nand \add_5_20_g13788/U$1 ( \640 , \635 , \637 , \638 , \639 );
nor \add_5_20_g13960/U$1 ( \641 , \c[4] , \d[4] );
nor \add_5_20_g13901/U$1 ( \642 , \c[5] , \d[5] );
nor \add_5_20_g13807/U$1 ( \643 , \641 , \642 );
nor \add_5_20_g13881/U$1 ( \644 , \c[9] , \d[9] );
nor \add_5_20_g45622/U$1 ( \645 , \c[8] , \d[8] );
nor \add_5_20_g13798/U$1 ( \646 , \644 , \645 );
nand \add_5_20_g13740/U$1 ( \647 , \643 , \646 );
nor \add_5_20_g13974/U$1 ( \648 , \c[10] , \d[10] );
not \add_5_20_g13973/U$1 ( \649 , \648 );
nor \add_5_20_g14009/U$1 ( \650 , \c[14] , \d[14] );
not \add_5_20_g13987/U$1 ( \651 , \650 );
nor \add_5_20_g13941/U$1 ( \652 , \c[6] , \d[6] );
not \add_5_20_g13940/U$1 ( \653 , \652 );
nor \add_5_20_g14010/U$1 ( \654 , \c[12] , \d[12] );
not \add_5_20_g13976/U$1 ( \655 , \654 );
nand \add_5_20_g13786/U$1 ( \656 , \649 , \651 , \653 , \655 );
nor \add_5_20_g13696/U$1 ( \657 , \640 , \647 , \656 );
nand \add_5_20_g13656/U$1 ( \658 , \633 , \657 );
nand \add_5_20_g13950/U$1 ( \659 , \c[12] , \d[12] );
not \add_5_20_g13949/U$1 ( \660 , \659 );
not \add_5_20_g13767/U$3 ( \661 , \660 );
not \add_5_20_g13767/U$4 ( \662 , \638 );
or \add_5_20_g13767/U$2 ( \663 , \661 , \662 );
nand \add_5_20_g13957/U$1 ( \664 , \c[13] , \d[13] );
nand \add_5_20_g13767/U$1 ( \665 , \663 , \664 );
not \add_5_20_g13893/U$1 ( \666 , \639 );
nor \add_5_20_g13850/U$1 ( \667 , \666 , \650 );
and \add_5_20_g13712/U$2 ( \668 , \665 , \667 );
nand \add_5_20_g13907/U$1 ( \669 , \c[14] , \d[14] );
or \add_5_20_g13779/U$2 ( \670 , \666 , \669 );
nand \add_5_20_g13904/U$1 ( \671 , \c[15] , \d[15] );
nand \add_5_20_g13779/U$1 ( \672 , \670 , \671 );
nor \add_5_20_g13712/U$1 ( \673 , \668 , \672 );
nand \add_5_20_g13936/U$1 ( \674 , \c[8] , \d[8] );
or \add_5_20_g13775/U$2 ( \675 , \674 , \644 );
nand \add_5_20_g13999/U$1 ( \676 , \c[9] , \d[9] );
nand \add_5_20_g13775/U$1 ( \677 , \675 , \676 );
not \add_5_20_g13708/U$3 ( \678 , \677 );
nor \add_5_20_g13838/U$1 ( \679 , \636 , \648 );
not \add_5_20_g13708/U$4 ( \680 , \679 );
or \add_5_20_g13708/U$2 ( \681 , \678 , \680 );
not \add_5_20_g13780/U$3 ( \682 , \636 );
nand \add_5_20_g45809/U$1 ( \683 , \c[10] , \d[10] );
not \add_5_20_g13780/U$4 ( \684 , \683 );
and \add_5_20_g13780/U$2 ( \685 , \682 , \684 );
nand \add_5_20_g13963/U$1 ( \686 , \c[11] , \d[11] );
not \add_5_20_g13962/U$1 ( \687 , \686 );
nor \add_5_20_g13780/U$1 ( \688 , \685 , \687 );
nand \add_5_20_g13708/U$1 ( \689 , \681 , \688 );
nand \add_5_20_g13849/U$1 ( \690 , \639 , \651 );
nand \add_5_20_g13865/U$1 ( \691 , \638 , \655 );
nor \add_5_20_g13754/U$1 ( \692 , \690 , \691 );
nand \add_5_20_g13683/U$1 ( \693 , \689 , \692 );
nand \add_5_20_g13955/U$1 ( \694 , \c[4] , \d[4] );
or \add_5_20_g13772/U$2 ( \695 , \642 , \694 );
nand \add_5_20_g13916/U$1 ( \696 , \c[5] , \d[5] );
nand \add_5_20_g13772/U$1 ( \697 , \695 , \696 );
not \add_5_20_g13715/U$3 ( \698 , \697 );
nor \add_5_20_g13851/U$1 ( \699 , \634 , \652 );
not \add_5_20_g13715/U$4 ( \700 , \699 );
or \add_5_20_g13715/U$2 ( \701 , \698 , \700 );
not \add_5_20_g13783/U$3 ( \702 , \634 );
nand \add_5_20_g13953/U$1 ( \703 , \c[6] , \d[6] );
not \add_5_20_g13783/U$4 ( \704 , \703 );
and \add_5_20_g13783/U$2 ( \705 , \702 , \704 );
nand \add_5_20_g13921/U$1 ( \706 , \c[7] , \d[7] );
not \add_5_20_g13920/U$1 ( \707 , \706 );
nor \add_5_20_g13783/U$1 ( \708 , \705 , \707 );
nand \add_5_20_g13715/U$1 ( \709 , \701 , \708 );
nand \add_5_20_g13784/U$1 ( \710 , \646 , \639 , \638 );
or \g45716/U$1 ( \711 , \636 , \654 , \648 , \650 );
nor \add_5_20_g13736/U$1 ( \712 , \710 , \711 );
nand \add_5_20_g13685/U$1 ( \713 , \709 , \712 );
and \add_5_20_g13643/U$1 ( \714 , \658 , \673 , \693 , \713 );
not \add_5_20_g13642/U$1 ( \715 , \714 );
not \add_5_20_g13616/U$4 ( \716 , \715 );
or \add_5_20_g13616/U$2 ( \717 , \614 , \716 );
not \add_5_20_g14012/U$3 ( \718 , \595 );
nand \add_5_20_g14003/U$1 ( \719 , \c[16] , \d[16] );
or \add_5_20_g13778/U$2 ( \720 , \585 , \719 );
nand \add_5_20_g13918/U$1 ( \721 , \c[17] , \d[17] );
nand \add_5_20_g13778/U$1 ( \722 , \720 , \721 );
not \add_5_20_g13702/U$3 ( \723 , \722 );
not \add_5_20_g13702/U$4 ( \724 , \584 );
or \add_5_20_g13702/U$2 ( \725 , \723 , \724 );
not \add_5_20_g13760/U$3 ( \726 , \582 );
nand \add_5_20_g13910/U$1 ( \727 , \c[18] , \d[18] );
not \add_5_20_g13760/U$4 ( \728 , \727 );
and \add_5_20_g13760/U$2 ( \729 , \726 , \728 );
and \add_5_20_g14015/U$1 ( \730 , \c[19] , \d[19] );
nor \add_5_20_g13760/U$1 ( \731 , \729 , \730 );
nand \add_5_20_g13702/U$1 ( \732 , \725 , \731 );
not \add_5_20_g14012/U$4 ( \733 , \732 );
or \add_5_20_g14012/U$2 ( \734 , \718 , \733 );
nand \add_5_20_g13888/U$1 ( \735 , \c[20] , \d[20] );
not \add_5_20_g13887/U$1 ( \736 , \735 );
not \add_5_20_g13764/U$3 ( \737 , \736 );
not \add_5_20_g13911/U$1 ( \738 , \589 );
not \add_5_20_g13764/U$4 ( \739 , \738 );
or \add_5_20_g13764/U$2 ( \740 , \737 , \739 );
nand \add_5_20_g14002/U$1 ( \741 , \c[21] , \d[21] );
nand \add_5_20_g13764/U$1 ( \742 , \740 , \741 );
and \g45855/U$2 ( \743 , \594 , \742 );
nand \add_5_20_g13913/U$1 ( \744 , \c[22] , \d[22] );
nor \add_5_20_g13830/U$1 ( \745 , \593 , \744 );
and \add_5_20_g13905/U$1 ( \746 , \c[23] , \d[23] );
nor \g45855/U$1 ( \747 , \743 , \745 , \746 );
nand \add_5_20_g14012/U$1 ( \748 , \734 , \747 );
and \add_5_20_g13657/U$2 ( \749 , \748 , \612 );
nand \add_5_20_g13968/U$1 ( \750 , \c[24] , \d[24] );
or \add_5_20_g13769/U$2 ( \751 , \607 , \750 );
nand \add_5_20_g13875/U$1 ( \752 , \c[25] , \d[25] );
nand \add_5_20_g13769/U$1 ( \753 , \751 , \752 );
not \add_5_20_g13710/U$3 ( \754 , \753 );
not \add_5_20_g13710/U$4 ( \755 , \606 );
or \add_5_20_g13710/U$2 ( \756 , \754 , \755 );
not \add_5_20_g13782/U$3 ( \757 , \604 );
nand \add_5_20_g13947/U$1 ( \758 , \c[26] , \d[26] );
not \add_5_20_g13782/U$4 ( \759 , \758 );
and \add_5_20_g13782/U$2 ( \760 , \757 , \759 );
and \add_5_20_g13874/U$1 ( \761 , \c[27] , \d[27] );
nor \add_5_20_g13782/U$1 ( \762 , \760 , \761 );
nand \add_5_20_g13710/U$1 ( \763 , \756 , \762 );
not \add_5_20_g13709/U$1 ( \764 , \763 );
or \add_5_20_g13679/U$2 ( \765 , \603 , \764 );
nand \add_5_20_g13934/U$1 ( \766 , \c[28] , \d[28] );
or \add_5_20_g13762/U$2 ( \767 , \600 , \766 );
nand \add_5_20_g13902/U$1 ( \768 , \c[29] , \d[29] );
nand \add_5_20_g13762/U$1 ( \769 , \767 , \768 );
not \add_5_20_g13761/U$1 ( \770 , \769 );
or \add_5_20_g13679/U$3 ( \771 , \598 , \770 );
nand \add_5_20_g13917/U$1 ( \772 , \c[30] , \d[30] );
nand \add_5_20_g13679/U$1 ( \773 , \765 , \771 , \772 );
nor \add_5_20_g13657/U$1 ( \774 , \749 , \773 );
nand \add_5_20_g13616/U$1 ( \775 , \717 , \774 );
not \add_5_20_g13867/U$3 ( \776 , \c[31] );
not \add_5_20_g13867/U$4 ( \777 , \d[31] );
and \add_5_20_g13867/U$2 ( \778 , \776 , \777 );
and \add_5_20_g13867/U$5 ( \779 , \c[31] , \d[31] );
nor \add_5_20_g13867/U$1 ( \780 , \778 , \779 );
xor \add_5_20_g14033/U$1 ( \781 , \775 , \780 );
and \g2878/U$3 ( \782 , \581 , \781 );
nor \g2878/U$1 ( \783 , \580 , \782 );
not \g2965/U$1 ( \784 , \243 );
not \g2964/U$1 ( \785 , \784 );
not \g2960/U$1 ( \786 , \291 );
not \g2959/U$1 ( \787 , \786 );
nand \g2956/U$1 ( \788 , \785 , \787 );
nand \g2957/U$1 ( \789 , \786 , \784 );
xor \g3027/U$1 ( \790 , \a[11] , \a[5] );
xor \g45561/U$1 ( \791 , \a[24] , \a[17] );
xnor \g2996/U$1 ( \792 , \790 , \791 );
not \g2978/U$3 ( \793 , \792 );
xor \g3023/U$1 ( \794 , \a[29] , \a[3] );
xor \g3014/U$1 ( \795 , \a[27] , \a[15] );
xor \g45559/U$1 ( \796 , \794 , \795 );
not \g2978/U$4 ( \797 , \796 );
or \g2978/U$2 ( \798 , \793 , \797 );
or \g2978/U$5 ( \799 , \792 , \796 );
nand \g2978/U$1 ( \800 , \798 , \799 );
not \g2968/U$3 ( \801 , \800 );
xor \g3032/U$1 ( \802 , \a[28] , \a[7] );
xor \g3034/U$1 ( \803 , \a[25] , \a[8] );
xor \g45545/U$1 ( \804 , \802 , \803 );
xor \g45713/U$1 ( \805 , \a[21] , \a[9] );
xnor \g2/U$1 ( \806 , \a[23] , \a[18] );
xnor \g45713/U$1_r1 ( \807 , \805 , \806 );
xnor \g3094/U$1 ( \808 , \804 , \807 );
not \g2968/U$4 ( \809 , \808 );
or \g2968/U$2 ( \810 , \801 , \809 );
or \g2968/U$5 ( \811 , \808 , \800 );
nand \g2968/U$1 ( \812 , \810 , \811 );
not \g2967/U$1 ( \813 , \812 );
xor \g45565/U$1 ( \814 , \a[22] , \a[4] );
xor \g3012/U$1 ( \815 , \a[12] , \a[6] );
xor \g45714/U$1 ( \816 , \814 , \815 );
xor \g45712/U$1 ( \817 , \a[26] , \a[16] );
xnor \g3097/U$1 ( \818 , \a[20] , \a[19] );
xnor \g45712/U$1_r1 ( \819 , \817 , \818 );
xnor \g45714/U$1_r1 ( \820 , \816 , \819 );
not \g2963/U$3 ( \821 , \820 );
xor \g3007/U$1 ( \822 , \a[30] , \a[1] );
xor \g3009/U$1 ( \823 , \a[10] , \a[2] );
xor \g2985/U$1 ( \824 , \822 , \823 );
xor \g45711/U$1 ( \825 , \a[31] , \a[0] );
xnor \g3080/U$1 ( \826 , \a[14] , \a[13] );
xnor \g45711/U$1_r1 ( \827 , \825 , \826 );
xor \g45543/U$1 ( \828 , \824 , \827 );
not \g2963/U$4 ( \829 , \828 );
and \g2963/U$2 ( \830 , \821 , \829 );
and \g2963/U$5 ( \831 , \820 , \828 );
nor \g2963/U$1 ( \832 , \830 , \831 );
not \g2962/U$1 ( \833 , \832 );
nand \g2955/U$1 ( \834 , \813 , \833 );
nand \g2958/U$1 ( \835 , \832 , \812 );
nand \g2865/U$1 ( \836 , \788 , \789 , \834 , \835 );
buf \fopt45604/U$1 ( \837 , \836 );
buf \fopt45603/U$1 ( \838 , \837 );
buf \fopt45602/U$1 ( \839 , \838 );
nand \g2804/U$1 ( \840 , \783 , \839 );
not \sub_5_33_g9319/U$2 ( \841 , \574 );
nand \sub_5_33_g9319/U$1 ( \842 , \841 , \334 );
not \sub_5_33_g9078/U$3 ( \843 , \842 );
nor \sub_5_33_g9217/U$1 ( \844 , \348 , \331 );
and \sub_5_33_g9176/U$1 ( \845 , \326 , \844 );
not \sub_5_33_g9087/U$3 ( \846 , \845 );
not \sub_5_33_g9087/U$4 ( \847 , \490 );
or \sub_5_33_g9087/U$2 ( \848 , \846 , \847 );
and \sub_5_33_g9135/U$2 ( \849 , \541 , \844 );
or \sub_5_33_g9156/U$2 ( \850 , \564 , \331 );
not \sub_5_33_g9242/U$1 ( \851 , \571 );
nand \sub_5_33_g9156/U$1 ( \852 , \850 , \851 );
nor \sub_5_33_g9135/U$1 ( \853 , \849 , \852 );
nand \sub_5_33_g9087/U$1 ( \854 , \848 , \853 );
not \sub_5_33_g9078/U$4 ( \855 , \854 );
or \sub_5_33_g9078/U$2 ( \856 , \843 , \855 );
or \sub_5_33_g9078/U$5 ( \857 , \854 , \842 );
nand \sub_5_33_g9078/U$1 ( \858 , \856 , \857 );
and \g2866/U$2 ( \859 , \298 , \858 );
and \add_5_20_g13728/U$1 ( \860 , \610 , \602 );
not \add_5_20_g13693/U$2 ( \861 , \860 );
nor \add_5_20_g13693/U$1 ( \862 , \861 , \596 );
not \add_5_20_g13629/U$3 ( \863 , \862 );
not \add_5_20_g13629/U$4 ( \864 , \715 );
or \add_5_20_g13629/U$2 ( \865 , \863 , \864 );
and \g45715/U$2 ( \866 , \763 , \602 );
and \g45715/U$3 ( \867 , \748 , \860 );
nor \g45715/U$1 ( \868 , \866 , \867 , \769 );
nand \add_5_20_g13629/U$1 ( \869 , \865 , \868 );
not \add_5_20_g13848/U$2 ( \870 , \598 );
nand \add_5_20_g13848/U$1 ( \871 , \870 , \772 );
xnor \add_5_20_g14030/U$1 ( \872 , \869 , \871 );
and \g2866/U$3 ( \873 , \872 , \297 );
nor \g2866/U$1 ( \874 , \859 , \873 );
nand \g2805/U$1 ( \875 , \874 , \839 );
nand \sub_5_33_g9327/U$1 ( \876 , \330 , \570 );
nand \sub_5_33_g9219/U$1 ( \877 , \347 , \328 );
nor \sub_5_33_g9177/U$1 ( \878 , \325 , \877 );
not \sub_5_33_g9088/U$3 ( \879 , \878 );
not \sub_5_33_g9088/U$4 ( \880 , \490 );
or \sub_5_33_g9088/U$2 ( \881 , \879 , \880 );
not \sub_5_33_g9218/U$1 ( \882 , \877 );
not \sub_5_33_g9137/U$3 ( \883 , \882 );
not \sub_5_33_g9137/U$4 ( \884 , \541 );
or \sub_5_33_g9137/U$2 ( \885 , \883 , \884 );
not \sub_5_33_g9158/U$3 ( \886 , \328 );
not \sub_5_33_g9158/U$4 ( \887 , \563 );
or \sub_5_33_g9158/U$2 ( \888 , \886 , \887 );
nand \sub_5_33_g9158/U$1 ( \889 , \888 , \567 );
not \sub_5_33_g9157/U$1 ( \890 , \889 );
nand \sub_5_33_g9137/U$1 ( \891 , \885 , \890 );
not \sub_5_33_g9136/U$1 ( \892 , \891 );
nand \sub_5_33_g9088/U$1 ( \893 , \881 , \892 );
xnor \g45535/U$1 ( \894 , \876 , \893 );
and \g2867/U$2 ( \895 , \894 , \298 );
not \add_5_20_g13927/U$1 ( \896 , \601 );
nand \add_5_20_g13730/U$1 ( \897 , \610 , \896 );
nor \add_5_20_g13690/U$1 ( \898 , \596 , \897 );
not \add_5_20_g13614/U$3 ( \899 , \898 );
not \add_5_20_g13614/U$4 ( \900 , \715 );
or \add_5_20_g13614/U$2 ( \901 , \899 , \900 );
not \add_5_20_g13729/U$1 ( \902 , \897 );
and \add_5_20_g13659/U$2 ( \903 , \748 , \902 );
or \add_5_20_g13672/U$2 ( \904 , \764 , \601 );
nand \add_5_20_g13672/U$1 ( \905 , \904 , \766 );
nor \add_5_20_g13659/U$1 ( \906 , \903 , \905 );
nand \add_5_20_g13614/U$1 ( \907 , \901 , \906 );
not \add_5_20_g13854/U$2 ( \908 , \768 );
nor \add_5_20_g13854/U$1 ( \909 , \908 , \600 );
xor \add_5_20_g14031/U$1 ( \910 , \907 , \909 );
and \g2867/U$3 ( \911 , \910 , \296 );
nor \g2867/U$1 ( \912 , \895 , \911 );
nand \g2806/U$1 ( \913 , \912 , \839 );
nor \add_5_20_g13692/U$1 ( \914 , \596 , \611 );
not \add_5_20_g13625/U$3 ( \915 , \914 );
not \add_5_20_g13625/U$4 ( \916 , \715 );
or \add_5_20_g13625/U$2 ( \917 , \915 , \916 );
not \add_5_20_g13655/U$3 ( \918 , \610 );
not \add_5_20_g13655/U$4 ( \919 , \748 );
or \add_5_20_g13655/U$2 ( \920 , \918 , \919 );
nand \add_5_20_g13655/U$1 ( \921 , \920 , \764 );
not \add_5_20_g13654/U$1 ( \922 , \921 );
nand \add_5_20_g13625/U$1 ( \923 , \917 , \922 );
nand \add_5_20_g13859/U$1 ( \924 , \896 , \766 );
xnor \add_5_20_g14032/U$1 ( \925 , \923 , \924 );
and \g2868/U$2 ( \926 , \297 , \925 );
not \g2868/U$4 ( \927 , \297 );
nor \sub_5_33_g9171/U$1 ( \928 , \325 , \348 );
not \sub_5_33_g9099/U$3 ( \929 , \928 );
not \sub_5_33_g9099/U$4 ( \930 , \490 );
or \sub_5_33_g9099/U$2 ( \931 , \929 , \930 );
not \sub_5_33_g9132/U$3 ( \932 , \347 );
not \sub_5_33_g9132/U$4 ( \933 , \541 );
or \sub_5_33_g9132/U$2 ( \934 , \932 , \933 );
nand \sub_5_33_g9132/U$1 ( \935 , \934 , \564 );
not \sub_5_33_g9131/U$1 ( \936 , \935 );
nand \sub_5_33_g9099/U$1 ( \937 , \931 , \936 );
nand \sub_5_33_g9286/U$1 ( \938 , \328 , \567 );
xnor \sub_5_33_g9538/U$1 ( \939 , \937 , \938 );
and \g2868/U$3 ( \940 , \927 , \939 );
nor \g2868/U$1 ( \941 , \926 , \940 );
nand \g2807/U$1 ( \942 , \941 , \839 );
nand \sub_5_33_g9280/U$1 ( \943 , \337 , \560 );
not \sub_5_33_g9064/U$3 ( \944 , \943 );
not \sub_5_33_g9283/U$1 ( \945 , \346 );
and \sub_5_33_g9221/U$1 ( \946 , \945 , \339 );
not \sub_5_33_g9532/U$2 ( \947 , \946 );
nor \sub_5_33_g9532/U$1 ( \948 , \947 , \325 );
not \sub_5_33_g9085/U$3 ( \949 , \948 );
not \sub_5_33_g9085/U$4 ( \950 , \489 );
or \sub_5_33_g9085/U$2 ( \951 , \949 , \950 );
and \g45709/U$2 ( \952 , \946 , \541 );
and \g45709/U$3 ( \953 , \550 , \339 );
nor \g45709/U$1 ( \954 , \952 , \953 , \555 );
nand \sub_5_33_g9085/U$1 ( \955 , \951 , \954 );
not \sub_5_33_g9064/U$4 ( \956 , \955 );
or \sub_5_33_g9064/U$2 ( \957 , \944 , \956 );
or \sub_5_33_g9064/U$5 ( \958 , \955 , \943 );
nand \sub_5_33_g9064/U$1 ( \959 , \957 , \958 );
not \g2923/U$1 ( \960 , \296 );
and \g2869/U$2 ( \961 , \959 , \960 );
not \add_5_20_g13929/U$1 ( \962 , \605 );
nand \add_5_20_g13739/U$1 ( \963 , \609 , \962 );
nor \add_5_20_g13694/U$1 ( \964 , \596 , \963 );
not \add_5_20_g13624/U$3 ( \965 , \964 );
not \add_5_20_g13624/U$4 ( \966 , \715 );
or \add_5_20_g13624/U$2 ( \967 , \965 , \966 );
not \add_5_20_g13738/U$1 ( \968 , \963 );
and \add_5_20_g13660/U$2 ( \969 , \748 , \968 );
not \add_5_20_g13697/U$3 ( \970 , \962 );
not \add_5_20_g13697/U$4 ( \971 , \753 );
or \add_5_20_g13697/U$2 ( \972 , \970 , \971 );
nand \add_5_20_g13697/U$1 ( \973 , \972 , \758 );
nor \add_5_20_g13660/U$1 ( \974 , \969 , \973 );
nand \add_5_20_g13624/U$1 ( \975 , \967 , \974 );
nor \add_5_20_g13791/U$1 ( \976 , \604 , \761 );
xor \add_5_20_g14016/U$1 ( \977 , \975 , \976 );
and \g2869/U$3 ( \978 , \297 , \977 );
nor \g2869/U$1 ( \979 , \961 , \978 );
nand \g2808/U$1 ( \980 , \979 , \839 );
buf \g2952/U$1 ( \981 , \292 );
not \g2950/U$1 ( \982 , \981 );
buf \g2943/U$1 ( \983 , \982 );
nor \add_5_20_g13689/U$1 ( \984 , \596 , \608 );
not \add_5_20_g13619/U$3 ( \985 , \984 );
not \add_5_20_g13619/U$4 ( \986 , \715 );
or \add_5_20_g13619/U$2 ( \987 , \985 , \986 );
not \add_5_20_g13870/U$1 ( \988 , \608 );
and \add_5_20_g13653/U$2 ( \989 , \748 , \988 );
not \add_5_20_g13967/U$1 ( \990 , \750 );
nor \add_5_20_g13653/U$1 ( \991 , \989 , \990 );
nand \add_5_20_g13619/U$1 ( \992 , \987 , \991 );
not \add_5_20_g13803/U$2 ( \993 , \752 );
nor \add_5_20_g13803/U$1 ( \994 , \993 , \607 );
xor \add_5_20_g14019/U$1 ( \995 , \992 , \994 );
and \g2872/U$2 ( \996 , \983 , \995 );
not \g2872/U$4 ( \997 , \983 );
not \sub_5_33_g9553/U$2 ( \998 , \345 );
nor \sub_5_33_g9553/U$1 ( \999 , \998 , \325 );
not \sub_5_33_g9091/U$3 ( \1000 , \999 );
not \sub_5_33_g9091/U$4 ( \1001 , \490 );
or \sub_5_33_g9091/U$2 ( \1002 , \1000 , \1001 );
not \sub_5_33_g9129/U$3 ( \1003 , \345 );
not \sub_5_33_g9129/U$4 ( \1004 , \541 );
or \sub_5_33_g9129/U$2 ( \1005 , \1003 , \1004 );
not \sub_5_33_g9450/U$1 ( \1006 , \545 );
nand \sub_5_33_g9129/U$1 ( \1007 , \1005 , \1006 );
not \sub_5_33_g9128/U$1 ( \1008 , \1007 );
nand \sub_5_33_g9091/U$1 ( \1009 , \1002 , \1008 );
nand \sub_5_33_g9291/U$1 ( \1010 , \343 , \549 );
not \sub_5_33_g9597/U$2 ( \1011 , \1010 );
xor \sub_5_33_g9597/U$1 ( \1012 , \1009 , \1011 );
and \g2872/U$3 ( \1013 , \997 , \1012 );
nor \g2872/U$1 ( \1014 , \996 , \1013 );
nand \g2810/U$1 ( \1015 , \1014 , \839 );
not \add_5_20_g13746/U$1 ( \1016 , \588 );
not \add_5_20_g13884/U$1 ( \1017 , \590 );
and \add_5_20_g13826/U$1 ( \1018 , \738 , \1017 );
not \add_5_20_g13990/U$1 ( \1019 , \592 );
nand \add_5_20_g13742/U$1 ( \1020 , \1018 , \1019 );
nor \add_5_20_g13734/U$1 ( \1021 , \1016 , \1020 );
not \add_5_20_g13621/U$3 ( \1022 , \1021 );
not \add_5_20_g13621/U$4 ( \1023 , \715 );
or \add_5_20_g13621/U$2 ( \1024 , \1022 , \1023 );
not \add_5_20_g13741/U$1 ( \1025 , \1020 );
and \add_5_20_g13681/U$2 ( \1026 , \732 , \1025 );
not \add_5_20_g13698/U$3 ( \1027 , \1019 );
not \add_5_20_g13698/U$4 ( \1028 , \742 );
or \add_5_20_g13698/U$2 ( \1029 , \1027 , \1028 );
nand \add_5_20_g13698/U$1 ( \1030 , \1029 , \744 );
nor \add_5_20_g13681/U$1 ( \1031 , \1026 , \1030 );
nand \add_5_20_g13621/U$1 ( \1032 , \1024 , \1031 );
nor \add_5_20_g13814/U$1 ( \1033 , \746 , \593 );
xor \add_5_20_g14022/U$1 ( \1034 , \1032 , \1033 );
and \g2873/U$2 ( \1035 , \983 , \1034 );
not \g2873/U$4 ( \1036 , \983 );
not \sub_5_33_g9385/U$1 ( \1037 , \322 );
nor \sub_5_33_g9224/U$1 ( \1038 , \318 , \1037 );
not \sub_5_33_g9533/U$2 ( \1039 , \1038 );
not \sub_5_33_g9350/U$1 ( \1040 , \310 );
nand \sub_5_33_g9241/U$1 ( \1041 , \304 , \1040 );
nor \sub_5_33_g9533/U$1 ( \1042 , \1039 , \1041 );
not \sub_5_33_g9086/U$3 ( \1043 , \1042 );
not \sub_5_33_g9086/U$4 ( \1044 , \489 );
or \sub_5_33_g9086/U$2 ( \1045 , \1043 , \1044 );
and \g45710/U$2 ( \1046 , \1038 , \514 );
and \g45710/U$3 ( \1047 , \527 , \322 );
nor \g45710/U$1 ( \1048 , \1046 , \1047 , \532 );
nand \sub_5_33_g9086/U$1 ( \1049 , \1045 , \1048 );
nand \sub_5_33_g9302/U$1 ( \1050 , \320 , \536 );
xnor \sub_5_33_g45888/U$1 ( \1051 , \1049 , \1050 );
and \g2873/U$3 ( \1052 , \1036 , \1051 );
nor \g2873/U$1 ( \1053 , \1035 , \1052 );
not \fopt45597/U$1 ( \1054 , \837 );
not \fopt45593/U$1 ( \1055 , \1054 );
nand \g2812/U$1 ( \1056 , \1053 , \1055 );
not \add_5_20_g14025/U$2 ( \1057 , \1018 );
nor \add_5_20_g14025/U$1 ( \1058 , \1057 , \1016 );
not \add_5_20_g13622/U$3 ( \1059 , \1058 );
not \add_5_20_g13622/U$4 ( \1060 , \715 );
or \add_5_20_g13622/U$2 ( \1061 , \1059 , \1060 );
and \add_5_20_g13667/U$2 ( \1062 , \732 , \1018 );
nor \add_5_20_g13667/U$1 ( \1063 , \1062 , \742 );
nand \add_5_20_g13622/U$1 ( \1064 , \1061 , \1063 );
nand \add_5_20_g13818/U$1 ( \1065 , \1019 , \744 );
xnor \add_5_20_g45815/U$1 ( \1066 , \1064 , \1065 );
and \g2874/U$2 ( \1067 , \983 , \1066 );
not \g2874/U$4 ( \1068 , \983 );
nor \sub_5_33_g9210/U$1 ( \1069 , \1041 , \318 );
not \sub_5_33_g9092/U$3 ( \1070 , \1069 );
not \sub_5_33_g9092/U$4 ( \1071 , \489 );
or \sub_5_33_g9092/U$2 ( \1072 , \1070 , \1071 );
not \sub_5_33_g9543/U$2 ( \1073 , \318 );
nand \sub_5_33_g9543/U$1 ( \1074 , \1073 , \514 );
not \sub_5_33_g9524/U$2 ( \1075 , \1074 );
nor \sub_5_33_g9524/U$1 ( \1076 , \1075 , \527 );
nand \sub_5_33_g9092/U$1 ( \1077 , \1072 , \1076 );
nor \sub_5_33_g9353/U$1 ( \1078 , \1037 , \532 );
xor \sub_5_33_g9550/U$1 ( \1079 , \1077 , \1078 );
and \g2874/U$3 ( \1080 , \1068 , \1079 );
nor \g2874/U$1 ( \1081 , \1067 , \1080 );
nand \g2813/U$1 ( \1082 , \1081 , \838 );
not \g2930/U$1 ( \1083 , \295 );
not \sub_5_33_g9554/U$2 ( \1084 , \317 );
nor \sub_5_33_g9554/U$1 ( \1085 , \1084 , \1041 );
not \sub_5_33_g9093/U$3 ( \1086 , \1085 );
not \sub_5_33_g9093/U$4 ( \1087 , \489 );
or \sub_5_33_g9093/U$2 ( \1088 , \1086 , \1087 );
nand \sub_5_33_g9164/U$1 ( \1089 , \514 , \317 );
not \sub_5_33_g9475/U$1 ( \1090 , \520 );
and \sub_5_33_g9525/U$1 ( \1091 , \1089 , \1090 );
nand \sub_5_33_g9093/U$1 ( \1092 , \1088 , \1091 );
nand \sub_5_33_g9305/U$1 ( \1093 , \522 , \526 );
xnor \sub_5_33_g45816/U$1 ( \1094 , \1092 , \1093 );
nand \g2884/U$1 ( \1095 , \1083 , \1094 );
nor \add_5_20_g13721/U$1 ( \1096 , \1016 , \590 );
not \add_5_20_g13615/U$3 ( \1097 , \1096 );
not \add_5_20_g13615/U$4 ( \1098 , \715 );
or \add_5_20_g13615/U$2 ( \1099 , \1097 , \1098 );
not \add_5_20_g13670/U$3 ( \1100 , \1017 );
not \add_5_20_g13670/U$4 ( \1101 , \732 );
or \add_5_20_g13670/U$2 ( \1102 , \1100 , \1101 );
nand \add_5_20_g13670/U$1 ( \1103 , \1102 , \735 );
not \add_5_20_g13669/U$1 ( \1104 , \1103 );
nand \add_5_20_g13615/U$1 ( \1105 , \1099 , \1104 );
nand \add_5_20_g13842/U$1 ( \1106 , \738 , \741 );
xnor \add_5_20_g14028/U$1 ( \1107 , \1105 , \1106 );
nand \g2883/U$1 ( \1108 , \296 , \1107 );
nand \g2814/U$1 ( \1109 , \1095 , \838 , \1108 );
not \g45325/U$2 ( \1110 , \983 );
nand \sub_5_33_g9310/U$1 ( \1111 , \317 , \1090 );
not \sub_5_33_g9101/U$3 ( \1112 , \311 );
not \sub_5_33_g9101/U$4 ( \1113 , \489 );
or \sub_5_33_g9101/U$2 ( \1114 , \1112 , \1113 );
not \sub_5_33_g9190/U$1 ( \1115 , \514 );
nand \sub_5_33_g9101/U$1 ( \1116 , \1114 , \1115 );
xnor \g45326/U$1 ( \1117 , \1111 , \1116 );
nand \g45325/U$1 ( \1118 , \1110 , \1117 );
nand \add_5_20_g13804/U$1 ( \1119 , \1017 , \735 );
not \add_5_20_g13627/U$3 ( \1120 , \588 );
not \add_5_20_g13627/U$4 ( \1121 , \715 );
or \add_5_20_g13627/U$2 ( \1122 , \1120 , \1121 );
not \add_5_20_g13700/U$1 ( \1123 , \732 );
nand \add_5_20_g13627/U$1 ( \1124 , \1122 , \1123 );
xnor \g45327/U$1 ( \1125 , \1119 , \1124 );
nand \g2885/U$1 ( \1126 , \296 , \1125 );
nand \g2815/U$1 ( \1127 , \1118 , \1126 , \1055 );
nand \sub_5_33_g9315/U$1 ( \1128 , \301 , \511 );
not \sub_5_33_g9229/U$2 ( \1129 , \303 );
nor \sub_5_33_g9229/U$1 ( \1130 , \1129 , \310 );
not \sub_5_33_g9094/U$3 ( \1131 , \1130 );
not \sub_5_33_g9094/U$4 ( \1132 , \489 );
or \sub_5_33_g9094/U$2 ( \1133 , \1131 , \1132 );
not \sub_5_33_g9181/U$3 ( \1134 , \303 );
not \sub_5_33_g9181/U$4 ( \1135 , \501 );
or \sub_5_33_g9181/U$2 ( \1136 , \1134 , \1135 );
not \sub_5_33_g9457/U$1 ( \1137 , \506 );
nand \sub_5_33_g9181/U$1 ( \1138 , \1136 , \1137 );
not \sub_5_33_g9180/U$1 ( \1139 , \1138 );
nand \sub_5_33_g9094/U$1 ( \1140 , \1133 , \1139 );
xnor \g45533/U$1 ( \1141 , \1128 , \1140 );
nand \g2888/U$1 ( \1142 , \1083 , \1141 );
or \add_5_20_g13789/U$1 ( \1143 , \582 , \730 );
not \add_5_20_g13597/U$3 ( \1144 , \1143 );
not \add_5_20_g13969/U$1 ( \1145 , \583 );
and \add_5_20_g13745/U$1 ( \1146 , \587 , \1145 );
not \add_5_20_g13628/U$3 ( \1147 , \1146 );
not \add_5_20_g13628/U$4 ( \1148 , \715 );
or \add_5_20_g13628/U$2 ( \1149 , \1147 , \1148 );
and \add_5_20_g13703/U$2 ( \1150 , \722 , \1145 );
not \add_5_20_g13908/U$1 ( \1151 , \727 );
nor \add_5_20_g13703/U$1 ( \1152 , \1150 , \1151 );
nand \add_5_20_g13628/U$1 ( \1153 , \1149 , \1152 );
not \add_5_20_g13597/U$4 ( \1154 , \1153 );
or \add_5_20_g13597/U$2 ( \1155 , \1144 , \1154 );
or \add_5_20_g13597/U$5 ( \1156 , \1153 , \1143 );
nand \add_5_20_g13597/U$1 ( \1157 , \1155 , \1156 );
nand \g2887/U$1 ( \1158 , \983 , \1157 );
nand \g2817/U$1 ( \1159 , \1142 , \1158 , \838 );
buf \g2816/U$1 ( \1160 , \1159 );
not \add_5_20_g13612/U$3 ( \1161 , \587 );
not \add_5_20_g13612/U$4 ( \1162 , \715 );
or \add_5_20_g13612/U$2 ( \1163 , \1161 , \1162 );
not \add_5_20_g13776/U$1 ( \1164 , \722 );
nand \add_5_20_g13612/U$1 ( \1165 , \1163 , \1164 );
nand \add_5_20_g13796/U$1 ( \1166 , \1145 , \727 );
not \add_5_20_g13795/U$1 ( \1167 , \1166 );
and \add_5_20_g13598/U$2 ( \1168 , \1165 , \1167 );
not \add_5_20_g13598/U$4 ( \1169 , \1165 );
and \add_5_20_g13598/U$3 ( \1170 , \1169 , \1166 );
nor \add_5_20_g13598/U$1 ( \1171 , \1168 , \1170 );
and \g2875/U$2 ( \1172 , \295 , \1171 );
not \g2875/U$4 ( \1173 , \295 );
not \sub_5_33_g9102/U$3 ( \1174 , \1040 );
nand \sub_5_33_g9120/U$1 ( \1175 , \488 , \463 , \434 , \377 );
not \sub_5_33_g9102/U$4 ( \1176 , \1175 );
or \sub_5_33_g9102/U$2 ( \1177 , \1174 , \1176 );
not \sub_5_33_g9261/U$1 ( \1178 , \501 );
nand \sub_5_33_g9102/U$1 ( \1179 , \1177 , \1178 );
nand \sub_5_33_g9336/U$1 ( \1180 , \303 , \1137 );
xnor \sub_5_33_g9548/U$1 ( \1181 , \1179 , \1180 );
and \g2875/U$3 ( \1182 , \1173 , \1181 );
nor \g2875/U$1 ( \1183 , \1172 , \1182 );
nand \g2818/U$1 ( \1184 , \1183 , \838 );
not \add_5_20_g13898/U$1 ( \1185 , \586 );
not \add_5_20_g13610/U$3 ( \1186 , \1185 );
not \add_5_20_g13706/U$1 ( \1187 , \689 );
not \add_5_20_g13661/U$3 ( \1188 , \1187 );
and \add_5_20_g13750/U$1 ( \1189 , \679 , \646 );
nand \add_5_20_g13682/U$1 ( \1190 , \709 , \1189 );
not \add_5_20_g13661/U$4 ( \1191 , \1190 );
or \add_5_20_g13661/U$2 ( \1192 , \1188 , \1191 );
nand \add_5_20_g13661/U$1 ( \1193 , \1192 , \692 );
nand \add_5_20_g13637/U$1 ( \1194 , \1193 , \658 , \673 );
not \add_5_20_g13610/U$4 ( \1195 , \1194 );
or \add_5_20_g13610/U$2 ( \1196 , \1186 , \1195 );
nand \add_5_20_g13610/U$1 ( \1197 , \1196 , \719 );
not \add_5_20_g13832/U$2 ( \1198 , \585 );
nand \add_5_20_g13832/U$1 ( \1199 , \1198 , \721 );
xnor \add_5_20_g13588/U$1 ( \1200 , \1197 , \1199 );
not \g2876/U$3 ( \1201 , \1200 );
buf \g2938/U$1 ( \1202 , \293 );
not \g2937/U$1 ( \1203 , \1202 );
not \g2876/U$4 ( \1204 , \1203 );
or \g2876/U$2 ( \1205 , \1201 , \1204 );
not \g2940/U$1 ( \1206 , \981 );
buf \g2945/U$1 ( \1207 , \1206 );
not \sub_5_33_g9103/U$3 ( \1208 , \309 );
not \sub_5_33_g9103/U$4 ( \1209 , \1175 );
or \sub_5_33_g9103/U$2 ( \1210 , \1208 , \1209 );
not \sub_5_33_g9359/U$1 ( \1211 , \496 );
nand \sub_5_33_g9103/U$1 ( \1212 , \1210 , \1211 );
nand \sub_5_33_g9321/U$1 ( \1213 , \307 , \500 );
xor \g45655/U$1 ( \1214 , \1212 , \1213 );
or \g2876/U$5 ( \1215 , \1207 , \1214 );
nand \g2876/U$1 ( \1216 , \1205 , \1215 );
nor \g2820/U$1 ( \1217 , \1216 , \1054 );
not \g2819/U$1 ( \1218 , \1217 );
nand \sub_5_33_g9322/U$1 ( \1219 , \309 , \1211 );
xnor \g45304/U$1 ( \1220 , \1219 , \489 );
nand \g45303/U$1 ( \1221 , \1083 , \1220 );
nand \add_5_20_g13834/U$1 ( \1222 , \1185 , \719 );
not \add_5_20_g13632/U$3 ( \1223 , \1222 );
not \add_5_20_g13632/U$4 ( \1224 , \715 );
or \add_5_20_g13632/U$2 ( \1225 , \1223 , \1224 );
or \add_5_20_g13632/U$5 ( \1226 , \715 , \1222 );
nand \add_5_20_g13632/U$1 ( \1227 , \1225 , \1226 );
nand \g2889/U$1 ( \1228 , \1227 , \295 );
nand \g2821/U$1 ( \1229 , \1221 , \1228 , \838 );
not \g2917/U$1 ( \1230 , \294 );
not \sub_5_33_g9551/U$2 ( \1231 , \374 );
nand \sub_5_33_g9551/U$1 ( \1232 , \1231 , \353 );
not \sub_5_33_g9075/U$3 ( \1233 , \1232 );
not \sub_5_33_g9234/U$2 ( \1234 , \437 );
nand \sub_5_33_g9234/U$1 ( \1235 , \1234 , \355 );
nor \sub_5_33_g9212/U$1 ( \1236 , \464 , \1235 );
not \sub_5_33_g9095/U$3 ( \1237 , \1236 );
not \sub_5_33_g9537/U$2 ( \1238 , \475 );
nor \sub_5_33_g9537/U$1 ( \1239 , \1238 , \392 );
not \sub_5_33_g9522/U$3 ( \1240 , \1239 );
not \sub_5_33_g9522/U$4 ( \1241 , \433 );
or \sub_5_33_g9522/U$2 ( \1242 , \1240 , \1241 );
not \sub_5_33_g9199/U$1 ( \1243 , \487 );
nand \sub_5_33_g9522/U$1 ( \1244 , \1242 , \1243 );
buf \fopt45583/U$1 ( \1245 , \1244 );
not \sub_5_33_g9095/U$4 ( \1246 , \1245 );
or \sub_5_33_g9095/U$2 ( \1247 , \1237 , \1246 );
not \sub_5_33_g9233/U$1 ( \1248 , \1235 );
and \sub_5_33_g9162/U$2 ( \1249 , \462 , \1248 );
not \sub_5_33_g9265/U$1 ( \1250 , \367 );
not \sub_5_33_g9432/U$1 ( \1251 , \355 );
or \sub_5_33_g9184/U$2 ( \1252 , \1250 , \1251 );
not \sub_5_33_g9395/U$1 ( \1253 , \371 );
nand \sub_5_33_g9184/U$1 ( \1254 , \1252 , \1253 );
nor \sub_5_33_g9162/U$1 ( \1255 , \1249 , \1254 );
nand \sub_5_33_g9095/U$1 ( \1256 , \1247 , \1255 );
not \sub_5_33_g9075/U$4 ( \1257 , \1256 );
or \sub_5_33_g9075/U$2 ( \1258 , \1233 , \1257 );
or \sub_5_33_g9075/U$5 ( \1259 , \1256 , \1232 );
nand \sub_5_33_g9075/U$1 ( \1260 , \1258 , \1259 );
nand \g2892/U$1 ( \1261 , \1230 , \1260 );
not \g2936/U$1 ( \1262 , \293 );
buf \g2935/U$1 ( \1263 , \1262 );
nand \add_5_20_g13835/U$1 ( \1264 , \639 , \671 );
not \add_5_20_g13861/U$1 ( \1265 , \691 );
nand \add_5_20_g13758/U$1 ( \1266 , \1265 , \651 );
not \add_5_20_g13749/U$1 ( \1267 , \1189 );
nor \add_5_20_g13733/U$1 ( \1268 , \1266 , \1267 );
not \add_5_20_g13623/U$3 ( \1269 , \1268 );
not \g45297/U$1 ( \1270 , \615 );
and \add_5_20_g13737/U$1 ( \1271 , \699 , \1270 , \643 );
not \add_5_20_g14011/U$3 ( \1272 , \1271 );
not \add_5_20_g13945/U$1 ( \1273 , \616 );
not \add_5_20_g13665/U$3 ( \1274 , \1273 );
not \add_5_20_g13665/U$4 ( \1275 , \623 );
or \add_5_20_g13665/U$2 ( \1276 , \1274 , \1275 );
and \add_5_20_g13846/U$1 ( \1277 , \630 , \627 );
nand \add_5_20_g13665/U$1 ( \1278 , \1276 , \1277 );
not \add_5_20_g14011/U$4 ( \1279 , \1278 );
or \add_5_20_g14011/U$2 ( \1280 , \1272 , \1279 );
not \add_5_20_g13714/U$1 ( \1281 , \709 );
nand \add_5_20_g14011/U$1 ( \1282 , \1280 , \1281 );
not \add_5_20_g13623/U$4 ( \1283 , \1282 );
or \add_5_20_g13623/U$2 ( \1284 , \1269 , \1283 );
not \add_5_20_g13757/U$1 ( \1285 , \1266 );
and \add_5_20_g13680/U$2 ( \1286 , \689 , \1285 );
not \add_5_20_g13704/U$3 ( \1287 , \651 );
not \add_5_20_g13704/U$4 ( \1288 , \665 );
or \add_5_20_g13704/U$2 ( \1289 , \1287 , \1288 );
nand \add_5_20_g13704/U$1 ( \1290 , \1289 , \669 );
nor \add_5_20_g13680/U$1 ( \1291 , \1286 , \1290 );
nand \add_5_20_g13623/U$1 ( \1292 , \1284 , \1291 );
xnor \g45329/U$1 ( \1293 , \1264 , \1292 );
nand \g2891/U$1 ( \1294 , \1263 , \1293 );
not \fopt45590/U$1 ( \1295 , \837 );
not \fopt45589/U$1 ( \1296 , \1295 );
nand \g2823/U$1 ( \1297 , \1261 , \1294 , \1296 );
buf \g2822/U$1 ( \1298 , \1297 );
not \g45323/U$2 ( \1299 , \1263 );
nand \sub_5_33_g9292/U$1 ( \1300 , \355 , \1253 );
nor \sub_5_33_g9213/U$1 ( \1301 , \464 , \437 );
not \sub_5_33_g9096/U$3 ( \1302 , \1301 );
not \sub_5_33_g9096/U$4 ( \1303 , \1244 );
or \sub_5_33_g9096/U$2 ( \1304 , \1302 , \1303 );
nand \sub_5_33_g9166/U$1 ( \1305 , \462 , \438 );
and \sub_5_33_g9526/U$1 ( \1306 , \1305 , \1250 );
nand \sub_5_33_g9096/U$1 ( \1307 , \1304 , \1306 );
xnor \g45324/U$1 ( \1308 , \1300 , \1307 );
nand \g45323/U$1 ( \1309 , \1299 , \1308 );
not \g45319/U$2 ( \1310 , \1230 );
nand \add_5_20_g13821/U$1 ( \1311 , \651 , \669 );
nor \add_5_20_g13731/U$1 ( \1312 , \1267 , \691 );
not \add_5_20_g13617/U$3 ( \1313 , \1312 );
not \add_5_20_g13617/U$4 ( \1314 , \1282 );
or \add_5_20_g13617/U$2 ( \1315 , \1313 , \1314 );
and \add_5_20_g13668/U$2 ( \1316 , \689 , \1265 );
nor \add_5_20_g13668/U$1 ( \1317 , \1316 , \665 );
nand \add_5_20_g13617/U$1 ( \1318 , \1315 , \1317 );
xnor \g45320/U$1 ( \1319 , \1311 , \1318 );
nand \g45319/U$1 ( \1320 , \1310 , \1319 );
nand \g2824/U$1 ( \1321 , \1309 , \838 , \1320 );
not \add_5_20_g14036/U$2 ( \1322 , \655 );
nor \add_5_20_g14036/U$1 ( \1323 , \1322 , \1267 );
not \add_5_20_g13620/U$3 ( \1324 , \1323 );
not \add_5_20_g13620/U$4 ( \1325 , \1282 );
or \add_5_20_g13620/U$2 ( \1326 , \1324 , \1325 );
not \add_5_20_g13674/U$3 ( \1327 , \655 );
not \add_5_20_g13674/U$4 ( \1328 , \689 );
or \add_5_20_g13674/U$2 ( \1329 , \1327 , \1328 );
nand \add_5_20_g13674/U$1 ( \1330 , \1329 , \659 );
not \add_5_20_g13673/U$1 ( \1331 , \1330 );
nand \add_5_20_g13620/U$1 ( \1332 , \1326 , \1331 );
nand \add_5_20_g13840/U$1 ( \1333 , \638 , \664 );
xnor \add_5_20_g14027/U$1 ( \1334 , \1332 , \1333 );
and \g3095/U$1 ( \1335 , \1206 , \1334 );
not \g2825/U$2 ( \1336 , \1335 );
nand \sub_5_33_g9341/U$1 ( \1337 , \359 , \366 );
not \sub_5_33_g9077/U$3 ( \1338 , \1337 );
not \sub_5_33_g9556/U$2 ( \1339 , \436 );
nor \sub_5_33_g9556/U$1 ( \1340 , \1339 , \464 );
not \sub_5_33_g9097/U$3 ( \1341 , \1340 );
not \sub_5_33_g9097/U$4 ( \1342 , \1244 );
or \sub_5_33_g9097/U$2 ( \1343 , \1341 , \1342 );
nand \sub_5_33_g9167/U$1 ( \1344 , \462 , \436 );
not \sub_5_33_g9469/U$1 ( \1345 , \362 );
and \sub_5_33_g9527/U$1 ( \1346 , \1344 , \1345 );
nand \sub_5_33_g9097/U$1 ( \1347 , \1343 , \1346 );
not \sub_5_33_g9077/U$4 ( \1348 , \1347 );
or \sub_5_33_g9077/U$2 ( \1349 , \1338 , \1348 );
or \sub_5_33_g9077/U$5 ( \1350 , \1347 , \1337 );
nand \sub_5_33_g9077/U$1 ( \1351 , \1349 , \1350 );
nand \g2896/U$1 ( \1352 , \1230 , \1351 );
nand \g2825/U$1 ( \1353 , \1336 , \1352 , \1055 );
nand \sub_5_33_g9337/U$1 ( \1354 , \436 , \1345 );
not \sub_5_33_g9235/U$1 ( \1355 , \464 );
not \sub_5_33_g9104/U$3 ( \1356 , \1355 );
not \sub_5_33_g9104/U$4 ( \1357 , \1244 );
or \sub_5_33_g9104/U$2 ( \1358 , \1356 , \1357 );
not \sub_5_33_g9194/U$1 ( \1359 , \462 );
nand \sub_5_33_g9104/U$1 ( \1360 , \1358 , \1359 );
xnor \g45534/U$1 ( \1361 , \1354 , \1360 );
nand \g2898/U$1 ( \1362 , \1083 , \1361 );
nand \add_5_20_g13857/U$1 ( \1363 , \655 , \659 );
not \add_5_20_g13630/U$3 ( \1364 , \1189 );
not \add_5_20_g13630/U$4 ( \1365 , \1282 );
or \add_5_20_g13630/U$2 ( \1366 , \1364 , \1365 );
nand \add_5_20_g13630/U$1 ( \1367 , \1366 , \1187 );
xnor \g45328/U$1 ( \1368 , \1363 , \1367 );
nand \g2897/U$1 ( \1369 , \295 , \1368 );
nand \g2826/U$1 ( \1370 , \1362 , \1369 , \1055 );
nand \add_5_20_g13822/U$1 ( \1371 , \637 , \686 );
and \add_5_20_g13759/U$1 ( \1372 , \646 , \649 );
not \add_5_20_g13626/U$3 ( \1373 , \1372 );
not \add_5_20_g13626/U$4 ( \1374 , \1282 );
or \add_5_20_g13626/U$2 ( \1375 , \1373 , \1374 );
and \add_5_20_g13713/U$2 ( \1376 , \677 , \649 );
not \add_5_20_g13931/U$1 ( \1377 , \683 );
nor \add_5_20_g13713/U$1 ( \1378 , \1376 , \1377 );
nand \add_5_20_g13626/U$1 ( \1379 , \1375 , \1378 );
xnor \g45330/U$1 ( \1380 , \1371 , \1379 );
nand \g2899/U$1 ( \1381 , \1262 , \1380 );
not \g2877/U$2 ( \1382 , \1381 );
and \sub_5_33_g9539/U$1 ( \1383 , \387 , \402 );
not \sub_5_33_g9098/U$3 ( \1384 , \1383 );
not \sub_5_33_g9098/U$4 ( \1385 , \1244 );
or \sub_5_33_g9098/U$2 ( \1386 , \1384 , \1385 );
nand \sub_5_33_g9215/U$1 ( \1387 , \450 , \402 );
not \sub_5_33_g9428/U$1 ( \1388 , \455 );
and \sub_5_33_g9528/U$1 ( \1389 , \1387 , \1388 );
nand \sub_5_33_g9098/U$1 ( \1390 , \1386 , \1389 );
nand \sub_5_33_g9339/U$1 ( \1391 , \459 , \381 );
xnor \sub_5_33_g45814/U$1 ( \1392 , \1390 , \1391 );
not \g3098/U$2 ( \1393 , \1392 );
nor \g3098/U$1 ( \1394 , \1393 , \1206 );
nor \g2877/U$1 ( \1395 , \1382 , \1394 );
nand \g2827/U$1 ( \1396 , \1395 , \838 );
nand \add_5_20_g13852/U$1 ( \1397 , \649 , \683 );
not \add_5_20_g13613/U$3 ( \1398 , \1282 );
not \add_5_20_g13613/U$4 ( \1399 , \646 );
or \add_5_20_g13613/U$2 ( \1400 , \1398 , \1399 );
not \add_5_20_g13773/U$1 ( \1401 , \677 );
nand \add_5_20_g13613/U$1 ( \1402 , \1400 , \1401 );
xor \g45875/U$1 ( \1403 , \1397 , \1402 );
nor \g45874/U$1 ( \1404 , \1403 , \981 );
not \g2828/U$2 ( \1405 , \1404 );
not \g45321/U$2 ( \1406 , \294 );
nand \sub_5_33_g9318/U$1 ( \1407 , \1388 , \402 );
not \sub_5_33_g9105/U$3 ( \1408 , \387 );
not \sub_5_33_g9105/U$4 ( \1409 , \1244 );
or \sub_5_33_g9105/U$2 ( \1410 , \1408 , \1409 );
not \sub_5_33_g9258/U$1 ( \1411 , \450 );
nand \sub_5_33_g9105/U$1 ( \1412 , \1410 , \1411 );
xnor \g45322/U$1 ( \1413 , \1407 , \1412 );
nand \g45321/U$1 ( \1414 , \1406 , \1413 );
nand \g2828/U$1 ( \1415 , \1405 , \1414 , \1296 );
not \sub_5_33_g9403/U$1 ( \1416 , \444 );
nand \sub_5_33_g9343/U$1 ( \1417 , \1416 , \386 );
not \sub_5_33_g9111/U$3 ( \1418 , \1417 );
not \sub_5_33_g9111/U$4 ( \1419 , \1245 );
or \sub_5_33_g9111/U$2 ( \1420 , \1418 , \1419 );
or \sub_5_33_g9111/U$5 ( \1421 , \1245 , \1417 );
nand \sub_5_33_g9111/U$1 ( \1422 , \1420 , \1421 );
not \g3099/U$2 ( \1423 , \1422 );
nor \g3099/U$1 ( \1424 , \1423 , \294 );
not \g2830/U$2 ( \1425 , \1424 );
not \g45702/U$2 ( \1426 , \645 );
nand \g45702/U$1 ( \1427 , \1426 , \674 );
not \add_5_20_g13633/U$3 ( \1428 , \1427 );
not \add_5_20_g13633/U$4 ( \1429 , \1282 );
or \add_5_20_g13633/U$2 ( \1430 , \1428 , \1429 );
or \add_5_20_g13633/U$5 ( \1431 , \1282 , \1427 );
nand \add_5_20_g13633/U$1 ( \1432 , \1430 , \1431 );
nand \g2906/U$1 ( \1433 , \982 , \1432 );
nand \g2830/U$1 ( \1434 , \1425 , \1433 , \837 );
nand \sub_5_33_g9326/U$1 ( \1435 , \379 , \484 );
not \sub_5_33_g9555/U$2 ( \1436 , \397 );
nor \sub_5_33_g9555/U$1 ( \1437 , \1436 , \392 );
not \sub_5_33_g9114/U$3 ( \1438 , \1437 );
not \sub_5_33_g9114/U$4 ( \1439 , \433 );
or \sub_5_33_g9114/U$2 ( \1440 , \1438 , \1439 );
and \sub_5_33_g9183/U$2 ( \1441 , \473 , \397 );
nor \sub_5_33_g9183/U$1 ( \1442 , \1441 , \479 );
nand \sub_5_33_g9114/U$1 ( \1443 , \1440 , \1442 );
xnor \g45536/U$1 ( \1444 , \1435 , \1443 );
nand \g2908/U$1 ( \1445 , \1444 , \981 );
nand \add_5_20_g13827/U$1 ( \1446 , \635 , \706 );
and \add_5_20_g13756/U$1 ( \1447 , \643 , \653 );
not \add_5_20_g13649/U$3 ( \1448 , \1447 );
not \add_5_20_g13649/U$4 ( \1449 , \633 );
or \add_5_20_g13649/U$2 ( \1450 , \1448 , \1449 );
and \add_5_20_g13716/U$2 ( \1451 , \697 , \653 );
not \add_5_20_g13951/U$1 ( \1452 , \703 );
nor \add_5_20_g13716/U$1 ( \1453 , \1451 , \1452 );
nand \add_5_20_g13649/U$1 ( \1454 , \1450 , \1453 );
xnor \g45310/U$1 ( \1455 , \1446 , \1454 );
nand \g45309/U$1 ( \1456 , \982 , \1455 );
and \g2832/U$1 ( \1457 , \1445 , \1456 , \837 );
not \g2831/U$1 ( \1458 , \1457 );
nand \add_5_20_g13816/U$1 ( \1459 , \653 , \703 );
not \add_5_20_g13647/U$3 ( \1460 , \643 );
not \add_5_20_g13647/U$4 ( \1461 , \633 );
or \add_5_20_g13647/U$2 ( \1462 , \1460 , \1461 );
not \add_5_20_g13770/U$1 ( \1463 , \697 );
nand \add_5_20_g13647/U$1 ( \1464 , \1462 , \1463 );
xnor \g45331/U$1 ( \1465 , \1459 , \1464 );
nand \g2910/U$1 ( \1466 , \1262 , \1465 );
not \sub_5_33_g9552/U$2 ( \1467 , \479 );
nand \sub_5_33_g9552/U$1 ( \1468 , \1467 , \397 );
not \sub_5_33_g9121/U$3 ( \1469 , \393 );
not \sub_5_33_g9121/U$4 ( \1470 , \433 );
or \sub_5_33_g9121/U$2 ( \1471 , \1469 , \1470 );
not \sub_5_33_g9247/U$1 ( \1472 , \473 );
nand \sub_5_33_g9121/U$1 ( \1473 , \1471 , \1472 );
xnor \g45537/U$1 ( \1474 , \1468 , \1473 );
nand \g2911/U$1 ( \1475 , \1474 , \981 );
and \g2834/U$1 ( \1476 , \1466 , \1475 , \837 );
nand \sub_5_33_g9317/U$1 ( \1477 , \389 , \472 );
not \sub_5_33_g9122/U$3 ( \1478 , \391 );
not \sub_5_33_g9122/U$4 ( \1479 , \433 );
or \sub_5_33_g9122/U$2 ( \1480 , \1478 , \1479 );
not \sub_5_33_g9378/U$1 ( \1481 , \468 );
nand \sub_5_33_g9122/U$1 ( \1482 , \1480 , \1481 );
xnor \g45538/U$1 ( \1483 , \1477 , \1482 );
not \g2879/U$3 ( \1484 , \1483 );
not \g2879/U$4 ( \1485 , \981 );
or \g2879/U$2 ( \1486 , \1484 , \1485 );
not \add_5_20_g13959/U$1 ( \1487 , \641 );
not \add_5_20_g13648/U$3 ( \1488 , \1487 );
not \add_5_20_g13648/U$4 ( \1489 , \633 );
or \add_5_20_g13648/U$2 ( \1490 , \1488 , \1489 );
nand \add_5_20_g13648/U$1 ( \1491 , \1490 , \694 );
not \add_5_20_g13801/U$2 ( \1492 , \696 );
nor \add_5_20_g13801/U$1 ( \1493 , \1492 , \642 );
xnor \g45652/U$1 ( \1494 , \1491 , \1493 );
or \g2879/U$5 ( \1495 , \981 , \1494 );
nand \g2879/U$1 ( \1496 , \1486 , \1495 );
not \fopt45591/U$1 ( \1497 , \837 );
nor \g2836/U$1 ( \1498 , \1496 , \1497 );
not \g2835/U$1 ( \1499 , \1498 );
nand \sub_5_33_g9340/U$1 ( \1500 , \391 , \1481 );
xnor \g45539/U$1 ( \1501 , \1500 , \433 );
nand \g2913/U$1 ( \1502 , \1202 , \1501 );
nand \add_5_20_g13792/U$1 ( \1503 , \1487 , \694 );
xnor \g45332/U$1 ( \1504 , \1503 , \633 );
nand \g2912/U$1 ( \1505 , \294 , \1504 );
and \g2838/U$1 ( \1506 , \1502 , \1505 , \837 );
not \g2837/U$1 ( \1507 , \1506 );
not \add_5_20_g13829/U$2 ( \1508 , \627 );
nor \add_5_20_g13829/U$1 ( \1509 , \1508 , \616 );
xnor \g45654/U$1 ( \1510 , \623 , \1509 );
or \g3073/U$2 ( \1511 , \1510 , \981 );
not \sub_5_33_g9473/U$1 ( \1512 , \425 );
nand \sub_5_33_g9356/U$1 ( \1513 , \420 , \1512 );
xnor \sub_5_33_g9523/U$1 ( \1514 , \415 , \1513 );
nand \g3074/U$1 ( \1515 , \293 , \1514 );
nand \g3073/U$1 ( \1516 , \1511 , \1515 );
nor \g2842/U$1 ( \1517 , \1516 , \1295 );
not \g2841/U$1 ( \1518 , \1517 );
not \add_5_20_g13812/U$2 ( \1519 , \622 );
nor \add_5_20_g13812/U$1 ( \1520 , \1519 , \619 );
xnor \g45333/U$1 ( \1521 , \620 , \1520 );
not \g2882/U$3 ( \1522 , \1521 );
not \g2947/U$1 ( \1523 , \981 );
not \g2882/U$4 ( \1524 , \1523 );
or \g2882/U$2 ( \1525 , \1522 , \1524 );
nand \sub_5_33_g9303/U$1 ( \1526 , \414 , \410 );
xor \g45656/U$1 ( \1527 , \1526 , \407 );
or \g2882/U$5 ( \1528 , \982 , \1527 );
nand \g2882/U$1 ( \1529 , \1525 , \1528 );
nor \g2844/U$1 ( \1530 , \1529 , \1054 );
not \g2843/U$1 ( \1531 , \1530 );
not \add_5_20_g14021/U$2 ( \1532 , \609 );
nor \add_5_20_g14021/U$1 ( \1533 , \1532 , \596 );
not \add_5_20_g13611/U$3 ( \1534 , \1533 );
not \add_5_20_g13611/U$4 ( \1535 , \715 );
or \add_5_20_g13611/U$2 ( \1536 , \1534 , \1535 );
and \add_5_20_g13652/U$2 ( \1537 , \748 , \609 );
nor \add_5_20_g13652/U$1 ( \1538 , \1537 , \753 );
nand \add_5_20_g13611/U$1 ( \1539 , \1536 , \1538 );
nand \add_5_20_g13794/U$1 ( \1540 , \962 , \758 );
xnor \add_5_20_g14017/U$1 ( \1541 , \1539 , \1540 );
and \g2870/U$2 ( \1542 , \297 , \1541 );
not \g2870/U$4 ( \1543 , \297 );
nor \sub_5_33_g9173/U$1 ( \1544 , \325 , \346 );
not \sub_5_33_g9090/U$3 ( \1545 , \1544 );
not \sub_5_33_g9090/U$4 ( \1546 , \490 );
or \sub_5_33_g9090/U$2 ( \1547 , \1545 , \1546 );
and \sub_5_33_g2/U$2 ( \1548 , \945 , \541 );
nor \sub_5_33_g2/U$1 ( \1549 , \1548 , \550 );
nand \sub_5_33_g9090/U$1 ( \1550 , \1547 , \1549 );
not \sub_5_33_g9279/U$2 ( \1551 , \555 );
nand \sub_5_33_g9279/U$1 ( \1552 , \1551 , \339 );
xnor \sub_5_33_g9536/U$1 ( \1553 , \1550 , \1552 );
and \g2870/U$3 ( \1554 , \1543 , \1553 );
nor \g2870/U$1 ( \1555 , \1542 , \1554 );
nand \sub_5_33_g9349/U$1 ( \1556 , \345 , \1006 );
not \sub_5_33_g9100/U$3 ( \1557 , \326 );
not \sub_5_33_g9100/U$4 ( \1558 , \489 );
or \sub_5_33_g9100/U$2 ( \1559 , \1557 , \1558 );
not \sub_5_33_g9153/U$1 ( \1560 , \541 );
nand \sub_5_33_g9100/U$1 ( \1561 , \1559 , \1560 );
xnor \g45532/U$1 ( \1562 , \1556 , \1561 );
and \g2871/U$2 ( \1563 , \960 , \1562 );
not \add_5_20_g13631/U$3 ( \1564 , \597 );
not \add_5_20_g13631/U$4 ( \1565 , \715 );
or \add_5_20_g13631/U$2 ( \1566 , \1564 , \1565 );
not \add_5_20_g13676/U$1 ( \1567 , \748 );
nand \add_5_20_g13631/U$1 ( \1568 , \1566 , \1567 );
nand \add_5_20_g13809/U$1 ( \1569 , \988 , \750 );
xnor \add_5_20_g14020/U$1 ( \1570 , \1568 , \1569 );
and \g2871/U$3 ( \1571 , \1570 , \983 );
nor \g2871/U$1 ( \1572 , \1563 , \1571 );
nand \sub_5_33_g9342/U$1 ( \1573 , \418 , \430 );
not \sub_5_33_g9141/U$3 ( \1574 , \420 );
not \sub_5_33_g9141/U$4 ( \1575 , \415 );
or \sub_5_33_g9141/U$2 ( \1576 , \1574 , \1575 );
nand \sub_5_33_g9141/U$1 ( \1577 , \1576 , \1512 );
xnor \g45540/U$1 ( \1578 , \1573 , \1577 );
not \g3069/U$3 ( \1579 , \1578 );
not \g3069/U$4 ( \1580 , \293 );
or \g3069/U$2 ( \1581 , \1579 , \1580 );
not \g3070/U$3 ( \1582 , \981 );
not \add_5_20_g13662/U$3 ( \1583 , \1273 );
not \add_5_20_g13662/U$4 ( \1584 , \623 );
or \add_5_20_g13662/U$2 ( \1585 , \1583 , \1584 );
nand \add_5_20_g13662/U$1 ( \1586 , \1585 , \627 );
not \add_5_20_g14035/U$2 ( \1587 , \630 );
nor \add_5_20_g14035/U$1 ( \1588 , \1587 , \615 );
xnor \g45653/U$1 ( \1589 , \1586 , \1588 );
not \g3070/U$4 ( \1590 , \1589 );
and \g3070/U$2 ( \1591 , \1582 , \1590 );
not \fopt45595/U$1 ( \1592 , \837 );
nor \g3070/U$1 ( \1593 , \1591 , \1592 );
nand \g3069/U$1 ( \1594 , \1581 , \1593 );
or \g45620/U$2 ( \1595 , \c[8] , \d[8] );
nand \g45620/U$1 ( \1596 , \1595 , \1282 );
nand \g45619/U$1 ( \1597 , \1596 , \674 );
not \add_5_20_g14034/U$2 ( \1598 , \676 );
nor \add_5_20_g14034/U$1 ( \1599 , \1598 , \644 );
xor \add_5_20_g14024/U$1 ( \1600 , \1597 , \1599 );
nor \add_6_14_g19606/U$1 ( \1601 , \a[27] , \b[27] );
not \add_6_14_g19477/U$2 ( \1602 , \1601 );
nand \add_6_14_g19605/U$1 ( \1603 , \a[27] , \b[27] );
nand \add_6_14_g19477/U$1 ( \1604 , \1602 , \1603 );
not \add_6_14_g19266/U$3 ( \1605 , \1604 );
nor \add_6_14_g19617/U$1 ( \1606 , \a[24] , \b[24] );
nor \add_6_14_g19651/U$1 ( \1607 , \a[25] , \b[25] );
nor \add_6_14_g19555/U$1 ( \1608 , \1606 , \1607 );
nor \add_6_14_g19585/U$1 ( \1609 , \a[26] , \b[26] );
not \add_6_14_g19584/U$1 ( \1610 , \1609 );
and \add_6_14_g19428/U$1 ( \1611 , \1608 , \1610 );
not \add_6_14_g19387/U$2 ( \1612 , \1611 );
nor \add_6_14_g19573/U$1 ( \1613 , \a[19] , \b[19] );
nor \add_6_14_g19604/U$1 ( \1614 , \a[18] , \b[18] );
nor \add_6_14_g19553/U$1 ( \1615 , \1613 , \1614 );
nor \add_6_14_g19629/U$1 ( \1616 , \a[16] , \b[16] );
nor \add_6_14_g19586/U$1 ( \1617 , \a[17] , \b[17] );
nor \add_6_14_g19556/U$1 ( \1618 , \1616 , \1617 );
and \add_6_14_g19440/U$1 ( \1619 , \1615 , \1618 );
nor \add_6_14_g19615/U$1 ( \1620 , \a[21] , \b[21] );
nor \add_6_14_g19626/U$1 ( \1621 , \a[20] , \b[20] );
nor \add_6_14_g19512/U$1 ( \1622 , \1620 , \1621 );
nor \add_6_14_g19588/U$1 ( \1623 , \a[22] , \b[22] );
nor \add_6_14_g19574/U$1 ( \1624 , \a[23] , \b[23] );
nor \add_6_14_g19521/U$1 ( \1625 , \1623 , \1624 );
and \add_6_14_g19436/U$1 ( \1626 , \1622 , \1625 );
and \add_6_14_g19420/U$1 ( \1627 , \1619 , \1626 );
not \add_6_14_g19419/U$1 ( \1628 , \1627 );
nor \add_6_14_g19387/U$1 ( \1629 , \1612 , \1628 );
not \add_6_14_g19301/U$3 ( \1630 , \1629 );
nor \add_6_14_g45823/U$1 ( \1631 , \a[9] , \b[9] );
nand \add_6_14_g19656/U$1 ( \1632 , \a[8] , \b[8] );
or \add_6_14_g19467/U$2 ( \1633 , \1631 , \1632 );
nand \add_6_14_g19646/U$1 ( \1634 , \a[9] , \b[9] );
nand \add_6_14_g19467/U$1 ( \1635 , \1633 , \1634 );
nor \add_6_14_g19640/U$1 ( \1636 , \a[11] , \b[11] );
nand \add_6_14_g19619/U$1 ( \1637 , \a[10] , \b[10] );
or \add_6_14_g19462/U$2 ( \1638 , \1636 , \1637 );
nand \add_6_14_g19608/U$1 ( \1639 , \a[11] , \b[11] );
nand \add_6_14_g19462/U$1 ( \1640 , \1638 , \1639 );
nor \add_6_14_g19418/U$1 ( \1641 , \1635 , \1640 );
not \g45821/U$3 ( \1642 , \a[9] );
not \g45821/U$4 ( \1643 , \b[9] );
and \g45821/U$2 ( \1644 , \1642 , \1643 );
nor \add_6_14_g45827/U$1 ( \1645 , \a[8] , \b[8] );
nor \g45821/U$1 ( \1646 , \1644 , \1645 );
nor \add_6_14_g19612/U$1 ( \1647 , \a[7] , \b[7] );
nand \add_6_14_g19643/U$1 ( \1648 , \a[6] , \b[6] );
or \add_6_14_g19469/U$2 ( \1649 , \1647 , \1648 );
nand \add_6_14_g19658/U$1 ( \1650 , \a[7] , \b[7] );
nand \add_6_14_g19469/U$1 ( \1651 , \1649 , \1650 );
nand \add_6_14_g19416/U$1 ( \1652 , \1646 , \1651 );
nor \add_6_14_g19592/U$1 ( \1653 , \a[9] , \b[9] );
nor \add_6_14_g19534/U$1 ( \1654 , \1653 , \1645 );
nand \add_6_14_g19634/U$1 ( \1655 , \a[5] , \b[5] );
not \add_6_14_g19633/U$1 ( \1656 , \1655 );
nand \add_6_14_g19446/U$1 ( \1657 , \1654 , \1656 );
nor \add_6_14_g19676/U$1 ( \1658 , \a[5] , \b[5] );
nand \add_6_14_g19602/U$1 ( \1659 , \a[4] , \b[4] );
nor \add_6_14_g19543/U$1 ( \1660 , \1658 , \1659 );
nand \add_6_14_g19447/U$1 ( \1661 , \1654 , \1660 );
nand \add_6_14_g19376/U$1 ( \1662 , \1641 , \1652 , \1657 , \1661 );
not \add_6_14_g19403/U$3 ( \1663 , \1640 );
nor \add_6_14_g19569/U$1 ( \1664 , \a[10] , \b[10] );
nor \add_6_14_g19641/U$1 ( \1665 , \a[11] , \b[11] );
nor \add_6_14_g19484/U$1 ( \1666 , \1664 , \1665 );
not \add_6_14_g19403/U$4 ( \1667 , \1666 );
and \add_6_14_g19403/U$2 ( \1668 , \1663 , \1667 );
or \g45665/U$1 ( \1669 , \a[13] , \b[13] );
not \add_6_14_g19706/U$2 ( \1670 , \1669 );
nor \add_6_14_g19650/U$1 ( \1671 , \a[12] , \b[12] );
nor \add_6_14_g19706/U$1 ( \1672 , \1670 , \1671 );
nor \add_6_14_g19670/U$1 ( \1673 , \a[15] , \b[15] );
nor \add_6_14_g19621/U$1 ( \1674 , \a[14] , \b[14] );
nor \add_6_14_g19560/U$1 ( \1675 , \1673 , \1674 );
nand \add_6_14_g19432/U$1 ( \1676 , \1672 , \1675 );
nor \add_6_14_g19403/U$1 ( \1677 , \1668 , \1676 );
not \add_6_14_g19409/U$2 ( \1678 , \1651 );
not \add_6_14_g19461/U$1 ( \1679 , \1640 );
not \add_6_14_g19466/U$1 ( \1680 , \1635 );
nor \add_6_14_g19594/U$1 ( \1681 , \a[6] , \b[6] );
nor \add_6_14_g19613/U$1 ( \1682 , \a[7] , \b[7] );
or \add_6_14_g19514/U$1 ( \1683 , \1681 , \1682 );
nand \add_6_14_g19409/U$1 ( \1684 , \1678 , \1679 , \1680 , \1683 );
nand \add_6_14_g19365/U$1 ( \1685 , \1662 , \1677 , \1684 );
nor \add_6_14_g19597/U$1 ( \1686 , \a[4] , \b[4] );
nor \add_6_14_g19519/U$1 ( \1687 , \1658 , \1686 );
nand \add_6_14_g19435/U$1 ( \1688 , \1646 , \1687 );
nor \add_6_14_g19540/U$1 ( \1689 , \1681 , \1671 );
nor \add_6_14_g19552/U$1 ( \1690 , \1664 , \1674 );
not \g45726/U$3 ( \1691 , \a[13] );
not \g45726/U$4 ( \1692 , \b[13] );
and \g45726/U$2 ( \1693 , \1691 , \1692 );
nor \g45726/U$1 ( \1694 , \1693 , \1647 );
nor \add_6_14_g19554/U$1 ( \1695 , \1673 , \1636 );
nand \add_6_14_g19426/U$1 ( \1696 , \1689 , \1690 , \1694 , \1695 );
nor \add_6_14_g19408/U$1 ( \1697 , \1688 , \1696 );
nor \add_6_14_g19662/U$1 ( \1698 , \a[3] , \b[3] );
nor \add_6_14_g19660/U$1 ( \1699 , \a[2] , \b[2] );
nor \add_6_14_g19488/U$1 ( \1700 , \1698 , \1699 );
not \g45725/U$3 ( \1701 , \1700 );
nand \add_6_14_g19599/U$1 ( \1702 , \a[3] , \b[3] );
not \add_6_14_g19598/U$1 ( \1703 , \1702 );
not \g45725/U$4 ( \1704 , \1703 );
and \g45725/U$2 ( \1705 , \1701 , \1704 );
nor \add_6_14_g19589/U$1 ( \1706 , \a[1] , \b[1] );
nand \g45805/U$2 ( \1707 , \a[0] , \b[0] );
nor \add_6_14_g19411/U$1 ( \1708 , \1706 , \1707 );
nand \add_6_14_g19638/U$1 ( \1709 , \a[2] , \b[2] );
nand \add_6_14_g19581/U$1 ( \1710 , \a[1] , \b[1] );
nand \add_6_14_g19475/U$1 ( \1711 , \1702 , \1709 , \1710 );
nor \add_6_14_g19392/U$1 ( \1712 , \1708 , \1711 );
nor \g45725/U$1 ( \1713 , \1705 , \1712 );
and \add_6_14_g19354/U$2 ( \1714 , \1697 , \1713 );
not \add_6_14_g19396/U$3 ( \1715 , \1675 );
and \add_6_14_g45828/U$1 ( \1716 , \a[12] , \b[12] );
not \add_6_14_g19474/U$3 ( \1717 , \1716 );
not \add_6_14_g19474/U$4 ( \1718 , \1669 );
or \add_6_14_g19474/U$2 ( \1719 , \1717 , \1718 );
nand \add_6_14_g19567/U$1 ( \1720 , \a[13] , \b[13] );
nand \add_6_14_g19474/U$1 ( \1721 , \1719 , \1720 );
not \add_6_14_g19396/U$4 ( \1722 , \1721 );
or \add_6_14_g19396/U$2 ( \1723 , \1715 , \1722 );
nor \add_6_14_g19671/U$1 ( \1724 , \a[15] , \b[15] );
nand \add_6_14_g19668/U$1 ( \1725 , \a[14] , \b[14] );
or \add_6_14_g19454/U$2 ( \1726 , \1724 , \1725 );
nand \add_6_14_g19609/U$1 ( \1727 , \a[15] , \b[15] );
nand \add_6_14_g19454/U$1 ( \1728 , \1726 , \1727 );
not \add_6_14_g19453/U$1 ( \1729 , \1728 );
nand \add_6_14_g19396/U$1 ( \1730 , \1723 , \1729 );
nor \add_6_14_g19354/U$1 ( \1731 , \1714 , \1730 );
nand \add_6_14_g19332/U$1 ( \1732 , \1685 , \1731 );
not \add_6_14_g19330/U$1 ( \1733 , \1732 );
not \add_6_14_g19328/U$1 ( \1734 , \1733 );
not \add_6_14_g19301/U$4 ( \1735 , \1734 );
or \add_6_14_g19301/U$2 ( \1736 , \1630 , \1735 );
not \add_6_14_g19367/U$3 ( \1737 , \1626 );
nand \add_6_14_g19653/U$1 ( \1738 , \a[16] , \b[16] );
or \add_6_14_g19459/U$2 ( \1739 , \1617 , \1738 );
nand \add_6_14_g19622/U$1 ( \1740 , \a[17] , \b[17] );
nand \add_6_14_g19459/U$1 ( \1741 , \1739 , \1740 );
not \add_6_14_g19400/U$3 ( \1742 , \1741 );
not \add_6_14_g19400/U$4 ( \1743 , \1615 );
or \add_6_14_g19400/U$2 ( \1744 , \1742 , \1743 );
not \add_6_14_g19572/U$1 ( \1745 , \1613 );
nand \add_6_14_g19645/U$1 ( \1746 , \a[18] , \b[18] );
not \add_6_14_g19644/U$1 ( \1747 , \1746 );
and \add_6_14_g19470/U$2 ( \1748 , \1745 , \1747 );
and \add_6_14_g19707/U$1 ( \1749 , \a[19] , \b[19] );
nor \add_6_14_g19470/U$1 ( \1750 , \1748 , \1749 );
nand \add_6_14_g19400/U$1 ( \1751 , \1744 , \1750 );
not \add_6_14_g19367/U$4 ( \1752 , \1751 );
or \add_6_14_g19367/U$2 ( \1753 , \1737 , \1752 );
nand \add_6_14_g19666/U$1 ( \1754 , \a[20] , \b[20] );
not \add_6_14_g19665/U$1 ( \1755 , \1754 );
not \add_6_14_g19452/U$3 ( \1756 , \1755 );
not \add_6_14_g19614/U$1 ( \1757 , \1620 );
not \add_6_14_g19452/U$4 ( \1758 , \1757 );
or \add_6_14_g19452/U$2 ( \1759 , \1756 , \1758 );
nand \add_6_14_g19657/U$1 ( \1760 , \a[21] , \b[21] );
nand \add_6_14_g19452/U$1 ( \1761 , \1759 , \1760 );
and \add_6_14_g19406/U$2 ( \1762 , \1761 , \1625 );
nand \add_6_14_g19623/U$1 ( \1763 , \a[22] , \b[22] );
or \add_6_14_g19471/U$2 ( \1764 , \1624 , \1763 );
nand \add_6_14_g19672/U$1 ( \1765 , \a[23] , \b[23] );
nand \add_6_14_g19471/U$1 ( \1766 , \1764 , \1765 );
nor \add_6_14_g19406/U$1 ( \1767 , \1762 , \1766 );
nand \add_6_14_g19367/U$1 ( \1768 , \1753 , \1767 );
and \add_6_14_g19346/U$2 ( \1769 , \1768 , \1611 );
not \add_6_14_g19394/U$3 ( \1770 , \1610 );
nand \add_6_14_g19611/U$1 ( \1771 , \a[24] , \b[24] );
or \add_6_14_g19455/U$2 ( \1772 , \1607 , \1771 );
nand \add_6_14_g19590/U$1 ( \1773 , \a[25] , \b[25] );
nand \add_6_14_g19455/U$1 ( \1774 , \1772 , \1773 );
not \add_6_14_g19394/U$4 ( \1775 , \1774 );
or \add_6_14_g19394/U$2 ( \1776 , \1770 , \1775 );
nand \add_6_14_g19630/U$1 ( \1777 , \a[26] , \b[26] );
nand \add_6_14_g19394/U$1 ( \1778 , \1776 , \1777 );
nor \add_6_14_g19346/U$1 ( \1779 , \1769 , \1778 );
nand \add_6_14_g19301/U$1 ( \1780 , \1736 , \1779 );
not \add_6_14_g19266/U$4 ( \1781 , \1780 );
or \add_6_14_g19266/U$2 ( \1782 , \1605 , \1781 );
or \add_6_14_g19266/U$5 ( \1783 , \1780 , \1604 );
nand \add_6_14_g19266/U$1 ( \1784 , \1782 , \1783 );
nor \add_6_14_g19635/U$1 ( \1785 , \a[29] , \b[29] );
and \add_6_14_g19639/U$1 ( \1786 , \a[29] , \b[29] );
or \add_6_14_g19559/U$1 ( \1787 , \1785 , \1786 );
not \add_6_14_g19278/U$3 ( \1788 , \1787 );
nor \add_6_14_g19509/U$1 ( \1789 , \1601 , \1609 );
nand \add_6_14_g19431/U$1 ( \1790 , \1789 , \1608 );
nor \add_6_14_g19669/U$1 ( \1791 , \a[28] , \b[28] );
nor \add_6_14_g19422/U$1 ( \1792 , \1790 , \1791 );
nand \g45719/U$1 ( \1793 , \1734 , \1627 , \1792 );
and \add_6_14_g19343/U$2 ( \1794 , \1768 , \1792 );
and \add_6_14_g19405/U$2 ( \1795 , \1789 , \1774 );
or \add_6_14_g19472/U$2 ( \1796 , \1601 , \1777 );
nand \add_6_14_g19472/U$1 ( \1797 , \1796 , \1603 );
nor \add_6_14_g19405/U$1 ( \1798 , \1795 , \1797 );
or \add_6_14_g19361/U$2 ( \1799 , \1798 , \1791 );
nand \add_6_14_g19627/U$1 ( \1800 , \a[28] , \b[28] );
nand \add_6_14_g19361/U$1 ( \1801 , \1799 , \1800 );
nor \add_6_14_g19343/U$1 ( \1802 , \1794 , \1801 );
nand \add_6_14_g19294/U$1 ( \1803 , \1793 , \1802 );
not \add_6_14_g19278/U$4 ( \1804 , \1803 );
or \add_6_14_g19278/U$2 ( \1805 , \1788 , \1804 );
or \add_6_14_g19278/U$5 ( \1806 , \1803 , \1787 );
nand \add_6_14_g19278/U$1 ( \1807 , \1805 , \1806 );
not \add_6_14_g19620/U$1 ( \1808 , \1674 );
nand \add_6_14_g19480/U$1 ( \1809 , \1808 , \1725 );
not \add_6_14_g19287/U$3 ( \1810 , \1809 );
not \add_6_14_g19686/U$2 ( \1811 , \1672 );
nand \add_6_14_g19443/U$1 ( \1812 , \1646 , \1666 );
nor \add_6_14_g19686/U$1 ( \1813 , \1811 , \1812 );
not \add_6_14_g19323/U$3 ( \1814 , \1813 );
not \add_6_14_g19693/U$2 ( \1815 , \1687 );
nor \add_6_14_g19693/U$1 ( \1816 , \1815 , \1683 );
not \add_6_14_g19352/U$3 ( \1817 , \1816 );
not \add_6_14_g19352/U$4 ( \1818 , \1713 );
or \add_6_14_g19352/U$2 ( \1819 , \1817 , \1818 );
not \add_6_14_g19698/U$2 ( \1820 , \1660 );
nand \add_6_14_g19698/U$1 ( \1821 , \1820 , \1655 );
not \add_6_14_g19513/U$1 ( \1822 , \1683 );
and \add_6_14_g19391/U$2 ( \1823 , \1821 , \1822 );
nor \add_6_14_g19391/U$1 ( \1824 , \1823 , \1651 );
nand \add_6_14_g19352/U$1 ( \1825 , \1819 , \1824 );
not \add_6_14_g19323/U$4 ( \1826 , \1825 );
or \add_6_14_g19323/U$2 ( \1827 , \1814 , \1826 );
not \add_6_14_g19390/U$3 ( \1828 , \1666 );
not \add_6_14_g19390/U$4 ( \1829 , \1635 );
or \add_6_14_g19390/U$2 ( \1830 , \1828 , \1829 );
nand \add_6_14_g19390/U$1 ( \1831 , \1830 , \1679 );
and \add_6_14_g19358/U$2 ( \1832 , \1831 , \1672 );
nor \add_6_14_g19358/U$1 ( \1833 , \1832 , \1721 );
nand \add_6_14_g19323/U$1 ( \1834 , \1827 , \1833 );
not \add_6_14_g19287/U$4 ( \1835 , \1834 );
or \add_6_14_g19287/U$2 ( \1836 , \1810 , \1835 );
or \add_6_14_g19287/U$5 ( \1837 , \1834 , \1809 );
nand \add_6_14_g19287/U$1 ( \1838 , \1836 , \1837 );
not \add_6_14_g19628/U$1 ( \1839 , \1616 );
not \add_6_14_g19289/U$3 ( \1840 , \1839 );
nand \add_6_14_g19325/U$1 ( \1841 , \1685 , \1731 );
not \add_6_14_g19289/U$4 ( \1842 , \1841 );
or \add_6_14_g19289/U$2 ( \1843 , \1840 , \1842 );
nand \add_6_14_g19289/U$1 ( \1844 , \1843 , \1738 );
not \add_6_14_g19320/U$3 ( \1845 , \1646 );
not \add_6_14_g19320/U$4 ( \1846 , \1825 );
or \add_6_14_g19320/U$2 ( \1847 , \1845 , \1846 );
nand \add_6_14_g19320/U$1 ( \1848 , \1847 , \1680 );
not \add_6_14_g19568/U$1 ( \1849 , \1664 );
nand \add_6_14_g19549/U$1 ( \1850 , \1849 , \1637 );
nand \add_6_14_g19290/U$1 ( \1851 , \1848 , \1850 );
nor \add_6_14_g19415/U$1 ( \1852 , \1812 , \1671 );
not \add_6_14_g19316/U$3 ( \1853 , \1852 );
not \add_6_14_g19316/U$4 ( \1854 , \1825 );
or \add_6_14_g19316/U$2 ( \1855 , \1853 , \1854 );
not \add_6_14_g19647/U$1 ( \1856 , \1671 );
and \add_6_14_g19359/U$2 ( \1857 , \1831 , \1856 );
nor \add_6_14_g19359/U$1 ( \1858 , \1857 , \1716 );
nand \add_6_14_g19316/U$1 ( \1859 , \1855 , \1858 );
nand \add_6_14_g19479/U$1 ( \1860 , \1669 , \1720 );
nand \add_6_14_g19291/U$1 ( \1861 , \1859 , \1860 );
not \add_6_14_g19292/U$3 ( \1862 , \1618 );
not \add_6_14_g19292/U$4 ( \1863 , \1732 );
or \add_6_14_g19292/U$2 ( \1864 , \1862 , \1863 );
not \add_6_14_g19457/U$1 ( \1865 , \1741 );
nand \add_6_14_g19292/U$1 ( \1866 , \1864 , \1865 );
and \add_6_14_g19379/U$1 ( \1867 , \1627 , \1608 );
not \add_6_14_g19295/U$3 ( \1868 , \1867 );
not \add_6_14_g19295/U$4 ( \1869 , \1734 );
or \add_6_14_g19295/U$2 ( \1870 , \1868 , \1869 );
and \add_6_14_g19333/U$2 ( \1871 , \1768 , \1608 );
nor \add_6_14_g19333/U$1 ( \1872 , \1871 , \1774 );
nand \add_6_14_g19295/U$1 ( \1873 , \1870 , \1872 );
nor \add_6_14_g19566/U$1 ( \1874 , \a[30] , \b[30] );
not \add_6_14_g19438/U$2 ( \1875 , \1874 );
nor \add_6_14_g19541/U$1 ( \1876 , \1785 , \1791 );
nand \add_6_14_g19438/U$1 ( \1877 , \1875 , \1876 );
nor \add_6_14_g19424/U$1 ( \1878 , \1790 , \1877 );
and \add_6_14_g19384/U$1 ( \1879 , \1627 , \1878 );
not \add_6_14_g19296/U$3 ( \1880 , \1879 );
not \add_6_14_g19296/U$4 ( \1881 , \1734 );
or \add_6_14_g19296/U$2 ( \1882 , \1880 , \1881 );
and \add_6_14_g19341/U$2 ( \1883 , \1768 , \1878 );
or \add_6_14_g19372/U$2 ( \1884 , \1798 , \1877 );
not \add_6_14_g19451/U$3 ( \1885 , \1785 );
not \add_6_14_g19451/U$4 ( \1886 , \1800 );
and \add_6_14_g19451/U$2 ( \1887 , \1885 , \1886 );
nor \add_6_14_g19451/U$1 ( \1888 , \1887 , \1786 );
or \add_6_14_g19372/U$3 ( \1889 , \1874 , \1888 );
nand \add_6_14_g19607/U$1 ( \1890 , \a[30] , \b[30] );
nand \add_6_14_g19372/U$1 ( \1891 , \1884 , \1889 , \1890 );
nor \add_6_14_g19341/U$1 ( \1892 , \1883 , \1891 );
nand \add_6_14_g19296/U$1 ( \1893 , \1882 , \1892 );
nor \add_6_14_g19380/U$1 ( \1894 , \1628 , \1606 );
not \add_6_14_g19297/U$3 ( \1895 , \1894 );
not \add_6_14_g19297/U$4 ( \1896 , \1734 );
or \add_6_14_g19297/U$2 ( \1897 , \1895 , \1896 );
not \add_6_14_g19616/U$1 ( \1898 , \1606 );
and \add_6_14_g19335/U$2 ( \1899 , \1768 , \1898 );
not \add_6_14_g19610/U$1 ( \1900 , \1771 );
nor \add_6_14_g19335/U$1 ( \1901 , \1899 , \1900 );
nand \add_6_14_g19297/U$1 ( \1902 , \1897 , \1901 );
not \add_6_14_g19587/U$1 ( \1903 , \1623 );
and \add_6_14_g19433/U$1 ( \1904 , \1622 , \1903 );
and \add_6_14_g19423/U$1 ( \1905 , \1619 , \1904 );
not \add_6_14_g19298/U$3 ( \1906 , \1905 );
not \add_6_14_g19298/U$4 ( \1907 , \1732 );
or \add_6_14_g19298/U$2 ( \1908 , \1906 , \1907 );
and \add_6_14_g19374/U$2 ( \1909 , \1751 , \1904 );
not \add_6_14_g19395/U$3 ( \1910 , \1903 );
not \add_6_14_g19395/U$4 ( \1911 , \1761 );
or \add_6_14_g19395/U$2 ( \1912 , \1910 , \1911 );
nand \add_6_14_g19395/U$1 ( \1913 , \1912 , \1763 );
nor \add_6_14_g19374/U$1 ( \1914 , \1909 , \1913 );
nand \add_6_14_g19298/U$1 ( \1915 , \1908 , \1914 );
not \add_6_14_g19692/U$2 ( \1916 , \1622 );
not \add_6_14_g19439/U$1 ( \1917 , \1619 );
nor \add_6_14_g19692/U$1 ( \1918 , \1916 , \1917 );
not \add_6_14_g19299/U$3 ( \1919 , \1918 );
not \add_6_14_g19299/U$4 ( \1920 , \1732 );
or \add_6_14_g19299/U$2 ( \1921 , \1919 , \1920 );
and \add_6_14_g19355/U$2 ( \1922 , \1751 , \1622 );
nor \add_6_14_g19355/U$1 ( \1923 , \1922 , \1761 );
nand \add_6_14_g19299/U$1 ( \1924 , \1921 , \1923 );
not \add_6_14_g19300/U$3 ( \1925 , \1619 );
not \add_6_14_g19300/U$4 ( \1926 , \1732 );
or \add_6_14_g19300/U$2 ( \1927 , \1925 , \1926 );
not \add_6_14_g19398/U$1 ( \1928 , \1751 );
nand \add_6_14_g19300/U$1 ( \1929 , \1927 , \1928 );
nor \add_6_14_g19385/U$1 ( \1930 , \1628 , \1790 );
not \add_6_14_g19302/U$3 ( \1931 , \1930 );
not \add_6_14_g19302/U$4 ( \1932 , \1734 );
or \add_6_14_g19302/U$2 ( \1933 , \1931 , \1932 );
not \add_6_14_g19430/U$1 ( \1934 , \1790 );
and \add_6_14_g19337/U$2 ( \1935 , \1768 , \1934 );
not \add_6_14_g19404/U$1 ( \1936 , \1798 );
nor \add_6_14_g19337/U$1 ( \1937 , \1935 , \1936 );
nand \add_6_14_g19302/U$1 ( \1938 , \1933 , \1937 );
not \add_6_14_g19603/U$1 ( \1939 , \1614 );
and \add_6_14_g19437/U$1 ( \1940 , \1618 , \1939 );
not \add_6_14_g19303/U$3 ( \1941 , \1940 );
not \add_6_14_g19303/U$4 ( \1942 , \1732 );
or \add_6_14_g19303/U$2 ( \1943 , \1941 , \1942 );
and \add_6_14_g19397/U$2 ( \1944 , \1741 , \1939 );
nor \add_6_14_g19397/U$1 ( \1945 , \1944 , \1747 );
nand \add_6_14_g19303/U$1 ( \1946 , \1943 , \1945 );
and \add_6_14_g19421/U$1 ( \1947 , \1934 , \1876 );
and \add_6_14_g19386/U$1 ( \1948 , \1627 , \1947 );
not \add_6_14_g19304/U$3 ( \1949 , \1948 );
not \add_6_14_g19304/U$4 ( \1950 , \1734 );
or \add_6_14_g19304/U$2 ( \1951 , \1949 , \1950 );
and \add_6_14_g19342/U$2 ( \1952 , \1768 , \1947 );
not \add_6_14_g19360/U$3 ( \1953 , \1876 );
not \add_6_14_g19360/U$4 ( \1954 , \1936 );
or \add_6_14_g19360/U$2 ( \1955 , \1953 , \1954 );
nand \add_6_14_g19360/U$1 ( \1956 , \1955 , \1888 );
nor \add_6_14_g19342/U$1 ( \1957 , \1952 , \1956 );
nand \add_6_14_g19304/U$1 ( \1958 , \1951 , \1957 );
not \add_6_14_g19305/U$3 ( \1959 , \1627 );
not \add_6_14_g19305/U$4 ( \1960 , \1732 );
or \add_6_14_g19305/U$2 ( \1961 , \1959 , \1960 );
not \add_6_14_g19366/U$1 ( \1962 , \1768 );
nand \add_6_14_g19305/U$1 ( \1963 , \1961 , \1962 );
nand \add_6_14_g19539/U$1 ( \1964 , \1839 , \1738 );
not \add_6_14_g19306/U$3 ( \1965 , \1964 );
not \add_6_14_g19306/U$4 ( \1966 , \1732 );
or \add_6_14_g19306/U$2 ( \1967 , \1965 , \1966 );
not \add_6_14_g19313/U$2 ( \1968 , \1964 );
nand \add_6_14_g19313/U$1 ( \1969 , \1968 , \1733 );
nand \add_6_14_g19306/U$1 ( \1970 , \1967 , \1969 );
not \add_6_14_g19538/U$2 ( \1971 , \1682 );
nand \add_6_14_g19538/U$1 ( \1972 , \1971 , \1650 );
not \add_6_14_g19308/U$3 ( \1973 , \1972 );
not \add_6_14_g19427/U$2 ( \1974 , \1687 );
nor \add_6_14_g19427/U$1 ( \1975 , \1974 , \1681 );
not \add_6_14_g19338/U$3 ( \1976 , \1975 );
not \add_6_14_g19680/U$2 ( \1977 , \1708 );
nand \add_6_14_g19680/U$1 ( \1978 , \1977 , \1710 );
nand \add_6_14_g19375/U$1 ( \1979 , \1978 , \1700 );
not \add_6_14_g19456/U$3 ( \1980 , \1698 );
not \add_6_14_g19456/U$4 ( \1981 , \1709 );
and \add_6_14_g19456/U$2 ( \1982 , \1980 , \1981 );
nor \add_6_14_g19456/U$1 ( \1983 , \1982 , \1703 );
nand \add_6_14_g19371/U$1 ( \1984 , \1979 , \1983 );
not \add_6_14_g19338/U$4 ( \1985 , \1984 );
or \add_6_14_g19338/U$2 ( \1986 , \1976 , \1985 );
not \add_6_14_g19444/U$1 ( \1987 , \1821 );
not \add_6_14_g19393/U$3 ( \1988 , \1987 );
not \add_6_14_g19393/U$4 ( \1989 , \1681 );
and \add_6_14_g19393/U$2 ( \1990 , \1988 , \1989 );
not \add_6_14_g19642/U$1 ( \1991 , \1648 );
nor \add_6_14_g19393/U$1 ( \1992 , \1990 , \1991 );
nand \add_6_14_g19338/U$1 ( \1993 , \1986 , \1992 );
not \add_6_14_g19308/U$4 ( \1994 , \1993 );
or \add_6_14_g19308/U$2 ( \1995 , \1973 , \1994 );
or \add_6_14_g19308/U$5 ( \1996 , \1993 , \1972 );
nand \add_6_14_g19308/U$1 ( \1997 , \1995 , \1996 );
buf \add_6_14_g19307/U$1 ( \1998 , \1997 );
not \add_6_14_g19595/U$1 ( \1999 , \1686 );
not \add_6_14_g19336/U$3 ( \2000 , \1999 );
not \add_6_14_g19336/U$4 ( \2001 , \1984 );
or \add_6_14_g19336/U$2 ( \2002 , \2000 , \2001 );
nand \add_6_14_g19336/U$1 ( \2003 , \2002 , \1659 );
nor \add_6_14_g19530/U$1 ( \2004 , \1656 , \1658 );
xor \add_6_14_g19696/U$1 ( \2005 , \2003 , \2004 );
buf \add_6_14_g19309/U$1 ( \2006 , \2005 );
not \add_6_14_g19441/U$1 ( \2007 , \1812 );
not \add_6_14_g19314/U$3 ( \2008 , \2007 );
not \add_6_14_g19314/U$4 ( \2009 , \1825 );
or \add_6_14_g19314/U$2 ( \2010 , \2008 , \2009 );
not \add_6_14_g19388/U$1 ( \2011 , \1831 );
nand \add_6_14_g19314/U$1 ( \2012 , \2010 , \2011 );
not \add_6_14_g19663/U$1 ( \2013 , \1645 );
not \add_6_14_g19317/U$3 ( \2014 , \2013 );
not \add_6_14_g19317/U$4 ( \2015 , \1825 );
or \add_6_14_g19317/U$2 ( \2016 , \2014 , \2015 );
nand \add_6_14_g19317/U$1 ( \2017 , \2016 , \1632 );
and \add_6_14_g19449/U$1 ( \2018 , \1672 , \1808 );
not \add_6_14_g19681/U$2 ( \2019 , \2018 );
nor \add_6_14_g19681/U$1 ( \2020 , \2019 , \1812 );
not \add_6_14_g19318/U$3 ( \2021 , \2020 );
not \add_6_14_g19318/U$4 ( \2022 , \1825 );
or \add_6_14_g19318/U$2 ( \2023 , \2021 , \2022 );
and \g45704/U$2 ( \2024 , \2018 , \1831 );
and \g45704/U$3 ( \2025 , \1721 , \1808 );
not \add_6_14_g19667/U$1 ( \2026 , \1725 );
nor \g45704/U$1 ( \2027 , \2024 , \2025 , \2026 );
nand \add_6_14_g19318/U$1 ( \2028 , \2023 , \2027 );
and \add_6_14_g19450/U$1 ( \2029 , \1646 , \1849 );
not \add_6_14_g19322/U$3 ( \2030 , \2029 );
not \add_6_14_g19322/U$4 ( \2031 , \1825 );
or \add_6_14_g19322/U$2 ( \2032 , \2030 , \2031 );
and \add_6_14_g19402/U$2 ( \2033 , \1635 , \1849 );
not \add_6_14_g19618/U$1 ( \2034 , \1637 );
nor \add_6_14_g19402/U$1 ( \2035 , \2033 , \2034 );
nand \add_6_14_g19322/U$1 ( \2036 , \2032 , \2035 );
not \add_6_14_g19340/U$3 ( \2037 , \1687 );
not \add_6_14_g19340/U$4 ( \2038 , \1984 );
or \add_6_14_g19340/U$2 ( \2039 , \2037 , \2038 );
nand \add_6_14_g19340/U$1 ( \2040 , \2039 , \1987 );
not \add_6_14_g19624/U$1 ( \2041 , \1621 );
not \add_6_14_g19357/U$3 ( \2042 , \2041 );
not \add_6_14_g19357/U$4 ( \2043 , \1751 );
or \add_6_14_g19357/U$2 ( \2044 , \2042 , \2043 );
nand \add_6_14_g19357/U$1 ( \2045 , \2044 , \1754 );
not \add_6_14_g19381/U$1 ( \2046 , \1978 );
or \add_6_14_g19363/U$2 ( \2047 , \2046 , \1699 );
nand \add_6_14_g19363/U$1 ( \2048 , \2047 , \1709 );
not \add_6_14_g19370/U$1 ( \2049 , \1984 );
not \add_6_14_g19407/U$3 ( \2050 , \1707 );
not \add_6_14_g19705/U$2 ( \2051 , \1710 );
nor \add_6_14_g19705/U$1 ( \2052 , \2051 , \1706 );
not \add_6_14_g19407/U$4 ( \2053 , \2052 );
or \add_6_14_g19407/U$2 ( \2054 , \2050 , \2053 );
or \add_6_14_g19425/U$1 ( \2055 , \2052 , \1707 );
nand \add_6_14_g19407/U$1 ( \2056 , \2054 , \2055 );
xor \g45805/U$1 ( \2057 , \a[0] , \b[0] );
buf \add_6_14_g19476/U$1 ( \2058 , \2057 );
nand \add_6_14_g19482/U$1 ( \2059 , \1610 , \1777 );
not \add_6_14_g19490/U$2 ( \2060 , \1890 );
nor \add_6_14_g19490/U$1 ( \2061 , \2060 , \1874 );
nand \add_6_14_g19492/U$1 ( \2062 , \1898 , \1771 );
not \add_6_14_g19498/U$2 ( \2063 , \1607 );
nand \add_6_14_g19498/U$1 ( \2064 , \2063 , \1773 );
not \add_6_14_g19500/U$2 ( \2065 , \1765 );
nor \add_6_14_g19500/U$1 ( \2066 , \2065 , \1624 );
nand \add_6_14_g19503/U$1 ( \2067 , \1903 , \1763 );
not \add_6_14_g19506/U$2 ( \2068 , \1740 );
nor \add_6_14_g19506/U$1 ( \2069 , \2068 , \1617 );
nand \add_6_14_g19508/U$1 ( \2070 , \1757 , \1760 );
not \add_6_14_g19515/U$2 ( \2071 , \1709 );
nor \add_6_14_g19515/U$1 ( \2072 , \2071 , \1699 );
nand \add_6_14_g19523/U$1 ( \2073 , \1939 , \1746 );
not \add_6_14_g19524/U$2 ( \2074 , \1659 );
nor \add_6_14_g19524/U$1 ( \2075 , \2074 , \1686 );
nor \add_6_14_g19526/U$1 ( \2076 , \1671 , \1716 );
not \add_6_14_g19537/U$2 ( \2077 , \1791 );
nand \add_6_14_g19537/U$1 ( \2078 , \2077 , \1800 );
not \add_6_14_g19545/U$2 ( \2079 , \1639 );
nor \add_6_14_g19545/U$1 ( \2080 , \2079 , \1665 );
not \add_6_14_g19547/U$2 ( \2081 , \1634 );
nor \add_6_14_g19547/U$1 ( \2082 , \2081 , \1653 );
not \add_6_14_g19551/U$2 ( \2083 , \1727 );
nor \add_6_14_g19551/U$1 ( \2084 , \2083 , \1724 );
nand \add_6_14_g19558/U$1 ( \2085 , \2041 , \1754 );
not \add_6_14_g19562/U$3 ( \2086 , \a[31] );
not \add_6_14_g19562/U$4 ( \2087 , \b[31] );
and \add_6_14_g19562/U$2 ( \2088 , \2086 , \2087 );
and \add_6_14_g19562/U$5 ( \2089 , \a[31] , \b[31] );
nor \add_6_14_g19562/U$1 ( \2090 , \2088 , \2089 );
or \add_6_14_g19678/U$2 ( \2091 , \1860 , \1859 );
nand \add_6_14_g19678/U$1 ( \2092 , \2091 , \1861 );
or \add_6_14_g19679/U$2 ( \2093 , \1850 , \1848 );
nand \add_6_14_g19679/U$1 ( \2094 , \2093 , \1851 );
xnor \add_6_14_g19682/U$1 ( \2095 , \1873 , \2059 );
xor \add_6_14_g19684/U$1 ( \2096 , \1958 , \2061 );
xnor \add_6_14_g19685/U$1 ( \2097 , \1963 , \2062 );
xnor \add_6_14_g19687/U$1 ( \2098 , \1902 , \2064 );
xor \add_6_14_g19688/U$1 ( \2099 , \1915 , \2066 );
xnor \add_6_14_g19689/U$1 ( \2100 , \1924 , \2067 );
xor \add_6_14_g19690/U$1 ( \2101 , \1844 , \2069 );
not \g45775/U$2 ( \2102 , \1732 );
nor \g45775/U$1 ( \2103 , \2102 , \1917 , \1621 );
or \g45774/U$1 ( \2104 , \2103 , \2045 );
xnor \add_6_14_g19691/U$1 ( \2105 , \2104 , \2070 );
xnor \add_6_14_g19694/U$1 ( \2106 , \1866 , \2073 );
xor \add_6_14_g19695/U$1 ( \2107 , \2012 , \2076 );
not \add_6_14_g19704/U$2 ( \2108 , \1745 );
nor \add_6_14_g19704/U$1 ( \2109 , \2108 , \1749 );
xor \add_6_14_g19697/U$1 ( \2110 , \1946 , \2109 );
xor \add_6_14_g19699/U$1 ( \2111 , \2036 , \2080 );
xor \add_6_14_g19700/U$1 ( \2112 , \2017 , \2082 );
xor \add_6_14_g19701/U$1 ( \2113 , \2028 , \2084 );
xnor \add_6_14_g19702/U$1 ( \2114 , \1929 , \2085 );
xor \add_6_14_g19703/U$1 ( \2115 , \1893 , \2090 );
not \mul_6_18_g44623/U$1 ( \2116 , \2058 );
not \mul_6_18_g44627/U$1 ( \2117 , \913 );
and \mul_6_18_g43892/U$2 ( \2118 , \2116 , \2117 );
not \mul_6_18_g43892/U$4 ( \2119 , \2116 );
and \mul_6_18_g43892/U$3 ( \2120 , \2119 , \913 );
nor \mul_6_18_g43892/U$1 ( \2121 , \2118 , \2120 );
not \mul_6_18_g43058/U$3 ( \2122 , \2121 );
not \mul_6_18_g44670/U$1 ( \2123 , \942 );
not \mul_6_18_g43865/U$3 ( \2124 , \2123 );
not \mul_6_18_g43865/U$4 ( \2125 , \980 );
or \mul_6_18_g43865/U$2 ( \2126 , \2124 , \2125 );
not \mul_6_18_g45249/U$2 ( \2127 , \980 );
nand \mul_6_18_g45249/U$1 ( \2128 , \2127 , \942 );
nand \mul_6_18_g43865/U$1 ( \2129 , \2126 , \2128 );
not \mul_6_18_g43739/U$3 ( \2130 , \2123 );
not \mul_6_18_g43739/U$4 ( \2131 , \2117 );
or \mul_6_18_g43739/U$2 ( \2132 , \2130 , \2131 );
nand \mul_6_18_g44160/U$1 ( \2133 , \913 , \942 );
nand \mul_6_18_g43739/U$1 ( \2134 , \2132 , \2133 );
nor \mul_6_18_g43701/U$1 ( \2135 , \2129 , \2134 );
not \mul_6_18_g43058/U$4 ( \2136 , \2135 );
or \mul_6_18_g43058/U$2 ( \2137 , \2122 , \2136 );
xor \mul_6_18_g45266/U$1 ( \2138 , \2056 , \913 );
nand \mul_6_18_g43584/U$1 ( \2139 , \2138 , \2129 );
nand \mul_6_18_g43058/U$1 ( \2140 , \2137 , \2139 );
and \g45858/U$2 ( \2141 , \2072 , \2046 );
not \g45858/U$4 ( \2142 , \2072 );
and \g45858/U$3 ( \2143 , \2142 , \1978 );
or \g45858/U$1 ( \2144 , \2141 , \2143 );
not \mul_6_18_g44571/U$1 ( \2145 , \2144 );
buf \mul_6_18_g44460/U$1 ( \2146 , \980 );
xnor \g45700/U$1 ( \2147 , \2145 , \2146 );
not \mul_6_18_g43066/U$3 ( \2148 , \2147 );
nand \g45626/U$1 ( \2149 , \1555 , \839 );
not \mul_6_18_g44406/U$1 ( \2150 , \1015 );
and \mul_6_18_g45268/U$2 ( \2151 , \2149 , \2150 );
not \mul_6_18_g45268/U$4 ( \2152 , \2149 );
and \mul_6_18_g45268/U$3 ( \2153 , \2152 , \1015 );
nor \mul_6_18_g45268/U$1 ( \2154 , \2151 , \2153 );
not \fopt45586/U$1 ( \2155 , \2154 );
and \g45625/U$1 ( \2156 , \1555 , \839 );
not \mul_6_18_g44668/U$1 ( \2157 , \2156 );
or \mul_6_18_g43734/U$2 ( \2158 , \2146 , \2157 );
not \mul_6_18_g44455/U$1 ( \2159 , \980 );
or \mul_6_18_g43734/U$3 ( \2160 , \2159 , \2156 );
nand \mul_6_18_g43734/U$1 ( \2161 , \2158 , \2160 );
nor \mul_6_18_g43698/U$1 ( \2162 , \2155 , \2161 );
not \mul_6_18_g43066/U$4 ( \2163 , \2162 );
or \mul_6_18_g43066/U$2 ( \2164 , \2148 , \2163 );
or \g45721/U$2 ( \2165 , \1703 , \1698 , \2048 );
or \g45723/U$2 ( \2166 , \1703 , \1698 );
nand \g45723/U$1 ( \2167 , \2166 , \2048 );
nand \g45721/U$1 ( \2168 , \2165 , \2167 );
and \g45614/U$2 ( \2169 , \2168 , \2159 );
not \g45614/U$4 ( \2170 , \2168 );
and \g45614/U$3 ( \2171 , \2170 , \2146 );
or \g45614/U$1 ( \2172 , \2169 , \2171 );
nand \mul_6_18_g43637/U$1 ( \2173 , \2172 , \2155 );
nand \mul_6_18_g43066/U$1 ( \2174 , \2164 , \2173 );
xor \mul_6_18_g42647/U$4 ( \2175 , \2140 , \2174 );
and \g45720/U$2 ( \2176 , \2075 , \2049 );
not \g45720/U$4 ( \2177 , \2075 );
and \g45720/U$3 ( \2178 , \2177 , \1984 );
or \g45720/U$1 ( \2179 , \2176 , \2178 );
not \mul_6_18_g44110/U$3 ( \2180 , \2179 );
buf \mul_6_18_g44413/U$1 ( \2181 , \1015 );
not \mul_6_18_g44412/U$1 ( \2182 , \2181 );
not \mul_6_18_g44110/U$4 ( \2183 , \2182 );
or \mul_6_18_g44110/U$2 ( \2184 , \2180 , \2183 );
not \mul_6_18_g44794/U$1 ( \2185 , \2179 );
nand \mul_6_18_g44277/U$1 ( \2186 , \2181 , \2185 );
nand \mul_6_18_g44110/U$1 ( \2187 , \2184 , \2186 );
not \mul_6_18_g43074/U$3 ( \2188 , \2187 );
nand \g45817/U$1 ( \2189 , \1572 , \839 );
not \mul_6_18_g44795/U$1 ( \2190 , \2189 );
and \g45773/U$2 ( \2191 , \2190 , \2150 );
not \g45773/U$4 ( \2192 , \2190 );
and \g45773/U$3 ( \2193 , \2192 , \1015 );
or \g45773/U$1 ( \2194 , \2191 , \2193 );
not \mul_6_18_g44793/U$1 ( \2195 , \1056 );
not \mul_6_18_g44789/U$1 ( \2196 , \2195 );
not \mul_6_18_g43842/U$3 ( \2197 , \2196 );
not \mul_6_18_g43842/U$4 ( \2198 , \2190 );
or \mul_6_18_g43842/U$2 ( \2199 , \2197 , \2198 );
nand \mul_6_18_g44187/U$1 ( \2200 , \2195 , \2189 );
nand \mul_6_18_g43842/U$1 ( \2201 , \2199 , \2200 );
nor \g45772/U$1 ( \2202 , \2194 , \2201 );
not \mul_6_18_g43074/U$4 ( \2203 , \2202 );
or \mul_6_18_g43074/U$2 ( \2204 , \2188 , \2203 );
and \mul_6_18_g44109/U$2 ( \2205 , \2006 , \2181 );
not \mul_6_18_g44109/U$4 ( \2206 , \2006 );
and \mul_6_18_g44109/U$3 ( \2207 , \2206 , \2182 );
nor \mul_6_18_g44109/U$1 ( \2208 , \2205 , \2207 );
not \mul_6_18_g43841/U$1 ( \2209 , \2201 );
not \mul_6_18_g43839/U$1 ( \2210 , \2209 );
nand \mul_6_18_g43453/U$1 ( \2211 , \2208 , \2210 );
nand \mul_6_18_g43074/U$1 ( \2212 , \2204 , \2211 );
and \mul_6_18_g42647/U$3 ( \2213 , \2175 , \2212 );
and \mul_6_18_g42647/U$5 ( \2214 , \2140 , \2174 );
or \mul_6_18_g42647/U$2 ( \2215 , \2213 , \2214 );
buf \mul_6_18_g44714/U$1 ( \2216 , \1531 );
not \mul_6_18_g44711/U$1 ( \2217 , \2216 );
xor \g45804/U$1 ( \2218 , \c[0] , \d[0] );
not \g45301/U$2 ( \2219 , \2218 );
nand \g45301/U$1 ( \2220 , \2219 , \838 );
nor \mul_6_18_g44394/U$1 ( \2221 , \2217 , \2220 );
buf \mul_6_18_g44393/U$1 ( \2222 , \2221 );
buf \mul_6_18_g44389/U$1 ( \2223 , \2222 );
not \mul_6_18_g44388/U$1 ( \2224 , \2223 );
buf \mul_6_18_g44691/U$1 ( \2225 , \1531 );
buf \mul_6_18_g44683/U$1 ( \2226 , \2225 );
and \mul_6_18_g43743/U$2 ( \2227 , \1807 , \2226 );
not \mul_6_18_g43743/U$4 ( \2228 , \1807 );
not \mul_6_18_g44682/U$1 ( \2229 , \2226 );
and \mul_6_18_g43743/U$3 ( \2230 , \2228 , \2229 );
nor \mul_6_18_g43743/U$1 ( \2231 , \2227 , \2230 );
not \mul_6_18_g43742/U$1 ( \2232 , \2231 );
or \mul_6_18_g43416/U$2 ( \2233 , \2224 , \2232 );
not \mul_6_18_g44475/U$1 ( \2234 , \2096 );
not \mul_6_18_g43741/U$3 ( \2235 , \2234 );
buf \mul_6_18_g44700/U$1 ( \2236 , \2216 );
not \mul_6_18_g43741/U$4 ( \2237 , \2236 );
or \mul_6_18_g43741/U$2 ( \2238 , \2235 , \2237 );
or \mul_6_18_g43741/U$5 ( \2239 , \2226 , \2234 );
nand \mul_6_18_g43741/U$1 ( \2240 , \2238 , \2239 );
not \mul_6_18_g43740/U$1 ( \2241 , \2240 );
not \mul_6_18_g44887/U$1 ( \2242 , \2220 );
buf \mul_6_18_g44886/U$1 ( \2243 , \2242 );
not \mul_6_18_g44883/U$1 ( \2244 , \2243 );
buf \mul_6_18_g44882/U$1 ( \2245 , \2244 );
not \mul_6_18_g44880/U$1 ( \2246 , \2245 );
or \mul_6_18_g43416/U$3 ( \2247 , \2241 , \2246 );
nand \mul_6_18_g43416/U$1 ( \2248 , \2233 , \2247 );
not \mul_6_18_g43875/U$3 ( \2249 , \2099 );
not \mul_6_18_g44962/U$1 ( \2250 , \1458 );
buf \mul_6_18_g44961/U$1 ( \2251 , \2250 );
not \mul_6_18_g44960/U$1 ( \2252 , \2251 );
not \mul_6_18_g44959/U$1 ( \2253 , \2252 );
not \mul_6_18_g43875/U$4 ( \2254 , \2253 );
or \mul_6_18_g43875/U$2 ( \2255 , \2249 , \2254 );
buf \mul_6_18_g44943/U$1 ( \2256 , \1458 );
not \mul_6_18_g44636/U$1 ( \2257 , \2099 );
nand \mul_6_18_g44205/U$1 ( \2258 , \2256 , \2257 );
nand \mul_6_18_g43875/U$1 ( \2259 , \2255 , \2258 );
not \mul_6_18_g43277/U$3 ( \2260 , \2259 );
nand \mul_6_18_g44176/U$1 ( \2261 , \1458 , \1476 );
not \mul_6_18_g43519/U$3 ( \2262 , \2261 );
not \fopt45607/U$1 ( \2263 , \1476 );
nand \mul_6_18_g44178/U$1 ( \2264 , \2250 , \2263 );
not \mul_6_18_g43519/U$4 ( \2265 , \2264 );
or \mul_6_18_g43519/U$2 ( \2266 , \2262 , \2265 );
and \mul_6_18_g43771/U$2 ( \2267 , \1499 , \1476 );
not \mul_6_18_g43771/U$4 ( \2268 , \1499 );
not \fopt45608/U$1 ( \2269 , \1476 );
and \mul_6_18_g43771/U$3 ( \2270 , \2268 , \2269 );
nor \mul_6_18_g43771/U$1 ( \2271 , \2267 , \2270 );
nand \mul_6_18_g43519/U$1 ( \2272 , \2266 , \2271 );
not \fopt45635/U$1 ( \2273 , \2272 );
buf \fopt45634/U$1 ( \2274 , \2273 );
not \mul_6_18_g43277/U$4 ( \2275 , \2274 );
or \mul_6_18_g43277/U$2 ( \2276 , \2260 , \2275 );
not \mul_6_18_g44942/U$1 ( \2277 , \2256 );
and \mul_6_18_g43861/U$2 ( \2278 , \2097 , \2277 );
not \mul_6_18_g43861/U$4 ( \2279 , \2097 );
not \mul_6_18_g44949/U$1 ( \2280 , \2251 );
and \mul_6_18_g43861/U$3 ( \2281 , \2279 , \2280 );
nor \mul_6_18_g43861/U$1 ( \2282 , \2278 , \2281 );
not \mul_6_18_g45234/U$2 ( \2283 , \2282 );
buf \mul_6_18_g43770/U$1 ( \2284 , \2271 );
not \mul_6_18_g43766/U$1 ( \2285 , \2284 );
nand \mul_6_18_g45234/U$1 ( \2286 , \2283 , \2285 );
nand \mul_6_18_g43277/U$1 ( \2287 , \2276 , \2286 );
xor \mul_6_18_g42650/U$1 ( \2288 , \2248 , \2287 );
not \mul_6_18_fopt45058/U$1 ( \2289 , \1353 );
and \mul_6_18_g43809/U$2 ( \2290 , \2289 , \1321 );
not \mul_6_18_g43809/U$4 ( \2291 , \2289 );
not \mul_6_18_g44398/U$1 ( \2292 , \1321 );
and \mul_6_18_g43809/U$3 ( \2293 , \2291 , \2292 );
nor \mul_6_18_g43809/U$1 ( \2294 , \2290 , \2293 );
not \mul_6_18_g44401/U$1 ( \2295 , \1321 );
not \mul_6_18_g44754/U$1 ( \2296 , \1298 );
and \mul_6_18_g43817/U$2 ( \2297 , \2295 , \2296 );
not \mul_6_18_g43817/U$4 ( \2298 , \2295 );
and \mul_6_18_g43817/U$3 ( \2299 , \2298 , \1298 );
nor \mul_6_18_g43817/U$1 ( \2300 , \2297 , \2299 );
nand \mul_6_18_g43463/U$1 ( \2301 , \2294 , \2300 );
not \mul_6_18_g43462/U$1 ( \2302 , \2301 );
buf \mul_6_18_g43461/U$1 ( \2303 , \2302 );
not \mul_6_18_g43458/U$1 ( \2304 , \2303 );
buf \mul_6_18_g44538/U$1 ( \2305 , \2113 );
not \mul_6_18_g43966/U$3 ( \2306 , \2305 );
buf \mul_6_18_g44752/U$1 ( \2307 , \1298 );
not \mul_6_18_g44768/U$1 ( \2308 , \2307 );
not \mul_6_18_g43966/U$4 ( \2309 , \2308 );
or \mul_6_18_g43966/U$2 ( \2310 , \2306 , \2309 );
buf \mul_6_18_g44761/U$1 ( \2311 , \2307 );
not \mul_6_18_g44537/U$1 ( \2312 , \2305 );
nand \mul_6_18_g44242/U$1 ( \2313 , \2311 , \2312 );
nand \mul_6_18_g43966/U$1 ( \2314 , \2310 , \2313 );
not \mul_6_18_g43965/U$1 ( \2315 , \2314 );
or \mul_6_18_g43171/U$2 ( \2316 , \2304 , \2315 );
not \mul_6_18_fopt45118/U$1 ( \2317 , \2294 );
buf \mul_6_18_fopt45117/U$1 ( \2318 , \2317 );
not \mul_6_18_fopt45114/U$1 ( \2319 , \2318 );
and \mul_6_18_g43942/U$2 ( \2320 , \2308 , \1970 );
not \mul_6_18_g44932/U$1 ( \2321 , \1970 );
and \mul_6_18_g43942/U$3 ( \2322 , \2307 , \2321 );
nor \mul_6_18_g43942/U$1 ( \2323 , \2320 , \2322 );
or \mul_6_18_g43171/U$3 ( \2324 , \2319 , \2323 );
nand \mul_6_18_g43171/U$1 ( \2325 , \2316 , \2324 );
xor \mul_6_18_g42650/U$1_r1 ( \2326 , \2288 , \2325 );
xor \mul_6_18_g42373/U$1 ( \2327 , \2215 , \2326 );
buf \mul_6_18_fopt45081/U$1 ( \2328 , \1353 );
buf \mul_6_18_fopt45074/U$1 ( \2329 , \2328 );
not \mul_6_18_fopt45073/U$1 ( \2330 , \2329 );
buf \mul_6_18_fopt45076/U$1 ( \2331 , \2330 );
not \mul_6_18_fopt45075/U$1 ( \2332 , \2331 );
and \mul_6_18_g43934/U$2 ( \2333 , \2101 , \2332 );
not \mul_6_18_g43934/U$4 ( \2334 , \2101 );
buf \mul_6_18_fopt45072/U$1 ( \2335 , \2329 );
not \mul_6_18_fopt45069/U$1 ( \2336 , \2335 );
and \mul_6_18_g43934/U$3 ( \2337 , \2334 , \2336 );
nor \mul_6_18_g43934/U$1 ( \2338 , \2333 , \2337 );
not \mul_6_18_g43174/U$3 ( \2339 , \2338 );
not \mul_6_18_fopt45057/U$1 ( \2340 , \1370 );
xor \g45495/U$1 ( \2341 , \2328 , \2340 );
not \mul_6_18_g43800/U$3 ( \2342 , \1396 );
not \mul_6_18_g43800/U$4 ( \2343 , \2340 );
or \mul_6_18_g43800/U$2 ( \2344 , \2342 , \2343 );
not \mul_6_18_g44545/U$1 ( \2345 , \1396 );
nand \mul_6_18_g44183/U$1 ( \2346 , \2345 , \1370 );
nand \mul_6_18_g43800/U$1 ( \2347 , \2344 , \2346 );
nor \mul_6_18_g43472/U$1 ( \2348 , \2341 , \2347 );
buf \mul_6_18_g43471/U$1 ( \2349 , \2348 );
not \mul_6_18_g43174/U$4 ( \2350 , \2349 );
or \mul_6_18_g43174/U$2 ( \2351 , \2339 , \2350 );
buf \mul_6_18_g44420/U$1 ( \2352 , \2106 );
and \mul_6_18_g43907/U$2 ( \2353 , \2336 , \2352 );
not \mul_6_18_g44419/U$1 ( \2354 , \2352 );
and \mul_6_18_g43907/U$3 ( \2355 , \2332 , \2354 );
nor \mul_6_18_g43907/U$1 ( \2356 , \2353 , \2355 );
not \mul_6_18_g43420/U$2 ( \2357 , \2356 );
buf \mul_6_18_fopt45134/U$1 ( \2358 , \2347 );
buf \mul_6_18_fopt45133/U$1 ( \2359 , \2358 );
nand \mul_6_18_g43420/U$1 ( \2360 , \2357 , \2359 );
nand \mul_6_18_g43174/U$1 ( \2361 , \2351 , \2360 );
not \mul_6_18_g43905/U$3 ( \2362 , \2110 );
buf \mul_6_18_g44558/U$1 ( \2363 , \1396 );
not \mul_6_18_g44547/U$1 ( \2364 , \2363 );
not \mul_6_18_g43905/U$4 ( \2365 , \2364 );
or \mul_6_18_g43905/U$2 ( \2366 , \2362 , \2365 );
not \mul_6_18_g44570/U$1 ( \2367 , \1396 );
not \mul_6_18_g44564/U$1 ( \2368 , \2367 );
not \mul_6_18_g44522/U$1 ( \2369 , \2110 );
nand \mul_6_18_g44225/U$1 ( \2370 , \2368 , \2369 );
nand \mul_6_18_g43905/U$1 ( \2371 , \2366 , \2370 );
not \mul_6_18_g43207/U$3 ( \2372 , \2371 );
not \sub_5_33_g9106/U$3 ( \2373 , \386 );
not \sub_5_33_g9106/U$4 ( \2374 , \1244 );
or \sub_5_33_g9106/U$2 ( \2375 , \2373 , \2374 );
nand \sub_5_33_g9106/U$1 ( \2376 , \2375 , \1416 );
nand \sub_5_33_g9312/U$1 ( \2377 , \384 , \449 );
xnor \sub_5_33_g9544/U$1 ( \2378 , \2376 , \2377 );
and \g45300/U$2 ( \2379 , \981 , \2378 );
not \g45300/U$4 ( \2380 , \981 );
and \g45300/U$3 ( \2381 , \2380 , \1600 );
nor \g45300/U$1 ( \2382 , \2379 , \2381 );
nand \g45299/U$1 ( \2383 , \2382 , \837 );
not \mul_6_18_g44835/U$1 ( \2384 , \2383 );
not \mul_6_18_g44834/U$1 ( \2385 , \2384 );
not \mul_6_18_g43794/U$3 ( \2386 , \2385 );
not \mul_6_18_g44891/U$1 ( \2387 , \1415 );
not \mul_6_18_g43794/U$4 ( \2388 , \2387 );
or \mul_6_18_g43794/U$2 ( \2389 , \2386 , \2388 );
nand \mul_6_18_g44181/U$1 ( \2390 , \2384 , \1415 );
nand \mul_6_18_g43794/U$1 ( \2391 , \2389 , \2390 );
not \mul_6_18_g43583/U$2 ( \2392 , \2391 );
not \mul_6_18_g43795/U$3 ( \2393 , \2387 );
not \mul_6_18_g43795/U$4 ( \2394 , \1396 );
or \mul_6_18_g43795/U$2 ( \2395 , \2393 , \2394 );
nand \mul_6_18_g44182/U$1 ( \2396 , \2345 , \1415 );
nand \mul_6_18_g43795/U$1 ( \2397 , \2395 , \2396 );
nand \mul_6_18_g43583/U$1 ( \2398 , \2392 , \2397 );
not \mul_6_18_g43582/U$1 ( \2399 , \2398 );
buf \mul_6_18_g43580/U$1 ( \2400 , \2399 );
not \mul_6_18_g43207/U$4 ( \2401 , \2400 );
or \mul_6_18_g43207/U$2 ( \2402 , \2372 , \2401 );
buf \mul_6_18_g43793/U$1 ( \2403 , \2391 );
not \mul_6_18_g44677/U$1 ( \2404 , \2114 );
not \mul_6_18_g44676/U$1 ( \2405 , \2404 );
xnor \g45617/U$1 ( \2406 , \2405 , \2364 );
nand \mul_6_18_g43423/U$1 ( \2407 , \2403 , \2406 );
nand \mul_6_18_g43207/U$1 ( \2408 , \2402 , \2407 );
xor \mul_6_18_g42522/U$1 ( \2409 , \2361 , \2408 );
not \mul_6_18_g43719/U$3 ( \2410 , \2116 );
not \mul_6_18_g43719/U$4 ( \2411 , \2123 );
or \mul_6_18_g43719/U$2 ( \2412 , \2410 , \2411 );
nand \mul_6_18_g43719/U$1 ( \2413 , \2412 , \2146 );
not \mul_6_18_g44632/U$1 ( \2414 , \2117 );
nand \mul_6_18_g44165/U$1 ( \2415 , \942 , \2058 );
and \mul_6_18_g43690/U$1 ( \2416 , \2413 , \2414 , \2415 );
buf \mul_6_18_g45008/U$1 ( \2417 , \1594 );
buf \mul_6_18_g45006/U$1 ( \2418 , \2417 );
not \mul_6_18_g45002/U$1 ( \2419 , \2418 );
and \mul_6_18_g43751/U$2 ( \2420 , \1784 , \2419 );
not \mul_6_18_g43751/U$4 ( \2421 , \1784 );
not \mul_6_18_g44991/U$1 ( \2422 , \1594 );
buf \mul_6_18_g44990/U$1 ( \2423 , \2422 );
not \mul_6_18_g44989/U$1 ( \2424 , \2423 );
and \mul_6_18_g43751/U$3 ( \2425 , \2421 , \2424 );
nor \mul_6_18_g43751/U$1 ( \2426 , \2420 , \2425 );
not \mul_6_18_g43750/U$1 ( \2427 , \2426 );
not \mul_6_18_g42925/U$3 ( \2428 , \2427 );
not \mul_6_18_g44530/U$1 ( \2429 , \1518 );
and \g45487/U$2 ( \2430 , \1531 , \2429 );
not \g45487/U$4 ( \2431 , \1531 );
and \g45487/U$3 ( \2432 , \2431 , \1518 );
or \g45487/U$1 ( \2433 , \2430 , \2432 );
buf \mul_6_18_g43397/U$1 ( \2434 , \2433 );
not \mul_6_18_g42925/U$4 ( \2435 , \2434 );
or \mul_6_18_g42925/U$2 ( \2436 , \2428 , \2435 );
and \mul_6_18_g43843/U$2 ( \2437 , \1531 , \2429 );
not \mul_6_18_g43843/U$4 ( \2438 , \1531 );
and \mul_6_18_g43843/U$3 ( \2439 , \2438 , \1518 );
nor \mul_6_18_g43843/U$1 ( \2440 , \2437 , \2439 );
not \mul_6_18_g43853/U$3 ( \2441 , \2429 );
not \mul_6_18_g43853/U$4 ( \2442 , \1594 );
or \mul_6_18_g43853/U$2 ( \2443 , \2441 , \2442 );
nand \mul_6_18_g44193/U$1 ( \2444 , \2422 , \1518 );
nand \mul_6_18_g43853/U$1 ( \2445 , \2443 , \2444 );
nand \mul_6_18_g45141/U$1 ( \2446 , \2440 , \2445 );
buf \mul_6_18_g43332/U$1 ( \2447 , \2446 );
not \mul_6_18_g43749/U$3 ( \2448 , \2095 );
not \mul_6_18_g43749/U$4 ( \2449 , \2423 );
or \mul_6_18_g43749/U$2 ( \2450 , \2448 , \2449 );
not \mul_6_18_g44773/U$1 ( \2451 , \2095 );
nand \mul_6_18_g44177/U$1 ( \2452 , \2424 , \2451 );
nand \mul_6_18_g43749/U$1 ( \2453 , \2450 , \2452 );
not \mul_6_18_g43748/U$1 ( \2454 , \2453 );
or \mul_6_18_g42925/U$5 ( \2455 , \2447 , \2454 );
nand \mul_6_18_g42925/U$1 ( \2456 , \2436 , \2455 );
and \mul_6_18_g42788/U$2 ( \2457 , \2416 , \2456 );
xor \mul_6_18_g42522/U$1_r1 ( \2458 , \2409 , \2457 );
xor \mul_6_18_g42373/U$1_r1 ( \2459 , \2327 , \2458 );
or \g45717/U$2 ( \2460 , \1681 , \1991 , \2040 );
or \g45728/U$2 ( \2461 , \1681 , \1991 );
nand \g45728/U$1 ( \2462 , \2461 , \2040 );
nand \g45717/U$1 ( \2463 , \2460 , \2462 );
not \mul_6_18_g44152/U$3 ( \2464 , \2463 );
not \mul_6_18_g44782/U$1 ( \2465 , \1056 );
not \mul_6_18_g44152/U$4 ( \2466 , \2465 );
or \mul_6_18_g44152/U$2 ( \2467 , \2464 , \2466 );
not \mul_6_18_g44473/U$1 ( \2468 , \2463 );
nand \mul_6_18_g44340/U$1 ( \2469 , \2196 , \2468 );
nand \mul_6_18_g44152/U$1 ( \2470 , \2467 , \2469 );
not \mul_6_18_g43076/U$3 ( \2471 , \2470 );
not \mul_6_18_g44446/U$1 ( \2472 , \1082 );
not \mul_6_18_g44445/U$1 ( \2473 , \2472 );
not \mul_6_18_g43737/U$3 ( \2474 , \2473 );
not \mul_6_18_g44779/U$1 ( \2475 , \2465 );
not \mul_6_18_g43737/U$4 ( \2476 , \2475 );
or \mul_6_18_g43737/U$2 ( \2477 , \2474 , \2476 );
nand \mul_6_18_g44159/U$1 ( \2478 , \2195 , \2472 );
nand \mul_6_18_g43737/U$1 ( \2479 , \2477 , \2478 );
xor \g45499/U$1 ( \2480 , \1109 , \1082 );
nor \mul_6_18_g43704/U$1 ( \2481 , \2479 , \2480 );
buf \mul_6_18_g43703/U$1 ( \2482 , \2481 );
not \mul_6_18_g43076/U$4 ( \2483 , \2482 );
or \mul_6_18_g43076/U$2 ( \2484 , \2471 , \2483 );
buf \mul_6_18_g43835/U$1 ( \2485 , \2480 );
not \mul_6_18_g44151/U$3 ( \2486 , \1998 );
not \mul_6_18_g44151/U$4 ( \2487 , \2465 );
or \mul_6_18_g44151/U$2 ( \2488 , \2486 , \2487 );
not \mul_6_18_g44836/U$1 ( \2489 , \1998 );
nand \mul_6_18_g44338/U$1 ( \2490 , \2475 , \2489 );
nand \mul_6_18_g44151/U$1 ( \2491 , \2488 , \2490 );
nand \mul_6_18_g43439/U$1 ( \2492 , \2485 , \2491 );
nand \mul_6_18_g43076/U$1 ( \2493 , \2484 , \2492 );
not \mul_6_18_g44071/U$3 ( \2494 , \2094 );
not \mul_6_18_fopt45101/U$1 ( \2495 , \1160 );
not \mul_6_18_fopt45098/U$1 ( \2496 , \2495 );
not \mul_6_18_fopt45096/U$1 ( \2497 , \2496 );
not \mul_6_18_g44071/U$4 ( \2498 , \2497 );
or \mul_6_18_g44071/U$2 ( \2499 , \2494 , \2498 );
not \mul_6_18_g44619/U$1 ( \2500 , \2094 );
nand \mul_6_18_g44280/U$1 ( \2501 , \2496 , \2500 );
nand \mul_6_18_g44071/U$1 ( \2502 , \2499 , \2501 );
not \mul_6_18_g43106/U$3 ( \2503 , \2502 );
xnor \mul_6_18_g45243/U$1 ( \2504 , \1218 , \1184 );
not \mul_6_18_g44404/U$1 ( \2505 , \1184 );
and \mul_6_18_g43738/U$2 ( \2506 , \2495 , \2505 );
and \mul_6_18_g43738/U$3 ( \2507 , \1184 , \1160 );
nor \mul_6_18_g43738/U$1 ( \2508 , \2506 , \2507 );
nand \mul_6_18_g43715/U$1 ( \2509 , \2504 , \2508 );
not \mul_6_18_g43714/U$1 ( \2510 , \2509 );
buf \mul_6_18_g43711/U$1 ( \2511 , \2510 );
not \mul_6_18_g43106/U$4 ( \2512 , \2511 );
or \mul_6_18_g43106/U$2 ( \2513 , \2503 , \2512 );
not \mul_6_18_g43823/U$1 ( \2514 , \2504 );
buf \mul_6_18_g43822/U$1 ( \2515 , \2514 );
and \mul_6_18_g44072/U$2 ( \2516 , \2111 , \2496 );
not \mul_6_18_g44072/U$4 ( \2517 , \2111 );
and \mul_6_18_g44072/U$3 ( \2518 , \2517 , \2497 );
nor \mul_6_18_g44072/U$1 ( \2519 , \2516 , \2518 );
nand \mul_6_18_g43430/U$1 ( \2520 , \2515 , \2519 );
nand \mul_6_18_g43106/U$1 ( \2521 , \2513 , \2520 );
xor \mul_6_18_g42574/U$1 ( \2522 , \2493 , \2521 );
xor \mul_6_18_g42788/U$1 ( \2523 , \2416 , \2456 );
xor \mul_6_18_g42574/U$1_r1 ( \2524 , \2522 , \2523 );
xor \g45611/U$1 ( \2525 , \2056 , \2146 );
not \mul_6_18_g43062/U$3 ( \2526 , \2525 );
buf \fopt45588/U$1 ( \2527 , \2162 );
not \mul_6_18_g43062/U$4 ( \2528 , \2527 );
or \mul_6_18_g43062/U$2 ( \2529 , \2526 , \2528 );
nand \mul_6_18_g43635/U$1 ( \2530 , \2147 , \2155 );
nand \mul_6_18_g43062/U$1 ( \2531 , \2529 , \2530 );
not \mul_6_18_g43720/U$3 ( \2532 , \2116 );
not \mul_6_18_g43720/U$4 ( \2533 , \2156 );
or \mul_6_18_g43720/U$2 ( \2534 , \2532 , \2533 );
nand \mul_6_18_g43720/U$1 ( \2535 , \2534 , \2181 );
not \mul_6_18_g45615/U$1 ( \2536 , \2159 );
nand \mul_6_18_g44167/U$1 ( \2537 , \2157 , \2058 );
nand \mul_6_18_g43689/U$1 ( \2538 , \2535 , \2536 , \2537 );
not \mul_6_18_g43688/U$1 ( \2539 , \2538 );
not \mul_6_18_g42756/U$3 ( \2540 , \2539 );
not \mul_6_18_g43746/U$3 ( \2541 , \2095 );
not \mul_6_18_g43746/U$4 ( \2542 , \2229 );
or \mul_6_18_g43746/U$2 ( \2543 , \2541 , \2542 );
nand \mul_6_18_g44188/U$1 ( \2544 , \2451 , \2216 );
nand \mul_6_18_g43746/U$1 ( \2545 , \2543 , \2544 );
not \mul_6_18_g43359/U$3 ( \2546 , \2545 );
not \mul_6_18_g43359/U$4 ( \2547 , \2223 );
or \mul_6_18_g43359/U$2 ( \2548 , \2546 , \2547 );
and \g45488/U$2 ( \2549 , \1784 , \2229 );
not \g45488/U$4 ( \2550 , \1784 );
and \g45488/U$3 ( \2551 , \2550 , \2225 );
or \g45488/U$1 ( \2552 , \2549 , \2551 );
nand \mul_6_18_g43487/U$1 ( \2553 , \2552 , \2245 );
nand \mul_6_18_g43359/U$1 ( \2554 , \2548 , \2553 );
not \mul_6_18_g42756/U$4 ( \2555 , \2554 );
or \mul_6_18_g42756/U$2 ( \2556 , \2540 , \2555 );
not \mul_6_18_g43885/U$3 ( \2557 , \2405 );
not \mul_6_18_g43885/U$4 ( \2558 , \2253 );
or \mul_6_18_g43885/U$2 ( \2559 , \2557 , \2558 );
nand \mul_6_18_g44210/U$1 ( \2560 , \2280 , \2404 );
nand \mul_6_18_g43885/U$1 ( \2561 , \2559 , \2560 );
not \mul_6_18_g43291/U$3 ( \2562 , \2561 );
not \mul_6_18_g43291/U$4 ( \2563 , \2274 );
or \mul_6_18_g43291/U$2 ( \2564 , \2562 , \2563 );
not \mul_6_18_g43886/U$3 ( \2565 , \2105 );
not \mul_6_18_g43886/U$4 ( \2566 , \2253 );
or \mul_6_18_g43886/U$2 ( \2567 , \2565 , \2566 );
not \mul_6_18_g44471/U$1 ( \2568 , \2105 );
nand \mul_6_18_g44208/U$1 ( \2569 , \2256 , \2568 );
nand \mul_6_18_g43886/U$1 ( \2570 , \2567 , \2569 );
nand \mul_6_18_g43627/U$1 ( \2571 , \2285 , \2570 );
nand \mul_6_18_g43291/U$1 ( \2572 , \2564 , \2571 );
not \mul_6_18_g43358/U$1 ( \2573 , \2554 );
nand \mul_6_18_g43017/U$1 ( \2574 , \2538 , \2573 );
nand \mul_6_18_g42798/U$1 ( \2575 , \2572 , \2574 );
nand \mul_6_18_g42756/U$1 ( \2576 , \2556 , \2575 );
xor \mul_6_18_g42417/U$4 ( \2577 , \2531 , \2576 );
and \mul_6_18_g43644/U$1 ( \2578 , \2129 , \2058 );
not \mul_6_18_g43850/U$3 ( \2579 , \2098 );
not \mul_6_18_g43850/U$4 ( \2580 , \2423 );
or \mul_6_18_g43850/U$2 ( \2581 , \2579 , \2580 );
not \mul_6_18_g44920/U$1 ( \2582 , \2098 );
nand \mul_6_18_g44196/U$1 ( \2583 , \2424 , \2582 );
nand \mul_6_18_g43850/U$1 ( \2584 , \2581 , \2583 );
not \mul_6_18_g42935/U$3 ( \2585 , \2584 );
not \mul_6_18_g43325/U$1 ( \2586 , \2447 );
not \mul_6_18_g42935/U$4 ( \2587 , \2586 );
or \mul_6_18_g42935/U$2 ( \2588 , \2585 , \2587 );
nand \mul_6_18_g43040/U$1 ( \2589 , \2434 , \2453 );
nand \mul_6_18_g42935/U$1 ( \2590 , \2588 , \2589 );
xor \mul_6_18_g42549/U$1 ( \2591 , \2578 , \2590 );
not \mul_6_18_g45007/U$1 ( \2592 , \2417 );
and \mul_6_18_g43852/U$2 ( \2593 , \1507 , \2592 );
not \mul_6_18_g43852/U$4 ( \2594 , \1507 );
and \mul_6_18_g43852/U$3 ( \2595 , \2594 , \2417 );
nor \mul_6_18_g43852/U$1 ( \2596 , \2593 , \2595 );
and \g45502/U$2 ( \2597 , \1499 , \1506 );
not \g45502/U$4 ( \2598 , \1499 );
and \g45502/U$3 ( \2599 , \2598 , \1507 );
or \g45502/U$1 ( \2600 , \2597 , \2599 );
nand \mul_6_18_g43350/U$1 ( \2601 , \2596 , \2600 );
buf \fopt45577/U$1 ( \2602 , \2601 );
not \fopt45570/U$1 ( \2603 , \2602 );
not \mul_6_18_g45223/U$3 ( \2604 , \2603 );
not \mul_6_18_g43874/U$3 ( \2605 , \2099 );
buf \mul_6_18_g44851/U$1 ( \2606 , \1499 );
not \mul_6_18_g44850/U$1 ( \2607 , \2606 );
not \mul_6_18_g43874/U$4 ( \2608 , \2607 );
or \mul_6_18_g43874/U$2 ( \2609 , \2605 , \2608 );
nand \mul_6_18_g44200/U$1 ( \2610 , \2606 , \2257 );
nand \mul_6_18_g43874/U$1 ( \2611 , \2609 , \2610 );
not \mul_6_18_g45223/U$4 ( \2612 , \2611 );
or \mul_6_18_g45223/U$2 ( \2613 , \2604 , \2612 );
not \mul_6_18_g44995/U$1 ( \2614 , \1594 );
not \mul_6_18_g43415/U$3 ( \2615 , \2614 );
not \mul_6_18_g43415/U$4 ( \2616 , \1507 );
or \mul_6_18_g43415/U$2 ( \2617 , \2615 , \2616 );
not \mul_6_18_g45289/U$2 ( \2618 , \2422 );
nand \mul_6_18_g45289/U$1 ( \2619 , \2618 , \1506 );
nand \mul_6_18_g43415/U$1 ( \2620 , \2617 , \2619 );
not \mul_6_18_g43414/U$1 ( \2621 , \2620 );
not \mul_6_18_g43412/U$1 ( \2622 , \2621 );
buf \mul_6_18_g43411/U$1 ( \2623 , \2622 );
not \mul_6_18_g43410/U$1 ( \2624 , \2623 );
not \mul_6_18_g44528/U$1 ( \2625 , \2097 );
buf \mul_6_18_g44866/U$1 ( \2626 , \1499 );
and \mul_6_18_g43858/U$2 ( \2627 , \2625 , \2626 );
not \mul_6_18_g43858/U$4 ( \2628 , \2625 );
not \mul_6_18_g44865/U$1 ( \2629 , \2626 );
and \mul_6_18_g43858/U$3 ( \2630 , \2628 , \2629 );
nor \mul_6_18_g43858/U$1 ( \2631 , \2627 , \2630 );
or \mul_6_18_g45223/U$5 ( \2632 , \2624 , \2631 );
nand \mul_6_18_g45223/U$1 ( \2633 , \2613 , \2632 );
xor \mul_6_18_g42549/U$1_r1 ( \2634 , \2591 , \2633 );
and \mul_6_18_g42417/U$3 ( \2635 , \2577 , \2634 );
and \mul_6_18_g42417/U$5 ( \2636 , \2531 , \2576 );
or \mul_6_18_g42417/U$2 ( \2637 , \2635 , \2636 );
xor \mul_6_18_g42199/U$4 ( \2638 , \2524 , \2637 );
not \mul_6_18_g44600/U$1 ( \2639 , \1838 );
not \mul_6_18_g44598/U$1 ( \2640 , \2639 );
not \mul_6_18_g43958/U$3 ( \2641 , \2640 );
not \mul_6_18_g43958/U$4 ( \2642 , \2336 );
or \mul_6_18_g43958/U$2 ( \2643 , \2641 , \2642 );
not \mul_6_18_fopt45064/U$1 ( \2644 , \2328 );
buf \mul_6_18_fopt45061/U$1 ( \2645 , \2644 );
not \mul_6_18_g45291/U$2 ( \2646 , \2645 );
nand \mul_6_18_g45291/U$1 ( \2647 , \2646 , \2639 );
nand \mul_6_18_g43958/U$1 ( \2648 , \2643 , \2647 );
not \mul_6_18_g43184/U$3 ( \2649 , \2648 );
not \mul_6_18_g43184/U$4 ( \2650 , \2349 );
or \mul_6_18_g43184/U$2 ( \2651 , \2649 , \2650 );
not \mul_6_18_g43957/U$3 ( \2652 , \2305 );
not \mul_6_18_g43957/U$4 ( \2653 , \2331 );
or \mul_6_18_g43957/U$2 ( \2654 , \2652 , \2653 );
nand \mul_6_18_g44246/U$1 ( \2655 , \2335 , \2312 );
nand \mul_6_18_g43957/U$1 ( \2656 , \2654 , \2655 );
nand \mul_6_18_g43421/U$1 ( \2657 , \2359 , \2656 );
nand \mul_6_18_g43184/U$1 ( \2658 , \2651 , \2657 );
not \g45794/U$3 ( \2659 , \2658 );
not \mul_6_18_g43925/U$3 ( \2660 , \1970 );
not \mul_6_18_g43925/U$4 ( \2661 , \2367 );
or \mul_6_18_g43925/U$2 ( \2662 , \2660 , \2661 );
buf \mul_6_18_g44551/U$1 ( \2663 , \2363 );
nand \mul_6_18_g44234/U$1 ( \2664 , \2663 , \2321 );
nand \mul_6_18_g43925/U$1 ( \2665 , \2662 , \2664 );
and \mul_6_18_g43216/U$2 ( \2666 , \2400 , \2665 );
not \mul_6_18_g43926/U$3 ( \2667 , \2101 );
not \mul_6_18_g43926/U$4 ( \2668 , \2367 );
or \mul_6_18_g43926/U$2 ( \2669 , \2667 , \2668 );
not \mul_6_18_g44578/U$1 ( \2670 , \2101 );
nand \mul_6_18_g44231/U$1 ( \2671 , \2368 , \2670 );
nand \mul_6_18_g43926/U$1 ( \2672 , \2669 , \2671 );
and \mul_6_18_g43216/U$3 ( \2673 , \2403 , \2672 );
nor \mul_6_18_g43216/U$1 ( \2674 , \2666 , \2673 );
not \mul_6_18_g43215/U$1 ( \2675 , \2674 );
not \g45794/U$4 ( \2676 , \2675 );
or \g45794/U$2 ( \2677 , \2659 , \2676 );
not \g45795/U$3 ( \2678 , \2674 );
not \mul_6_18_g43183/U$1 ( \2679 , \2658 );
not \g45795/U$4 ( \2680 , \2679 );
or \g45795/U$2 ( \2681 , \2678 , \2680 );
xor \g45497/U$1 ( \2682 , \1127 , \1160 );
not \mul_6_18_g43832/U$1 ( \2683 , \2682 );
buf \mul_6_18_g44443/U$1 ( \2684 , \1109 );
and \mul_6_18_g43735/U$2 ( \2685 , \1127 , \2684 );
not \mul_6_18_g43735/U$4 ( \2686 , \1127 );
not \mul_6_18_g44442/U$1 ( \2687 , \2684 );
and \mul_6_18_g43735/U$3 ( \2688 , \2686 , \2687 );
nor \mul_6_18_g43735/U$1 ( \2689 , \2685 , \2688 );
nand \mul_6_18_g43695/U$1 ( \2690 , \2683 , \2689 );
not \mul_6_18_g43694/U$1 ( \2691 , \2690 );
buf \mul_6_18_g43693/U$1 ( \2692 , \2691 );
not \mul_6_18_g44131/U$3 ( \2693 , \2463 );
not \mul_6_18_g44432/U$1 ( \2694 , \2684 );
not \mul_6_18_g44131/U$4 ( \2695 , \2694 );
or \mul_6_18_g44131/U$2 ( \2696 , \2693 , \2695 );
buf \mul_6_18_g44440/U$1 ( \2697 , \2684 );
nand \mul_6_18_g44320/U$1 ( \2698 , \2697 , \2468 );
nand \mul_6_18_g44131/U$1 ( \2699 , \2696 , \2698 );
and \mul_6_18_g43099/U$2 ( \2700 , \2692 , \2699 );
not \mul_6_18_g43831/U$1 ( \2701 , \2683 );
not \mul_6_18_g44133/U$3 ( \2702 , \1998 );
not \mul_6_18_g44133/U$4 ( \2703 , \2694 );
or \mul_6_18_g44133/U$2 ( \2704 , \2702 , \2703 );
not \mul_6_18_g44431/U$1 ( \2705 , \2694 );
nand \mul_6_18_g44317/U$1 ( \2706 , \2705 , \2489 );
nand \mul_6_18_g44133/U$1 ( \2707 , \2704 , \2706 );
and \mul_6_18_g43099/U$3 ( \2708 , \2701 , \2707 );
nor \mul_6_18_g43099/U$1 ( \2709 , \2700 , \2708 );
not \mul_6_18_g43097/U$1 ( \2710 , \2709 );
nand \g45795/U$1 ( \2711 , \2681 , \2710 );
nand \g45794/U$1 ( \2712 , \2677 , \2711 );
not \mul_6_18_g43903/U$3 ( \2713 , \2352 );
buf \mul_6_18_g44833/U$1 ( \2714 , \2385 );
not \mul_6_18_g44826/U$1 ( \2715 , \2714 );
not \mul_6_18_g43903/U$4 ( \2716 , \2715 );
or \mul_6_18_g43903/U$2 ( \2717 , \2713 , \2716 );
buf \mul_6_18_g44813/U$1 ( \2718 , \2384 );
not \mul_6_18_g44808/U$1 ( \2719 , \2718 );
nand \mul_6_18_g44222/U$1 ( \2720 , \2719 , \2354 );
nand \mul_6_18_g43903/U$1 ( \2721 , \2717 , \2720 );
not \mul_6_18_g43261/U$3 ( \2722 , \2721 );
xor \g45494/U$1 ( \2723 , \1458 , \1434 );
and \mul_6_18_g43785/U$2 ( \2724 , \1434 , \2384 );
not \mul_6_18_g43785/U$4 ( \2725 , \1434 );
and \mul_6_18_g43785/U$3 ( \2726 , \2725 , \2385 );
nor \mul_6_18_g43785/U$1 ( \2727 , \2724 , \2726 );
nor \mul_6_18_g43599/U$1 ( \2728 , \2723 , \2727 );
buf \mul_6_18_g43589/U$1 ( \2729 , \2728 );
not \mul_6_18_g43261/U$4 ( \2730 , \2729 );
or \mul_6_18_g43261/U$2 ( \2731 , \2722 , \2730 );
not \mul_6_18_g43783/U$1 ( \2732 , \2723 );
not \mul_6_18_g43774/U$1 ( \2733 , \2732 );
not \mul_6_18_g43902/U$3 ( \2734 , \2110 );
not \mul_6_18_g43902/U$4 ( \2735 , \2715 );
or \mul_6_18_g43902/U$2 ( \2736 , \2734 , \2735 );
nand \mul_6_18_g44227/U$1 ( \2737 , \2714 , \2369 );
nand \mul_6_18_g43902/U$1 ( \2738 , \2736 , \2737 );
nand \mul_6_18_g43555/U$1 ( \2739 , \2733 , \2738 );
nand \mul_6_18_g43261/U$1 ( \2740 , \2731 , \2739 );
not \mul_6_18_g43994/U$3 ( \2741 , \2107 );
not \mul_6_18_g44759/U$1 ( \2742 , \2311 );
not \mul_6_18_g43994/U$4 ( \2743 , \2742 );
or \mul_6_18_g43994/U$2 ( \2744 , \2741 , \2743 );
not \mul_6_18_g44589/U$1 ( \2745 , \2107 );
nand \mul_6_18_g44262/U$1 ( \2746 , \2311 , \2745 );
nand \mul_6_18_g43994/U$1 ( \2747 , \2744 , \2746 );
not \mul_6_18_g43163/U$3 ( \2748 , \2747 );
not \mul_6_18_g43163/U$4 ( \2749 , \2303 );
or \mul_6_18_g43163/U$2 ( \2750 , \2748 , \2749 );
not \mul_6_18_g43995/U$3 ( \2751 , \2092 );
not \mul_6_18_g43995/U$4 ( \2752 , \2742 );
or \mul_6_18_g43995/U$2 ( \2753 , \2751 , \2752 );
not \mul_6_18_g44772/U$1 ( \2754 , \2092 );
nand \mul_6_18_g44264/U$1 ( \2755 , \2311 , \2754 );
nand \mul_6_18_g43995/U$1 ( \2756 , \2753 , \2755 );
nand \mul_6_18_g43521/U$1 ( \2757 , \2318 , \2756 );
nand \mul_6_18_g43163/U$1 ( \2758 , \2750 , \2757 );
xor \mul_6_18_g42718/U$4 ( \2759 , \2740 , \2758 );
not \mul_6_18_g44052/U$3 ( \2760 , \2094 );
buf \mul_6_18_g44503/U$1 ( \2761 , \1218 );
not \mul_6_18_g44497/U$1 ( \2762 , \2761 );
not \mul_6_18_g44052/U$4 ( \2763 , \2762 );
or \mul_6_18_g44052/U$2 ( \2764 , \2760 , \2763 );
not \mul_6_18_g44495/U$1 ( \2765 , \2762 );
nand \mul_6_18_g44279/U$1 ( \2766 , \2765 , \2500 );
nand \mul_6_18_g44052/U$1 ( \2767 , \2764 , \2766 );
not \mul_6_18_g43144/U$3 ( \2768 , \2767 );
xor \g45496/U$1 ( \2769 , \1229 , \1218 );
xnor \mul_6_18_g45275/U$1 ( \2770 , \1298 , \1229 );
and \mul_6_18_g43621/U$1 ( \2771 , \2769 , \2770 );
not \mul_6_18_g43620/U$1 ( \2772 , \2771 );
not \mul_6_18_g43619/U$1 ( \2773 , \2772 );
not \mul_6_18_g43144/U$4 ( \2774 , \2773 );
or \mul_6_18_g43144/U$2 ( \2775 , \2768 , \2774 );
not \mul_6_18_g44053/U$3 ( \2776 , \2111 );
not \mul_6_18_g44053/U$4 ( \2777 , \2762 );
or \mul_6_18_g44053/U$2 ( \2778 , \2776 , \2777 );
not \mul_6_18_g44924/U$1 ( \2779 , \2111 );
nand \mul_6_18_g44289/U$1 ( \2780 , \2765 , \2779 );
nand \mul_6_18_g44053/U$1 ( \2781 , \2778 , \2780 );
buf \mul_6_18_g43815/U$1 ( \2782 , \2770 );
not \mul_6_18_g43811/U$1 ( \2783 , \2782 );
buf \mul_6_18_g43810/U$1 ( \2784 , \2783 );
nand \mul_6_18_g43568/U$1 ( \2785 , \2781 , \2784 );
nand \mul_6_18_g43144/U$1 ( \2786 , \2775 , \2785 );
and \mul_6_18_g42718/U$3 ( \2787 , \2759 , \2786 );
and \mul_6_18_g42718/U$5 ( \2788 , \2740 , \2758 );
or \mul_6_18_g42718/U$2 ( \2789 , \2787 , \2788 );
xor \mul_6_18_g42422/U$4 ( \2790 , \2712 , \2789 );
not \mul_6_18_g43079/U$3 ( \2791 , \2485 );
not \mul_6_18_g44144/U$3 ( \2792 , \2006 );
not \mul_6_18_g44144/U$4 ( \2793 , \2195 );
or \mul_6_18_g44144/U$2 ( \2794 , \2792 , \2793 );
not \mul_6_18_g44901/U$1 ( \2795 , \2006 );
nand \mul_6_18_g44321/U$1 ( \2796 , \2196 , \2795 );
nand \mul_6_18_g44144/U$1 ( \2797 , \2794 , \2796 );
not \mul_6_18_g43079/U$4 ( \2798 , \2797 );
or \mul_6_18_g43079/U$2 ( \2799 , \2791 , \2798 );
not \mul_6_18_g44143/U$3 ( \2800 , \2179 );
not \mul_6_18_g44143/U$4 ( \2801 , \2465 );
or \mul_6_18_g44143/U$2 ( \2802 , \2800 , \2801 );
nand \mul_6_18_g44327/U$1 ( \2803 , \2475 , \2185 );
nand \mul_6_18_g44143/U$1 ( \2804 , \2802 , \2803 );
nand \mul_6_18_g43316/U$1 ( \2805 , \2481 , \2804 );
nand \mul_6_18_g43079/U$1 ( \2806 , \2799 , \2805 );
not \mul_6_18_g43078/U$1 ( \2807 , \2806 );
not \mul_6_18_g42676/U$3 ( \2808 , \2807 );
and \g45338/U$1 ( \2809 , \2013 , \1632 );
xor \g45337/U$1 ( \2810 , \2809 , \1825 );
not \mul_6_18_g44913/U$1 ( \2811 , \2810 );
not \mul_6_18_g44910/U$1 ( \2812 , \2811 );
not \mul_6_18_g44098/U$3 ( \2813 , \2812 );
not \mul_6_18_g44098/U$4 ( \2814 , \2497 );
or \mul_6_18_g44098/U$2 ( \2815 , \2813 , \2814 );
not \mul_6_18_fopt45107/U$1 ( \2816 , \1160 );
not \mul_6_18_fopt45103/U$1 ( \2817 , \2816 );
nand \mul_6_18_g44298/U$1 ( \2818 , \2817 , \2811 );
nand \mul_6_18_g44098/U$1 ( \2819 , \2815 , \2818 );
and \mul_6_18_g43122/U$2 ( \2820 , \2511 , \2819 );
not \mul_6_18_g44097/U$3 ( \2821 , \2112 );
not \mul_6_18_g44097/U$4 ( \2822 , \2497 );
or \mul_6_18_g44097/U$2 ( \2823 , \2821 , \2822 );
not \mul_6_18_g44479/U$1 ( \2824 , \2112 );
nand \mul_6_18_g44294/U$1 ( \2825 , \2817 , \2824 );
nand \mul_6_18_g44097/U$1 ( \2826 , \2823 , \2825 );
and \mul_6_18_g43122/U$3 ( \2827 , \2515 , \2826 );
nor \mul_6_18_g43122/U$1 ( \2828 , \2820 , \2827 );
not \mul_6_18_g42676/U$4 ( \2829 , \2828 );
or \mul_6_18_g42676/U$2 ( \2830 , \2808 , \2829 );
not \mul_6_18_g44899/U$1 ( \2831 , \2100 );
not \mul_6_18_g44896/U$1 ( \2832 , \2831 );
not \mul_6_18_g43872/U$3 ( \2833 , \2832 );
not \mul_6_18_g44848/U$1 ( \2834 , \2606 );
not \mul_6_18_g43872/U$4 ( \2835 , \2834 );
or \mul_6_18_g43872/U$2 ( \2836 , \2833 , \2835 );
nand \mul_6_18_g44201/U$1 ( \2837 , \2626 , \2831 );
nand \mul_6_18_g43872/U$1 ( \2838 , \2836 , \2837 );
not \mul_6_18_g42966/U$3 ( \2839 , \2838 );
not \mul_6_18_g42966/U$4 ( \2840 , \2603 );
or \mul_6_18_g42966/U$2 ( \2841 , \2839 , \2840 );
buf \mul_6_18_g43408/U$1 ( \2842 , \2620 );
nand \mul_6_18_g43010/U$1 ( \2843 , \2842 , \2611 );
nand \mul_6_18_g42966/U$1 ( \2844 , \2841 , \2843 );
not \mul_6_18_g43851/U$3 ( \2845 , \2097 );
not \mul_6_18_g43851/U$4 ( \2846 , \2423 );
or \mul_6_18_g43851/U$2 ( \2847 , \2845 , \2846 );
not \mul_6_18_g44997/U$1 ( \2848 , \2419 );
nand \mul_6_18_g44191/U$1 ( \2849 , \2848 , \2625 );
nand \mul_6_18_g43851/U$1 ( \2850 , \2847 , \2849 );
not \mul_6_18_g42961/U$3 ( \2851 , \2850 );
not \mul_6_18_g42961/U$4 ( \2852 , \2586 );
or \mul_6_18_g42961/U$2 ( \2853 , \2851 , \2852 );
nand \mul_6_18_g43048/U$1 ( \2854 , \2434 , \2584 );
nand \mul_6_18_g42961/U$1 ( \2855 , \2853 , \2854 );
xnor \g45479/U$1 ( \2856 , \2844 , \2855 );
not \mul_6_18_g42777/U$1 ( \2857 , \2856 );
nand \mul_6_18_g42676/U$1 ( \2858 , \2830 , \2857 );
not \mul_6_18_g45214/U$2 ( \2859 , \2828 );
nand \mul_6_18_g45214/U$1 ( \2860 , \2859 , \2806 );
nand \mul_6_18_g42605/U$1 ( \2861 , \2858 , \2860 );
and \mul_6_18_g42422/U$3 ( \2862 , \2790 , \2861 );
and \mul_6_18_g42422/U$5 ( \2863 , \2712 , \2789 );
or \mul_6_18_g42422/U$2 ( \2864 , \2862 , \2863 );
and \mul_6_18_g42199/U$3 ( \2865 , \2638 , \2864 );
and \mul_6_18_g42199/U$5 ( \2866 , \2524 , \2637 );
or \mul_6_18_g42199/U$2 ( \2867 , \2865 , \2866 );
xor \mul_6_18_g42068/U$1 ( \2868 , \2459 , \2867 );
not \fopt45587/U$1 ( \2869 , \2527 );
not \mul_6_18_g44014/U$1 ( \2870 , \2172 );
or \mul_6_18_g43061/U$2 ( \2871 , \2869 , \2870 );
and \mul_6_18_g44039/U$2 ( \2872 , \2179 , \2159 );
not \mul_6_18_g44039/U$4 ( \2873 , \2179 );
and \mul_6_18_g44039/U$3 ( \2874 , \2873 , \2146 );
nor \mul_6_18_g44039/U$1 ( \2875 , \2872 , \2874 );
or \mul_6_18_g43061/U$3 ( \2876 , \2875 , \2154 );
nand \mul_6_18_g43061/U$1 ( \2877 , \2871 , \2876 );
not \mul_6_18_g43057/U$3 ( \2878 , \2138 );
buf \mul_6_18_g43700/U$1 ( \2879 , \2135 );
not \mul_6_18_g43057/U$4 ( \2880 , \2879 );
or \mul_6_18_g43057/U$2 ( \2881 , \2878 , \2880 );
not \mul_6_18_g43944/U$3 ( \2882 , \2144 );
not \mul_6_18_g43944/U$4 ( \2883 , \2117 );
or \mul_6_18_g43944/U$2 ( \2884 , \2882 , \2883 );
nand \mul_6_18_g44226/U$1 ( \2885 , \2414 , \2145 );
nand \mul_6_18_g43944/U$1 ( \2886 , \2884 , \2885 );
nand \mul_6_18_g43443/U$1 ( \2887 , \2886 , \2129 );
nand \mul_6_18_g43057/U$1 ( \2888 , \2881 , \2887 );
xor \mul_6_18_g42450/U$1 ( \2889 , \2877 , \2888 );
xnor \g45334/U$1 ( \2890 , \2078 , \1938 );
and \g45754/U$2 ( \2891 , \2890 , \2423 );
not \g45754/U$4 ( \2892 , \2890 );
and \g45754/U$3 ( \2893 , \2892 , \2848 );
or \g45754/U$1 ( \2894 , \2891 , \2893 );
not \mul_6_18_g43002/U$3 ( \2895 , \2894 );
not \mul_6_18_g43002/U$4 ( \2896 , \2434 );
or \mul_6_18_g43002/U$2 ( \2897 , \2895 , \2896 );
or \mul_6_18_g43002/U$5 ( \2898 , \2447 , \2426 );
nand \mul_6_18_g43002/U$1 ( \2899 , \2897 , \2898 );
and \g45755/U$2 ( \2900 , \2117 , \875 );
not \g45755/U$4 ( \2901 , \2117 );
not \mul_6_18_g44544/U$1 ( \2902 , \875 );
and \g45755/U$3 ( \2903 , \2901 , \2902 );
or \g45755/U$1 ( \2904 , \2900 , \2903 );
and \mul_6_18_g43450/U$1 ( \2905 , \2904 , \2058 );
xor \mul_6_18_g42583/U$1 ( \2906 , \2899 , \2905 );
not \fopt45576/U$1 ( \2907 , \2602 );
not \fopt45573/U$1 ( \2908 , \2907 );
not \mul_6_18_g44854/U$1 ( \2909 , \2626 );
and \mul_6_18_g43855/U$2 ( \2910 , \2098 , \2909 );
not \mul_6_18_g43855/U$4 ( \2911 , \2098 );
and \mul_6_18_g43855/U$3 ( \2912 , \2911 , \2606 );
nor \mul_6_18_g43855/U$1 ( \2913 , \2910 , \2912 );
or \mul_6_18_g42965/U$2 ( \2914 , \2908 , \2913 );
and \mul_6_18_g43755/U$2 ( \2915 , \2095 , \2834 );
and \mul_6_18_g43755/U$3 ( \2916 , \2626 , \2451 );
nor \mul_6_18_g43755/U$1 ( \2917 , \2915 , \2916 );
or \mul_6_18_g42965/U$3 ( \2918 , \2624 , \2917 );
nand \mul_6_18_g42965/U$1 ( \2919 , \2914 , \2918 );
xor \mul_6_18_g42583/U$1_r1 ( \2920 , \2906 , \2919 );
xor \mul_6_18_g42450/U$1_r1 ( \2921 , \2889 , \2920 );
xor \mul_6_18_g42549/U$4 ( \2922 , \2578 , \2590 );
and \mul_6_18_g42549/U$3 ( \2923 , \2922 , \2633 );
and \mul_6_18_g42549/U$5 ( \2924 , \2578 , \2590 );
or \mul_6_18_g42549/U$2 ( \2925 , \2923 , \2924 );
not \mul_6_18_g43419/U$3 ( \2926 , \2222 );
not \mul_6_18_g43419/U$4 ( \2927 , \2552 );
or \mul_6_18_g43419/U$2 ( \2928 , \2926 , \2927 );
not \mul_6_18_g44699/U$1 ( \2929 , \2236 );
and \g45489/U$2 ( \2930 , \2890 , \2929 );
not \g45489/U$4 ( \2931 , \2890 );
and \g45489/U$3 ( \2932 , \2931 , \2226 );
or \g45489/U$1 ( \2933 , \2930 , \2932 );
not \mul_6_18_g44871/U$1 ( \2934 , \2243 );
nand \mul_6_18_g43654/U$1 ( \2935 , \2933 , \2934 );
nand \mul_6_18_g43419/U$1 ( \2936 , \2928 , \2935 );
not \mul_6_18_g43282/U$3 ( \2937 , \2570 );
not \fopt45631/U$1 ( \2938 , \2272 );
not \mul_6_18_g43282/U$4 ( \2939 , \2938 );
or \mul_6_18_g43282/U$2 ( \2940 , \2937 , \2939 );
not \mul_6_18_g43876/U$3 ( \2941 , \2832 );
not \mul_6_18_g43876/U$4 ( \2942 , \2251 );
or \mul_6_18_g43876/U$2 ( \2943 , \2941 , \2942 );
nand \mul_6_18_g44202/U$1 ( \2944 , \2256 , \2831 );
nand \mul_6_18_g43876/U$1 ( \2945 , \2943 , \2944 );
nand \mul_6_18_g43422/U$1 ( \2946 , \2285 , \2945 );
nand \mul_6_18_g43282/U$1 ( \2947 , \2940 , \2946 );
xor \mul_6_18_g42629/U$4 ( \2948 , \2936 , \2947 );
not \mul_6_18_g43170/U$3 ( \2949 , \2756 );
not \mul_6_18_g43170/U$4 ( \2950 , \2303 );
or \mul_6_18_g43170/U$2 ( \2951 , \2949 , \2950 );
not \mul_6_18_g43964/U$3 ( \2952 , \2640 );
not \mul_6_18_g43964/U$4 ( \2953 , \2308 );
or \mul_6_18_g43964/U$2 ( \2954 , \2952 , \2953 );
nand \mul_6_18_g44245/U$1 ( \2955 , \2311 , \2639 );
nand \mul_6_18_g43964/U$1 ( \2956 , \2954 , \2955 );
nand \mul_6_18_g43425/U$1 ( \2957 , \2318 , \2956 );
nand \mul_6_18_g43170/U$1 ( \2958 , \2951 , \2957 );
and \mul_6_18_g42629/U$3 ( \2959 , \2948 , \2958 );
and \mul_6_18_g42629/U$5 ( \2960 , \2936 , \2947 );
or \mul_6_18_g42629/U$2 ( \2961 , \2959 , \2960 );
xor \mul_6_18_g42360/U$4 ( \2962 , \2925 , \2961 );
not \mul_6_18_g43260/U$3 ( \2963 , \2738 );
not \mul_6_18_g43598/U$1 ( \2964 , \2728 );
not \mul_6_18_g43597/U$1 ( \2965 , \2964 );
not \mul_6_18_g43260/U$4 ( \2966 , \2965 );
or \mul_6_18_g43260/U$2 ( \2967 , \2963 , \2966 );
not \mul_6_18_g43888/U$3 ( \2968 , \2405 );
buf \mul_6_18_g44825/U$1 ( \2969 , \2715 );
not \mul_6_18_g43888/U$4 ( \2970 , \2969 );
or \mul_6_18_g43888/U$2 ( \2971 , \2968 , \2970 );
not \mul_6_18_g44803/U$1 ( \2972 , \2718 );
nand \mul_6_18_g44209/U$1 ( \2973 , \2972 , \2404 );
nand \mul_6_18_g43888/U$1 ( \2974 , \2971 , \2973 );
nand \mul_6_18_g43446/U$1 ( \2975 , \2733 , \2974 );
nand \mul_6_18_g43260/U$1 ( \2976 , \2967 , \2975 );
not \mul_6_18_g43140/U$3 ( \2977 , \2781 );
not \mul_6_18_g43140/U$4 ( \2978 , \2773 );
or \mul_6_18_g43140/U$2 ( \2979 , \2977 , \2978 );
not \mul_6_18_g44010/U$3 ( \2980 , \2107 );
not \mul_6_18_g44010/U$4 ( \2981 , \2762 );
or \mul_6_18_g44010/U$2 ( \2982 , \2980 , \2981 );
nand \mul_6_18_g44260/U$1 ( \2983 , \2765 , \2745 );
nand \mul_6_18_g44010/U$1 ( \2984 , \2982 , \2983 );
nand \mul_6_18_g43636/U$1 ( \2985 , \2984 , \2784 );
nand \mul_6_18_g43140/U$1 ( \2986 , \2979 , \2985 );
xor \mul_6_18_g42725/U$4 ( \2987 , \2976 , \2986 );
not \mul_6_18_g43095/U$3 ( \2988 , \2707 );
not \mul_6_18_g43095/U$4 ( \2989 , \2692 );
or \mul_6_18_g43095/U$2 ( \2990 , \2988 , \2989 );
and \mul_6_18_g44119/U$2 ( \2991 , \2812 , \2697 );
not \mul_6_18_g44119/U$4 ( \2992 , \2812 );
not \mul_6_18_g44439/U$1 ( \2993 , \2697 );
and \mul_6_18_g44119/U$3 ( \2994 , \2992 , \2993 );
nor \mul_6_18_g44119/U$1 ( \2995 , \2991 , \2994 );
nand \mul_6_18_g43428/U$1 ( \2996 , \2701 , \2995 );
nand \mul_6_18_g43095/U$1 ( \2997 , \2990 , \2996 );
and \mul_6_18_g42725/U$3 ( \2998 , \2987 , \2997 );
and \mul_6_18_g42725/U$5 ( \2999 , \2976 , \2986 );
or \mul_6_18_g42725/U$2 ( \3000 , \2998 , \2999 );
and \mul_6_18_g42360/U$3 ( \3001 , \2962 , \3000 );
and \mul_6_18_g42360/U$5 ( \3002 , \2925 , \2961 );
or \mul_6_18_g42360/U$2 ( \3003 , \3001 , \3002 );
xor \mul_6_18_g42202/U$1 ( \3004 , \2921 , \3003 );
not \mul_6_18_g43418/U$3 ( \3005 , \2933 );
not \mul_6_18_g43418/U$4 ( \3006 , \2223 );
or \mul_6_18_g43418/U$2 ( \3007 , \3005 , \3006 );
nand \mul_6_18_g43650/U$1 ( \3008 , \2231 , \2245 );
nand \mul_6_18_g43418/U$1 ( \3009 , \3007 , \3008 );
not \mul_6_18_g42656/U$3 ( \3010 , \3009 );
not \mul_6_18_g43857/U$1 ( \3011 , \2631 );
not \mul_6_18_g42989/U$3 ( \3012 , \3011 );
not \fopt45572/U$1 ( \3013 , \2908 );
not \mul_6_18_g42989/U$4 ( \3014 , \3013 );
or \mul_6_18_g42989/U$2 ( \3015 , \3012 , \3014 );
not \mul_6_18_g45233/U$2 ( \3016 , \2913 );
nand \mul_6_18_g45233/U$1 ( \3017 , \3016 , \2842 );
nand \mul_6_18_g42989/U$1 ( \3018 , \3015 , \3017 );
not \mul_6_18_g42656/U$4 ( \3019 , \3018 );
or \mul_6_18_g42656/U$2 ( \3020 , \3010 , \3019 );
or \mul_6_18_g42684/U$2 ( \3021 , \3018 , \3009 );
not \mul_6_18_g43306/U$3 ( \3022 , \2945 );
not \mul_6_18_g43306/U$4 ( \3023 , \2274 );
or \mul_6_18_g43306/U$2 ( \3024 , \3022 , \3023 );
nand \mul_6_18_g43570/U$1 ( \3025 , \2285 , \2259 );
nand \mul_6_18_g43306/U$1 ( \3026 , \3024 , \3025 );
nand \mul_6_18_g42684/U$1 ( \3027 , \3021 , \3026 );
nand \mul_6_18_g42656/U$1 ( \3028 , \3020 , \3027 );
not \mul_6_18_g43904/U$3 ( \3029 , \2352 );
not \mul_6_18_g43904/U$4 ( \3030 , \2367 );
or \mul_6_18_g43904/U$2 ( \3031 , \3029 , \3030 );
nand \mul_6_18_g44218/U$1 ( \3032 , \2368 , \2354 );
nand \mul_6_18_g43904/U$1 ( \3033 , \3031 , \3032 );
not \mul_6_18_g43238/U$3 ( \3034 , \3033 );
not \mul_6_18_g43238/U$4 ( \3035 , \2400 );
or \mul_6_18_g43238/U$2 ( \3036 , \3034 , \3035 );
nand \mul_6_18_g43610/U$1 ( \3037 , \2403 , \2371 );
nand \mul_6_18_g43238/U$1 ( \3038 , \3036 , \3037 );
not \mul_6_18_g43933/U$3 ( \3039 , \1970 );
not \mul_6_18_g43933/U$4 ( \3040 , \2331 );
or \mul_6_18_g43933/U$2 ( \3041 , \3039 , \3040 );
nand \mul_6_18_g44233/U$1 ( \3042 , \2335 , \2321 );
nand \mul_6_18_g43933/U$1 ( \3043 , \3041 , \3042 );
not \mul_6_18_g43193/U$3 ( \3044 , \3043 );
not \mul_6_18_g43193/U$4 ( \3045 , \2349 );
or \mul_6_18_g43193/U$2 ( \3046 , \3044 , \3045 );
nand \mul_6_18_g43544/U$1 ( \3047 , \2359 , \2338 );
nand \mul_6_18_g43193/U$1 ( \3048 , \3046 , \3047 );
xor \mul_6_18_g42731/U$4 ( \3049 , \3038 , \3048 );
not \mul_6_18_g43096/U$3 ( \3050 , \2692 );
not \mul_6_18_g43096/U$4 ( \3051 , \2995 );
or \mul_6_18_g43096/U$2 ( \3052 , \3050 , \3051 );
and \mul_6_18_g44118/U$2 ( \3053 , \2112 , \2705 );
not \mul_6_18_g44118/U$4 ( \3054 , \2112 );
and \mul_6_18_g44118/U$3 ( \3055 , \3054 , \2993 );
nor \mul_6_18_g44118/U$1 ( \3056 , \3053 , \3055 );
nand \mul_6_18_g43609/U$1 ( \3057 , \2701 , \3056 );
nand \mul_6_18_g43096/U$1 ( \3058 , \3052 , \3057 );
and \mul_6_18_g42731/U$3 ( \3059 , \3049 , \3058 );
and \mul_6_18_g42731/U$5 ( \3060 , \3038 , \3048 );
or \mul_6_18_g42731/U$2 ( \3061 , \3059 , \3060 );
xor \mul_6_18_g42372/U$1 ( \3062 , \3028 , \3061 );
not \mul_6_18_g43167/U$3 ( \3063 , \2956 );
not \mul_6_18_g43167/U$4 ( \3064 , \2303 );
or \mul_6_18_g43167/U$2 ( \3065 , \3063 , \3064 );
nand \mul_6_18_g43607/U$1 ( \3066 , \2318 , \2314 );
nand \mul_6_18_g43167/U$1 ( \3067 , \3065 , \3066 );
not \mul_6_18_g43143/U$3 ( \3068 , \2984 );
not \mul_6_18_g43143/U$4 ( \3069 , \2773 );
or \mul_6_18_g43143/U$2 ( \3070 , \3068 , \3069 );
not \mul_6_18_g44011/U$3 ( \3071 , \2092 );
not \mul_6_18_g44011/U$4 ( \3072 , \2762 );
or \mul_6_18_g44011/U$2 ( \3073 , \3071 , \3072 );
nand \mul_6_18_g44255/U$1 ( \3074 , \2765 , \2754 );
nand \mul_6_18_g44011/U$1 ( \3075 , \3073 , \3074 );
nand \mul_6_18_g43465/U$1 ( \3076 , \2784 , \3075 );
nand \mul_6_18_g43143/U$1 ( \3077 , \3070 , \3076 );
xor \mul_6_18_g42717/U$4 ( \3078 , \3067 , \3077 );
not \mul_6_18_g43593/U$1 ( \3079 , \2965 );
not \mul_6_18_g43887/U$1 ( \3080 , \2974 );
or \mul_6_18_g43275/U$2 ( \3081 , \3079 , \3080 );
and \mul_6_18_g43889/U$2 ( \3082 , \2969 , \2105 );
not \mul_6_18_g44821/U$1 ( \3083 , \2969 );
and \mul_6_18_g43889/U$3 ( \3084 , \3083 , \2568 );
nor \mul_6_18_g43889/U$1 ( \3085 , \3082 , \3084 );
not \mul_6_18_g43772/U$1 ( \3086 , \2733 );
or \mul_6_18_g43275/U$3 ( \3087 , \3085 , \3086 );
nand \mul_6_18_g43275/U$1 ( \3088 , \3081 , \3087 );
and \mul_6_18_g42717/U$3 ( \3089 , \3078 , \3088 );
and \mul_6_18_g42717/U$5 ( \3090 , \3067 , \3077 );
or \mul_6_18_g42717/U$2 ( \3091 , \3089 , \3090 );
xor \mul_6_18_g42372/U$1_r1 ( \3092 , \3062 , \3091 );
xor \mul_6_18_g42202/U$1_r1 ( \3093 , \3004 , \3092 );
xor \mul_6_18_g42068/U$1_r1 ( \3094 , \2868 , \3093 );
xor \mul_6_18_g42199/U$1 ( \3095 , \2524 , \2637 );
xor \mul_6_18_g42199/U$1_r1 ( \3096 , \3095 , \2864 );
xor \mul_6_18_g42360/U$1 ( \3097 , \2925 , \2961 );
xor \mul_6_18_g42360/U$1_r1 ( \3098 , \3097 , \3000 );
xor \mul_6_18_g42629/U$1 ( \3099 , \2936 , \2947 );
xor \mul_6_18_g42629/U$1_r1 ( \3100 , \3099 , \2958 );
not \mul_6_18_g43178/U$3 ( \3101 , \2656 );
not \mul_6_18_g43178/U$4 ( \3102 , \2349 );
or \mul_6_18_g43178/U$2 ( \3103 , \3101 , \3102 );
nand \mul_6_18_g43643/U$1 ( \3104 , \2359 , \3043 );
nand \mul_6_18_g43178/U$1 ( \3105 , \3103 , \3104 );
not \mul_6_18_g43212/U$3 ( \3106 , \2672 );
not \mul_6_18_g43212/U$4 ( \3107 , \2400 );
or \mul_6_18_g43212/U$2 ( \3108 , \3106 , \3107 );
nand \mul_6_18_g43437/U$1 ( \3109 , \2403 , \3033 );
nand \mul_6_18_g43212/U$1 ( \3110 , \3108 , \3109 );
xor \mul_6_18_g42578/U$1 ( \3111 , \3105 , \3110 );
and \mul_6_18_g42850/U$1 ( \3112 , \2844 , \2855 );
xor \mul_6_18_g42578/U$1_r1 ( \3113 , \3111 , \3112 );
xor \mul_6_18_g42413/U$4 ( \3114 , \3100 , \3113 );
xor \mul_6_18_g42725/U$1 ( \3115 , \2976 , \2986 );
xor \mul_6_18_g42725/U$1_r1 ( \3116 , \3115 , \2997 );
and \mul_6_18_g42413/U$3 ( \3117 , \3114 , \3116 );
and \mul_6_18_g42413/U$5 ( \3118 , \3100 , \3113 );
or \mul_6_18_g42413/U$2 ( \3119 , \3117 , \3118 );
xor \mul_6_18_g42196/U$1 ( \3120 , \3098 , \3119 );
xor \mul_6_18_g42647/U$1 ( \3121 , \2140 , \2174 );
xor \mul_6_18_g42647/U$1_r1 ( \3122 , \3121 , \2212 );
xor \mul_6_18_g42717/U$1 ( \3123 , \3067 , \3077 );
xor \mul_6_18_g42717/U$1_r1 ( \3124 , \3123 , \3088 );
xor \mul_6_18_g42405/U$1 ( \3125 , \3122 , \3124 );
xor \mul_6_18_g42731/U$1 ( \3126 , \3038 , \3048 );
xor \mul_6_18_g42731/U$1_r1 ( \3127 , \3126 , \3058 );
xor \mul_6_18_g42405/U$1_r1 ( \3128 , \3125 , \3127 );
xor \mul_6_18_g42196/U$1_r1 ( \3129 , \3120 , \3128 );
xor \mul_6_18_g42045/U$4 ( \3130 , \3096 , \3129 );
xor \mul_6_18_g42413/U$1 ( \3131 , \3100 , \3113 );
xor \mul_6_18_g42413/U$1_r1 ( \3132 , \3131 , \3116 );
not \mul_6_18_g45174/U$2 ( \3133 , \3132 );
not \mul_6_18_g43000/U$3 ( \3134 , \2573 );
not \mul_6_18_g43000/U$4 ( \3135 , \2539 );
or \mul_6_18_g43000/U$2 ( \3136 , \3134 , \3135 );
nand \mul_6_18_g43050/U$1 ( \3137 , \2538 , \2554 );
nand \mul_6_18_g43000/U$1 ( \3138 , \3136 , \3137 );
xnor \mul_6_18_g45219/U$1 ( \3139 , \3138 , \2572 );
xor \mul_6_18_g42660/U$1 ( \3140 , \2806 , \2828 );
xnor \mul_6_18_g42660/U$1_r1 ( \3141 , \3140 , \2856 );
xor \mul_6_18_g42251/U$4 ( \3142 , \3139 , \3141 );
not \mul_6_18_g44095/U$3 ( \3143 , \2144 );
not \mul_6_18_g44095/U$4 ( \3144 , \2182 );
or \mul_6_18_g44095/U$2 ( \3145 , \3143 , \3144 );
nand \mul_6_18_g44284/U$1 ( \3146 , \2181 , \2145 );
nand \mul_6_18_g44095/U$1 ( \3147 , \3145 , \3146 );
not \mul_6_18_g43070/U$3 ( \3148 , \3147 );
not \mul_6_18_g43070/U$4 ( \3149 , \2202 );
or \mul_6_18_g43070/U$2 ( \3150 , \3148 , \3149 );
not \mul_6_18_g44093/U$3 ( \3151 , \2168 );
not \mul_6_18_g44093/U$4 ( \3152 , \2182 );
or \mul_6_18_g44093/U$2 ( \3153 , \3151 , \3152 );
not \mul_6_18_g44529/U$1 ( \3154 , \2168 );
nand \mul_6_18_g44285/U$1 ( \3155 , \2181 , \3154 );
nand \mul_6_18_g44093/U$1 ( \3156 , \3153 , \3155 );
nand \mul_6_18_g43475/U$1 ( \3157 , \3156 , \2210 );
nand \mul_6_18_g43070/U$1 ( \3158 , \3150 , \3157 );
and \mul_6_18_g43923/U$2 ( \3159 , \2116 , \2159 );
not \mul_6_18_g43923/U$4 ( \3160 , \2116 );
and \mul_6_18_g43923/U$3 ( \3161 , \3160 , \2146 );
nor \mul_6_18_g43923/U$1 ( \3162 , \3159 , \3161 );
not \mul_6_18_g43065/U$3 ( \3163 , \3162 );
not \mul_6_18_g43065/U$4 ( \3164 , \2162 );
or \mul_6_18_g43065/U$2 ( \3165 , \3163 , \3164 );
nand \mul_6_18_g43563/U$1 ( \3166 , \2525 , \2155 );
nand \mul_6_18_g43065/U$1 ( \3167 , \3165 , \3166 );
and \mul_6_18_g42865/U$2 ( \3168 , \3158 , \3167 );
not \mul_6_18_g42865/U$4 ( \3169 , \3158 );
not \fopt45609/U$1 ( \3170 , \3167 );
and \mul_6_18_g42865/U$3 ( \3171 , \3169 , \3170 );
nor \mul_6_18_g42865/U$1 ( \3172 , \3168 , \3171 );
nor \mul_6_18_g43645/U$1 ( \3173 , \2154 , \2116 );
not \mul_6_18_g43870/U$3 ( \3174 , \2099 );
not \mul_6_18_g43870/U$4 ( \3175 , \2423 );
or \mul_6_18_g43870/U$2 ( \3176 , \3174 , \3175 );
nand \mul_6_18_g44199/U$1 ( \3177 , \2848 , \2257 );
nand \mul_6_18_g43870/U$1 ( \3178 , \3176 , \3177 );
not \mul_6_18_g42924/U$3 ( \3179 , \3178 );
not \mul_6_18_g42924/U$4 ( \3180 , \2586 );
or \mul_6_18_g42924/U$2 ( \3181 , \3179 , \3180 );
nand \mul_6_18_g43009/U$1 ( \3182 , \2434 , \2850 );
nand \mul_6_18_g42924/U$1 ( \3183 , \3181 , \3182 );
xor \mul_6_18_g42561/U$4 ( \3184 , \3173 , \3183 );
not \mul_6_18_g43883/U$3 ( \3185 , \2105 );
not \mul_6_18_g44859/U$1 ( \3186 , \2626 );
not \mul_6_18_g43883/U$4 ( \3187 , \3186 );
or \mul_6_18_g43883/U$2 ( \3188 , \3185 , \3187 );
nand \mul_6_18_g44213/U$1 ( \3189 , \2626 , \2568 );
nand \mul_6_18_g43883/U$1 ( \3190 , \3188 , \3189 );
not \mul_6_18_g42967/U$3 ( \3191 , \3190 );
not \mul_6_18_g42967/U$4 ( \3192 , \2907 );
or \mul_6_18_g42967/U$2 ( \3193 , \3191 , \3192 );
nand \mul_6_18_g43011/U$1 ( \3194 , \2623 , \2838 );
nand \mul_6_18_g42967/U$1 ( \3195 , \3193 , \3194 );
and \mul_6_18_g42561/U$3 ( \3196 , \3184 , \3195 );
and \mul_6_18_g42561/U$5 ( \3197 , \3173 , \3183 );
or \mul_6_18_g42561/U$2 ( \3198 , \3196 , \3197 );
not \mul_6_18_g42560/U$1 ( \3199 , \3198 );
and \mul_6_18_g42492/U$2 ( \3200 , \3172 , \3199 );
not \mul_6_18_g42492/U$4 ( \3201 , \3172 );
and \mul_6_18_g42492/U$3 ( \3202 , \3201 , \3198 );
nor \mul_6_18_g42492/U$1 ( \3203 , \3200 , \3202 );
and \mul_6_18_g42251/U$3 ( \3204 , \3142 , \3203 );
and \mul_6_18_g42251/U$5 ( \3205 , \3139 , \3141 );
or \mul_6_18_g42251/U$2 ( \3206 , \3204 , \3205 );
nand \mul_6_18_g45174/U$1 ( \3207 , \3133 , \3206 );
not \mul_6_18_g42127/U$3 ( \3208 , \3207 );
xor \mul_6_18_g42561/U$1 ( \3209 , \3173 , \3183 );
xor \mul_6_18_g42561/U$1_r1 ( \3210 , \3209 , \3195 );
not \mul_6_18_g44713/U$1 ( \3211 , \2216 );
and \g45501/U$2 ( \3212 , \2098 , \3211 );
not \g45501/U$4 ( \3213 , \2098 );
not \mul_6_18_g44702/U$1 ( \3214 , \2216 );
not \mul_6_18_g44701/U$1 ( \3215 , \3214 );
and \g45501/U$3 ( \3216 , \3213 , \3215 );
or \g45501/U$1 ( \3217 , \3212 , \3216 );
not \mul_6_18_g43363/U$3 ( \3218 , \3217 );
not \mul_6_18_g43363/U$4 ( \3219 , \2222 );
or \mul_6_18_g43363/U$2 ( \3220 , \3218 , \3219 );
nand \mul_6_18_g43496/U$1 ( \3221 , \2545 , \2934 );
nand \mul_6_18_g43363/U$1 ( \3222 , \3220 , \3221 );
not \mul_6_18_g43900/U$3 ( \3223 , \2110 );
not \mul_6_18_g44971/U$1 ( \3224 , \2256 );
not \mul_6_18_g43900/U$4 ( \3225 , \3224 );
or \mul_6_18_g43900/U$2 ( \3226 , \3223 , \3225 );
nand \mul_6_18_g44228/U$1 ( \3227 , \2256 , \2369 );
nand \mul_6_18_g43900/U$1 ( \3228 , \3226 , \3227 );
not \mul_6_18_g43286/U$3 ( \3229 , \3228 );
not \mul_6_18_g43286/U$4 ( \3230 , \2938 );
or \mul_6_18_g43286/U$2 ( \3231 , \3229 , \3230 );
not \mul_6_18_g43757/U$1 ( \3232 , \2284 );
nand \mul_6_18_g43499/U$1 ( \3233 , \3232 , \2561 );
nand \mul_6_18_g43286/U$1 ( \3234 , \3231 , \3233 );
xor \mul_6_18_g42622/U$1 ( \3235 , \3222 , \3234 );
not \mul_6_18_g44025/U$3 ( \3236 , \2111 );
not \mul_6_18_g44756/U$1 ( \3237 , \2307 );
not \mul_6_18_g44025/U$4 ( \3238 , \3237 );
or \mul_6_18_g44025/U$2 ( \3239 , \3236 , \3238 );
nand \mul_6_18_g44283/U$1 ( \3240 , \2311 , \2779 );
nand \mul_6_18_g44025/U$1 ( \3241 , \3239 , \3240 );
not \mul_6_18_g43156/U$3 ( \3242 , \3241 );
not \mul_6_18_g43156/U$4 ( \3243 , \2303 );
or \mul_6_18_g43156/U$2 ( \3244 , \3242 , \3243 );
nand \mul_6_18_g43531/U$1 ( \3245 , \2318 , \2747 );
nand \mul_6_18_g43156/U$1 ( \3246 , \3244 , \3245 );
xor \mul_6_18_g42622/U$1_r1 ( \3247 , \3235 , \3246 );
xor \mul_6_18_g42370/U$4 ( \3248 , \3210 , \3247 );
not \mul_6_18_g44115/U$3 ( \3249 , \2463 );
not \mul_6_18_g44115/U$4 ( \3250 , \2495 );
or \mul_6_18_g44115/U$2 ( \3251 , \3249 , \3250 );
nand \mul_6_18_g44329/U$1 ( \3252 , \2496 , \2468 );
nand \mul_6_18_g44115/U$1 ( \3253 , \3251 , \3252 );
not \mul_6_18_g43105/U$3 ( \3254 , \3253 );
not \mul_6_18_g43105/U$4 ( \3255 , \2511 );
or \mul_6_18_g43105/U$2 ( \3256 , \3254 , \3255 );
buf \mul_6_18_fopt45112/U$1 ( \3257 , \1160 );
and \mul_6_18_g44116/U$2 ( \3258 , \1998 , \3257 );
not \mul_6_18_g44116/U$4 ( \3259 , \1998 );
and \mul_6_18_g44116/U$3 ( \3260 , \3259 , \2495 );
nor \mul_6_18_g44116/U$1 ( \3261 , \3258 , \3260 );
nand \mul_6_18_g43504/U$1 ( \3262 , \2515 , \3261 );
nand \mul_6_18_g43105/U$1 ( \3263 , \3256 , \3262 );
not \mul_6_18_g44132/U$3 ( \3264 , \2144 );
not \mul_6_18_g44132/U$4 ( \3265 , \2465 );
or \mul_6_18_g44132/U$2 ( \3266 , \3264 , \3265 );
nand \mul_6_18_g44325/U$1 ( \3267 , \2475 , \2145 );
nand \mul_6_18_g44132/U$1 ( \3268 , \3266 , \3267 );
not \mul_6_18_g43082/U$3 ( \3269 , \3268 );
nor \mul_6_18_g43705/U$1 ( \3270 , \2480 , \2479 );
not \mul_6_18_g43082/U$4 ( \3271 , \3270 );
or \mul_6_18_g43082/U$2 ( \3272 , \3269 , \3271 );
not \mul_6_18_g44130/U$3 ( \3273 , \2168 );
not \mul_6_18_g44130/U$4 ( \3274 , \2465 );
or \mul_6_18_g44130/U$2 ( \3275 , \3273 , \3274 );
nand \mul_6_18_g44328/U$1 ( \3276 , \2475 , \3154 );
nand \mul_6_18_g44130/U$1 ( \3277 , \3275 , \3276 );
nand \mul_6_18_g43573/U$1 ( \3278 , \3277 , \2480 );
nand \mul_6_18_g43082/U$1 ( \3279 , \3272 , \3278 );
or \mul_6_18_g45211/U$1 ( \3280 , \3263 , \3279 );
not \g45553/U$3 ( \3281 , \3280 );
not \mul_6_18_g43871/U$3 ( \3282 , \2832 );
not \mul_6_18_g43871/U$4 ( \3283 , \2423 );
or \mul_6_18_g43871/U$2 ( \3284 , \3282 , \3283 );
nand \mul_6_18_g44203/U$1 ( \3285 , \2418 , \2831 );
nand \mul_6_18_g43871/U$1 ( \3286 , \3284 , \3285 );
not \mul_6_18_g42933/U$3 ( \3287 , \3286 );
not \mul_6_18_g42933/U$4 ( \3288 , \2586 );
or \mul_6_18_g42933/U$2 ( \3289 , \3287 , \3288 );
nand \mul_6_18_g43022/U$1 ( \3290 , \2434 , \3178 );
nand \mul_6_18_g42933/U$1 ( \3291 , \3289 , \3290 );
not \mul_6_18_g43884/U$3 ( \3292 , \2405 );
not \mul_6_18_g43884/U$4 ( \3293 , \2629 );
or \mul_6_18_g43884/U$2 ( \3294 , \3292 , \3293 );
nand \mul_6_18_g44212/U$1 ( \3295 , \2606 , \2404 );
nand \mul_6_18_g43884/U$1 ( \3296 , \3294 , \3295 );
not \mul_6_18_g42976/U$3 ( \3297 , \3296 );
not \mul_6_18_g42976/U$4 ( \3298 , \2907 );
or \mul_6_18_g42976/U$2 ( \3299 , \3297 , \3298 );
nand \mul_6_18_g43023/U$1 ( \3300 , \2623 , \3190 );
nand \mul_6_18_g42976/U$1 ( \3301 , \3299 , \3300 );
xor \mul_6_18_g42787/U$1 ( \3302 , \3291 , \3301 );
not \g45553/U$4 ( \3303 , \3302 );
or \g45553/U$2 ( \3304 , \3281 , \3303 );
nand \mul_6_18_g42911/U$1 ( \3305 , \3263 , \3279 );
nand \g45553/U$1 ( \3306 , \3304 , \3305 );
and \mul_6_18_g42370/U$3 ( \3307 , \3248 , \3306 );
and \mul_6_18_g42370/U$5 ( \3308 , \3210 , \3247 );
or \mul_6_18_g42370/U$2 ( \3309 , \3307 , \3308 );
not \mul_6_18_g42369/U$1 ( \3310 , \3309 );
not \mul_6_18_g42368/U$1 ( \3311 , \3310 );
xor \mul_6_18_g42622/U$4 ( \3312 , \3222 , \3234 );
and \mul_6_18_g42622/U$3 ( \3313 , \3312 , \3246 );
and \mul_6_18_g42622/U$5 ( \3314 , \3222 , \3234 );
or \mul_6_18_g42622/U$2 ( \3315 , \3313 , \3314 );
not \mul_6_18_g43922/U$3 ( \3316 , \2972 );
not \mul_6_18_g43922/U$4 ( \3317 , \2670 );
and \mul_6_18_g43922/U$2 ( \3318 , \3316 , \3317 );
and \mul_6_18_g43922/U$5 ( \3319 , \2719 , \2670 );
nor \mul_6_18_g43922/U$1 ( \3320 , \3318 , \3319 );
not \mul_6_18_g43921/U$1 ( \3321 , \3320 );
not \mul_6_18_g43259/U$3 ( \3322 , \3321 );
not \mul_6_18_g43591/U$1 ( \3323 , \2964 );
not \mul_6_18_g43259/U$4 ( \3324 , \3323 );
or \mul_6_18_g43259/U$2 ( \3325 , \3322 , \3324 );
not \mul_6_18_g43782/U$1 ( \3326 , \2732 );
nand \mul_6_18_g43530/U$1 ( \3327 , \3326 , \2721 );
nand \mul_6_18_g43259/U$1 ( \3328 , \3325 , \3327 );
not \mul_6_18_g44079/U$3 ( \3329 , \2112 );
buf \mul_6_18_g44508/U$1 ( \3330 , \1218 );
not \mul_6_18_g44510/U$1 ( \3331 , \3330 );
not \mul_6_18_g44079/U$4 ( \3332 , \3331 );
or \mul_6_18_g44079/U$2 ( \3333 , \3329 , \3332 );
nand \mul_6_18_g44312/U$1 ( \3334 , \3330 , \2824 );
nand \mul_6_18_g44079/U$1 ( \3335 , \3333 , \3334 );
not \mul_6_18_g43145/U$3 ( \3336 , \3335 );
not \mul_6_18_g43145/U$4 ( \3337 , \2773 );
or \mul_6_18_g43145/U$2 ( \3338 , \3336 , \3337 );
nand \mul_6_18_g43613/U$1 ( \3339 , \2784 , \2767 );
nand \mul_6_18_g43145/U$1 ( \3340 , \3338 , \3339 );
xor \mul_6_18_g42623/U$4 ( \3341 , \3328 , \3340 );
and \mul_6_18_g44146/U$2 ( \3342 , \2006 , \2684 );
not \mul_6_18_g44146/U$4 ( \3343 , \2006 );
and \mul_6_18_g44146/U$3 ( \3344 , \3343 , \2993 );
nor \mul_6_18_g44146/U$1 ( \3345 , \3342 , \3344 );
not \mul_6_18_g43102/U$3 ( \3346 , \3345 );
not \mul_6_18_g43102/U$4 ( \3347 , \2692 );
or \mul_6_18_g43102/U$2 ( \3348 , \3346 , \3347 );
nand \mul_6_18_g43533/U$1 ( \3349 , \2701 , \2699 );
nand \mul_6_18_g43102/U$1 ( \3350 , \3348 , \3349 );
and \mul_6_18_g42623/U$3 ( \3351 , \3341 , \3350 );
and \mul_6_18_g42623/U$5 ( \3352 , \3328 , \3340 );
or \mul_6_18_g42623/U$2 ( \3353 , \3351 , \3352 );
xor \mul_6_18_g42424/U$1 ( \3354 , \3315 , \3353 );
not \mul_6_18_g43085/U$3 ( \3355 , \3277 );
not \mul_6_18_g43085/U$4 ( \3356 , \2481 );
or \mul_6_18_g43085/U$2 ( \3357 , \3355 , \3356 );
nand \mul_6_18_g43527/U$1 ( \3358 , \2804 , \2480 );
nand \mul_6_18_g43085/U$1 ( \3359 , \3357 , \3358 );
not \mul_6_18_g44474/U$1 ( \3360 , \2056 );
and \mul_6_18_g44085/U$2 ( \3361 , \3360 , \2182 );
not \mul_6_18_g44085/U$4 ( \3362 , \3360 );
and \mul_6_18_g44085/U$3 ( \3363 , \3362 , \2181 );
nor \mul_6_18_g44085/U$1 ( \3364 , \3361 , \3363 );
not \mul_6_18_g43072/U$3 ( \3365 , \3364 );
not \mul_6_18_g43072/U$4 ( \3366 , \2202 );
or \mul_6_18_g43072/U$2 ( \3367 , \3365 , \3366 );
nand \mul_6_18_g43523/U$1 ( \3368 , \3147 , \2210 );
nand \mul_6_18_g43072/U$1 ( \3369 , \3367 , \3368 );
xor \mul_6_18_g42585/U$4 ( \3370 , \3359 , \3369 );
and \mul_6_18_g42787/U$2 ( \3371 , \3291 , \3301 );
and \mul_6_18_g42585/U$3 ( \3372 , \3370 , \3371 );
and \mul_6_18_g42585/U$5 ( \3373 , \3359 , \3369 );
or \mul_6_18_g42585/U$2 ( \3374 , \3372 , \3373 );
xor \mul_6_18_g42424/U$1_r1 ( \3375 , \3354 , \3374 );
or \mul_6_18_g42283/U$2 ( \3376 , \3311 , \3375 );
not \mul_6_18_g43984/U$3 ( \3377 , \2107 );
not \mul_6_18_g43984/U$4 ( \3378 , \2644 );
or \mul_6_18_g43984/U$2 ( \3379 , \3377 , \3378 );
not \mul_6_18_fopt45059/U$1 ( \3380 , \2644 );
nand \mul_6_18_g44263/U$1 ( \3381 , \3380 , \2745 );
nand \mul_6_18_g43984/U$1 ( \3382 , \3379 , \3381 );
not \mul_6_18_g43194/U$3 ( \3383 , \3382 );
not \mul_6_18_g43194/U$4 ( \3384 , \2349 );
or \mul_6_18_g43194/U$2 ( \3385 , \3383 , \3384 );
not \mul_6_18_g43985/U$3 ( \3386 , \2092 );
not \mul_6_18_g43985/U$4 ( \3387 , \2645 );
or \mul_6_18_g43985/U$2 ( \3388 , \3386 , \3387 );
nand \mul_6_18_g45807/U$1 ( \3389 , \2335 , \2754 );
nand \mul_6_18_g43985/U$1 ( \3390 , \3388 , \3389 );
nand \mul_6_18_g43552/U$1 ( \3391 , \2359 , \3390 );
nand \mul_6_18_g43194/U$1 ( \3392 , \3385 , \3391 );
not \mul_6_18_g43953/U$3 ( \3393 , \2640 );
not \mul_6_18_g44550/U$1 ( \3394 , \2663 );
not \mul_6_18_g43953/U$4 ( \3395 , \3394 );
or \mul_6_18_g43953/U$2 ( \3396 , \3393 , \3395 );
nand \mul_6_18_g44247/U$1 ( \3397 , \2368 , \2639 );
nand \mul_6_18_g43953/U$1 ( \3398 , \3396 , \3397 );
not \mul_6_18_g43243/U$3 ( \3399 , \3398 );
not \mul_6_18_g43243/U$4 ( \3400 , \2400 );
or \mul_6_18_g43243/U$2 ( \3401 , \3399 , \3400 );
not \mul_6_18_g43954/U$3 ( \3402 , \2305 );
not \mul_6_18_g43954/U$4 ( \3403 , \2367 );
or \mul_6_18_g43954/U$2 ( \3404 , \3402 , \3403 );
nand \mul_6_18_g44250/U$1 ( \3405 , \2663 , \2312 );
nand \mul_6_18_g43954/U$1 ( \3406 , \3404 , \3405 );
nand \mul_6_18_g43556/U$1 ( \3407 , \2403 , \3406 );
nand \mul_6_18_g43243/U$1 ( \3408 , \3401 , \3407 );
xor \mul_6_18_g42730/U$4 ( \3409 , \3392 , \3408 );
and \mul_6_18_g44147/U$2 ( \3410 , \2179 , \2697 );
not \mul_6_18_g44147/U$4 ( \3411 , \2179 );
and \mul_6_18_g44147/U$3 ( \3412 , \3411 , \2993 );
nor \mul_6_18_g44147/U$1 ( \3413 , \3410 , \3412 );
not \mul_6_18_g43101/U$3 ( \3414 , \3413 );
not \mul_6_18_g43101/U$4 ( \3415 , \2691 );
or \mul_6_18_g43101/U$2 ( \3416 , \3414 , \3415 );
nand \mul_6_18_g43632/U$1 ( \3417 , \2701 , \3345 );
nand \mul_6_18_g43101/U$1 ( \3418 , \3416 , \3417 );
and \mul_6_18_g42730/U$3 ( \3419 , \3409 , \3418 );
and \mul_6_18_g42730/U$5 ( \3420 , \3392 , \3408 );
or \mul_6_18_g42730/U$2 ( \3421 , \3419 , \3420 );
not \mul_6_18_g44688/U$1 ( \3422 , \2225 );
and \g45500/U$2 ( \3423 , \2097 , \3422 );
not \g45500/U$4 ( \3424 , \2097 );
and \g45500/U$3 ( \3425 , \3424 , \2225 );
or \g45500/U$1 ( \3426 , \3423 , \3425 );
not \mul_6_18_g43371/U$3 ( \3427 , \3426 );
not \mul_6_18_g43371/U$4 ( \3428 , \2222 );
or \mul_6_18_g43371/U$2 ( \3429 , \3427 , \3428 );
not \mul_6_18_g44878/U$1 ( \3430 , \2243 );
nand \mul_6_18_g43545/U$1 ( \3431 , \3217 , \3430 );
nand \mul_6_18_g43371/U$1 ( \3432 , \3429 , \3431 );
nand \mul_6_18_g44163/U$1 ( \3433 , \2190 , \2116 );
and \mul_6_18_g43687/U$2 ( \3434 , \2475 , \3433 );
not \mul_6_18_g43726/U$3 ( \3435 , \2058 );
not \mul_6_18_g43726/U$4 ( \3436 , \2189 );
or \mul_6_18_g43726/U$2 ( \3437 , \3435 , \3436 );
nand \mul_6_18_g43726/U$1 ( \3438 , \3437 , \1015 );
nor \mul_6_18_g43687/U$1 ( \3439 , \3434 , \3438 );
xor \mul_6_18_g42713/U$4 ( \3440 , \3432 , \3439 );
not \mul_6_18_g43901/U$3 ( \3441 , \2352 );
not \mul_6_18_g43901/U$4 ( \3442 , \3224 );
or \mul_6_18_g43901/U$2 ( \3443 , \3441 , \3442 );
nand \mul_6_18_g44216/U$1 ( \3444 , \2280 , \2354 );
nand \mul_6_18_g43901/U$1 ( \3445 , \3443 , \3444 );
not \mul_6_18_g43302/U$3 ( \3446 , \3445 );
not \mul_6_18_g43302/U$4 ( \3447 , \2273 );
or \mul_6_18_g43302/U$2 ( \3448 , \3446 , \3447 );
not \mul_6_18_g43768/U$1 ( \3449 , \2284 );
nand \mul_6_18_g43559/U$1 ( \3450 , \3449 , \3228 );
nand \mul_6_18_g43302/U$1 ( \3451 , \3448 , \3450 );
and \mul_6_18_g42713/U$3 ( \3452 , \3440 , \3451 );
and \mul_6_18_g42713/U$5 ( \3453 , \3432 , \3439 );
or \mul_6_18_g42713/U$2 ( \3454 , \3452 , \3453 );
or \mul_6_18_g42541/U$2 ( \3455 , \3421 , \3454 );
not \mul_6_18_g44026/U$3 ( \3456 , \2094 );
not \mul_6_18_g44026/U$4 ( \3457 , \3237 );
or \mul_6_18_g44026/U$2 ( \3458 , \3456 , \3457 );
nand \mul_6_18_g44275/U$1 ( \3459 , \2307 , \2500 );
nand \mul_6_18_g44026/U$1 ( \3460 , \3458 , \3459 );
not \mul_6_18_g43166/U$3 ( \3461 , \3460 );
not \mul_6_18_g43166/U$4 ( \3462 , \2303 );
or \mul_6_18_g43166/U$2 ( \3463 , \3461 , \3462 );
nand \mul_6_18_g43605/U$1 ( \3464 , \2318 , \3241 );
nand \mul_6_18_g43166/U$1 ( \3465 , \3463 , \3464 );
not \mul_6_18_g42693/U$3 ( \3466 , \3465 );
not \mul_6_18_g44831/U$1 ( \3467 , \2715 );
and \mul_6_18_g43920/U$2 ( \3468 , \2321 , \3467 );
not \mul_6_18_g43920/U$4 ( \3469 , \2321 );
and \mul_6_18_g43920/U$3 ( \3470 , \3469 , \2718 );
nor \mul_6_18_g43920/U$1 ( \3471 , \3468 , \3470 );
or \mul_6_18_g43248/U$2 ( \3472 , \2964 , \3471 );
not \mul_6_18_g43781/U$1 ( \3473 , \3326 );
or \mul_6_18_g43248/U$3 ( \3474 , \3473 , \3320 );
nand \mul_6_18_g43248/U$1 ( \3475 , \3472 , \3474 );
not \mul_6_18_g42693/U$4 ( \3476 , \3475 );
or \mul_6_18_g42693/U$2 ( \3477 , \3466 , \3476 );
or \mul_6_18_g42747/U$2 ( \3478 , \3475 , \3465 );
not \mul_6_18_g44078/U$3 ( \3479 , \2812 );
not \mul_6_18_g44078/U$4 ( \3480 , \3331 );
or \mul_6_18_g44078/U$2 ( \3481 , \3479 , \3480 );
nand \mul_6_18_g44302/U$1 ( \3482 , \3330 , \2811 );
nand \mul_6_18_g44078/U$1 ( \3483 , \3481 , \3482 );
not \mul_6_18_g43139/U$3 ( \3484 , \3483 );
not \mul_6_18_g43139/U$4 ( \3485 , \2773 );
or \mul_6_18_g43139/U$2 ( \3486 , \3484 , \3485 );
nand \mul_6_18_g43566/U$1 ( \3487 , \2784 , \3335 );
nand \mul_6_18_g43139/U$1 ( \3488 , \3486 , \3487 );
nand \mul_6_18_g42747/U$1 ( \3489 , \3478 , \3488 );
nand \mul_6_18_g42693/U$1 ( \3490 , \3477 , \3489 );
nand \mul_6_18_g42541/U$1 ( \3491 , \3455 , \3490 );
nand \mul_6_18_g42589/U$1 ( \3492 , \3421 , \3454 );
nand \mul_6_18_g42519/U$1 ( \3493 , \3491 , \3492 );
nand \mul_6_18_g42283/U$1 ( \3494 , \3376 , \3493 );
nand \mul_6_18_g42309/U$1 ( \3495 , \3311 , \3375 );
nand \mul_6_18_g42244/U$1 ( \3496 , \3494 , \3495 );
not \mul_6_18_g42127/U$4 ( \3497 , \3496 );
or \mul_6_18_g42127/U$2 ( \3498 , \3208 , \3497 );
not \mul_6_18_g42250/U$1 ( \3499 , \3206 );
nand \mul_6_18_g42219/U$1 ( \3500 , \3132 , \3499 );
nand \mul_6_18_g42127/U$1 ( \3501 , \3498 , \3500 );
and \mul_6_18_g42045/U$3 ( \3502 , \3130 , \3501 );
and \mul_6_18_g42045/U$5 ( \3503 , \3096 , \3129 );
or \mul_6_18_g42045/U$2 ( \3504 , \3502 , \3503 );
xor \mul_6_18_g41910/U$1 ( \3505 , \3094 , \3504 );
xor \mul_6_18_g42196/U$4 ( \3506 , \3098 , \3119 );
and \mul_6_18_g42196/U$3 ( \3507 , \3506 , \3128 );
and \mul_6_18_g42196/U$5 ( \3508 , \3098 , \3119 );
or \mul_6_18_g42196/U$2 ( \3509 , \3507 , \3508 );
xor \mul_6_18_g42578/U$4 ( \3510 , \3105 , \3110 );
and \mul_6_18_g42578/U$3 ( \3511 , \3510 , \3112 );
and \mul_6_18_g42578/U$5 ( \3512 , \3105 , \3110 );
or \mul_6_18_g42578/U$2 ( \3513 , \3511 , \3512 );
not \mul_6_18_g42577/U$1 ( \3514 , \3513 );
not \mul_6_18_g42460/U$3 ( \3515 , \3514 );
xor \mul_6_18_g42657/U$1 ( \3516 , \3009 , \3018 );
xnor \mul_6_18_g42657/U$1_r1 ( \3517 , \3516 , \3026 );
not \mul_6_18_g42460/U$4 ( \3518 , \3517 );
or \mul_6_18_g42460/U$2 ( \3519 , \3515 , \3518 );
not \mul_6_18_g43068/U$3 ( \3520 , \3156 );
not \mul_6_18_g43068/U$4 ( \3521 , \2202 );
or \mul_6_18_g43068/U$2 ( \3522 , \3520 , \3521 );
nand \mul_6_18_g43476/U$1 ( \3523 , \2187 , \2210 );
nand \mul_6_18_g43068/U$1 ( \3524 , \3522 , \3523 );
not \mul_6_18_g42896/U$2 ( \3525 , \3524 );
and \mul_6_18_g43128/U$2 ( \3526 , \2511 , \2826 );
and \mul_6_18_g43128/U$3 ( \3527 , \2502 , \2515 );
nor \mul_6_18_g43128/U$1 ( \3528 , \3526 , \3527 );
nand \mul_6_18_g42896/U$1 ( \3529 , \3525 , \3528 );
and \mul_6_18_g43084/U$2 ( \3530 , \2482 , \2797 );
and \mul_6_18_g43084/U$3 ( \3531 , \2485 , \2470 );
nor \mul_6_18_g43084/U$1 ( \3532 , \3530 , \3531 );
not \mul_6_18_g43083/U$1 ( \3533 , \3532 );
and \mul_6_18_g42810/U$2 ( \3534 , \3529 , \3533 );
not \mul_6_18_g42900/U$2 ( \3535 , \3524 );
nor \mul_6_18_g42900/U$1 ( \3536 , \3535 , \3528 );
nor \mul_6_18_g42810/U$1 ( \3537 , \3534 , \3536 );
not \mul_6_18_g42720/U$1 ( \3538 , \3537 );
nand \mul_6_18_g42460/U$1 ( \3539 , \3519 , \3538 );
not \mul_6_18_g45185/U$2 ( \3540 , \3517 );
nand \mul_6_18_g45185/U$1 ( \3541 , \3540 , \3513 );
nand \mul_6_18_g42440/U$1 ( \3542 , \3539 , \3541 );
xor \mul_6_18_g42405/U$4 ( \3543 , \3122 , \3124 );
and \mul_6_18_g42405/U$3 ( \3544 , \3543 , \3127 );
and \mul_6_18_g42405/U$5 ( \3545 , \3122 , \3124 );
or \mul_6_18_g42405/U$2 ( \3546 , \3544 , \3545 );
xor \mul_6_18_g42203/U$1 ( \3547 , \3542 , \3546 );
xor \mul_6_18_g42574/U$4 ( \3548 , \2493 , \2521 );
and \mul_6_18_g42574/U$3 ( \3549 , \3548 , \2523 );
and \mul_6_18_g42574/U$5 ( \3550 , \2493 , \2521 );
or \mul_6_18_g42574/U$2 ( \3551 , \3549 , \3550 );
or \mul_6_18_g43274/U$2 ( \3552 , \3079 , \3085 );
and \mul_6_18_g43878/U$2 ( \3553 , \2969 , \2832 );
and \mul_6_18_g43878/U$3 ( \3554 , \3083 , \2831 );
nor \mul_6_18_g43878/U$1 ( \3555 , \3553 , \3554 );
or \mul_6_18_g43274/U$3 ( \3556 , \3086 , \3555 );
nand \mul_6_18_g43274/U$1 ( \3557 , \3552 , \3556 );
not \mul_6_18_g43129/U$3 ( \3558 , \3075 );
not \mul_6_18_g43129/U$4 ( \3559 , \2773 );
or \mul_6_18_g43129/U$2 ( \3560 , \3558 , \3559 );
and \mul_6_18_g43980/U$2 ( \3561 , \2640 , \2765 );
not \mul_6_18_g43980/U$4 ( \3562 , \2640 );
and \mul_6_18_g43980/U$3 ( \3563 , \3562 , \2762 );
nor \mul_6_18_g43980/U$1 ( \3564 , \3561 , \3563 );
nand \mul_6_18_g43454/U$1 ( \3565 , \2784 , \3564 );
nand \mul_6_18_g43129/U$1 ( \3566 , \3560 , \3565 );
xor \mul_6_18_g42704/U$1 ( \3567 , \3557 , \3566 );
not \mul_6_18_g43103/U$3 ( \3568 , \3056 );
not \mul_6_18_g43103/U$4 ( \3569 , \2692 );
or \mul_6_18_g43103/U$2 ( \3570 , \3568 , \3569 );
or \mul_6_18_g44096/U$2 ( \3571 , \2705 , \2500 );
or \mul_6_18_g44096/U$3 ( \3572 , \2694 , \2094 );
nand \mul_6_18_g44096/U$1 ( \3573 , \3571 , \3572 );
nand \mul_6_18_g43641/U$1 ( \3574 , \2701 , \3573 );
nand \mul_6_18_g43103/U$1 ( \3575 , \3570 , \3574 );
xor \mul_6_18_g42704/U$1_r1 ( \3576 , \3567 , \3575 );
xor \mul_6_18_g42374/U$1 ( \3577 , \3551 , \3576 );
not \mul_6_18_g43088/U$3 ( \3578 , \2485 );
not \mul_6_18_g44138/U$3 ( \3579 , \2812 );
not \mul_6_18_g44138/U$4 ( \3580 , \2195 );
or \mul_6_18_g44138/U$2 ( \3581 , \3579 , \3580 );
nand \mul_6_18_g44293/U$1 ( \3582 , \2196 , \2811 );
nand \mul_6_18_g44138/U$1 ( \3583 , \3581 , \3582 );
not \mul_6_18_g43088/U$4 ( \3584 , \3583 );
or \mul_6_18_g43088/U$2 ( \3585 , \3578 , \3584 );
nand \mul_6_18_g43318/U$1 ( \3586 , \2482 , \2491 );
nand \mul_6_18_g43088/U$1 ( \3587 , \3585 , \3586 );
not \mul_6_18_g43067/U$3 ( \3588 , \2208 );
not \mul_6_18_g43067/U$4 ( \3589 , \2202 );
or \mul_6_18_g43067/U$2 ( \3590 , \3588 , \3589 );
and \mul_6_18_g44121/U$2 ( \3591 , \2468 , \2182 );
not \mul_6_18_g44121/U$4 ( \3592 , \2468 );
and \mul_6_18_g44121/U$3 ( \3593 , \3592 , \2181 );
nor \mul_6_18_g44121/U$1 ( \3594 , \3591 , \3593 );
nand \mul_6_18_g43571/U$1 ( \3595 , \3594 , \2210 );
nand \mul_6_18_g43067/U$1 ( \3596 , \3590 , \3595 );
xor \mul_6_18_g42715/U$1 ( \3597 , \3587 , \3596 );
not \mul_6_18_g43117/U$3 ( \3598 , \2519 );
not \mul_6_18_g43117/U$4 ( \3599 , \2511 );
or \mul_6_18_g43117/U$2 ( \3600 , \3598 , \3599 );
and \mul_6_18_g44034/U$2 ( \3601 , \2745 , \2496 );
not \mul_6_18_g44034/U$4 ( \3602 , \2745 );
and \mul_6_18_g44034/U$3 ( \3603 , \3602 , \2497 );
nor \mul_6_18_g44034/U$1 ( \3604 , \3601 , \3603 );
not \mul_6_18_g43626/U$2 ( \3605 , \3604 );
nand \mul_6_18_g43626/U$1 ( \3606 , \3605 , \2515 );
nand \mul_6_18_g43117/U$1 ( \3607 , \3600 , \3606 );
xor \mul_6_18_g42715/U$1_r1 ( \3608 , \3597 , \3607 );
xor \mul_6_18_g42374/U$1_r1 ( \3609 , \3577 , \3608 );
xor \mul_6_18_g42203/U$1_r1 ( \3610 , \3547 , \3609 );
xor \mul_6_18_g42027/U$1 ( \3611 , \3509 , \3610 );
xor \mul_6_18_g42424/U$4 ( \3612 , \3315 , \3353 );
and \mul_6_18_g42424/U$3 ( \3613 , \3612 , \3374 );
and \mul_6_18_g42424/U$5 ( \3614 , \3315 , \3353 );
or \mul_6_18_g42424/U$2 ( \3615 , \3613 , \3614 );
not \mul_6_18_g43242/U$3 ( \3616 , \3406 );
not \mul_6_18_g43242/U$4 ( \3617 , \2400 );
or \mul_6_18_g43242/U$2 ( \3618 , \3616 , \3617 );
nand \mul_6_18_g43615/U$1 ( \3619 , \2403 , \2665 );
nand \mul_6_18_g43242/U$1 ( \3620 , \3618 , \3619 );
not \mul_6_18_g43241/U$1 ( \3621 , \3620 );
not \mul_6_18_g42749/U$3 ( \3622 , \3621 );
not \mul_6_18_g43205/U$3 ( \3623 , \3390 );
not \mul_6_18_g43205/U$4 ( \3624 , \2349 );
or \mul_6_18_g43205/U$2 ( \3625 , \3623 , \3624 );
nand \mul_6_18_g43445/U$1 ( \3626 , \2359 , \2648 );
nand \mul_6_18_g43205/U$1 ( \3627 , \3625 , \3626 );
not \mul_6_18_g43204/U$1 ( \3628 , \3627 );
not \mul_6_18_g42749/U$4 ( \3629 , \3628 );
or \mul_6_18_g42749/U$2 ( \3630 , \3622 , \3629 );
not \mul_6_18_g43124/U$3 ( \3631 , \3261 );
not \mul_6_18_g43124/U$4 ( \3632 , \2511 );
or \mul_6_18_g43124/U$2 ( \3633 , \3631 , \3632 );
nand \mul_6_18_g43543/U$1 ( \3634 , \2515 , \2819 );
nand \mul_6_18_g43124/U$1 ( \3635 , \3633 , \3634 );
nand \mul_6_18_g42749/U$1 ( \3636 , \3630 , \3635 );
nand \mul_6_18_g42912/U$1 ( \3637 , \3627 , \3620 );
and \mul_6_18_g42695/U$1 ( \3638 , \3636 , \3637 );
not \mul_6_18_g42651/U$1 ( \3639 , \3638 );
not \mul_6_18_g42397/U$3 ( \3640 , \3639 );
xor \mul_6_18_g42718/U$1 ( \3641 , \2740 , \2758 );
xor \mul_6_18_g42718/U$1_r1 ( \3642 , \3641 , \2786 );
not \mul_6_18_g42397/U$4 ( \3643 , \3642 );
or \mul_6_18_g42397/U$2 ( \3644 , \3640 , \3643 );
or \mul_6_18_g42435/U$2 ( \3645 , \3642 , \3639 );
not \mul_6_18_g42878/U$3 ( \3646 , \2679 );
not \mul_6_18_g42878/U$4 ( \3647 , \2710 );
or \mul_6_18_g42878/U$2 ( \3648 , \3646 , \3647 );
nand \mul_6_18_g42893/U$1 ( \3649 , \2709 , \2658 );
nand \mul_6_18_g42878/U$1 ( \3650 , \3648 , \3649 );
and \mul_6_18_g42789/U$2 ( \3651 , \3650 , \2675 );
not \mul_6_18_g42789/U$4 ( \3652 , \3650 );
and \mul_6_18_g42789/U$3 ( \3653 , \3652 , \2674 );
nor \mul_6_18_g42789/U$1 ( \3654 , \3651 , \3653 );
nand \mul_6_18_g42435/U$1 ( \3655 , \3645 , \3654 );
nand \mul_6_18_g42397/U$1 ( \3656 , \3644 , \3655 );
xor \mul_6_18_g42195/U$4 ( \3657 , \3615 , \3656 );
xor \mul_6_18_g42422/U$1 ( \3658 , \2712 , \2789 );
xor \mul_6_18_g42422/U$1_r1 ( \3659 , \3658 , \2861 );
and \mul_6_18_g42195/U$3 ( \3660 , \3657 , \3659 );
and \mul_6_18_g42195/U$5 ( \3661 , \3615 , \3656 );
or \mul_6_18_g42195/U$2 ( \3662 , \3660 , \3661 );
not \g45623/U$3 ( \3663 , \3662 );
not \mul_6_18_g42466/U$3 ( \3664 , \3198 );
not \mul_6_18_g45210/U$2 ( \3665 , \3158 );
nand \mul_6_18_g45210/U$1 ( \3666 , \3665 , \3170 );
not \mul_6_18_g42466/U$4 ( \3667 , \3666 );
or \mul_6_18_g42466/U$2 ( \3668 , \3664 , \3667 );
nand \mul_6_18_g42910/U$1 ( \3669 , \3158 , \3167 );
nand \mul_6_18_g42466/U$1 ( \3670 , \3668 , \3669 );
not \mul_6_18_g42862/U$3 ( \3671 , \3524 );
not \mul_6_18_g42862/U$4 ( \3672 , \3532 );
and \mul_6_18_g42862/U$2 ( \3673 , \3671 , \3672 );
and \mul_6_18_g42862/U$5 ( \3674 , \3524 , \3532 );
nor \mul_6_18_g42862/U$1 ( \3675 , \3673 , \3674 );
xor \g45462/U$1 ( \3676 , \3528 , \3675 );
xor \mul_6_18_g42236/U$4 ( \3677 , \3670 , \3676 );
xor \mul_6_18_g42417/U$1 ( \3678 , \2531 , \2576 );
xor \mul_6_18_g42417/U$1_r1 ( \3679 , \3678 , \2634 );
and \mul_6_18_g42236/U$3 ( \3680 , \3677 , \3679 );
and \mul_6_18_g42236/U$5 ( \3681 , \3670 , \3676 );
or \mul_6_18_g42236/U$2 ( \3682 , \3680 , \3681 );
not \mul_6_18_g45159/U$2 ( \3683 , \3682 );
not \mul_6_18_g42486/U$3 ( \3684 , \3514 );
not \mul_6_18_g42486/U$4 ( \3685 , \3538 );
or \mul_6_18_g42486/U$2 ( \3686 , \3684 , \3685 );
nand \mul_6_18_g42501/U$1 ( \3687 , \3537 , \3513 );
nand \mul_6_18_g42486/U$1 ( \3688 , \3686 , \3687 );
not \mul_6_18_g42429/U$3 ( \3689 , \3688 );
buf \fopt45639/U$1 ( \3690 , \3517 );
not \mul_6_18_g42429/U$4 ( \3691 , \3690 );
and \mul_6_18_g42429/U$2 ( \3692 , \3689 , \3691 );
and \mul_6_18_g42429/U$5 ( \3693 , \3688 , \3690 );
nor \mul_6_18_g42429/U$1 ( \3694 , \3692 , \3693 );
nand \mul_6_18_g45159/U$1 ( \3695 , \3683 , \3694 );
not \g45623/U$4 ( \3696 , \3695 );
or \g45623/U$2 ( \3697 , \3663 , \3696 );
not \g45624/U$2 ( \3698 , \3694 );
nand \g45624/U$1 ( \3699 , \3698 , \3682 );
nand \g45623/U$1 ( \3700 , \3697 , \3699 );
xor \mul_6_18_g42027/U$1_r1 ( \3701 , \3611 , \3700 );
xor \mul_6_18_g41910/U$1_r1 ( \3702 , \3505 , \3701 );
not \mul_6_18_g42179/U$3 ( \3703 , \3694 );
not \mul_6_18_g42179/U$4 ( \3704 , \3682 );
or \mul_6_18_g42179/U$2 ( \3705 , \3703 , \3704 );
or \mul_6_18_g42179/U$5 ( \3706 , \3682 , \3694 );
nand \mul_6_18_g42179/U$1 ( \3707 , \3705 , \3706 );
and \mul_6_18_g42111/U$2 ( \3708 , \3707 , \3662 );
not \mul_6_18_g42111/U$4 ( \3709 , \3707 );
not \fopt45550/U$1 ( \3710 , \3662 );
and \mul_6_18_g42111/U$3 ( \3711 , \3709 , \3710 );
nor \mul_6_18_g42111/U$1 ( \3712 , \3708 , \3711 );
xor \mul_6_18_g42236/U$1 ( \3713 , \3670 , \3676 );
xor \mul_6_18_g42236/U$1_r1 ( \3714 , \3713 , \3679 );
not \mul_6_18_g42078/U$3 ( \3715 , \3714 );
xor \mul_6_18_g42195/U$1 ( \3716 , \3615 , \3656 );
xor \mul_6_18_g42195/U$1_r1 ( \3717 , \3716 , \3659 );
not \mul_6_18_g42078/U$4 ( \3718 , \3717 );
or \mul_6_18_g42078/U$2 ( \3719 , \3715 , \3718 );
or \mul_6_18_g42095/U$2 ( \3720 , \3717 , \3714 );
xor \g45413/U$1 ( \3721 , \3638 , \3642 );
xor \g45413/U$1_r1 ( \3722 , \3721 , \3654 );
not \mul_6_18_g42376/U$1 ( \3723 , \3722 );
not \mul_6_18_g42171/U$3 ( \3724 , \3723 );
xor \mul_6_18_g42251/U$1 ( \3725 , \3139 , \3141 );
xor \mul_6_18_g42251/U$1_r1 ( \3726 , \3725 , \3203 );
not \mul_6_18_g42249/U$1 ( \3727 , \3726 );
not \mul_6_18_g42171/U$4 ( \3728 , \3727 );
or \mul_6_18_g42171/U$2 ( \3729 , \3724 , \3728 );
not \mul_6_18_g42188/U$3 ( \3730 , \3722 );
not \mul_6_18_g42188/U$4 ( \3731 , \3726 );
or \mul_6_18_g42188/U$2 ( \3732 , \3730 , \3731 );
not \mul_6_18_g42875/U$3 ( \3733 , \3620 );
not \mul_6_18_g42875/U$4 ( \3734 , \3628 );
or \mul_6_18_g42875/U$2 ( \3735 , \3733 , \3734 );
nand \mul_6_18_g42892/U$1 ( \3736 , \3627 , \3621 );
nand \mul_6_18_g42875/U$1 ( \3737 , \3735 , \3736 );
and \mul_6_18_g42739/U$2 ( \3738 , \3737 , \3635 );
not \mul_6_18_g42739/U$4 ( \3739 , \3737 );
not \mul_6_18_g43123/U$1 ( \3740 , \3635 );
and \mul_6_18_g42739/U$3 ( \3741 , \3739 , \3740 );
nor \mul_6_18_g42739/U$1 ( \3742 , \3738 , \3741 );
xor \mul_6_18_g42623/U$1 ( \3743 , \3328 , \3340 );
xor \mul_6_18_g42623/U$1_r1 ( \3744 , \3743 , \3350 );
xor \mul_6_18_g42421/U$4 ( \3745 , \3742 , \3744 );
xor \mul_6_18_g42585/U$1 ( \3746 , \3359 , \3369 );
xor \mul_6_18_g42585/U$1_r1 ( \3747 , \3746 , \3371 );
and \mul_6_18_g42421/U$3 ( \3748 , \3745 , \3747 );
and \mul_6_18_g42421/U$5 ( \3749 , \3742 , \3744 );
or \mul_6_18_g42421/U$2 ( \3750 , \3748 , \3749 );
nand \mul_6_18_g42188/U$1 ( \3751 , \3732 , \3750 );
nand \mul_6_18_g42171/U$1 ( \3752 , \3729 , \3751 );
nand \mul_6_18_g42095/U$1 ( \3753 , \3720 , \3752 );
nand \mul_6_18_g42078/U$1 ( \3754 , \3719 , \3753 );
xor \mul_6_18_g41970/U$4 ( \3755 , \3712 , \3754 );
xor \mul_6_18_g42045/U$1 ( \3756 , \3096 , \3129 );
xor \mul_6_18_g42045/U$1_r1 ( \3757 , \3756 , \3501 );
and \mul_6_18_g41970/U$3 ( \3758 , \3755 , \3757 );
and \mul_6_18_g41970/U$5 ( \3759 , \3712 , \3754 );
or \mul_6_18_g41970/U$2 ( \3760 , \3758 , \3759 );
nor \mul_6_18_g41873/U$1 ( \3761 , \3702 , \3760 );
xor \mul_6_18_g41970/U$1 ( \3762 , \3712 , \3754 );
xor \mul_6_18_g41970/U$1_r1 ( \3763 , \3762 , \3757 );
not \mul_6_18_g41937/U$2 ( \3764 , \3763 );
and \mul_6_18_g42207/U$2 ( \3765 , \3132 , \3499 );
not \mul_6_18_g42207/U$4 ( \3766 , \3132 );
and \mul_6_18_g42207/U$3 ( \3767 , \3766 , \3206 );
nor \mul_6_18_g42207/U$1 ( \3768 , \3765 , \3767 );
not \mul_6_18_g42228/U$1 ( \3769 , \3496 );
and \mul_6_18_g42137/U$2 ( \3770 , \3768 , \3769 );
not \mul_6_18_g42137/U$4 ( \3771 , \3768 );
and \mul_6_18_g42137/U$3 ( \3772 , \3771 , \3496 );
nor \mul_6_18_g42137/U$1 ( \3773 , \3770 , \3772 );
and \mul_6_18_g43959/U$2 ( \3774 , \2116 , \2182 );
not \mul_6_18_g43959/U$4 ( \3775 , \2116 );
and \mul_6_18_g43959/U$3 ( \3776 , \3775 , \2181 );
nor \mul_6_18_g43959/U$1 ( \3777 , \3774 , \3776 );
not \mul_6_18_g43073/U$3 ( \3778 , \3777 );
not \mul_6_18_g43073/U$4 ( \3779 , \2202 );
or \mul_6_18_g43073/U$2 ( \3780 , \3778 , \3779 );
nand \mul_6_18_g43630/U$1 ( \3781 , \3364 , \2210 );
nand \mul_6_18_g43073/U$1 ( \3782 , \3780 , \3781 );
not \mul_6_18_g43372/U$3 ( \3783 , \2244 );
not \mul_6_18_g43372/U$4 ( \3784 , \3426 );
or \mul_6_18_g43372/U$2 ( \3785 , \3783 , \3784 );
not \mul_6_18_g43866/U$3 ( \3786 , \2099 );
not \mul_6_18_g43866/U$4 ( \3787 , \2217 );
or \mul_6_18_g43866/U$2 ( \3788 , \3786 , \3787 );
not \mul_6_18_g45267/U$2 ( \3789 , \2099 );
nand \mul_6_18_g45267/U$1 ( \3790 , \3789 , \2216 );
nand \mul_6_18_g43866/U$1 ( \3791 , \3788 , \3790 );
nand \mul_6_18_g43608/U$1 ( \3792 , \2222 , \3791 );
nand \mul_6_18_g43372/U$1 ( \3793 , \3785 , \3792 );
and \mul_6_18_g43916/U$2 ( \3794 , \2670 , \2256 );
not \mul_6_18_g43916/U$4 ( \3795 , \2670 );
and \mul_6_18_g43916/U$3 ( \3796 , \3795 , \2277 );
nor \mul_6_18_g43916/U$1 ( \3797 , \3794 , \3796 );
not \mul_6_18_g43915/U$1 ( \3798 , \3797 );
not \mul_6_18_g43301/U$3 ( \3799 , \3798 );
not \mul_6_18_g43301/U$4 ( \3800 , \2273 );
or \mul_6_18_g43301/U$2 ( \3801 , \3799 , \3800 );
nand \mul_6_18_g43546/U$1 ( \3802 , \3445 , \3449 );
nand \mul_6_18_g43301/U$1 ( \3803 , \3801 , \3802 );
xor \mul_6_18_g42655/U$4 ( \3804 , \3793 , \3803 );
not \mul_6_18_g44060/U$3 ( \3805 , \2112 );
not \mul_6_18_g44060/U$4 ( \3806 , \3237 );
or \mul_6_18_g44060/U$2 ( \3807 , \3805 , \3806 );
nand \mul_6_18_g44303/U$1 ( \3808 , \2307 , \2824 );
nand \mul_6_18_g44060/U$1 ( \3809 , \3807 , \3808 );
not \mul_6_18_g43164/U$3 ( \3810 , \3809 );
not \mul_6_18_g43164/U$4 ( \3811 , \2303 );
or \mul_6_18_g43164/U$2 ( \3812 , \3810 , \3811 );
nand \mul_6_18_g43547/U$1 ( \3813 , \3460 , \2318 );
nand \mul_6_18_g43164/U$1 ( \3814 , \3812 , \3813 );
and \mul_6_18_g42655/U$3 ( \3815 , \3804 , \3814 );
and \mul_6_18_g42655/U$5 ( \3816 , \3793 , \3803 );
or \mul_6_18_g42655/U$2 ( \3817 , \3815 , \3816 );
xor \mul_6_18_g42380/U$4 ( \3818 , \3782 , \3817 );
and \mul_6_18_g43646/U$1 ( \3819 , \2201 , \2058 );
not \mul_6_18_g43899/U$3 ( \3820 , \2110 );
not \mul_6_18_g43899/U$4 ( \3821 , \2909 );
or \mul_6_18_g43899/U$2 ( \3822 , \3820 , \3821 );
nand \mul_6_18_g44221/U$1 ( \3823 , \2606 , \2369 );
nand \mul_6_18_g43899/U$1 ( \3824 , \3822 , \3823 );
not \mul_6_18_g42982/U$3 ( \3825 , \3824 );
not \fopt45569/U$1 ( \3826 , \2602 );
not \mul_6_18_g42982/U$4 ( \3827 , \3826 );
or \mul_6_18_g42982/U$2 ( \3828 , \3825 , \3827 );
nand \mul_6_18_g43030/U$1 ( \3829 , \3296 , \2842 );
nand \mul_6_18_g42982/U$1 ( \3830 , \3828 , \3829 );
xor \mul_6_18_g42548/U$4 ( \3831 , \3819 , \3830 );
not \mul_6_18_g43882/U$3 ( \3832 , \2105 );
not \mul_6_18_g43882/U$4 ( \3833 , \2423 );
or \mul_6_18_g43882/U$2 ( \3834 , \3832 , \3833 );
nand \mul_6_18_g44207/U$1 ( \3835 , \2424 , \2568 );
nand \mul_6_18_g43882/U$1 ( \3836 , \3834 , \3835 );
not \mul_6_18_g42937/U$3 ( \3837 , \3836 );
not \mul_6_18_g42937/U$4 ( \3838 , \2586 );
or \mul_6_18_g42937/U$2 ( \3839 , \3837 , \3838 );
nand \mul_6_18_g43029/U$1 ( \3840 , \2434 , \3286 );
nand \mul_6_18_g42937/U$1 ( \3841 , \3839 , \3840 );
and \mul_6_18_g42548/U$3 ( \3842 , \3831 , \3841 );
and \mul_6_18_g42548/U$5 ( \3843 , \3819 , \3830 );
or \mul_6_18_g42548/U$2 ( \3844 , \3842 , \3843 );
and \mul_6_18_g42380/U$3 ( \3845 , \3818 , \3844 );
and \mul_6_18_g42380/U$5 ( \3846 , \3782 , \3817 );
or \mul_6_18_g42380/U$2 ( \3847 , \3845 , \3846 );
not \fopt45638/U$1 ( \3848 , \3847 );
not \mul_6_18_g42285/U$3 ( \3849 , \3848 );
xor \mul_6_18_g42455/U$1 ( \3850 , \3454 , \3490 );
xnor \mul_6_18_g42455/U$1_r1 ( \3851 , \3850 , \3421 );
not \mul_6_18_g42285/U$4 ( \3852 , \3851 );
or \mul_6_18_g42285/U$2 ( \3853 , \3849 , \3852 );
xor \mul_6_18_g42713/U$1 ( \3854 , \3432 , \3439 );
xor \mul_6_18_g42713/U$1_r1 ( \3855 , \3854 , \3451 );
not \mul_6_18_g43975/U$3 ( \3856 , \2092 );
not \mul_6_18_g43975/U$4 ( \3857 , \2364 );
or \mul_6_18_g43975/U$2 ( \3858 , \3856 , \3857 );
nand \mul_6_18_g44256/U$1 ( \3859 , \2363 , \2754 );
nand \mul_6_18_g43975/U$1 ( \3860 , \3858 , \3859 );
and \mul_6_18_g43228/U$2 ( \3861 , \2400 , \3860 );
and \mul_6_18_g43228/U$3 ( \3862 , \2403 , \3398 );
nor \mul_6_18_g43228/U$1 ( \3863 , \3861 , \3862 );
not \mul_6_18_g43227/U$1 ( \3864 , \3863 );
not \mul_6_18_g42692/U$3 ( \3865 , \3864 );
not \mul_6_18_g44008/U$3 ( \3866 , \2111 );
not \mul_6_18_g44008/U$4 ( \3867 , \2330 );
or \mul_6_18_g44008/U$2 ( \3868 , \3866 , \3867 );
nand \mul_6_18_g44288/U$1 ( \3869 , \2329 , \2779 );
nand \mul_6_18_g44008/U$1 ( \3870 , \3868 , \3869 );
not \mul_6_18_g43191/U$3 ( \3871 , \3870 );
not \mul_6_18_g43191/U$4 ( \3872 , \2349 );
or \mul_6_18_g43191/U$2 ( \3873 , \3871 , \3872 );
nand \mul_6_18_g43554/U$1 ( \3874 , \2359 , \3382 );
nand \mul_6_18_g43191/U$1 ( \3875 , \3873 , \3874 );
not \mul_6_18_g42692/U$4 ( \3876 , \3875 );
or \mul_6_18_g42692/U$2 ( \3877 , \3865 , \3876 );
not \mul_6_18_g42746/U$3 ( \3878 , \3863 );
not \mul_6_18_g43190/U$1 ( \3879 , \3875 );
not \mul_6_18_g42746/U$4 ( \3880 , \3879 );
or \mul_6_18_g42746/U$2 ( \3881 , \3878 , \3880 );
not \mul_6_18_g44127/U$3 ( \3882 , \2006 );
not \mul_6_18_fopt45110/U$1 ( \3883 , \3257 );
not \mul_6_18_g44127/U$4 ( \3884 , \3883 );
or \mul_6_18_g44127/U$2 ( \3885 , \3882 , \3884 );
nand \mul_6_18_g44356/U$1 ( \3886 , \2817 , \2795 );
nand \mul_6_18_g44127/U$1 ( \3887 , \3885 , \3886 );
not \mul_6_18_g43116/U$3 ( \3888 , \3887 );
not \mul_6_18_g43116/U$4 ( \3889 , \2511 );
or \mul_6_18_g43116/U$2 ( \3890 , \3888 , \3889 );
nand \mul_6_18_g43434/U$1 ( \3891 , \2515 , \3253 );
nand \mul_6_18_g43116/U$1 ( \3892 , \3890 , \3891 );
nand \mul_6_18_g42746/U$1 ( \3893 , \3881 , \3892 );
nand \mul_6_18_g42692/U$1 ( \3894 , \3877 , \3893 );
xor \mul_6_18_g42402/U$4 ( \3895 , \3855 , \3894 );
not \mul_6_18_g43947/U$3 ( \3896 , \2305 );
not \mul_6_18_g43947/U$4 ( \3897 , \2715 );
or \mul_6_18_g43947/U$2 ( \3898 , \3896 , \3897 );
not \mul_6_18_g44541/U$1 ( \3899 , \2113 );
nand \mul_6_18_g44249/U$1 ( \3900 , \2714 , \3899 );
nand \mul_6_18_g43947/U$1 ( \3901 , \3898 , \3900 );
not \mul_6_18_g43263/U$3 ( \3902 , \3901 );
not \mul_6_18_g43263/U$4 ( \3903 , \2729 );
or \mul_6_18_g43263/U$2 ( \3904 , \3902 , \3903 );
not \mul_6_18_g43919/U$1 ( \3905 , \3471 );
nand \mul_6_18_g43490/U$1 ( \3906 , \3905 , \2733 );
nand \mul_6_18_g43263/U$1 ( \3907 , \3904 , \3906 );
not \mul_6_18_g44155/U$3 ( \3908 , \2168 );
not \mul_6_18_g44155/U$4 ( \3909 , \2993 );
or \mul_6_18_g44155/U$2 ( \3910 , \3908 , \3909 );
nand \mul_6_18_g44366/U$1 ( \3911 , \2697 , \3154 );
nand \mul_6_18_g44155/U$1 ( \3912 , \3910 , \3911 );
not \mul_6_18_g43100/U$3 ( \3913 , \3912 );
not \mul_6_18_g43100/U$4 ( \3914 , \2691 );
or \mul_6_18_g43100/U$2 ( \3915 , \3913 , \3914 );
nand \mul_6_18_g43561/U$1 ( \3916 , \3413 , \2701 );
nand \mul_6_18_g43100/U$1 ( \3917 , \3915 , \3916 );
xor \mul_6_18_g42648/U$4 ( \3918 , \3907 , \3917 );
not \mul_6_18_g44100/U$3 ( \3919 , \1998 );
not \mul_6_18_g44502/U$1 ( \3920 , \2761 );
not \mul_6_18_g44100/U$4 ( \3921 , \3920 );
or \mul_6_18_g44100/U$2 ( \3922 , \3919 , \3921 );
nand \mul_6_18_g44315/U$1 ( \3923 , \3330 , \2489 );
nand \mul_6_18_g44100/U$1 ( \3924 , \3922 , \3923 );
not \mul_6_18_g43137/U$3 ( \3925 , \3924 );
not \mul_6_18_g43137/U$4 ( \3926 , \2773 );
or \mul_6_18_g43137/U$2 ( \3927 , \3925 , \3926 );
nand \mul_6_18_g43551/U$1 ( \3928 , \2784 , \3483 );
nand \mul_6_18_g43137/U$1 ( \3929 , \3927 , \3928 );
and \mul_6_18_g42648/U$3 ( \3930 , \3918 , \3929 );
and \mul_6_18_g42648/U$5 ( \3931 , \3907 , \3917 );
or \mul_6_18_g42648/U$2 ( \3932 , \3930 , \3931 );
and \mul_6_18_g42402/U$3 ( \3933 , \3895 , \3932 );
and \mul_6_18_g42402/U$5 ( \3934 , \3855 , \3894 );
or \mul_6_18_g42402/U$2 ( \3935 , \3933 , \3934 );
nand \mul_6_18_g42285/U$1 ( \3936 , \3853 , \3935 );
not \mul_6_18_g45175/U$2 ( \3937 , \3851 );
not \fopt45637/U$1 ( \3938 , \3848 );
nand \mul_6_18_g45175/U$1 ( \3939 , \3937 , \3938 );
and \mul_6_18_g42245/U$1 ( \3940 , \3936 , \3939 );
xor \mul_6_18_g45176/U$1 ( \3941 , \3493 , \3310 );
xor \mul_6_18_g45176/U$1_r1 ( \3942 , \3941 , \3375 );
xor \mul_6_18_g42081/U$4 ( \3943 , \3940 , \3942 );
xor \mul_6_18_g42421/U$1 ( \3944 , \3742 , \3744 );
xor \mul_6_18_g42421/U$1_r1 ( \3945 , \3944 , \3747 );
not \mul_6_18_g42419/U$1 ( \3946 , \3945 );
xor \mul_6_18_g42662/U$1 ( \3947 , \3279 , \3263 );
xnor \mul_6_18_g42662/U$1_r1 ( \3948 , \3947 , \3302 );
xor \mul_6_18_g42730/U$1 ( \3949 , \3392 , \3408 );
xor \mul_6_18_g42730/U$1_r1 ( \3950 , \3949 , \3418 );
not \mul_6_18_g42729/U$1 ( \3951 , \3950 );
nand \mul_6_18_g42499/U$1 ( \3952 , \3948 , \3951 );
not \mul_6_18_g42874/U$3 ( \3953 , \3475 );
not \mul_6_18_g43165/U$1 ( \3954 , \3465 );
not \mul_6_18_g42874/U$4 ( \3955 , \3954 );
or \mul_6_18_g42874/U$2 ( \3956 , \3953 , \3955 );
not \mul_6_18_g42880/U$2 ( \3957 , \3475 );
nand \mul_6_18_g42880/U$1 ( \3958 , \3957 , \3465 );
nand \mul_6_18_g42874/U$1 ( \3959 , \3956 , \3958 );
not \mul_6_18_g43138/U$1 ( \3960 , \3488 );
and \mul_6_18_g42740/U$2 ( \3961 , \3959 , \3960 );
not \mul_6_18_g42740/U$4 ( \3962 , \3959 );
and \mul_6_18_g42740/U$3 ( \3963 , \3962 , \3488 );
nor \mul_6_18_g42740/U$1 ( \3964 , \3961 , \3963 );
not \mul_6_18_g42638/U$1 ( \3965 , \3964 );
and \mul_6_18_g42439/U$2 ( \3966 , \3952 , \3965 );
nor \mul_6_18_g42498/U$1 ( \3967 , \3948 , \3951 );
nor \mul_6_18_g42439/U$1 ( \3968 , \3966 , \3967 );
buf \mul_6_18_g42403/U$1 ( \3969 , \3968 );
nand \mul_6_18_g42345/U$1 ( \3970 , \3946 , \3969 );
xor \mul_6_18_g42370/U$1 ( \3971 , \3210 , \3247 );
xor \mul_6_18_g42370/U$1_r1 ( \3972 , \3971 , \3306 );
and \mul_6_18_g42295/U$2 ( \3973 , \3970 , \3972 );
nor \mul_6_18_g42344/U$1 ( \3974 , \3946 , \3969 );
nor \mul_6_18_g42295/U$1 ( \3975 , \3973 , \3974 );
and \mul_6_18_g42081/U$3 ( \3976 , \3943 , \3975 );
and \mul_6_18_g42081/U$5 ( \3977 , \3940 , \3942 );
or \mul_6_18_g42081/U$2 ( \3978 , \3976 , \3977 );
xor \mul_6_18_g41991/U$4 ( \3979 , \3773 , \3978 );
xor \mul_6_18_g42089/U$1 ( \3980 , \3714 , \3717 );
xnor \mul_6_18_g42089/U$1_r1 ( \3981 , \3980 , \3752 );
and \mul_6_18_g41991/U$3 ( \3982 , \3979 , \3981 );
and \mul_6_18_g41991/U$5 ( \3983 , \3773 , \3978 );
or \mul_6_18_g41991/U$2 ( \3984 , \3982 , \3983 );
nand \mul_6_18_g41937/U$1 ( \3985 , \3764 , \3984 );
xor \mul_6_18_g41991/U$1 ( \3986 , \3773 , \3978 );
xor \mul_6_18_g41991/U$1_r1 ( \3987 , \3986 , \3981 );
not \mul_6_18_g42304/U$3 ( \3988 , \3750 );
not \mul_6_18_g42304/U$4 ( \3989 , \3722 );
or \mul_6_18_g42304/U$2 ( \3990 , \3988 , \3989 );
or \mul_6_18_g42304/U$5 ( \3991 , \3750 , \3722 );
nand \mul_6_18_g42304/U$1 ( \3992 , \3990 , \3991 );
and \mul_6_18_g42211/U$2 ( \3993 , \3992 , \3726 );
not \mul_6_18_g42211/U$4 ( \3994 , \3992 );
and \mul_6_18_g42211/U$3 ( \3995 , \3994 , \3727 );
nor \mul_6_18_g42211/U$1 ( \3996 , \3993 , \3995 );
and \g45514/U$2 ( \3997 , \2106 , \3186 );
not \g45514/U$4 ( \3998 , \2106 );
and \g45514/U$3 ( \3999 , \3998 , \2606 );
or \g45514/U$1 ( \4000 , \3997 , \3999 );
not \mul_6_18_g42988/U$3 ( \4001 , \4000 );
not \fopt45580/U$1 ( \4002 , \2601 );
not \mul_6_18_g42988/U$4 ( \4003 , \4002 );
or \mul_6_18_g42988/U$2 ( \4004 , \4001 , \4003 );
not \mul_6_18_g43409/U$1 ( \4005 , \2621 );
nand \mul_6_18_g43035/U$1 ( \4006 , \4005 , \3824 );
nand \mul_6_18_g42988/U$1 ( \4007 , \4004 , \4006 );
not \mul_6_18_g45005/U$1 ( \4008 , \2418 );
and \g45870/U$2 ( \4009 , \2114 , \4008 );
not \g45870/U$4 ( \4010 , \2114 );
and \g45870/U$3 ( \4011 , \4010 , \2418 );
or \g45870/U$1 ( \4012 , \4009 , \4011 );
not \mul_6_18_g42941/U$3 ( \4013 , \4012 );
not \mul_6_18_g43329/U$1 ( \4014 , \2447 );
not \mul_6_18_g42941/U$4 ( \4015 , \4014 );
or \mul_6_18_g42941/U$2 ( \4016 , \4013 , \4015 );
nand \mul_6_18_g43036/U$1 ( \4017 , \2434 , \3836 );
nand \mul_6_18_g42941/U$1 ( \4018 , \4016 , \4017 );
nand \mul_6_18_g42852/U$1 ( \4019 , \4007 , \4018 );
not \mul_6_18_g44123/U$3 ( \4020 , \3360 );
not \mul_6_18_g44123/U$4 ( \4021 , \2475 );
or \mul_6_18_g44123/U$2 ( \4022 , \4020 , \4021 );
nand \mul_6_18_g44334/U$1 ( \4023 , \2195 , \2056 );
nand \mul_6_18_g44123/U$1 ( \4024 , \4022 , \4023 );
and \mul_6_18_g43087/U$2 ( \4025 , \2481 , \4024 );
and \mul_6_18_g43087/U$3 ( \4026 , \3268 , \2480 );
nor \mul_6_18_g43087/U$1 ( \4027 , \4025 , \4026 );
nand \mul_6_18_g42666/U$1 ( \4028 , \4019 , \4027 );
not \mul_6_18_g42461/U$3 ( \4029 , \4028 );
not \mul_6_18_g43946/U$3 ( \4030 , \2640 );
not \mul_6_18_g43946/U$4 ( \4031 , \2715 );
or \mul_6_18_g43946/U$2 ( \4032 , \4030 , \4031 );
nand \mul_6_18_g44252/U$1 ( \4033 , \2714 , \2639 );
nand \mul_6_18_g43946/U$1 ( \4034 , \4032 , \4033 );
not \mul_6_18_g43267/U$3 ( \4035 , \4034 );
not \mul_6_18_g43267/U$4 ( \4036 , \2965 );
or \mul_6_18_g43267/U$2 ( \4037 , \4035 , \4036 );
nand \mul_6_18_g43529/U$1 ( \4038 , \3326 , \3901 );
nand \mul_6_18_g43267/U$1 ( \4039 , \4037 , \4038 );
not \mul_6_18_g43266/U$1 ( \4040 , \4039 );
not \mul_6_18_g42750/U$3 ( \4041 , \4040 );
not \mul_6_18_g44061/U$3 ( \4042 , \2812 );
not \mul_6_18_g44061/U$4 ( \4043 , \3237 );
or \mul_6_18_g44061/U$2 ( \4044 , \4042 , \4043 );
not \mul_6_18_g45274/U$2 ( \4045 , \2296 );
nand \mul_6_18_g45274/U$1 ( \4046 , \4045 , \2811 );
nand \mul_6_18_g44061/U$1 ( \4047 , \4044 , \4046 );
not \mul_6_18_g43169/U$3 ( \4048 , \4047 );
not \mul_6_18_g43457/U$1 ( \4049 , \2301 );
not \mul_6_18_g43169/U$4 ( \4050 , \4049 );
or \mul_6_18_g43169/U$2 ( \4051 , \4048 , \4050 );
nand \mul_6_18_g43586/U$1 ( \4052 , \2317 , \3809 );
nand \mul_6_18_g43169/U$1 ( \4053 , \4051 , \4052 );
not \mul_6_18_g43168/U$1 ( \4054 , \4053 );
not \mul_6_18_g42750/U$4 ( \4055 , \4054 );
or \mul_6_18_g42750/U$2 ( \4056 , \4041 , \4055 );
not \mul_6_18_g44101/U$3 ( \4057 , \2463 );
not \mul_6_18_g44101/U$4 ( \4058 , \3920 );
or \mul_6_18_g44101/U$2 ( \4059 , \4057 , \4058 );
nand \mul_6_18_g44323/U$1 ( \4060 , \3330 , \2468 );
nand \mul_6_18_g44101/U$1 ( \4061 , \4059 , \4060 );
not \mul_6_18_g43141/U$3 ( \4062 , \4061 );
not \mul_6_18_g43141/U$4 ( \4063 , \2771 );
or \mul_6_18_g43141/U$2 ( \4064 , \4062 , \4063 );
nand \mul_6_18_g43562/U$1 ( \4065 , \3924 , \2783 );
nand \mul_6_18_g43141/U$1 ( \4066 , \4064 , \4065 );
nand \mul_6_18_g42750/U$1 ( \4067 , \4056 , \4066 );
nand \mul_6_18_g42913/U$1 ( \4068 , \4039 , \4053 );
nand \mul_6_18_g42694/U$1 ( \4069 , \4067 , \4068 );
not \mul_6_18_g42461/U$4 ( \4070 , \4069 );
or \mul_6_18_g42461/U$2 ( \4071 , \4029 , \4070 );
not \mul_6_18_g45212/U$2 ( \4072 , \4027 );
not \mul_6_18_g42775/U$1 ( \4073 , \4019 );
nand \mul_6_18_g45212/U$1 ( \4074 , \4072 , \4073 );
nand \mul_6_18_g42461/U$1 ( \4075 , \4071 , \4074 );
and \mul_6_18_g44395/U$1 ( \4076 , \2242 , \2216 );
not \mul_6_18_g43379/U$3 ( \4077 , \4076 );
and \g45507/U$2 ( \4078 , \2100 , \3211 );
not \g45507/U$4 ( \4079 , \2100 );
and \g45507/U$3 ( \4080 , \4079 , \2216 );
or \g45507/U$1 ( \4081 , \4078 , \4080 );
not \mul_6_18_g43379/U$4 ( \4082 , \4081 );
or \mul_6_18_g43379/U$2 ( \4083 , \4077 , \4082 );
nand \mul_6_18_g43606/U$1 ( \4084 , \3791 , \2934 );
nand \mul_6_18_g43379/U$1 ( \4085 , \4083 , \4084 );
nor \mul_6_18_g44170/U$1 ( \4086 , \2473 , \2058 );
not \mul_6_18_g43685/U$3 ( \4087 , \4086 );
not \mul_6_18_g43685/U$4 ( \4088 , \2694 );
and \mul_6_18_g43685/U$2 ( \4089 , \4087 , \4088 );
not \mul_6_18_g43730/U$3 ( \4090 , \2058 );
not \mul_6_18_g43730/U$4 ( \4091 , \2473 );
or \mul_6_18_g43730/U$2 ( \4092 , \4090 , \4091 );
nand \mul_6_18_g43730/U$1 ( \4093 , \4092 , \2196 );
nor \mul_6_18_g43685/U$1 ( \4094 , \4089 , \4093 );
xor \mul_6_18_g42703/U$4 ( \4095 , \4085 , \4094 );
and \g45517/U$2 ( \4096 , \1970 , \2251 );
not \g45517/U$4 ( \4097 , \1970 );
and \g45517/U$3 ( \4098 , \4097 , \2256 );
or \g45517/U$1 ( \4099 , \4096 , \4098 );
not \g5/U$3 ( \4100 , \4099 );
not \g5/U$4 ( \4101 , \2273 );
or \g5/U$2 ( \4102 , \4100 , \4101 );
or \g6/U$1 ( \4103 , \3797 , \2284 );
nand \g5/U$1 ( \4104 , \4102 , \4103 );
and \mul_6_18_g42703/U$3 ( \4105 , \4095 , \4104 );
and \mul_6_18_g42703/U$5 ( \4106 , \4085 , \4094 );
or \mul_6_18_g42703/U$2 ( \4107 , \4105 , \4106 );
not \mul_6_18_g43973/U$3 ( \4108 , \2107 );
not \mul_6_18_g43973/U$4 ( \4109 , \2367 );
or \mul_6_18_g43973/U$2 ( \4110 , \4108 , \4109 );
nand \mul_6_18_g44267/U$1 ( \4111 , \2363 , \2745 );
nand \mul_6_18_g43973/U$1 ( \4112 , \4110 , \4111 );
not \mul_6_18_g43237/U$3 ( \4113 , \4112 );
not \mul_6_18_g43237/U$4 ( \4114 , \2399 );
or \mul_6_18_g43237/U$2 ( \4115 , \4113 , \4114 );
nand \mul_6_18_g43452/U$1 ( \4116 , \2403 , \3860 );
nand \mul_6_18_g43237/U$1 ( \4117 , \4115 , \4116 );
not \mul_6_18_g43236/U$1 ( \4118 , \4117 );
not \mul_6_18_g42858/U$3 ( \4119 , \4118 );
nor \mul_6_18_g43473/U$1 ( \4120 , \2341 , \2347 );
not \mul_6_18_g44009/U$3 ( \4121 , \2094 );
not \mul_6_18_g44009/U$4 ( \4122 , \2644 );
or \mul_6_18_g44009/U$2 ( \4123 , \4121 , \4122 );
nand \mul_6_18_g44286/U$1 ( \4124 , \2329 , \2500 );
nand \mul_6_18_g44009/U$1 ( \4125 , \4123 , \4124 );
and \mul_6_18_g43201/U$2 ( \4126 , \4120 , \4125 );
and \mul_6_18_g43201/U$3 ( \4127 , \2358 , \3870 );
nor \mul_6_18_g43201/U$1 ( \4128 , \4126 , \4127 );
not \mul_6_18_g42858/U$4 ( \4129 , \4128 );
or \mul_6_18_g42858/U$2 ( \4130 , \4119 , \4129 );
not \mul_6_18_g44154/U$3 ( \4131 , \2144 );
not \mul_6_18_g44154/U$4 ( \4132 , \2687 );
or \mul_6_18_g44154/U$2 ( \4133 , \4131 , \4132 );
nand \mul_6_18_g44362/U$1 ( \4134 , \2697 , \2145 );
nand \mul_6_18_g44154/U$1 ( \4135 , \4133 , \4134 );
not \mul_6_18_g43092/U$3 ( \4136 , \4135 );
not \mul_6_18_g43092/U$4 ( \4137 , \2691 );
or \mul_6_18_g43092/U$2 ( \4138 , \4136 , \4137 );
nand \mul_6_18_g43441/U$1 ( \4139 , \2701 , \3912 );
nand \mul_6_18_g43092/U$1 ( \4140 , \4138 , \4139 );
nand \mul_6_18_g42858/U$1 ( \4141 , \4130 , \4140 );
not \mul_6_18_g45216/U$2 ( \4142 , \4118 );
not \mul_6_18_g43200/U$1 ( \4143 , \4128 );
nand \mul_6_18_g45216/U$1 ( \4144 , \4142 , \4143 );
nand \mul_6_18_g42809/U$1 ( \4145 , \4141 , \4144 );
xor \mul_6_18_g42326/U$4 ( \4146 , \4107 , \4145 );
xor \mul_6_18_g42548/U$1 ( \4147 , \3819 , \3830 );
xor \mul_6_18_g42548/U$1_r1 ( \4148 , \4147 , \3841 );
and \mul_6_18_g42326/U$3 ( \4149 , \4146 , \4148 );
and \mul_6_18_g42326/U$5 ( \4150 , \4107 , \4145 );
or \mul_6_18_g42326/U$2 ( \4151 , \4149 , \4150 );
xor \mul_6_18_g42172/U$4 ( \4152 , \4075 , \4151 );
xor \mul_6_18_g42380/U$1 ( \4153 , \3782 , \3817 );
xor \mul_6_18_g42380/U$1_r1 ( \4154 , \4153 , \3844 );
and \mul_6_18_g42172/U$3 ( \4155 , \4152 , \4154 );
and \mul_6_18_g42172/U$5 ( \4156 , \4075 , \4151 );
or \mul_6_18_g42172/U$2 ( \4157 , \4155 , \4156 );
xor \mul_6_18_g42237/U$1 ( \4158 , \3847 , \3935 );
xnor \mul_6_18_g42237/U$1_r1 ( \4159 , \4158 , \3851 );
xor \mul_6_18_g42048/U$4 ( \4160 , \4157 , \4159 );
xor \mul_6_18_g42402/U$1 ( \4161 , \3855 , \3894 );
xor \mul_6_18_g42402/U$1_r1 ( \4162 , \4161 , \3932 );
xor \mul_6_18_g42655/U$1 ( \4163 , \3793 , \3803 );
xor \mul_6_18_g42655/U$1_r1 ( \4164 , \4163 , \3814 );
xor \mul_6_18_g42648/U$1 ( \4165 , \3907 , \3917 );
xor \mul_6_18_g42648/U$1_r1 ( \4166 , \4165 , \3929 );
xor \mul_6_18_g42410/U$4 ( \4167 , \4164 , \4166 );
xor \g45744/U$1 ( \4168 , \3864 , \3879 );
xnor \g45744/U$1_r1 ( \4169 , \4168 , \3892 );
and \mul_6_18_g42410/U$3 ( \4170 , \4167 , \4169 );
and \mul_6_18_g42410/U$5 ( \4171 , \4164 , \4166 );
or \mul_6_18_g42410/U$2 ( \4172 , \4170 , \4171 );
xor \mul_6_18_g42229/U$4 ( \4173 , \4162 , \4172 );
not \mul_6_18_g42527/U$3 ( \4174 , \3951 );
not \mul_6_18_g42527/U$4 ( \4175 , \3965 );
or \mul_6_18_g42527/U$2 ( \4176 , \4174 , \4175 );
nand \mul_6_18_g42537/U$1 ( \4177 , \3950 , \3964 );
nand \mul_6_18_g42527/U$1 ( \4178 , \4176 , \4177 );
not \mul_6_18_g42581/U$1 ( \4179 , \3948 );
and \mul_6_18_g42456/U$2 ( \4180 , \4178 , \4179 );
not \mul_6_18_g42456/U$4 ( \4181 , \4178 );
and \mul_6_18_g42456/U$3 ( \4182 , \4181 , \3948 );
nor \mul_6_18_g42456/U$1 ( \4183 , \4180 , \4182 );
and \mul_6_18_g42229/U$3 ( \4184 , \4173 , \4183 );
and \mul_6_18_g42229/U$5 ( \4185 , \4162 , \4172 );
or \mul_6_18_g42229/U$2 ( \4186 , \4184 , \4185 );
and \mul_6_18_g42048/U$3 ( \4187 , \4160 , \4186 );
and \mul_6_18_g42048/U$5 ( \4188 , \4157 , \4159 );
or \mul_6_18_g42048/U$2 ( \4189 , \4187 , \4188 );
not \mul_6_18_g42047/U$1 ( \4190 , \4189 );
xor \mul_6_18_g41948/U$4 ( \4191 , \3996 , \4190 );
xor \mul_6_18_g42081/U$1 ( \4192 , \3940 , \3942 );
xor \mul_6_18_g42081/U$1_r1 ( \4193 , \4192 , \3975 );
and \mul_6_18_g41948/U$3 ( \4194 , \4191 , \4193 );
and \mul_6_18_g41948/U$5 ( \4195 , \3996 , \4190 );
or \mul_6_18_g41948/U$2 ( \4196 , \4194 , \4195 );
nand \mul_6_18_g41920/U$1 ( \4197 , \3987 , \4196 );
nand \mul_6_18_g41904/U$1 ( \4198 , \3985 , \4197 );
nor \mul_6_18_g41862/U$1 ( \4199 , \3761 , \4198 );
not \mul_6_18_g41837/U$3 ( \4200 , \4199 );
xor \mul_6_18_g41948/U$1 ( \4201 , \3996 , \4190 );
xor \mul_6_18_g41948/U$1_r1 ( \4202 , \4201 , \4193 );
xor \mul_6_18_g42048/U$1 ( \4203 , \4157 , \4159 );
xor \mul_6_18_g42048/U$1_r1 ( \4204 , \4203 , \4186 );
not \mul_6_18_g42046/U$1 ( \4205 , \4204 );
or \g45681/U$2 ( \4206 , \3968 , \3972 );
nand \mul_6_18_g42315/U$1 ( \4207 , \3972 , \3968 );
nand \g45681/U$1 ( \4208 , \4206 , \4207 );
xnor \mul_6_18_g42238/U$1 ( \4209 , \4208 , \3945 );
buf \mul_6_18_fopt45113/U$1 ( \4210 , \4209 );
nand \mul_6_18_g42010/U$1 ( \4211 , \4205 , \4210 );
xor \g45521/U$1 ( \4212 , \2058 , \2196 );
not \mul_6_18_g43090/U$3 ( \4213 , \4212 );
not \mul_6_18_g43090/U$4 ( \4214 , \3270 );
or \mul_6_18_g43090/U$2 ( \4215 , \4213 , \4214 );
nand \mul_6_18_g43440/U$1 ( \4216 , \4024 , \2480 );
nand \mul_6_18_g43090/U$1 ( \4217 , \4215 , \4216 );
not \mul_6_18_g42607/U$3 ( \4218 , \4217 );
not \mul_6_18_g44128/U$3 ( \4219 , \2179 );
not \mul_6_18_g44128/U$4 ( \4220 , \3883 );
or \mul_6_18_g44128/U$2 ( \4221 , \4219 , \4220 );
nand \mul_6_18_g44349/U$1 ( \4222 , \2496 , \2185 );
nand \mul_6_18_g44128/U$1 ( \4223 , \4221 , \4222 );
not \mul_6_18_g43126/U$3 ( \4224 , \4223 );
not \mul_6_18_g43126/U$4 ( \4225 , \2510 );
or \mul_6_18_g43126/U$2 ( \4226 , \4224 , \4225 );
nand \mul_6_18_g43624/U$1 ( \4227 , \2514 , \3887 );
nand \mul_6_18_g43126/U$1 ( \4228 , \4226 , \4227 );
not \mul_6_18_g42607/U$4 ( \4229 , \4228 );
or \mul_6_18_g42607/U$2 ( \4230 , \4218 , \4229 );
not \mul_6_18_g43089/U$1 ( \4231 , \4217 );
not \mul_6_18_g42675/U$3 ( \4232 , \4231 );
not \mul_6_18_g43125/U$1 ( \4233 , \4228 );
not \mul_6_18_g42675/U$4 ( \4234 , \4233 );
or \mul_6_18_g42675/U$2 ( \4235 , \4232 , \4234 );
xor \g45478/U$1 ( \4236 , \4007 , \4018 );
nand \mul_6_18_g42675/U$1 ( \4237 , \4235 , \4236 );
nand \mul_6_18_g42607/U$1 ( \4238 , \4230 , \4237 );
not \mul_6_18_g42473/U$3 ( \4239 , \4069 );
not \mul_6_18_g42611/U$3 ( \4240 , \4073 );
not \mul_6_18_g42611/U$4 ( \4241 , \4027 );
and \mul_6_18_g42611/U$2 ( \4242 , \4240 , \4241 );
and \mul_6_18_g42611/U$5 ( \4243 , \4073 , \4027 );
nor \mul_6_18_g42611/U$1 ( \4244 , \4242 , \4243 );
not \mul_6_18_g42473/U$4 ( \4245 , \4244 );
or \mul_6_18_g42473/U$2 ( \4246 , \4239 , \4245 );
or \mul_6_18_g42473/U$5 ( \4247 , \4069 , \4244 );
nand \mul_6_18_g42473/U$1 ( \4248 , \4246 , \4247 );
xor \mul_6_18_g42233/U$4 ( \4249 , \4238 , \4248 );
and \g45516/U$2 ( \4250 , \2101 , \3186 );
not \g45516/U$4 ( \4251 , \2101 );
and \g45516/U$3 ( \4252 , \4251 , \2626 );
or \g45516/U$1 ( \4253 , \4250 , \4252 );
not \mul_6_18_g42992/U$3 ( \4254 , \4253 );
nand \mul_6_18_g43351/U$1 ( \4255 , \2596 , \2600 );
not \mul_6_18_g43349/U$1 ( \4256 , \4255 );
not \mul_6_18_g42992/U$4 ( \4257 , \4256 );
or \mul_6_18_g42992/U$2 ( \4258 , \4254 , \4257 );
nand \mul_6_18_g43028/U$1 ( \4259 , \2622 , \4000 );
nand \mul_6_18_g42992/U$1 ( \4260 , \4258 , \4259 );
not \g45800/U$3 ( \4261 , \2434 );
not \g45800/U$4 ( \4262 , \4012 );
or \g45800/U$2 ( \4263 , \4261 , \4262 );
not \mul_6_18_g43321/U$1 ( \4264 , \2446 );
not \mul_6_18_g43319/U$1 ( \4265 , \4264 );
not \g45801/U$2 ( \4266 , \4265 );
and \g45757/U$2 ( \4267 , \2110 , \2614 );
not \g45757/U$4 ( \4268 , \2110 );
and \g45757/U$3 ( \4269 , \4268 , \2418 );
or \g45757/U$1 ( \4270 , \4267 , \4269 );
nand \g45801/U$1 ( \4271 , \4266 , \4270 );
nand \g45800/U$1 ( \4272 , \4263 , \4271 );
xor \mul_6_18_g42635/U$4 ( \4273 , \4260 , \4272 );
and \mul_6_18_g43647/U$1 ( \4274 , \2480 , \2058 );
and \mul_6_18_g42635/U$3 ( \4275 , \4273 , \4274 );
and \mul_6_18_g42635/U$5 ( \4276 , \4260 , \4272 );
or \mul_6_18_g42635/U$2 ( \4277 , \4275 , \4276 );
not \mul_6_18_g44084/U$3 ( \4278 , \1998 );
not \mul_6_18_g44084/U$4 ( \4279 , \2308 );
or \mul_6_18_g44084/U$2 ( \4280 , \4278 , \4279 );
nand \mul_6_18_g44318/U$1 ( \4281 , \2307 , \2489 );
nand \mul_6_18_g44084/U$1 ( \4282 , \4280 , \4281 );
not \mul_6_18_g43173/U$3 ( \4283 , \4282 );
not \mul_6_18_g43173/U$4 ( \4284 , \4049 );
or \mul_6_18_g43173/U$2 ( \4285 , \4283 , \4284 );
buf \mul_6_18_fopt45121/U$1 ( \4286 , \2294 );
not \mul_6_18_fopt45120/U$1 ( \4287 , \4286 );
nand \mul_6_18_g43548/U$1 ( \4288 , \4287 , \4047 );
nand \mul_6_18_g43173/U$1 ( \4289 , \4285 , \4288 );
not \g45766/U$3 ( \4290 , \4289 );
and \g45519/U$2 ( \4291 , \2113 , \2251 );
not \g45519/U$4 ( \4292 , \2113 );
and \g45519/U$3 ( \4293 , \4292 , \2256 );
or \g45519/U$1 ( \4294 , \4291 , \4293 );
not \mul_6_18_g43296/U$3 ( \4295 , \4294 );
not \mul_6_18_g43296/U$4 ( \4296 , \2273 );
or \mul_6_18_g43296/U$2 ( \4297 , \4295 , \4296 );
nand \mul_6_18_g43481/U$1 ( \4298 , \4099 , \3232 );
nand \mul_6_18_g43296/U$1 ( \4299 , \4297 , \4298 );
not \mul_6_18_g43295/U$1 ( \4300 , \4299 );
not \mul_6_18_g43879/U$3 ( \4301 , \2105 );
not \mul_6_18_g43879/U$4 ( \4302 , \3211 );
or \mul_6_18_g43879/U$2 ( \4303 , \4301 , \4302 );
not \mul_6_18_g45250/U$2 ( \4304 , \2105 );
nand \mul_6_18_g45250/U$1 ( \4305 , \4304 , \2225 );
nand \mul_6_18_g43879/U$1 ( \4306 , \4303 , \4305 );
not \mul_6_18_g43355/U$3 ( \4307 , \4306 );
not \mul_6_18_g43355/U$4 ( \4308 , \4076 );
or \mul_6_18_g43355/U$2 ( \4309 , \4307 , \4308 );
nand \mul_6_18_g43549/U$1 ( \4310 , \4081 , \2244 );
nand \mul_6_18_g43355/U$1 ( \4311 , \4309 , \4310 );
not \mul_6_18_g43354/U$1 ( \4312 , \4311 );
nand \mul_6_18_g42890/U$1 ( \4313 , \4300 , \4312 );
not \g45766/U$4 ( \4314 , \4313 );
or \g45766/U$2 ( \4315 , \4290 , \4314 );
or \g45766/U$5 ( \4316 , \4312 , \4300 );
nand \g45766/U$1 ( \4317 , \4315 , \4316 );
xor \mul_6_18_g42411/U$4 ( \4318 , \4277 , \4317 );
and \mul_6_18_g43970/U$2 ( \4319 , \2092 , \2718 );
not \mul_6_18_g43970/U$4 ( \4320 , \2092 );
and \mul_6_18_g43970/U$3 ( \4321 , \4320 , \2719 );
nor \mul_6_18_g43970/U$1 ( \4322 , \4319 , \4321 );
not \mul_6_18_g43969/U$1 ( \4323 , \4322 );
not \mul_6_18_g43254/U$3 ( \4324 , \4323 );
not \mul_6_18_g43254/U$4 ( \4325 , \2965 );
or \mul_6_18_g43254/U$2 ( \4326 , \4324 , \4325 );
not \mul_6_18_g43775/U$1 ( \4327 , \2732 );
nand \mul_6_18_g43539/U$1 ( \4328 , \4327 , \4034 );
nand \mul_6_18_g43254/U$1 ( \4329 , \4326 , \4328 );
and \mul_6_18_g44148/U$2 ( \4330 , \2056 , \2705 );
not \mul_6_18_g44148/U$4 ( \4331 , \2056 );
and \mul_6_18_g44148/U$3 ( \4332 , \4331 , \2687 );
nor \mul_6_18_g44148/U$1 ( \4333 , \4330 , \4332 );
not \mul_6_18_g43094/U$3 ( \4334 , \4333 );
not \mul_6_18_g43094/U$4 ( \4335 , \2691 );
or \mul_6_18_g43094/U$2 ( \4336 , \4334 , \4335 );
nand \mul_6_18_g43572/U$1 ( \4337 , \2701 , \4135 );
nand \mul_6_18_g43094/U$1 ( \4338 , \4336 , \4337 );
xor \mul_6_18_g42637/U$4 ( \4339 , \4329 , \4338 );
not \mul_6_18_g44111/U$3 ( \4340 , \2006 );
not \mul_6_18_g44111/U$4 ( \4341 , \3331 );
or \mul_6_18_g44111/U$2 ( \4342 , \4340 , \4341 );
nand \mul_6_18_g44358/U$1 ( \4343 , \3330 , \2795 );
nand \mul_6_18_g44111/U$1 ( \4344 , \4342 , \4343 );
not \mul_6_18_g43142/U$3 ( \4345 , \4344 );
not \mul_6_18_g43142/U$4 ( \4346 , \2771 );
or \mul_6_18_g43142/U$2 ( \4347 , \4345 , \4346 );
nand \mul_6_18_g43585/U$1 ( \4348 , \2783 , \4061 );
nand \mul_6_18_g43142/U$1 ( \4349 , \4347 , \4348 );
and \mul_6_18_g42637/U$3 ( \4350 , \4339 , \4349 );
and \mul_6_18_g42637/U$5 ( \4351 , \4329 , \4338 );
or \mul_6_18_g42637/U$2 ( \4352 , \4350 , \4351 );
and \mul_6_18_g42411/U$3 ( \4353 , \4318 , \4352 );
and \mul_6_18_g42411/U$5 ( \4354 , \4277 , \4317 );
or \mul_6_18_g42411/U$2 ( \4355 , \4353 , \4354 );
and \mul_6_18_g42233/U$3 ( \4356 , \4249 , \4355 );
and \mul_6_18_g42233/U$5 ( \4357 , \4238 , \4248 );
or \mul_6_18_g42233/U$2 ( \4358 , \4356 , \4357 );
xor \mul_6_18_g42172/U$1 ( \4359 , \4075 , \4151 );
xor \mul_6_18_g42172/U$1_r1 ( \4360 , \4359 , \4154 );
xor \mul_6_18_g42050/U$4 ( \4361 , \4358 , \4360 );
xor \mul_6_18_g42326/U$1 ( \4362 , \4107 , \4145 );
xor \mul_6_18_g42326/U$1_r1 ( \4363 , \4362 , \4148 );
not \mul_6_18_g42879/U$3 ( \4364 , \4053 );
not \mul_6_18_g42879/U$4 ( \4365 , \4040 );
or \mul_6_18_g42879/U$2 ( \4366 , \4364 , \4365 );
or \mul_6_18_g42879/U$5 ( \4367 , \4040 , \4053 );
nand \mul_6_18_g42879/U$1 ( \4368 , \4366 , \4367 );
xor \mul_6_18_g42742/U$1 ( \4369 , \4368 , \4066 );
not \mul_6_18_g44044/U$3 ( \4370 , \2112 );
not \mul_6_18_g44044/U$4 ( \4371 , \2330 );
or \mul_6_18_g44044/U$2 ( \4372 , \4370 , \4371 );
nand \mul_6_18_g45806/U$1 ( \4373 , \2329 , \2824 );
nand \mul_6_18_g44044/U$1 ( \4374 , \4372 , \4373 );
not \mul_6_18_g43206/U$3 ( \4375 , \4374 );
not \mul_6_18_g43206/U$4 ( \4376 , \4120 );
or \mul_6_18_g43206/U$2 ( \4377 , \4375 , \4376 );
nand \mul_6_18_g43474/U$1 ( \4378 , \2358 , \4125 );
nand \mul_6_18_g43206/U$1 ( \4379 , \4377 , \4378 );
not \mul_6_18_g43999/U$3 ( \4380 , \2111 );
not \mul_6_18_g43999/U$4 ( \4381 , \2364 );
or \mul_6_18_g43999/U$2 ( \4382 , \4380 , \4381 );
nand \mul_6_18_g44290/U$1 ( \4383 , \2368 , \2779 );
nand \mul_6_18_g43999/U$1 ( \4384 , \4382 , \4383 );
not \mul_6_18_g43244/U$3 ( \4385 , \4384 );
not \mul_6_18_g43244/U$4 ( \4386 , \2399 );
or \mul_6_18_g43244/U$2 ( \4387 , \4385 , \4386 );
nand \mul_6_18_g43541/U$1 ( \4388 , \2403 , \4112 );
nand \mul_6_18_g43244/U$1 ( \4389 , \4387 , \4388 );
xor \mul_6_18_g42643/U$4 ( \4390 , \4379 , \4389 );
and \mul_6_18_g45293/U$2 ( \4391 , \3154 , \2495 );
not \mul_6_18_g45293/U$4 ( \4392 , \3154 );
and \mul_6_18_g45293/U$3 ( \4393 , \4392 , \3257 );
or \mul_6_18_g45293/U$1 ( \4394 , \4391 , \4393 );
not \mul_6_18_g44141/U$1 ( \4395 , \4394 );
not \mul_6_18_g43113/U$3 ( \4396 , \4395 );
not \mul_6_18_g43113/U$4 ( \4397 , \2510 );
or \mul_6_18_g43113/U$2 ( \4398 , \4396 , \4397 );
nand \mul_6_18_g43480/U$1 ( \4399 , \2515 , \4223 );
nand \mul_6_18_g43113/U$1 ( \4400 , \4398 , \4399 );
and \mul_6_18_g42643/U$3 ( \4401 , \4390 , \4400 );
and \mul_6_18_g42643/U$5 ( \4402 , \4379 , \4389 );
or \mul_6_18_g42643/U$2 ( \4403 , \4401 , \4402 );
or \mul_6_18_g42517/U$2 ( \4404 , \4369 , \4403 );
xor \mul_6_18_g42796/U$1 ( \4405 , \4117 , \4143 );
xor \mul_6_18_g42796/U$1_r1 ( \4406 , \4405 , \4140 );
nand \mul_6_18_g42517/U$1 ( \4407 , \4404 , \4406 );
nand \mul_6_18_g42539/U$1 ( \4408 , \4369 , \4403 );
nand \mul_6_18_g42472/U$1 ( \4409 , \4407 , \4408 );
xor \mul_6_18_g42177/U$4 ( \4410 , \4363 , \4409 );
xor \mul_6_18_g42410/U$1 ( \4411 , \4164 , \4166 );
xor \mul_6_18_g42410/U$1_r1 ( \4412 , \4411 , \4169 );
and \mul_6_18_g42177/U$3 ( \4413 , \4410 , \4412 );
and \mul_6_18_g42177/U$5 ( \4414 , \4363 , \4409 );
or \mul_6_18_g42177/U$2 ( \4415 , \4413 , \4414 );
and \mul_6_18_g42050/U$3 ( \4416 , \4361 , \4415 );
and \mul_6_18_g42050/U$5 ( \4417 , \4358 , \4360 );
or \mul_6_18_g42050/U$2 ( \4418 , \4416 , \4417 );
buf \mul_6_18_g42049/U$1 ( \4419 , \4418 );
and \mul_6_18_g41988/U$2 ( \4420 , \4211 , \4419 );
nor \mul_6_18_g42011/U$1 ( \4421 , \4205 , \4210 );
nor \mul_6_18_g41988/U$1 ( \4422 , \4420 , \4421 );
nand \mul_6_18_g41917/U$1 ( \4423 , \4202 , \4422 );
not \mul_6_18_g41842/U$3 ( \4424 , \4423 );
not \mul_6_18_g41971/U$3 ( \4425 , \4204 );
not \mul_6_18_g42006/U$3 ( \4426 , \4418 );
not \mul_6_18_g42006/U$4 ( \4427 , \4209 );
and \mul_6_18_g42006/U$2 ( \4428 , \4426 , \4427 );
and \mul_6_18_g42006/U$5 ( \4429 , \4418 , \4209 );
nor \mul_6_18_g42006/U$1 ( \4430 , \4428 , \4429 );
not \mul_6_18_g41971/U$4 ( \4431 , \4430 );
or \mul_6_18_g41971/U$2 ( \4432 , \4425 , \4431 );
or \mul_6_18_g41971/U$5 ( \4433 , \4430 , \4204 );
nand \mul_6_18_g41971/U$1 ( \4434 , \4432 , \4433 );
xor \mul_6_18_g42229/U$1 ( \4435 , \4162 , \4172 );
xor \mul_6_18_g42229/U$1_r1 ( \4436 , \4435 , \4183 );
xor \mul_6_18_g42703/U$1 ( \4437 , \4085 , \4094 );
xor \mul_6_18_g42703/U$1_r1 ( \4438 , \4437 , \4104 );
not \mul_6_18_g42494/U$2 ( \4439 , \4438 );
not \mul_6_18_g42861/U$3 ( \4440 , \4231 );
not \mul_6_18_g42861/U$4 ( \4441 , \4228 );
or \mul_6_18_g42861/U$2 ( \4442 , \4440 , \4441 );
nand \mul_6_18_g42884/U$1 ( \4443 , \4233 , \4217 );
nand \mul_6_18_g42861/U$1 ( \4444 , \4442 , \4443 );
not \mul_6_18_g42772/U$1 ( \4445 , \4236 );
and \mul_6_18_g42659/U$2 ( \4446 , \4444 , \4445 );
not \mul_6_18_g42659/U$4 ( \4447 , \4444 );
and \mul_6_18_g42659/U$3 ( \4448 , \4447 , \4236 );
nor \mul_6_18_g42659/U$1 ( \4449 , \4446 , \4448 );
nand \mul_6_18_g42494/U$1 ( \4450 , \4439 , \4449 );
not \mul_6_18_g43682/U$3 ( \4451 , \2495 );
nor \mul_6_18_g44162/U$1 ( \4452 , \1127 , \2058 );
not \mul_6_18_g43682/U$4 ( \4453 , \4452 );
and \mul_6_18_g43682/U$2 ( \4454 , \4451 , \4453 );
not \mul_6_18_g43727/U$3 ( \4455 , \2058 );
not \mul_6_18_g43727/U$4 ( \4456 , \1127 );
or \mul_6_18_g43727/U$2 ( \4457 , \4455 , \4456 );
nand \mul_6_18_g43727/U$1 ( \4458 , \4457 , \2684 );
nor \mul_6_18_g43682/U$1 ( \4459 , \4454 , \4458 );
and \g45756/U$2 ( \4460 , \2106 , \2423 );
not \g45756/U$4 ( \4461 , \2106 );
and \g45756/U$3 ( \4462 , \4461 , \2418 );
or \g45756/U$1 ( \4463 , \4460 , \4462 );
not \mul_6_18_g42916/U$3 ( \4464 , \4463 );
not \mul_6_18_g42916/U$4 ( \4465 , \4264 );
or \mul_6_18_g42916/U$2 ( \4466 , \4464 , \4465 );
nand \mul_6_18_g43003/U$1 ( \4467 , \2434 , \4270 );
nand \mul_6_18_g42916/U$1 ( \4468 , \4466 , \4467 );
and \mul_6_18_g42776/U$2 ( \4469 , \4459 , \4468 );
not \mul_6_18_g43247/U$3 ( \4470 , \2964 );
and \g45854/U$2 ( \4471 , \2107 , \2718 );
not \g45854/U$4 ( \4472 , \2107 );
and \g45854/U$3 ( \4473 , \4472 , \2719 );
nor \g45854/U$1 ( \4474 , \4471 , \4473 );
not \mul_6_18_g43247/U$4 ( \4475 , \4474 );
and \mul_6_18_g43247/U$2 ( \4476 , \4470 , \4475 );
nor \mul_6_18_g43442/U$1 ( \4477 , \4322 , \2732 );
nor \mul_6_18_g43247/U$1 ( \4478 , \4476 , \4477 );
not \mul_6_18_g43246/U$1 ( \4479 , \4478 );
not \mul_6_18_g42691/U$3 ( \4480 , \4479 );
not \mul_6_18_g44083/U$3 ( \4481 , \2463 );
not \mul_6_18_g44083/U$4 ( \4482 , \2296 );
or \mul_6_18_g44083/U$2 ( \4483 , \4481 , \4482 );
nand \mul_6_18_g44314/U$1 ( \4484 , \2307 , \2468 );
nand \mul_6_18_g44083/U$1 ( \4485 , \4483 , \4484 );
not \mul_6_18_g43147/U$3 ( \4486 , \4485 );
not \mul_6_18_g43147/U$4 ( \4487 , \2302 );
or \mul_6_18_g43147/U$2 ( \4488 , \4486 , \4487 );
nand \mul_6_18_g43485/U$1 ( \4489 , \4282 , \2317 );
nand \mul_6_18_g43147/U$1 ( \4490 , \4488 , \4489 );
buf \mul_6_18_g43146/U$1 ( \4491 , \4490 );
not \mul_6_18_g42691/U$4 ( \4492 , \4491 );
or \mul_6_18_g42691/U$2 ( \4493 , \4480 , \4492 );
or \mul_6_18_g42743/U$2 ( \4494 , \4491 , \4479 );
not \mul_6_18_g44112/U$3 ( \4495 , \2179 );
not \mul_6_18_g44112/U$4 ( \4496 , \2762 );
or \mul_6_18_g44112/U$2 ( \4497 , \4495 , \4496 );
nand \mul_6_18_g44360/U$1 ( \4498 , \3330 , \2185 );
nand \mul_6_18_g44112/U$1 ( \4499 , \4497 , \4498 );
not \mul_6_18_g43136/U$3 ( \4500 , \4499 );
not \mul_6_18_g43136/U$4 ( \4501 , \2771 );
or \mul_6_18_g43136/U$2 ( \4502 , \4500 , \4501 );
nand \mul_6_18_g43524/U$1 ( \4503 , \4344 , \2783 );
nand \mul_6_18_g43136/U$1 ( \4504 , \4502 , \4503 );
nand \mul_6_18_g42743/U$1 ( \4505 , \4494 , \4504 );
nand \mul_6_18_g42691/U$1 ( \4506 , \4493 , \4505 );
xor \mul_6_18_g42416/U$4 ( \4507 , \4469 , \4506 );
and \g45522/U$2 ( \4508 , \2094 , \2367 );
not \g45522/U$4 ( \4509 , \2094 );
and \g45522/U$3 ( \4510 , \4509 , \2363 );
or \g45522/U$1 ( \4511 , \4508 , \4510 );
not \mul_6_18_g43208/U$3 ( \4512 , \4511 );
not \mul_6_18_g43208/U$4 ( \4513 , \2399 );
or \mul_6_18_g43208/U$2 ( \4514 , \4512 , \4513 );
nand \mul_6_18_g43484/U$1 ( \4515 , \4384 , \2403 );
nand \mul_6_18_g43208/U$1 ( \4516 , \4514 , \4515 );
not \mul_6_18_g44045/U$3 ( \4517 , \2812 );
not \mul_6_18_g44045/U$4 ( \4518 , \2645 );
or \mul_6_18_g44045/U$2 ( \4519 , \4517 , \4518 );
nand \mul_6_18_g44300/U$1 ( \4520 , \3380 , \2811 );
nand \mul_6_18_g44045/U$1 ( \4521 , \4519 , \4520 );
not \mul_6_18_g43175/U$3 ( \4522 , \4521 );
not \mul_6_18_g43175/U$4 ( \4523 , \2349 );
or \mul_6_18_g43175/U$2 ( \4524 , \4522 , \4523 );
nand \mul_6_18_g43424/U$1 ( \4525 , \2358 , \4374 );
nand \mul_6_18_g43175/U$1 ( \4526 , \4524 , \4525 );
xor \mul_6_18_g42719/U$4 ( \4527 , \4516 , \4526 );
and \mul_6_18_g44036/U$2 ( \4528 , \2116 , \2993 );
not \mul_6_18_g44036/U$4 ( \4529 , \2116 );
and \mul_6_18_g44036/U$3 ( \4530 , \4529 , \2697 );
nor \mul_6_18_g44036/U$1 ( \4531 , \4528 , \4530 );
not \mul_6_18_g43091/U$3 ( \4532 , \4531 );
not \mul_6_18_g43091/U$4 ( \4533 , \2691 );
or \mul_6_18_g43091/U$2 ( \4534 , \4532 , \4533 );
nand \mul_6_18_g43528/U$1 ( \4535 , \4333 , \2701 );
nand \mul_6_18_g43091/U$1 ( \4536 , \4534 , \4535 );
and \mul_6_18_g42719/U$3 ( \4537 , \4527 , \4536 );
and \mul_6_18_g42719/U$5 ( \4538 , \4516 , \4526 );
or \mul_6_18_g42719/U$2 ( \4539 , \4537 , \4538 );
and \mul_6_18_g42416/U$3 ( \4540 , \4507 , \4539 );
and \mul_6_18_g42416/U$5 ( \4541 , \4469 , \4506 );
or \mul_6_18_g42416/U$2 ( \4542 , \4540 , \4541 );
and \mul_6_18_g42320/U$2 ( \4543 , \4450 , \4542 );
not \mul_6_18_g45194/U$2 ( \4544 , \4438 );
nor \mul_6_18_g45194/U$1 ( \4545 , \4544 , \4449 );
nor \mul_6_18_g42320/U$1 ( \4546 , \4543 , \4545 );
buf \mul_6_18_g42299/U$1 ( \4547 , \4546 );
not \mul_6_18_g42094/U$3 ( \4548 , \4547 );
and \g45508/U$2 ( \4549 , \2114 , \3211 );
not \g45508/U$4 ( \4550 , \2114 );
and \g45508/U$3 ( \4551 , \4550 , \2225 );
or \g45508/U$1 ( \4552 , \4549 , \4551 );
not \mul_6_18_g43352/U$3 ( \4553 , \4552 );
not \mul_6_18_g43352/U$4 ( \4554 , \4076 );
or \mul_6_18_g43352/U$2 ( \4555 , \4553 , \4554 );
nand \mul_6_18_g43550/U$1 ( \4556 , \4306 , \3430 );
nand \mul_6_18_g43352/U$1 ( \4557 , \4555 , \4556 );
and \g45515/U$2 ( \4558 , \1970 , \2607 );
not \g45515/U$4 ( \4559 , \1970 );
and \g45515/U$3 ( \4560 , \4559 , \2626 );
or \g45515/U$1 ( \4561 , \4558 , \4560 );
not \mul_6_18_g42962/U$3 ( \4562 , \4561 );
not \mul_6_18_g42962/U$4 ( \4563 , \4256 );
or \mul_6_18_g42962/U$2 ( \4564 , \4562 , \4563 );
nand \mul_6_18_g43004/U$1 ( \4565 , \2842 , \4253 );
nand \mul_6_18_g42962/U$1 ( \4566 , \4564 , \4565 );
xor \mul_6_18_g42569/U$4 ( \4567 , \4557 , \4566 );
not \mul_6_18_g43938/U$3 ( \4568 , \2640 );
not \mul_6_18_g43938/U$4 ( \4569 , \2251 );
or \mul_6_18_g43938/U$2 ( \4570 , \4568 , \4569 );
nand \mul_6_18_g44238/U$1 ( \4571 , \2256 , \2639 );
nand \mul_6_18_g43938/U$1 ( \4572 , \4570 , \4571 );
not \mul_6_18_g43276/U$3 ( \4573 , \4572 );
not \mul_6_18_g43276/U$4 ( \4574 , \2273 );
or \mul_6_18_g43276/U$2 ( \4575 , \4573 , \4574 );
nand \mul_6_18_g43431/U$1 ( \4576 , \3449 , \4294 );
nand \mul_6_18_g43276/U$1 ( \4577 , \4575 , \4576 );
and \mul_6_18_g42569/U$3 ( \4578 , \4567 , \4577 );
and \mul_6_18_g42569/U$5 ( \4579 , \4557 , \4566 );
or \mul_6_18_g42569/U$2 ( \4580 , \4578 , \4579 );
not \mul_6_18_g42568/U$1 ( \4581 , \4580 );
not \mul_6_18_g42567/U$1 ( \4582 , \4581 );
not \mul_6_18_g42348/U$3 ( \4583 , \4582 );
xor \mul_6_18_g42635/U$1 ( \4584 , \4260 , \4272 );
xor \mul_6_18_g42635/U$1_r1 ( \4585 , \4584 , \4274 );
not \mul_6_18_g42348/U$4 ( \4586 , \4585 );
or \mul_6_18_g42348/U$2 ( \4587 , \4583 , \4586 );
xor \mul_6_18_g42637/U$1 ( \4588 , \4329 , \4338 );
xor \mul_6_18_g42637/U$1_r1 ( \4589 , \4588 , \4349 );
not \mul_6_18_g45191/U$2 ( \4590 , \4585 );
nand \mul_6_18_g45191/U$1 ( \4591 , \4590 , \4581 );
nand \mul_6_18_g42391/U$1 ( \4592 , \4589 , \4591 );
nand \mul_6_18_g42348/U$1 ( \4593 , \4587 , \4592 );
not \mul_6_18_g42169/U$3 ( \4594 , \4593 );
xor \mul_6_18_g42411/U$1 ( \4595 , \4277 , \4317 );
xor \mul_6_18_g42411/U$1_r1 ( \4596 , \4595 , \4352 );
not \mul_6_18_g42169/U$4 ( \4597 , \4596 );
or \mul_6_18_g42169/U$2 ( \4598 , \4594 , \4597 );
or \mul_6_18_g42187/U$2 ( \4599 , \4596 , \4593 );
xor \mul_6_18_g42643/U$1 ( \4600 , \4379 , \4389 );
xor \mul_6_18_g42643/U$1_r1 ( \4601 , \4600 , \4400 );
buf \mul_6_18_g42641/U$1 ( \4602 , \4601 );
xor \mul_6_18_g42734/U$1 ( \4603 , \4311 , \4299 );
xnor \mul_6_18_g42734/U$1_r1 ( \4604 , \4603 , \4289 );
not \mul_6_18_g42636/U$1 ( \4605 , \4604 );
or \mul_6_18_g42392/U$2 ( \4606 , \4602 , \4605 );
not \mul_6_18_g43108/U$3 ( \4607 , \2509 );
and \mul_6_18_g44140/U$2 ( \4608 , \2145 , \3257 );
not \mul_6_18_g44140/U$4 ( \4609 , \2145 );
and \mul_6_18_g44140/U$3 ( \4610 , \4609 , \2816 );
nor \mul_6_18_g44140/U$1 ( \4611 , \4608 , \4610 );
not \mul_6_18_g43108/U$4 ( \4612 , \4611 );
and \mul_6_18_g43108/U$2 ( \4613 , \4607 , \4612 );
nor \mul_6_18_g43438/U$1 ( \4614 , \2504 , \4394 );
nor \mul_6_18_g43108/U$1 ( \4615 , \4613 , \4614 );
not \mul_6_18_g43107/U$1 ( \4616 , \4615 );
not \mul_6_18_g42464/U$3 ( \4617 , \4616 );
xor \mul_6_18_g42776/U$1 ( \4618 , \4459 , \4468 );
not \mul_6_18_g42464/U$4 ( \4619 , \4618 );
or \mul_6_18_g42464/U$2 ( \4620 , \4617 , \4619 );
or \mul_6_18_g42512/U$2 ( \4621 , \4616 , \4618 );
nand \mul_6_18_g43649/U$1 ( \4622 , \2682 , \2058 );
not \mul_6_18_g43648/U$1 ( \4623 , \4622 );
not \mul_6_18_g42598/U$3 ( \4624 , \4623 );
and \g45758/U$2 ( \4625 , \2101 , \2423 );
not \g45758/U$4 ( \4626 , \2101 );
and \g45758/U$3 ( \4627 , \4626 , \2418 );
or \g45758/U$1 ( \4628 , \4625 , \4627 );
not \mul_6_18_g42918/U$3 ( \4629 , \4628 );
not \mul_6_18_g42918/U$4 ( \4630 , \4264 );
or \mul_6_18_g42918/U$2 ( \4631 , \4629 , \4630 );
nand \mul_6_18_g43005/U$1 ( \4632 , \2434 , \4463 );
nand \mul_6_18_g42918/U$1 ( \4633 , \4631 , \4632 );
not \mul_6_18_g42598/U$4 ( \4634 , \4633 );
or \mul_6_18_g42598/U$2 ( \4635 , \4624 , \4634 );
or \mul_6_18_g42677/U$2 ( \4636 , \4633 , \4623 );
and \g45760/U$2 ( \4637 , \2113 , \2834 );
not \g45760/U$4 ( \4638 , \2113 );
and \g45760/U$3 ( \4639 , \4638 , \2626 );
or \g45760/U$1 ( \4640 , \4637 , \4639 );
not \mul_6_18_g42964/U$3 ( \4641 , \4640 );
not \mul_6_18_g42964/U$4 ( \4642 , \4256 );
or \mul_6_18_g42964/U$2 ( \4643 , \4641 , \4642 );
nand \mul_6_18_g43006/U$1 ( \4644 , \2842 , \4561 );
nand \mul_6_18_g42964/U$1 ( \4645 , \4643 , \4644 );
nand \mul_6_18_g42677/U$1 ( \4646 , \4636 , \4645 );
nand \mul_6_18_g42598/U$1 ( \4647 , \4635 , \4646 );
nand \mul_6_18_g42512/U$1 ( \4648 , \4621 , \4647 );
nand \mul_6_18_g42464/U$1 ( \4649 , \4620 , \4648 );
buf \mul_6_18_g42452/U$1 ( \4650 , \4649 );
nand \mul_6_18_g42392/U$1 ( \4651 , \4606 , \4650 );
nand \mul_6_18_g42528/U$1 ( \4652 , \4602 , \4605 );
nand \mul_6_18_g42354/U$1 ( \4653 , \4651 , \4652 );
nand \mul_6_18_g42187/U$1 ( \4654 , \4599 , \4653 );
nand \mul_6_18_g42169/U$1 ( \4655 , \4598 , \4654 );
not \mul_6_18_g42161/U$1 ( \4656 , \4655 );
not \mul_6_18_g42094/U$4 ( \4657 , \4656 );
or \mul_6_18_g42094/U$2 ( \4658 , \4548 , \4657 );
xor \mul_6_18_g42233/U$1 ( \4659 , \4238 , \4248 );
xor \mul_6_18_g42233/U$1_r1 ( \4660 , \4659 , \4355 );
nand \mul_6_18_g42094/U$1 ( \4661 , \4658 , \4660 );
not \mul_6_18_g45165/U$2 ( \4662 , \4547 );
nand \mul_6_18_g45165/U$1 ( \4663 , \4662 , \4655 );
nand \mul_6_18_g42079/U$1 ( \4664 , \4661 , \4663 );
xor \mul_6_18_g41931/U$4 ( \4665 , \4436 , \4664 );
xor \mul_6_18_g42050/U$1 ( \4666 , \4358 , \4360 );
xor \mul_6_18_g42050/U$1_r1 ( \4667 , \4666 , \4415 );
and \mul_6_18_g41931/U$3 ( \4668 , \4665 , \4667 );
and \mul_6_18_g41931/U$5 ( \4669 , \4436 , \4664 );
or \mul_6_18_g41931/U$2 ( \4670 , \4668 , \4669 );
nor \mul_6_18_g41898/U$1 ( \4671 , \4434 , \4670 );
xor \mul_6_18_g42177/U$1 ( \4672 , \4363 , \4409 );
xor \mul_6_18_g42177/U$1_r1 ( \4673 , \4672 , \4412 );
xor \mul_6_18_g45812/U$1 ( \4674 , \4403 , \4406 );
xor \mul_6_18_g45812/U$1_r1 ( \4675 , \4674 , \4369 );
xor \mul_6_18_g42341/U$1 ( \4676 , \4438 , \4449 );
xnor \mul_6_18_g42341/U$1_r1 ( \4677 , \4676 , \4542 );
xor \mul_6_18_g42069/U$4 ( \4678 , \4675 , \4677 );
and \g45509/U$2 ( \4679 , \2110 , \3422 );
not \g45509/U$4 ( \4680 , \2110 );
and \g45509/U$3 ( \4681 , \4680 , \2225 );
or \g45509/U$1 ( \4682 , \4679 , \4681 );
not \mul_6_18_g43356/U$3 ( \4683 , \4682 );
not \mul_6_18_g43356/U$4 ( \4684 , \2222 );
or \mul_6_18_g43356/U$2 ( \4685 , \4683 , \4684 );
nand \mul_6_18_g43447/U$1 ( \4686 , \4552 , \3430 );
nand \mul_6_18_g43356/U$1 ( \4687 , \4685 , \4686 );
not \mul_6_18_g44024/U$3 ( \4688 , \2112 );
not \mul_6_18_g44024/U$4 ( \4689 , \2364 );
or \mul_6_18_g44024/U$2 ( \4690 , \4688 , \4689 );
not \mul_6_18_g44567/U$1 ( \4691 , \2367 );
nand \mul_6_18_g44296/U$1 ( \4692 , \4691 , \2824 );
nand \mul_6_18_g44024/U$1 ( \4693 , \4690 , \4692 );
not \mul_6_18_g43211/U$3 ( \4694 , \4693 );
not \mul_6_18_g43211/U$4 ( \4695 , \2399 );
or \mul_6_18_g43211/U$2 ( \4696 , \4694 , \4695 );
nand \mul_6_18_g43448/U$1 ( \4697 , \2403 , \4511 );
nand \mul_6_18_g43211/U$1 ( \4698 , \4696 , \4697 );
xor \mul_6_18_g42711/U$4 ( \4699 , \4687 , \4698 );
not \g45751/U$3 ( \4700 , \2729 );
not \mul_6_18_g43993/U$3 ( \4701 , \2111 );
not \mul_6_18_g43993/U$4 ( \4702 , \2715 );
or \mul_6_18_g43993/U$2 ( \4703 , \4701 , \4702 );
nand \mul_6_18_g44272/U$1 ( \4704 , \2972 , \2779 );
nand \mul_6_18_g43993/U$1 ( \4705 , \4703 , \4704 );
not \g45751/U$4 ( \4706 , \4705 );
or \g45751/U$2 ( \4707 , \4700 , \4706 );
not \mul_6_18_g45235/U$2 ( \4708 , \4474 );
nand \mul_6_18_g45235/U$1 ( \4709 , \4708 , \3326 );
nand \g45751/U$1 ( \4710 , \4707 , \4709 );
and \mul_6_18_g42711/U$3 ( \4711 , \4699 , \4710 );
and \mul_6_18_g42711/U$5 ( \4712 , \4687 , \4698 );
or \mul_6_18_g42711/U$2 ( \4713 , \4711 , \4712 );
not \mul_6_18_g44102/U$3 ( \4714 , \2006 );
not \mul_6_18_g44102/U$4 ( \4715 , \3237 );
or \mul_6_18_g44102/U$2 ( \4716 , \4714 , \4715 );
nand \mul_6_18_g44353/U$1 ( \4717 , \2307 , \2795 );
nand \mul_6_18_g44102/U$1 ( \4718 , \4716 , \4717 );
not \mul_6_18_g43149/U$3 ( \4719 , \4718 );
not \mul_6_18_g43149/U$4 ( \4720 , \2302 );
or \mul_6_18_g43149/U$2 ( \4721 , \4719 , \4720 );
nand \mul_6_18_g43492/U$1 ( \4722 , \4485 , \2317 );
nand \mul_6_18_g43149/U$1 ( \4723 , \4721 , \4722 );
not \mul_6_18_g43961/U$3 ( \4724 , \2092 );
not \mul_6_18_g43961/U$4 ( \4725 , \2277 );
or \mul_6_18_g43961/U$2 ( \4726 , \4724 , \4725 );
nand \mul_6_18_g44257/U$1 ( \4727 , \2256 , \2754 );
nand \mul_6_18_g43961/U$1 ( \4728 , \4726 , \4727 );
not \mul_6_18_g43300/U$3 ( \4729 , \4728 );
not \mul_6_18_g43300/U$4 ( \4730 , \2273 );
or \mul_6_18_g43300/U$2 ( \4731 , \4729 , \4730 );
nand \mul_6_18_g43501/U$1 ( \4732 , \4572 , \3449 );
nand \mul_6_18_g43300/U$1 ( \4733 , \4731 , \4732 );
or \mul_6_18_g42854/U$2 ( \4734 , \4723 , \4733 );
and \mul_6_18_g44126/U$2 ( \4735 , \3154 , \2762 );
not \mul_6_18_g44126/U$4 ( \4736 , \3154 );
and \mul_6_18_g44126/U$3 ( \4737 , \4736 , \3330 );
nor \mul_6_18_g44126/U$1 ( \4738 , \4735 , \4737 );
not \mul_6_18_g43130/U$3 ( \4739 , \4738 );
not \mul_6_18_g43130/U$4 ( \4740 , \2771 );
or \mul_6_18_g43130/U$2 ( \4741 , \4739 , \4740 );
nand \mul_6_18_g43426/U$1 ( \4742 , \4499 , \2783 );
nand \mul_6_18_g43130/U$1 ( \4743 , \4741 , \4742 );
nand \mul_6_18_g42854/U$1 ( \4744 , \4734 , \4743 );
nand \mul_6_18_g42881/U$1 ( \4745 , \4723 , \4733 );
nand \mul_6_18_g42804/U$1 ( \4746 , \4744 , \4745 );
xor \mul_6_18_g42418/U$4 ( \4747 , \4713 , \4746 );
xor \mul_6_18_g42719/U$1 ( \4748 , \4516 , \4526 );
xor \mul_6_18_g42719/U$1_r1 ( \4749 , \4748 , \4536 );
and \mul_6_18_g42418/U$3 ( \4750 , \4747 , \4749 );
and \mul_6_18_g42418/U$5 ( \4751 , \4713 , \4746 );
or \mul_6_18_g42418/U$2 ( \4752 , \4750 , \4751 );
xor \mul_6_18_g42416/U$1 ( \4753 , \4469 , \4506 );
xor \mul_6_18_g42416/U$1_r1 ( \4754 , \4753 , \4539 );
or \mul_6_18_g42220/U$2 ( \4755 , \4752 , \4754 );
xor \mul_6_18_g42569/U$1 ( \4756 , \4557 , \4566 );
xor \mul_6_18_g42569/U$1_r1 ( \4757 , \4756 , \4577 );
and \mul_6_18_g42863/U$2 ( \4758 , \4490 , \4479 );
not \mul_6_18_g42863/U$4 ( \4759 , \4490 );
and \mul_6_18_g42863/U$3 ( \4760 , \4759 , \4478 );
nor \mul_6_18_g42863/U$1 ( \4761 , \4758 , \4760 );
and \mul_6_18_g42738/U$2 ( \4762 , \4761 , \4504 );
not \mul_6_18_g42738/U$4 ( \4763 , \4761 );
not \mul_6_18_g43135/U$1 ( \4764 , \4504 );
and \mul_6_18_g42738/U$3 ( \4765 , \4763 , \4764 );
nor \mul_6_18_g42738/U$1 ( \4766 , \4762 , \4765 );
xor \mul_6_18_g42261/U$4 ( \4767 , \4757 , \4766 );
and \mul_6_18_g44150/U$2 ( \4768 , \2056 , \2496 );
not \mul_6_18_g44150/U$4 ( \4769 , \2056 );
and \mul_6_18_g44150/U$3 ( \4770 , \4769 , \3883 );
nor \mul_6_18_g44150/U$1 ( \4771 , \4768 , \4770 );
not \mul_6_18_g43110/U$3 ( \4772 , \4771 );
not \mul_6_18_g43110/U$4 ( \4773 , \2511 );
or \mul_6_18_g43110/U$2 ( \4774 , \4772 , \4773 );
not \mul_6_18_g45241/U$2 ( \4775 , \4611 );
nand \mul_6_18_g45241/U$1 ( \4776 , \4775 , \2515 );
nand \mul_6_18_g43110/U$1 ( \4777 , \4774 , \4776 );
not \mul_6_18_g44067/U$3 ( \4778 , \1998 );
not \mul_6_18_g44067/U$4 ( \4779 , \2644 );
or \mul_6_18_g44067/U$2 ( \4780 , \4778 , \4779 );
nand \mul_6_18_g44339/U$1 ( \4781 , \2335 , \2489 );
nand \mul_6_18_g44067/U$1 ( \4782 , \4780 , \4781 );
not \mul_6_18_g43182/U$3 ( \4783 , \4782 );
not \mul_6_18_g43182/U$4 ( \4784 , \2349 );
or \mul_6_18_g43182/U$2 ( \4785 , \4783 , \4784 );
nand \mul_6_18_g43628/U$1 ( \4786 , \2359 , \4521 );
nand \mul_6_18_g43182/U$1 ( \4787 , \4785 , \4786 );
nor \mul_6_18_g42883/U$1 ( \4788 , \4777 , \4787 );
and \g45759/U$2 ( \4789 , \1970 , \2423 );
not \g45759/U$4 ( \4790 , \1970 );
and \g45759/U$3 ( \4791 , \4790 , \2418 );
or \g45759/U$1 ( \4792 , \4789 , \4791 );
not \mul_6_18_g42923/U$3 ( \4793 , \4792 );
not \mul_6_18_g42923/U$4 ( \4794 , \4014 );
or \mul_6_18_g42923/U$2 ( \4795 , \4793 , \4794 );
nand \mul_6_18_g45644/U$1 ( \4796 , \2434 , \4628 );
nand \mul_6_18_g42923/U$1 ( \4797 , \4795 , \4796 );
nand \mul_6_18_g44169/U$1 ( \4798 , \2505 , \2116 );
and \mul_6_18_g43680/U$2 ( \4799 , \4798 , \2761 );
not \mul_6_18_g43728/U$3 ( \4800 , \2058 );
not \mul_6_18_g44403/U$1 ( \4801 , \2505 );
not \mul_6_18_g43728/U$4 ( \4802 , \4801 );
or \mul_6_18_g43728/U$2 ( \4803 , \4800 , \4802 );
nand \mul_6_18_g43728/U$1 ( \4804 , \4803 , \2817 );
nor \mul_6_18_g43680/U$1 ( \4805 , \4799 , \4804 );
nand \mul_6_18_g42839/U$1 ( \4806 , \4797 , \4805 );
or \mul_6_18_g42600/U$2 ( \4807 , \4788 , \4806 );
nand \mul_6_18_g42882/U$1 ( \4808 , \4777 , \4787 );
nand \mul_6_18_g42600/U$1 ( \4809 , \4807 , \4808 );
and \mul_6_18_g42261/U$3 ( \4810 , \4767 , \4809 );
and \mul_6_18_g42261/U$5 ( \4811 , \4757 , \4766 );
or \mul_6_18_g42261/U$2 ( \4812 , \4810 , \4811 );
nand \mul_6_18_g42220/U$1 ( \4813 , \4755 , \4812 );
nand \mul_6_18_g42343/U$1 ( \4814 , \4752 , \4754 );
nand \mul_6_18_g42192/U$1 ( \4815 , \4813 , \4814 );
and \mul_6_18_g42069/U$3 ( \4816 , \4678 , \4815 );
and \mul_6_18_g42069/U$5 ( \4817 , \4675 , \4677 );
or \mul_6_18_g42069/U$2 ( \4818 , \4816 , \4817 );
xor \mul_6_18_g41950/U$1 ( \4819 , \4673 , \4818 );
xor \mul_6_18_g42110/U$1 ( \4820 , \4546 , \4660 );
xnor \mul_6_18_g42110/U$1_r1 ( \4821 , \4820 , \4655 );
xor \mul_6_18_g41950/U$1_r1 ( \4822 , \4819 , \4821 );
xor \g45377/U$1 ( \4823 , \4596 , \4593 );
and \mul_6_18_g42180/U$2 ( \4824 , \4823 , \4653 );
not \mul_6_18_g42180/U$4 ( \4825 , \4823 );
not \mul_6_18_g42257/U$1 ( \4826 , \4653 );
and \mul_6_18_g42180/U$3 ( \4827 , \4825 , \4826 );
nor \mul_6_18_g42180/U$1 ( \4828 , \4824 , \4827 );
xor \mul_6_18_g45542/U$1 ( \4829 , \4604 , \4649 );
xor \mul_6_18_g45542/U$1_r1 ( \4830 , \4829 , \4601 );
not \mul_6_18_g42256/U$1 ( \4831 , \4830 );
not \mul_6_18_g45162/U$2 ( \4832 , \4831 );
xor \mul_6_18_g42384/U$1 ( \4833 , \4580 , \4585 );
xnor \mul_6_18_g42384/U$1_r1 ( \4834 , \4833 , \4589 );
nand \mul_6_18_g45162/U$1 ( \4835 , \4832 , \4834 );
not \mul_6_18_g42128/U$3 ( \4836 , \4835 );
not \mul_6_18_g42490/U$3 ( \4837 , \4647 );
not \mul_6_18_g42621/U$3 ( \4838 , \4618 );
not \mul_6_18_g42621/U$4 ( \4839 , \4615 );
and \mul_6_18_g42621/U$2 ( \4840 , \4838 , \4839 );
and \mul_6_18_g42621/U$5 ( \4841 , \4618 , \4615 );
nor \mul_6_18_g42621/U$1 ( \4842 , \4840 , \4841 );
not \mul_6_18_g42490/U$4 ( \4843 , \4842 );
or \mul_6_18_g42490/U$2 ( \4844 , \4837 , \4843 );
or \mul_6_18_g42490/U$5 ( \4845 , \4842 , \4647 );
nand \mul_6_18_g42490/U$1 ( \4846 , \4844 , \4845 );
not \mul_6_18_g43894/U$3 ( \4847 , \2106 );
not \mul_6_18_g43894/U$4 ( \4848 , \3422 );
or \mul_6_18_g43894/U$2 ( \4849 , \4847 , \4848 );
not \mul_6_18_g45245/U$2 ( \4850 , \2106 );
nand \mul_6_18_g45245/U$1 ( \4851 , \4850 , \2216 );
nand \mul_6_18_g43894/U$1 ( \4852 , \4849 , \4851 );
not \mul_6_18_g43380/U$3 ( \4853 , \4852 );
not \mul_6_18_g43380/U$4 ( \4854 , \2222 );
or \mul_6_18_g43380/U$2 ( \4855 , \4853 , \4854 );
nand \mul_6_18_g43477/U$1 ( \4856 , \4682 , \2934 );
nand \mul_6_18_g43380/U$1 ( \4857 , \4855 , \4856 );
not \mul_6_18_g43992/U$3 ( \4858 , \2094 );
not \mul_6_18_g43992/U$4 ( \4859 , \2715 );
or \mul_6_18_g43992/U$2 ( \4860 , \4858 , \4859 );
not \mul_6_18_g45263/U$2 ( \4861 , \2094 );
nand \mul_6_18_g45263/U$1 ( \4862 , \4861 , \2719 );
nand \mul_6_18_g43992/U$1 ( \4863 , \4860 , \4862 );
not \mul_6_18_g43250/U$3 ( \4864 , \4863 );
not \mul_6_18_g43250/U$4 ( \4865 , \2965 );
or \mul_6_18_g43250/U$2 ( \4866 , \4864 , \4865 );
nand \mul_6_18_g43432/U$1 ( \4867 , \4327 , \4705 );
nand \mul_6_18_g43250/U$1 ( \4868 , \4866 , \4867 );
xor \mul_6_18_g42728/U$4 ( \4869 , \4857 , \4868 );
not \mul_6_18_g44125/U$3 ( \4870 , \2144 );
not \mul_6_18_g44125/U$4 ( \4871 , \3920 );
or \mul_6_18_g44125/U$2 ( \4872 , \4870 , \4871 );
nand \mul_6_18_g44376/U$1 ( \4873 , \3330 , \2145 );
nand \mul_6_18_g44125/U$1 ( \4874 , \4872 , \4873 );
not \mul_6_18_g43131/U$3 ( \4875 , \4874 );
not \mul_6_18_g43131/U$4 ( \4876 , \2771 );
or \mul_6_18_g43131/U$2 ( \4877 , \4875 , \4876 );
nand \mul_6_18_g43478/U$1 ( \4878 , \4738 , \2783 );
nand \mul_6_18_g43131/U$1 ( \4879 , \4877 , \4878 );
and \mul_6_18_g42728/U$3 ( \4880 , \4869 , \4879 );
and \mul_6_18_g42728/U$5 ( \4881 , \4857 , \4868 );
or \mul_6_18_g42728/U$2 ( \4882 , \4880 , \4881 );
xnor \g45761/U$1 ( \4883 , \2107 , \2251 );
not \mul_6_18_g43280/U$3 ( \4884 , \4883 );
not \mul_6_18_g43280/U$4 ( \4885 , \2938 );
or \mul_6_18_g43280/U$2 ( \4886 , \4884 , \4885 );
nand \mul_6_18_g43498/U$1 ( \4887 , \4728 , \3232 );
nand \mul_6_18_g43280/U$1 ( \4888 , \4886 , \4887 );
not \mul_6_18_g43936/U$3 ( \4889 , \2640 );
not \mul_6_18_g43936/U$4 ( \4890 , \2607 );
or \mul_6_18_g43936/U$2 ( \4891 , \4889 , \4890 );
nand \mul_6_18_g44248/U$1 ( \4892 , \2626 , \2639 );
nand \mul_6_18_g43936/U$1 ( \4893 , \4891 , \4892 );
not \mul_6_18_g42969/U$3 ( \4894 , \4893 );
not \mul_6_18_g42969/U$4 ( \4895 , \4256 );
or \mul_6_18_g42969/U$2 ( \4896 , \4894 , \4895 );
nand \mul_6_18_g43013/U$1 ( \4897 , \4005 , \4640 );
nand \mul_6_18_g42969/U$1 ( \4898 , \4896 , \4897 );
or \mul_6_18_g45206/U$2 ( \4899 , \4888 , \4898 );
not \mul_6_18_g44103/U$3 ( \4900 , \2179 );
not \mul_6_18_g44103/U$4 ( \4901 , \2296 );
or \mul_6_18_g44103/U$2 ( \4902 , \4900 , \4901 );
nand \mul_6_18_g44341/U$1 ( \4903 , \2307 , \2185 );
nand \mul_6_18_g44103/U$1 ( \4904 , \4902 , \4903 );
not \mul_6_18_g43151/U$3 ( \4905 , \4904 );
not \mul_6_18_g43151/U$4 ( \4906 , \2303 );
or \mul_6_18_g43151/U$2 ( \4907 , \4905 , \4906 );
nand \mul_6_18_g43558/U$1 ( \4908 , \4287 , \4718 );
nand \mul_6_18_g43151/U$1 ( \4909 , \4907 , \4908 );
nand \mul_6_18_g45206/U$1 ( \4910 , \4899 , \4909 );
nand \mul_6_18_g42827/U$1 ( \4911 , \4898 , \4888 );
nand \mul_6_18_g42757/U$1 ( \4912 , \4910 , \4911 );
nor \mul_6_18_g42530/U$1 ( \4913 , \4882 , \4912 );
not \mul_6_18_g42813/U$3 ( \4914 , \4623 );
not \mul_6_18_g42917/U$1 ( \4915 , \4633 );
not \mul_6_18_g42813/U$4 ( \4916 , \4915 );
or \mul_6_18_g42813/U$2 ( \4917 , \4914 , \4916 );
nand \mul_6_18_g42832/U$1 ( \4918 , \4633 , \4622 );
nand \mul_6_18_g42813/U$1 ( \4919 , \4917 , \4918 );
not \mul_6_18_g42963/U$1 ( \4920 , \4645 );
and \mul_6_18_g42620/U$2 ( \4921 , \4919 , \4920 );
not \mul_6_18_g42620/U$4 ( \4922 , \4919 );
and \mul_6_18_g42620/U$3 ( \4923 , \4922 , \4645 );
nor \mul_6_18_g42620/U$1 ( \4924 , \4921 , \4923 );
buf \mul_6_18_g42572/U$1 ( \4925 , \4924 );
or \mul_6_18_g42468/U$2 ( \4926 , \4913 , \4925 );
nand \mul_6_18_g42529/U$1 ( \4927 , \4882 , \4912 );
nand \mul_6_18_g42468/U$1 ( \4928 , \4926 , \4927 );
xor \mul_6_18_g42206/U$4 ( \4929 , \4846 , \4928 );
xor \mul_6_18_g42418/U$1 ( \4930 , \4713 , \4746 );
xor \mul_6_18_g42418/U$1_r1 ( \4931 , \4930 , \4749 );
and \mul_6_18_g42206/U$3 ( \4932 , \4929 , \4931 );
and \mul_6_18_g42206/U$5 ( \4933 , \4846 , \4928 );
or \mul_6_18_g42206/U$2 ( \4934 , \4932 , \4933 );
not \mul_6_18_g42128/U$4 ( \4935 , \4934 );
or \mul_6_18_g42128/U$2 ( \4936 , \4836 , \4935 );
not \mul_6_18_g45168/U$2 ( \4937 , \4834 );
nand \mul_6_18_g45168/U$1 ( \4938 , \4937 , \4831 );
nand \mul_6_18_g42128/U$1 ( \4939 , \4936 , \4938 );
xor \mul_6_18_g41953/U$4 ( \4940 , \4828 , \4939 );
xor \mul_6_18_g42069/U$1 ( \4941 , \4675 , \4677 );
xor \mul_6_18_g42069/U$1_r1 ( \4942 , \4941 , \4815 );
and \mul_6_18_g41953/U$3 ( \4943 , \4940 , \4942 );
and \mul_6_18_g41953/U$5 ( \4944 , \4828 , \4939 );
or \mul_6_18_g41953/U$2 ( \4945 , \4943 , \4944 );
nand \mul_6_18_g41915/U$1 ( \4946 , \4822 , \4945 );
xor \mul_6_18_g41931/U$1 ( \4947 , \4436 , \4664 );
xor \mul_6_18_g41931/U$1_r1 ( \4948 , \4947 , \4667 );
xor \mul_6_18_g41950/U$4 ( \4949 , \4673 , \4818 );
and \mul_6_18_g41950/U$3 ( \4950 , \4949 , \4821 );
and \mul_6_18_g41950/U$5 ( \4951 , \4673 , \4818 );
or \mul_6_18_g41950/U$2 ( \4952 , \4950 , \4951 );
nand \mul_6_18_g41902/U$1 ( \4953 , \4948 , \4952 );
nand \mul_6_18_g41871/U$1 ( \4954 , \4946 , \4953 );
not \mul_6_18_g41930/U$1 ( \4955 , \4948 );
not \mul_6_18_g41949/U$1 ( \4956 , \4952 );
nand \mul_6_18_g41900/U$1 ( \4957 , \4955 , \4956 );
nand \mul_6_18_g41864/U$1 ( \4958 , \4954 , \4957 );
nor \mul_6_18_g41852/U$1 ( \4959 , \4671 , \4958 );
nand \mul_6_18_g41908/U$1 ( \4960 , \4434 , \4670 );
not \mul_6_18_g41907/U$1 ( \4961 , \4960 );
nor \mul_6_18_g41850/U$1 ( \4962 , \4959 , \4961 );
not \mul_6_18_g41946/U$1 ( \4963 , \4202 );
not \mul_6_18_g41954/U$1 ( \4964 , \4422 );
nand \mul_6_18_g41916/U$1 ( \4965 , \4963 , \4964 );
nand \mul_6_18_g41847/U$1 ( \4966 , \4962 , \4965 );
not \mul_6_18_g41842/U$4 ( \4967 , \4966 );
or \mul_6_18_g41842/U$2 ( \4968 , \4424 , \4967 );
and \g45523/U$2 ( \4969 , \2810 , \2277 );
not \g45523/U$4 ( \4970 , \2810 );
and \g45523/U$3 ( \4971 , \4970 , \2256 );
or \g45523/U$1 ( \4972 , \4969 , \4971 );
not \mul_6_18_g43298/U$3 ( \4973 , \4972 );
not \mul_6_18_g43298/U$4 ( \4974 , \2273 );
or \mul_6_18_g43298/U$2 ( \4975 , \4973 , \4974 );
and \g45524/U$2 ( \4976 , \2112 , \2277 );
not \g45524/U$4 ( \4977 , \2112 );
and \g45524/U$3 ( \4978 , \4977 , \2256 );
or \g45524/U$1 ( \4979 , \4976 , \4978 );
nand \mul_6_18_g43526/U$1 ( \4980 , \4979 , \3449 );
nand \mul_6_18_g43298/U$1 ( \4981 , \4975 , \4980 );
not \mul_6_18_g43297/U$1 ( \4982 , \4981 );
not \mul_6_18_g42873/U$3 ( \4983 , \4982 );
not \mul_6_18_g44076/U$3 ( \4984 , \2179 );
not \mul_6_18_g44076/U$4 ( \4985 , \2367 );
or \mul_6_18_g44076/U$2 ( \4986 , \4984 , \4985 );
nand \mul_6_18_g44347/U$1 ( \4987 , \4691 , \2185 );
nand \mul_6_18_g44076/U$1 ( \4988 , \4986 , \4987 );
not \mul_6_18_g43223/U$3 ( \4989 , \4988 );
not \mul_6_18_g43223/U$4 ( \4990 , \2399 );
or \mul_6_18_g43223/U$2 ( \4991 , \4989 , \4990 );
not \mul_6_18_g44077/U$3 ( \4992 , \2006 );
not \mul_6_18_g44077/U$4 ( \4993 , \2367 );
or \mul_6_18_g44077/U$2 ( \4994 , \4992 , \4993 );
nand \mul_6_18_g44359/U$1 ( \4995 , \2363 , \2795 );
nand \mul_6_18_g44077/U$1 ( \4996 , \4994 , \4995 );
nand \mul_6_18_g43427/U$1 ( \4997 , \2403 , \4996 );
nand \mul_6_18_g43223/U$1 ( \4998 , \4991 , \4997 );
not \mul_6_18_g42873/U$4 ( \4999 , \4998 );
or \mul_6_18_g42873/U$2 ( \5000 , \4983 , \4999 );
or \mul_6_18_g42873/U$5 ( \5001 , \4998 , \4982 );
nand \mul_6_18_g42873/U$1 ( \5002 , \5000 , \5001 );
not \mul_6_18_g43587/U$1 ( \5003 , \2729 );
not \mul_6_18_g43258/U$3 ( \5004 , \5003 );
and \mul_6_18_g44043/U$2 ( \5005 , \2468 , \2714 );
not \mul_6_18_g44043/U$4 ( \5006 , \2468 );
and \mul_6_18_g44043/U$3 ( \5007 , \5006 , \2718 );
nor \mul_6_18_g44043/U$1 ( \5008 , \5005 , \5007 );
not \mul_6_18_g43258/U$4 ( \5009 , \5008 );
and \mul_6_18_g43258/U$2 ( \5010 , \5004 , \5009 );
not \mul_6_18_g44041/U$3 ( \5011 , \1998 );
not \mul_6_18_g44041/U$4 ( \5012 , \2715 );
or \mul_6_18_g44041/U$2 ( \5013 , \5011 , \5012 );
nand \mul_6_18_g44331/U$1 ( \5014 , \2972 , \2489 );
nand \mul_6_18_g44041/U$1 ( \5015 , \5013 , \5014 );
not \mul_6_18_g45238/U$2 ( \5016 , \5015 );
nor \mul_6_18_g45238/U$1 ( \5017 , \5016 , \3473 );
nor \mul_6_18_g43258/U$1 ( \5018 , \5010 , \5017 );
and \mul_6_18_g42793/U$2 ( \5019 , \5002 , \5018 );
not \mul_6_18_g42793/U$4 ( \5020 , \5002 );
not \mul_6_18_g43257/U$1 ( \5021 , \5018 );
and \mul_6_18_g42793/U$3 ( \5022 , \5020 , \5021 );
nor \mul_6_18_g42793/U$1 ( \5023 , \5019 , \5022 );
and \g45518/U$2 ( \5024 , \1838 , \3214 );
not \g45518/U$4 ( \5025 , \1838 );
and \g45518/U$3 ( \5026 , \5025 , \2225 );
or \g45518/U$1 ( \5027 , \5024 , \5026 );
not \mul_6_18_g43366/U$3 ( \5028 , \5027 );
not \mul_6_18_g43366/U$4 ( \5029 , \2222 );
or \mul_6_18_g43366/U$2 ( \5030 , \5028 , \5029 );
not \mul_6_18_g43927/U$3 ( \5031 , \2113 );
not \mul_6_18_g43927/U$4 ( \5032 , \3214 );
or \mul_6_18_g43927/U$2 ( \5033 , \5031 , \5032 );
nand \mul_6_18_g44243/U$1 ( \5034 , \2225 , \3899 );
nand \mul_6_18_g43927/U$1 ( \5035 , \5033 , \5034 );
nand \mul_6_18_g43436/U$1 ( \5036 , \5035 , \2934 );
nand \mul_6_18_g43366/U$1 ( \5037 , \5030 , \5036 );
not \g45750/U$3 ( \5038 , \4005 );
not \mul_6_18_g43977/U$3 ( \5039 , \2111 );
not \mul_6_18_g43977/U$4 ( \5040 , \2607 );
or \mul_6_18_g43977/U$2 ( \5041 , \5039 , \5040 );
nand \mul_6_18_g44281/U$1 ( \5042 , \2626 , \2779 );
nand \mul_6_18_g43977/U$1 ( \5043 , \5041 , \5042 );
not \g45750/U$4 ( \5044 , \5043 );
or \g45750/U$2 ( \5045 , \5038 , \5044 );
not \fopt45578/U$1 ( \5046 , \4002 );
and \mul_6_18_g43979/U$2 ( \5047 , \2500 , \2606 );
not \mul_6_18_g43979/U$4 ( \5048 , \2500 );
and \mul_6_18_g43979/U$3 ( \5049 , \5048 , \2834 );
nor \mul_6_18_g43979/U$1 ( \5050 , \5047 , \5049 );
or \g45750/U$5 ( \5051 , \5046 , \5050 );
nand \g45750/U$1 ( \5052 , \5045 , \5051 );
xor \mul_6_18_g42550/U$1 ( \5053 , \5037 , \5052 );
and \mul_6_18_g44108/U$2 ( \5054 , \2058 , \2311 );
not \mul_6_18_g44108/U$4 ( \5055 , \2058 );
and \mul_6_18_g44108/U$3 ( \5056 , \5055 , \2308 );
nor \mul_6_18_g44108/U$1 ( \5057 , \5054 , \5056 );
not \mul_6_18_g43162/U$3 ( \5058 , \5057 );
not \mul_6_18_g43162/U$4 ( \5059 , \2303 );
or \mul_6_18_g43162/U$2 ( \5060 , \5058 , \5059 );
not \mul_6_18_g44124/U$3 ( \5061 , \2056 );
not \mul_6_18_g44124/U$4 ( \5062 , \3237 );
or \mul_6_18_g44124/U$2 ( \5063 , \5061 , \5062 );
nand \mul_6_18_g44387/U$1 ( \5064 , \2307 , \3360 );
nand \mul_6_18_g44124/U$1 ( \5065 , \5063 , \5064 );
nand \mul_6_18_g43639/U$1 ( \5066 , \2318 , \5065 );
nand \mul_6_18_g43162/U$1 ( \5067 , \5060 , \5066 );
xor \mul_6_18_g42550/U$1_r1 ( \5068 , \5053 , \5067 );
not \mul_6_18_g43949/U$3 ( \5069 , \2092 );
not \mul_6_18_g43949/U$4 ( \5070 , \3422 );
or \mul_6_18_g43949/U$2 ( \5071 , \5069 , \5070 );
nand \mul_6_18_g44258/U$1 ( \5072 , \2225 , \2754 );
nand \mul_6_18_g43949/U$1 ( \5073 , \5071 , \5072 );
not \mul_6_18_g43373/U$3 ( \5074 , \5073 );
not \mul_6_18_g43373/U$4 ( \5075 , \4076 );
or \mul_6_18_g43373/U$2 ( \5076 , \5074 , \5075 );
not \mul_6_18_g45278/U$2 ( \5077 , \2243 );
nand \mul_6_18_g45278/U$1 ( \5078 , \5077 , \5027 );
nand \mul_6_18_g43373/U$1 ( \5079 , \5076 , \5078 );
not \mul_6_18_g44028/U$3 ( \5080 , \1998 );
not \mul_6_18_g44028/U$4 ( \5081 , \2251 );
or \mul_6_18_g44028/U$2 ( \5082 , \5080 , \5081 );
nand \mul_6_18_g44336/U$1 ( \5083 , \2256 , \2489 );
nand \mul_6_18_g44028/U$1 ( \5084 , \5082 , \5083 );
not \mul_6_18_g43303/U$3 ( \5085 , \5084 );
not \mul_6_18_g43303/U$4 ( \5086 , \2273 );
or \mul_6_18_g43303/U$2 ( \5087 , \5085 , \5086 );
nand \mul_6_18_g43611/U$1 ( \5088 , \3449 , \4972 );
nand \mul_6_18_g43303/U$1 ( \5089 , \5087 , \5088 );
xor \mul_6_18_g42631/U$4 ( \5090 , \5079 , \5089 );
not \mul_6_18_g44064/U$3 ( \5091 , \2006 );
not \mul_6_18_g44064/U$4 ( \5092 , \2715 );
or \mul_6_18_g44064/U$2 ( \5093 , \5091 , \5092 );
nand \mul_6_18_g44357/U$1 ( \5094 , \2972 , \2795 );
nand \mul_6_18_g44064/U$1 ( \5095 , \5093 , \5094 );
not \mul_6_18_g43262/U$3 ( \5096 , \5095 );
not \mul_6_18_g43262/U$4 ( \5097 , \3323 );
or \mul_6_18_g43262/U$2 ( \5098 , \5096 , \5097 );
not \mul_6_18_g45239/U$2 ( \5099 , \5008 );
nand \mul_6_18_g45239/U$1 ( \5100 , \5099 , \4327 );
nand \mul_6_18_g43262/U$1 ( \5101 , \5098 , \5100 );
and \mul_6_18_g42631/U$3 ( \5102 , \5090 , \5101 );
and \mul_6_18_g42631/U$5 ( \5103 , \5079 , \5089 );
or \mul_6_18_g42631/U$2 ( \5104 , \5102 , \5103 );
and \mul_6_18_g42485/U$2 ( \5105 , \5068 , \5104 );
not \mul_6_18_g42485/U$4 ( \5106 , \5068 );
not \mul_6_18_g42630/U$1 ( \5107 , \5104 );
and \mul_6_18_g42485/U$3 ( \5108 , \5106 , \5107 );
nor \mul_6_18_g42485/U$1 ( \5109 , \5105 , \5108 );
not \g45549/U$2 ( \5110 , \5109 );
xor \g45549/U$1 ( \5111 , \5023 , \5110 );
xor \mul_6_18_g42631/U$1 ( \5112 , \5079 , \5089 );
xor \mul_6_18_g42631/U$1_r1 ( \5113 , \5112 , \5101 );
not \mul_6_18_g44117/U$3 ( \5114 , \2056 );
not \mul_6_18_g44117/U$4 ( \5115 , \2645 );
or \mul_6_18_g44117/U$2 ( \5116 , \5114 , \5115 );
nand \mul_6_18_g44380/U$1 ( \5117 , \2335 , \3360 );
nand \mul_6_18_g44117/U$1 ( \5118 , \5116 , \5117 );
not \mul_6_18_g43177/U$3 ( \5119 , \5118 );
not \mul_6_18_g43177/U$4 ( \5120 , \2349 );
or \mul_6_18_g43177/U$2 ( \5121 , \5119 , \5120 );
not \mul_6_18_g44106/U$3 ( \5122 , \2144 );
not \mul_6_18_g44106/U$4 ( \5123 , \2336 );
or \mul_6_18_g44106/U$2 ( \5124 , \5122 , \5123 );
nand \mul_6_18_g44373/U$1 ( \5125 , \3380 , \2145 );
nand \mul_6_18_g44106/U$1 ( \5126 , \5124 , \5125 );
nand \mul_6_18_g43522/U$1 ( \5127 , \2359 , \5126 );
nand \mul_6_18_g43177/U$1 ( \5128 , \5121 , \5127 );
not \mul_6_18_g43176/U$1 ( \5129 , \5128 );
not \mul_6_18_g42610/U$3 ( \5130 , \5129 );
not \mul_6_18_g43972/U$3 ( \5131 , \2094 );
not \mul_6_18_g43972/U$4 ( \5132 , \2419 );
or \mul_6_18_g43972/U$2 ( \5133 , \5131 , \5132 );
nand \mul_6_18_g44292/U$1 ( \5134 , \2848 , \2500 );
nand \mul_6_18_g43972/U$1 ( \5135 , \5133 , \5134 );
not \mul_6_18_g42930/U$3 ( \5136 , \5135 );
not \mul_6_18_g42930/U$4 ( \5137 , \4014 );
or \mul_6_18_g42930/U$2 ( \5138 , \5136 , \5137 );
not \mul_6_18_g43971/U$3 ( \5139 , \2111 );
not \mul_6_18_g44993/U$1 ( \5140 , \2614 );
not \mul_6_18_g44992/U$1 ( \5141 , \5140 );
not \mul_6_18_g43971/U$4 ( \5142 , \5141 );
or \mul_6_18_g43971/U$2 ( \5143 , \5139 , \5142 );
not \g45695/U$2 ( \5144 , \4008 );
nand \g45695/U$1 ( \5145 , \5144 , \2779 );
nand \mul_6_18_g43971/U$1 ( \5146 , \5143 , \5145 );
nand \mul_6_18_g43044/U$1 ( \5147 , \2434 , \5146 );
nand \mul_6_18_g42930/U$1 ( \5148 , \5138 , \5147 );
not \mul_6_18_g43723/U$3 ( \5149 , \2116 );
not \mul_6_18_g43723/U$4 ( \5150 , \2340 );
or \mul_6_18_g43723/U$2 ( \5151 , \5149 , \5150 );
nand \mul_6_18_g43723/U$1 ( \5152 , \5151 , \2663 );
not \mul_6_18_g45290/U$2 ( \5153 , \2340 );
nand \mul_6_18_g45290/U$1 ( \5154 , \5153 , \2058 );
nand \mul_6_18_g43676/U$1 ( \5155 , \5152 , \2335 , \5154 );
not \mul_6_18_g43675/U$1 ( \5156 , \5155 );
and \mul_6_18_g45145/U$1 ( \5157 , \5148 , \5156 );
not \mul_6_18_g42610/U$4 ( \5158 , \5157 );
or \mul_6_18_g42610/U$2 ( \5159 , \5130 , \5158 );
or \mul_6_18_g42610/U$5 ( \5160 , \5157 , \5129 );
nand \mul_6_18_g42610/U$1 ( \5161 , \5159 , \5160 );
not \mul_6_18_g44091/U$3 ( \5162 , \2168 );
not \mul_6_18_g44091/U$4 ( \5163 , \2367 );
or \mul_6_18_g44091/U$2 ( \5164 , \5162 , \5163 );
not \mul_6_18_g44562/U$1 ( \5165 , \2367 );
nand \mul_6_18_g44361/U$1 ( \5166 , \5165 , \3154 );
nand \mul_6_18_g44091/U$1 ( \5167 , \5164 , \5166 );
and \mul_6_18_g43233/U$2 ( \5168 , \2400 , \5167 );
and \mul_6_18_g43233/U$3 ( \5169 , \2403 , \4988 );
nor \mul_6_18_g43233/U$1 ( \5170 , \5168 , \5169 );
not \mul_6_18_g43231/U$1 ( \5171 , \5170 );
xor \mul_6_18_g42521/U$1 ( \5172 , \5161 , \5171 );
xor \mul_6_18_g42201/U$4 ( \5173 , \5113 , \5172 );
and \mul_6_18_g42816/U$2 ( \5174 , \5148 , \5156 );
not \mul_6_18_g42816/U$4 ( \5175 , \5148 );
and \mul_6_18_g42816/U$3 ( \5176 , \5175 , \5155 );
nor \mul_6_18_g42816/U$1 ( \5177 , \5174 , \5176 );
not \mul_6_18_g42347/U$3 ( \5178 , \5177 );
nand \mul_6_18_g43659/U$1 ( \5179 , \2358 , \2058 );
not \mul_6_18_g43658/U$1 ( \5180 , \5179 );
not \mul_6_18_g42595/U$3 ( \5181 , \5180 );
not \mul_6_18_g42955/U$3 ( \5182 , \2447 );
not \mul_6_18_g43990/U$3 ( \5183 , \2112 );
not \mul_6_18_g43990/U$4 ( \5184 , \4008 );
or \mul_6_18_g43990/U$2 ( \5185 , \5183 , \5184 );
not \mul_6_18_g45252/U$2 ( \5186 , \2112 );
nand \mul_6_18_g45252/U$1 ( \5187 , \5186 , \2418 );
nand \mul_6_18_g43990/U$1 ( \5188 , \5185 , \5187 );
not \mul_6_18_g43989/U$1 ( \5189 , \5188 );
not \mul_6_18_g42955/U$4 ( \5190 , \5189 );
and \mul_6_18_g42955/U$2 ( \5191 , \5182 , \5190 );
and \mul_6_18_g42955/U$5 ( \5192 , \2434 , \5135 );
nor \mul_6_18_g42955/U$1 ( \5193 , \5191 , \5192 );
not \mul_6_18_g42954/U$1 ( \5194 , \5193 );
not \mul_6_18_g42595/U$4 ( \5195 , \5194 );
or \mul_6_18_g42595/U$2 ( \5196 , \5181 , \5195 );
or \mul_6_18_g42679/U$2 ( \5197 , \5194 , \5180 );
not \mul_6_18_g44019/U$3 ( \5198 , \1998 );
not \mul_6_18_g44019/U$4 ( \5199 , \2607 );
or \mul_6_18_g44019/U$2 ( \5200 , \5198 , \5199 );
nand \mul_6_18_g44330/U$1 ( \5201 , \2626 , \2489 );
nand \mul_6_18_g44019/U$1 ( \5202 , \5200 , \5201 );
not \mul_6_18_g42986/U$3 ( \5203 , \5202 );
not \mul_6_18_g42986/U$4 ( \5204 , \2603 );
or \mul_6_18_g42986/U$2 ( \5205 , \5203 , \5204 );
not \mul_6_18_g43997/U$3 ( \5206 , \2812 );
not \mul_6_18_g43997/U$4 ( \5207 , \2629 );
or \mul_6_18_g43997/U$2 ( \5208 , \5206 , \5207 );
nand \mul_6_18_g44308/U$1 ( \5209 , \2606 , \2811 );
nand \mul_6_18_g43997/U$1 ( \5210 , \5208 , \5209 );
nand \mul_6_18_g43033/U$1 ( \5211 , \2842 , \5210 );
nand \mul_6_18_g42986/U$1 ( \5212 , \5205 , \5211 );
nand \mul_6_18_g42679/U$1 ( \5213 , \5197 , \5212 );
nand \mul_6_18_g42595/U$1 ( \5214 , \5196 , \5213 );
not \mul_6_18_g42347/U$4 ( \5215 , \5214 );
or \mul_6_18_g42347/U$2 ( \5216 , \5178 , \5215 );
or \g45738/U$2 ( \5217 , \5214 , \5177 );
not \mul_6_18_g43963/U$3 ( \5218 , \2111 );
not \mul_6_18_g43963/U$4 ( \5219 , \2929 );
or \mul_6_18_g43963/U$2 ( \5220 , \5218 , \5219 );
nand \mul_6_18_g44291/U$1 ( \5221 , \2236 , \2779 );
nand \mul_6_18_g43963/U$1 ( \5222 , \5220 , \5221 );
not \mul_6_18_g43369/U$3 ( \5223 , \5222 );
not \mul_6_18_g43369/U$4 ( \5224 , \2222 );
or \mul_6_18_g43369/U$2 ( \5225 , \5223 , \5224 );
not \mul_6_18_g43948/U$3 ( \5226 , \2107 );
not \mul_6_18_g43948/U$4 ( \5227 , \2217 );
or \mul_6_18_g43948/U$2 ( \5228 , \5226 , \5227 );
not \mul_6_18_g44593/U$1 ( \5229 , \2107 );
nand \mul_6_18_g44265/U$1 ( \5230 , \2236 , \5229 );
nand \mul_6_18_g43948/U$1 ( \5231 , \5228 , \5230 );
nand \mul_6_18_g43569/U$1 ( \5232 , \5231 , \2934 );
nand \mul_6_18_g43369/U$1 ( \5233 , \5225 , \5232 );
not \mul_6_18_g42688/U$3 ( \5234 , \5233 );
not \mul_6_18_g44057/U$3 ( \5235 , \2006 );
not \mul_6_18_g44057/U$4 ( \5236 , \3224 );
or \mul_6_18_g44057/U$2 ( \5237 , \5235 , \5236 );
nand \mul_6_18_g44351/U$1 ( \5238 , \2256 , \2795 );
nand \mul_6_18_g44057/U$1 ( \5239 , \5237 , \5238 );
not \mul_6_18_g43305/U$3 ( \5240 , \5239 );
not \mul_6_18_g43305/U$4 ( \5241 , \2938 );
or \mul_6_18_g43305/U$2 ( \5242 , \5240 , \5241 );
not \mul_6_18_g44030/U$3 ( \5243 , \2463 );
not \mul_6_18_g44030/U$4 ( \5244 , \2251 );
or \mul_6_18_g44030/U$2 ( \5245 , \5243 , \5244 );
nand \mul_6_18_g44324/U$1 ( \5246 , \2256 , \2468 );
nand \mul_6_18_g44030/U$1 ( \5247 , \5245 , \5246 );
nand \mul_6_18_g43464/U$1 ( \5248 , \5247 , \3232 );
nand \mul_6_18_g43305/U$1 ( \5249 , \5242 , \5248 );
not \mul_6_18_g42688/U$4 ( \5250 , \5249 );
or \mul_6_18_g42688/U$2 ( \5251 , \5234 , \5250 );
or \g45745/U$2 ( \5252 , \5249 , \5233 );
not \mul_6_18_g44081/U$3 ( \5253 , \2168 );
not \mul_6_18_g44081/U$4 ( \5254 , \2715 );
or \mul_6_18_g44081/U$2 ( \5255 , \5253 , \5254 );
nand \mul_6_18_g44363/U$1 ( \5256 , \2972 , \3154 );
nand \mul_6_18_g44081/U$1 ( \5257 , \5255 , \5256 );
not \mul_6_18_g43265/U$3 ( \5258 , \5257 );
not \mul_6_18_g43265/U$4 ( \5259 , \3323 );
or \mul_6_18_g43265/U$2 ( \5260 , \5258 , \5259 );
not \mul_6_18_g44065/U$3 ( \5261 , \2179 );
not \mul_6_18_g44065/U$4 ( \5262 , \2715 );
or \mul_6_18_g44065/U$2 ( \5263 , \5261 , \5262 );
nand \mul_6_18_g44348/U$1 ( \5264 , \2972 , \2185 );
nand \mul_6_18_g44065/U$1 ( \5265 , \5263 , \5264 );
nand \mul_6_18_g43634/U$1 ( \5266 , \2733 , \5265 );
nand \mul_6_18_g43265/U$1 ( \5267 , \5260 , \5266 );
nand \g45745/U$1 ( \5268 , \5252 , \5267 );
nand \mul_6_18_g42688/U$1 ( \5269 , \5251 , \5268 );
nand \g45738/U$1 ( \5270 , \5217 , \5269 );
nand \mul_6_18_g42347/U$1 ( \5271 , \5216 , \5270 );
and \mul_6_18_g42201/U$3 ( \5272 , \5173 , \5271 );
and \mul_6_18_g42201/U$5 ( \5273 , \5113 , \5172 );
or \mul_6_18_g42201/U$2 ( \5274 , \5272 , \5273 );
xor \mul_6_18_g42085/U$1 ( \5275 , \5111 , \5274 );
not \mul_6_18_g42685/U$3 ( \5276 , \5170 );
not \mul_6_18_g42685/U$4 ( \5277 , \5129 );
or \mul_6_18_g42685/U$2 ( \5278 , \5276 , \5277 );
nand \mul_6_18_g42685/U$1 ( \5279 , \5278 , \5157 );
nand \mul_6_18_g42897/U$1 ( \5280 , \5128 , \5171 );
nand \mul_6_18_g42599/U$1 ( \5281 , \5279 , \5280 );
not \mul_6_18_g43195/U$3 ( \5282 , \5126 );
not \mul_6_18_g43195/U$4 ( \5283 , \2349 );
or \mul_6_18_g43195/U$2 ( \5284 , \5282 , \5283 );
and \mul_6_18_g44105/U$2 ( \5285 , \3154 , \2330 );
not \mul_6_18_g44105/U$4 ( \5286 , \3154 );
and \mul_6_18_g44105/U$3 ( \5287 , \5286 , \2329 );
nor \mul_6_18_g44105/U$1 ( \5288 , \5285 , \5287 );
nand \mul_6_18_g43537/U$1 ( \5289 , \2359 , \5288 );
nand \mul_6_18_g43195/U$1 ( \5290 , \5284 , \5289 );
not \mul_6_18_g43722/U$3 ( \5291 , \2116 );
not \mul_6_18_g43722/U$4 ( \5292 , \2295 );
or \mul_6_18_g43722/U$2 ( \5293 , \5291 , \5292 );
nand \mul_6_18_g43722/U$1 ( \5294 , \5293 , \2329 );
not \mul_6_18_g45242/U$2 ( \5295 , \2295 );
nand \mul_6_18_g45242/U$1 ( \5296 , \5295 , \2058 );
and \mul_6_18_g43677/U$1 ( \5297 , \5294 , \2311 , \5296 );
not \mul_6_18_g43952/U$3 ( \5298 , \2107 );
not \mul_6_18_g43952/U$4 ( \5299 , \2423 );
or \mul_6_18_g43952/U$2 ( \5300 , \5298 , \5299 );
nand \mul_6_18_g44259/U$1 ( \5301 , \2424 , \2745 );
nand \mul_6_18_g43952/U$1 ( \5302 , \5300 , \5301 );
not \mul_6_18_g42934/U$3 ( \5303 , \5302 );
not \mul_6_18_g42934/U$4 ( \5304 , \2586 );
or \mul_6_18_g42934/U$2 ( \5305 , \5303 , \5304 );
not \mul_6_18_g43951/U$3 ( \5306 , \2092 );
not \mul_6_18_g43951/U$4 ( \5307 , \2423 );
or \mul_6_18_g43951/U$2 ( \5308 , \5306 , \5307 );
nand \mul_6_18_g44269/U$1 ( \5309 , \5140 , \2754 );
nand \mul_6_18_g43951/U$1 ( \5310 , \5308 , \5309 );
nand \mul_6_18_g43024/U$1 ( \5311 , \2434 , \5310 );
nand \mul_6_18_g42934/U$1 ( \5312 , \5305 , \5311 );
xor \mul_6_18_g42771/U$1 ( \5313 , \5297 , \5312 );
xor \mul_6_18_g42446/U$1 ( \5314 , \5290 , \5313 );
nand \mul_6_18_g43657/U$1 ( \5315 , \4287 , \2058 );
not \mul_6_18_g42682/U$3 ( \5316 , \5315 );
not \mul_6_18_g42939/U$3 ( \5317 , \5146 );
not \mul_6_18_g42939/U$4 ( \5318 , \2586 );
or \mul_6_18_g42939/U$2 ( \5319 , \5317 , \5318 );
nand \mul_6_18_g45643/U$1 ( \5320 , \2434 , \5302 );
nand \mul_6_18_g42939/U$1 ( \5321 , \5319 , \5320 );
not \mul_6_18_g42938/U$1 ( \5322 , \5321 );
not \mul_6_18_g42682/U$4 ( \5323 , \5322 );
or \mul_6_18_g42682/U$2 ( \5324 , \5316 , \5323 );
not \mul_6_18_g43998/U$3 ( \5325 , \2112 );
not \mul_6_18_g43998/U$4 ( \5326 , \2834 );
or \mul_6_18_g43998/U$2 ( \5327 , \5325 , \5326 );
nand \mul_6_18_g44301/U$1 ( \5328 , \2606 , \2824 );
nand \mul_6_18_g43998/U$1 ( \5329 , \5327 , \5328 );
not \mul_6_18_g42998/U$3 ( \5330 , \5329 );
not \mul_6_18_g42998/U$4 ( \5331 , \2907 );
or \mul_6_18_g42998/U$2 ( \5332 , \5330 , \5331 );
not \mul_6_18_g45236/U$2 ( \5333 , \5050 );
nand \mul_6_18_g45236/U$1 ( \5334 , \5333 , \2842 );
nand \mul_6_18_g42998/U$1 ( \5335 , \5332 , \5334 );
nand \mul_6_18_g42682/U$1 ( \5336 , \5324 , \5335 );
not \mul_6_18_g45231/U$2 ( \5337 , \5315 );
nand \mul_6_18_g45231/U$1 ( \5338 , \5337 , \5321 );
nand \mul_6_18_g42596/U$1 ( \5339 , \5336 , \5338 );
xor \mul_6_18_g42446/U$1_r1 ( \5340 , \5314 , \5339 );
xor \mul_6_18_g42269/U$1 ( \5341 , \5281 , \5340 );
not \mul_6_18_g43264/U$3 ( \5342 , \5265 );
not \mul_6_18_g43264/U$4 ( \5343 , \2729 );
or \mul_6_18_g43264/U$2 ( \5344 , \5342 , \5343 );
nand \mul_6_18_g43538/U$1 ( \5345 , \4327 , \5095 );
nand \mul_6_18_g43264/U$1 ( \5346 , \5344 , \5345 );
not \mul_6_18_g42895/U$2 ( \5347 , \5346 );
and \g45529/U$2 ( \5348 , \2364 , \2144 );
not \g45529/U$4 ( \5349 , \2364 );
and \g45529/U$3 ( \5350 , \5349 , \2145 );
or \g45529/U$1 ( \5351 , \5348 , \5350 );
and \mul_6_18_g43230/U$2 ( \5352 , \2400 , \5351 );
and \mul_6_18_g43230/U$3 ( \5353 , \2403 , \5167 );
nor \mul_6_18_g43230/U$1 ( \5354 , \5352 , \5353 );
nand \mul_6_18_g42895/U$1 ( \5355 , \5347 , \5354 );
and \mul_6_18_g44120/U$2 ( \5356 , \2058 , \2335 );
not \mul_6_18_g44120/U$4 ( \5357 , \2058 );
and \mul_6_18_g44120/U$3 ( \5358 , \5357 , \2330 );
nor \mul_6_18_g44120/U$1 ( \5359 , \5356 , \5358 );
not \mul_6_18_g43198/U$3 ( \5360 , \5359 );
not \mul_6_18_g43198/U$4 ( \5361 , \2349 );
or \mul_6_18_g43198/U$2 ( \5362 , \5360 , \5361 );
nand \mul_6_18_g43564/U$1 ( \5363 , \2359 , \5118 );
nand \mul_6_18_g43198/U$1 ( \5364 , \5362 , \5363 );
and \mul_6_18_g42808/U$2 ( \5365 , \5355 , \5364 );
not \mul_6_18_g42894/U$2 ( \5366 , \5346 );
nor \mul_6_18_g42894/U$1 ( \5367 , \5366 , \5354 );
nor \mul_6_18_g42808/U$1 ( \5368 , \5365 , \5367 );
not \mul_6_18_g42724/U$1 ( \5369 , \5368 );
not \g45788/U$3 ( \5370 , \5369 );
and \g45708/U$2 ( \5371 , \5231 , \2222 );
and \g45708/U$3 ( \5372 , \5073 , \3430 );
nor \g45708/U$1 ( \5373 , \5371 , \5372 );
and \g45706/U$2 ( \5374 , \5210 , \4002 );
and \g45706/U$3 ( \5375 , \2842 , \5329 );
nor \g45706/U$1 ( \5376 , \5374 , \5375 );
xor \mul_6_18_g42552/U$4 ( \5377 , \5373 , \5376 );
and \g45752/U$2 ( \5378 , \2274 , \5247 );
not \mul_6_18_g45237/U$2 ( \5379 , \5084 );
nor \mul_6_18_g45237/U$1 ( \5380 , \5379 , \2284 );
nor \g45752/U$1 ( \5381 , \5378 , \5380 );
and \mul_6_18_g42552/U$3 ( \5382 , \5377 , \5381 );
and \mul_6_18_g42552/U$5 ( \5383 , \5373 , \5376 );
or \mul_6_18_g42552/U$2 ( \5384 , \5382 , \5383 );
not \mul_6_18_g42551/U$1 ( \5385 , \5384 );
not \g45788/U$4 ( \5386 , \5385 );
or \g45788/U$2 ( \5387 , \5370 , \5386 );
not \g45789/U$3 ( \5388 , \5368 );
not \g45789/U$4 ( \5389 , \5384 );
or \g45789/U$2 ( \5390 , \5388 , \5389 );
xor \mul_6_18_g42617/U$1 ( \5391 , \5315 , \5321 );
xor \mul_6_18_g42617/U$1_r1 ( \5392 , \5391 , \5335 );
not \mul_6_18_g42579/U$1 ( \5393 , \5392 );
nand \g45789/U$1 ( \5394 , \5390 , \5393 );
nand \g45788/U$1 ( \5395 , \5387 , \5394 );
xor \mul_6_18_g42269/U$1_r1 ( \5396 , \5341 , \5395 );
xor \mul_6_18_g42085/U$1_r1 ( \5397 , \5275 , \5396 );
not \mul_6_18_g42083/U$1 ( \5398 , \5397 );
not \mul_6_18_g42487/U$3 ( \5399 , \5384 );
not \mul_6_18_g42487/U$4 ( \5400 , \5393 );
or \mul_6_18_g42487/U$2 ( \5401 , \5399 , \5400 );
nand \mul_6_18_g42493/U$1 ( \5402 , \5392 , \5385 );
nand \mul_6_18_g42487/U$1 ( \5403 , \5401 , \5402 );
and \mul_6_18_g42430/U$2 ( \5404 , \5403 , \5369 );
not \mul_6_18_g42430/U$4 ( \5405 , \5403 );
and \mul_6_18_g42430/U$3 ( \5406 , \5405 , \5368 );
nor \mul_6_18_g42430/U$1 ( \5407 , \5404 , \5406 );
not \mul_6_18_g42357/U$1 ( \5408 , \5407 );
not \mul_6_18_g42168/U$3 ( \5409 , \5408 );
xor \mul_6_18_g42552/U$1 ( \5410 , \5373 , \5376 );
xor \mul_6_18_g42552/U$1_r1 ( \5411 , \5410 , \5381 );
xor \g45869/U$1 ( \5412 , \5346 , \5364 );
xor \g45869/U$1_r1 ( \5413 , \5412 , \5354 );
xor \mul_6_18_g42332/U$4 ( \5414 , \5411 , \5413 );
not \mul_6_18_g43962/U$3 ( \5415 , \2094 );
not \mul_6_18_g44705/U$1 ( \5416 , \2236 );
not \mul_6_18_g43962/U$4 ( \5417 , \5416 );
or \mul_6_18_g43962/U$2 ( \5418 , \5415 , \5417 );
nand \mul_6_18_g44274/U$1 ( \5419 , \2226 , \2500 );
nand \mul_6_18_g43962/U$1 ( \5420 , \5418 , \5419 );
not \mul_6_18_g43357/U$3 ( \5421 , \5420 );
not \mul_6_18_g43357/U$4 ( \5422 , \2222 );
or \mul_6_18_g43357/U$2 ( \5423 , \5421 , \5422 );
nand \mul_6_18_g43602/U$1 ( \5424 , \5222 , \2934 );
nand \mul_6_18_g43357/U$1 ( \5425 , \5423 , \5424 );
buf \fopt45575/U$1 ( \5426 , \2907 );
not \mul_6_18_g45224/U$3 ( \5427 , \5426 );
not \mul_6_18_g44018/U$3 ( \5428 , \2463 );
not \mul_6_18_g44018/U$4 ( \5429 , \2629 );
or \mul_6_18_g44018/U$2 ( \5430 , \5428 , \5429 );
nand \mul_6_18_g44332/U$1 ( \5431 , \2468 , \2606 );
nand \mul_6_18_g44018/U$1 ( \5432 , \5430 , \5431 );
not \mul_6_18_g45224/U$4 ( \5433 , \5432 );
or \mul_6_18_g45224/U$2 ( \5434 , \5427 , \5433 );
nand \mul_6_18_g43039/U$1 ( \5435 , \2842 , \5202 );
nand \mul_6_18_g45224/U$1 ( \5436 , \5434 , \5435 );
xor \mul_6_18_g42559/U$4 ( \5437 , \5425 , \5436 );
not \mul_6_18_g44056/U$3 ( \5438 , \2179 );
not \mul_6_18_g44056/U$4 ( \5439 , \2277 );
or \mul_6_18_g44056/U$2 ( \5440 , \5438 , \5439 );
nand \mul_6_18_g44352/U$1 ( \5441 , \2252 , \2185 );
nand \mul_6_18_g44056/U$1 ( \5442 , \5440 , \5441 );
not \mul_6_18_g43307/U$3 ( \5443 , \5442 );
not \mul_6_18_g43307/U$4 ( \5444 , \2274 );
or \mul_6_18_g43307/U$2 ( \5445 , \5443 , \5444 );
nand \mul_6_18_g43466/U$1 ( \5446 , \2285 , \5239 );
nand \mul_6_18_g43307/U$1 ( \5447 , \5445 , \5446 );
and \mul_6_18_g42559/U$3 ( \5448 , \5437 , \5447 );
and \mul_6_18_g42559/U$5 ( \5449 , \5425 , \5436 );
or \mul_6_18_g42559/U$2 ( \5450 , \5448 , \5449 );
not \mul_6_18_g43991/U$3 ( \5451 , \2810 );
not \mul_6_18_g43991/U$4 ( \5452 , \4008 );
or \mul_6_18_g43991/U$2 ( \5453 , \5451 , \5452 );
nand \mul_6_18_g44304/U$1 ( \5454 , \2418 , \2811 );
nand \mul_6_18_g43991/U$1 ( \5455 , \5453 , \5454 );
not \mul_6_18_g42943/U$3 ( \5456 , \5455 );
not \mul_6_18_g42943/U$4 ( \5457 , \2586 );
or \mul_6_18_g42943/U$2 ( \5458 , \5456 , \5457 );
nand \mul_6_18_g43027/U$1 ( \5459 , \2434 , \5188 );
nand \mul_6_18_g42943/U$1 ( \5460 , \5458 , \5459 );
not \mul_6_18_g43724/U$3 ( \5461 , \2116 );
not \mul_6_18_g43724/U$4 ( \5462 , \2387 );
or \mul_6_18_g43724/U$2 ( \5463 , \5461 , \5462 );
nand \mul_6_18_g43724/U$1 ( \5464 , \5463 , \2714 );
not \mul_6_18_g45279/U$2 ( \5465 , \2387 );
nand \mul_6_18_g45279/U$1 ( \5466 , \5465 , \2058 );
nand \mul_6_18_g43674/U$1 ( \5467 , \5464 , \2663 , \5466 );
not \mul_6_18_g43673/U$1 ( \5468 , \5467 );
nand \mul_6_18_g45142/U$1 ( \5469 , \5460 , \5468 );
not \mul_6_18_g44107/U$3 ( \5470 , \2056 );
not \mul_6_18_g44107/U$4 ( \5471 , \2367 );
or \mul_6_18_g44107/U$2 ( \5472 , \5470 , \5471 );
nand \mul_6_18_g44383/U$1 ( \5473 , \2663 , \3360 );
nand \mul_6_18_g44107/U$1 ( \5474 , \5472 , \5473 );
not \mul_6_18_g43210/U$3 ( \5475 , \5474 );
not \mul_6_18_g43210/U$4 ( \5476 , \2400 );
or \mul_6_18_g43210/U$2 ( \5477 , \5475 , \5476 );
nand \mul_6_18_g43444/U$1 ( \5478 , \2403 , \5351 );
nand \mul_6_18_g43210/U$1 ( \5479 , \5477 , \5478 );
not \mul_6_18_g43209/U$1 ( \5480 , \5479 );
nand \mul_6_18_g42668/U$1 ( \5481 , \5469 , \5480 );
and \mul_6_18_g42462/U$2 ( \5482 , \5450 , \5481 );
nor \mul_6_18_g42667/U$1 ( \5483 , \5469 , \5480 );
nor \mul_6_18_g42462/U$1 ( \5484 , \5482 , \5483 );
and \mul_6_18_g42332/U$3 ( \5485 , \5414 , \5484 );
and \mul_6_18_g42332/U$5 ( \5486 , \5411 , \5413 );
or \mul_6_18_g42332/U$2 ( \5487 , \5485 , \5486 );
not \mul_6_18_g42168/U$4 ( \5488 , \5487 );
or \mul_6_18_g42168/U$2 ( \5489 , \5409 , \5488 );
xor \mul_6_18_g42201/U$1 ( \5490 , \5113 , \5172 );
xor \mul_6_18_g42201/U$1_r1 ( \5491 , \5490 , \5271 );
nand \mul_6_18_g42168/U$1 ( \5492 , \5489 , \5491 );
or \mul_6_18_g45167/U$1 ( \5493 , \5487 , \5408 );
nand \mul_6_18_g42152/U$1 ( \5494 , \5492 , \5493 );
not \mul_6_18_g42132/U$1 ( \5495 , \5494 );
nand \mul_6_18_g42057/U$1 ( \5496 , \5398 , \5495 );
and \mul_6_18_g42265/U$2 ( \5497 , \5487 , \5408 );
not \mul_6_18_g42265/U$4 ( \5498 , \5487 );
and \mul_6_18_g42265/U$3 ( \5499 , \5498 , \5407 );
nor \mul_6_18_g42265/U$1 ( \5500 , \5497 , \5499 );
not \mul_6_18_g42200/U$1 ( \5501 , \5491 );
and \mul_6_18_g42164/U$2 ( \5502 , \5500 , \5501 );
not \mul_6_18_g42164/U$4 ( \5503 , \5500 );
and \mul_6_18_g42164/U$3 ( \5504 , \5503 , \5491 );
nor \mul_6_18_g42164/U$1 ( \5505 , \5502 , \5504 );
xor \mul_6_18_g42332/U$1 ( \5506 , \5411 , \5413 );
xor \mul_6_18_g42332/U$1_r1 ( \5507 , \5506 , \5484 );
xor \mul_6_18_g42383/U$1 ( \5508 , \5177 , \5214 );
xnor \mul_6_18_g42383/U$1_r1 ( \5509 , \5508 , \5269 );
nand \mul_6_18_g42279/U$1 ( \5510 , \5507 , \5509 );
xor \mul_6_18_g45207/U$1 ( \5511 , \5179 , \5194 );
xor \mul_6_18_g45207/U$1_r1 ( \5512 , \5511 , \5212 );
not \mul_6_18_g42395/U$3 ( \5513 , \5512 );
xor \mul_6_18_g42736/U$1 ( \5514 , \5233 , \5249 );
xnor \mul_6_18_g42736/U$1_r1 ( \5515 , \5514 , \5267 );
not \mul_6_18_g42395/U$4 ( \5516 , \5515 );
or \mul_6_18_g42395/U$2 ( \5517 , \5513 , \5516 );
not \mul_6_18_g44082/U$3 ( \5518 , \2144 );
not \mul_6_18_g44082/U$4 ( \5519 , \2715 );
or \mul_6_18_g44082/U$2 ( \5520 , \5518 , \5519 );
nand \mul_6_18_g44374/U$1 ( \5521 , \2972 , \2145 );
nand \mul_6_18_g44082/U$1 ( \5522 , \5520 , \5521 );
not \mul_6_18_g43268/U$3 ( \5523 , \5522 );
not \mul_6_18_g43268/U$4 ( \5524 , \3323 );
or \mul_6_18_g43268/U$2 ( \5525 , \5523 , \5524 );
nand \mul_6_18_g43536/U$1 ( \5526 , \4327 , \5257 );
nand \mul_6_18_g43268/U$1 ( \5527 , \5525 , \5526 );
not \mul_6_18_g44129/U$3 ( \5528 , \2058 );
not \mul_6_18_g44129/U$4 ( \5529 , \2367 );
or \mul_6_18_g44129/U$2 ( \5530 , \5528 , \5529 );
nand \mul_6_18_g44396/U$1 ( \5531 , \5165 , \2116 );
nand \mul_6_18_g44129/U$1 ( \5532 , \5530 , \5531 );
not \mul_6_18_g43234/U$3 ( \5533 , \5532 );
not \mul_6_18_g43234/U$4 ( \5534 , \2400 );
or \mul_6_18_g43234/U$2 ( \5535 , \5533 , \5534 );
nand \mul_6_18_g43540/U$1 ( \5536 , \2403 , \5474 );
nand \mul_6_18_g43234/U$1 ( \5537 , \5535 , \5536 );
xor \mul_6_18_g42480/U$4 ( \5538 , \5527 , \5537 );
and \mul_6_18_g42817/U$2 ( \5539 , \5460 , \5468 );
not \mul_6_18_g42817/U$4 ( \5540 , \5460 );
and \mul_6_18_g42817/U$3 ( \5541 , \5540 , \5467 );
nor \mul_6_18_g42817/U$1 ( \5542 , \5539 , \5541 );
and \mul_6_18_g42480/U$3 ( \5543 , \5538 , \5542 );
and \mul_6_18_g42480/U$5 ( \5544 , \5527 , \5537 );
or \mul_6_18_g42480/U$2 ( \5545 , \5543 , \5544 );
nand \mul_6_18_g42395/U$1 ( \5546 , \5517 , \5545 );
not \mul_6_18_g42632/U$1 ( \5547 , \5515 );
not \mul_6_18_g42555/U$1 ( \5548 , \5512 );
nand \mul_6_18_g42515/U$1 ( \5549 , \5547 , \5548 );
nand \mul_6_18_g42350/U$1 ( \5550 , \5546 , \5549 );
and \mul_6_18_g42227/U$2 ( \5551 , \5510 , \5550 );
nor \mul_6_18_g42278/U$1 ( \5552 , \5507 , \5509 );
nor \mul_6_18_g42227/U$1 ( \5553 , \5551 , \5552 );
nand \mul_6_18_g42092/U$1 ( \5554 , \5505 , \5553 );
and \mul_6_18_g42039/U$1 ( \5555 , \5496 , \5554 );
not \mul_6_18_g41969/U$3 ( \5556 , \5555 );
nand \mul_6_18_g43662/U$1 ( \5557 , \2403 , \2058 );
not \mul_6_18_g44006/U$3 ( \5558 , \1998 );
not \mul_6_18_g44006/U$4 ( \5559 , \2423 );
or \mul_6_18_g44006/U$2 ( \5560 , \5558 , \5559 );
not \mul_6_18_g44978/U$1 ( \5561 , \2423 );
nand \mul_6_18_g44319/U$1 ( \5562 , \5561 , \2489 );
nand \mul_6_18_g44006/U$1 ( \5563 , \5560 , \5562 );
not \mul_6_18_g42949/U$3 ( \5564 , \5563 );
not \mul_6_18_g42949/U$4 ( \5565 , \4264 );
or \mul_6_18_g42949/U$2 ( \5566 , \5564 , \5565 );
nand \mul_6_18_g43007/U$1 ( \5567 , \2434 , \5455 );
nand \mul_6_18_g42949/U$1 ( \5568 , \5566 , \5567 );
xor \mul_6_18_g42615/U$1 ( \5569 , \5557 , \5568 );
not \mul_6_18_g44047/U$3 ( \5570 , \2006 );
not \mul_6_18_g44047/U$4 ( \5571 , \2629 );
or \mul_6_18_g44047/U$2 ( \5572 , \5570 , \5571 );
nand \mul_6_18_g44342/U$1 ( \5573 , \2606 , \2795 );
nand \mul_6_18_g44047/U$1 ( \5574 , \5572 , \5573 );
not \mul_6_18_g42978/U$3 ( \5575 , \5574 );
not \mul_6_18_g42978/U$4 ( \5576 , \2603 );
or \mul_6_18_g42978/U$2 ( \5577 , \5575 , \5576 );
nand \mul_6_18_g43041/U$1 ( \5578 , \2842 , \5432 );
nand \mul_6_18_g42978/U$1 ( \5579 , \5577 , \5578 );
xor \mul_6_18_g42615/U$1_r1 ( \5580 , \5569 , \5579 );
not \mul_6_18_g44007/U$3 ( \5581 , \2463 );
not \mul_6_18_g44007/U$4 ( \5582 , \2419 );
or \mul_6_18_g44007/U$2 ( \5583 , \5581 , \5582 );
nand \mul_6_18_g44333/U$1 ( \5584 , \5140 , \2468 );
nand \mul_6_18_g44007/U$1 ( \5585 , \5583 , \5584 );
not \mul_6_18_g42946/U$3 ( \5586 , \5585 );
not \mul_6_18_g42946/U$4 ( \5587 , \2586 );
or \mul_6_18_g42946/U$2 ( \5588 , \5586 , \5587 );
nand \mul_6_18_g43026/U$1 ( \5589 , \2434 , \5563 );
nand \mul_6_18_g42946/U$1 ( \5590 , \5588 , \5589 );
not \mul_6_18_g45248/U$2 ( \5591 , \1434 );
nand \mul_6_18_g45248/U$1 ( \5592 , \5591 , \2116 );
and \mul_6_18_g43671/U$2 ( \5593 , \2280 , \5592 );
not \mul_6_18_g43731/U$3 ( \5594 , \2058 );
not \mul_6_18_g43731/U$4 ( \5595 , \1434 );
or \mul_6_18_g43731/U$2 ( \5596 , \5594 , \5595 );
nand \mul_6_18_g43731/U$1 ( \5597 , \5596 , \2714 );
nor \mul_6_18_g43671/U$1 ( \5598 , \5593 , \5597 );
nand \mul_6_18_g45651/U$1 ( \5599 , \5590 , \5598 );
nand \mul_6_18_g42503/U$1 ( \5600 , \5580 , \5599 );
not \mul_6_18_g43987/U$3 ( \5601 , \2810 );
not \mul_6_18_g43987/U$4 ( \5602 , \2929 );
or \mul_6_18_g43987/U$2 ( \5603 , \5601 , \5602 );
nand \mul_6_18_g44295/U$1 ( \5604 , \2236 , \2811 );
nand \mul_6_18_g43987/U$1 ( \5605 , \5603 , \5604 );
not \mul_6_18_g43382/U$3 ( \5606 , \5605 );
not \mul_6_18_g43382/U$4 ( \5607 , \2222 );
or \mul_6_18_g43382/U$2 ( \5608 , \5606 , \5607 );
not \mul_6_18_g43988/U$3 ( \5609 , \2112 );
not \mul_6_18_g43988/U$4 ( \5610 , \2217 );
or \mul_6_18_g43988/U$2 ( \5611 , \5609 , \5610 );
nand \mul_6_18_g44297/U$1 ( \5612 , \3215 , \2824 );
nand \mul_6_18_g43988/U$1 ( \5613 , \5611 , \5612 );
nand \mul_6_18_g43623/U$1 ( \5614 , \5613 , \3430 );
nand \mul_6_18_g43382/U$1 ( \5615 , \5608 , \5614 );
not \mul_6_18_g44046/U$3 ( \5616 , \2179 );
not \mul_6_18_g44046/U$4 ( \5617 , \2629 );
or \mul_6_18_g44046/U$2 ( \5618 , \5616 , \5617 );
nand \mul_6_18_g44343/U$1 ( \5619 , \2606 , \2185 );
nand \mul_6_18_g44046/U$1 ( \5620 , \5618 , \5619 );
not \mul_6_18_g42991/U$3 ( \5621 , \5620 );
not \mul_6_18_g42991/U$4 ( \5622 , \2907 );
or \mul_6_18_g42991/U$2 ( \5623 , \5621 , \5622 );
nand \mul_6_18_g43014/U$1 ( \5624 , \2623 , \5574 );
nand \mul_6_18_g42991/U$1 ( \5625 , \5623 , \5624 );
xor \mul_6_18_g42563/U$4 ( \5626 , \5615 , \5625 );
not \mul_6_18_g44073/U$3 ( \5627 , \2144 );
not \mul_6_18_g44073/U$4 ( \5628 , \2251 );
or \mul_6_18_g44073/U$2 ( \5629 , \5627 , \5628 );
nand \mul_6_18_g44370/U$1 ( \5630 , \2256 , \2145 );
nand \mul_6_18_g44073/U$1 ( \5631 , \5629 , \5630 );
not \mul_6_18_g43308/U$3 ( \5632 , \5631 );
not \mul_6_18_g43308/U$4 ( \5633 , \2274 );
or \mul_6_18_g43308/U$2 ( \5634 , \5632 , \5633 );
not \mul_6_18_g44074/U$3 ( \5635 , \2168 );
not \mul_6_18_g44074/U$4 ( \5636 , \2277 );
or \mul_6_18_g44074/U$2 ( \5637 , \5635 , \5636 );
nand \mul_6_18_g44368/U$1 ( \5638 , \2256 , \3154 );
nand \mul_6_18_g44074/U$1 ( \5639 , \5637 , \5638 );
nand \mul_6_18_g43629/U$1 ( \5640 , \3232 , \5639 );
nand \mul_6_18_g43308/U$1 ( \5641 , \5634 , \5640 );
and \mul_6_18_g42563/U$3 ( \5642 , \5626 , \5641 );
and \mul_6_18_g42563/U$5 ( \5643 , \5615 , \5625 );
or \mul_6_18_g42563/U$2 ( \5644 , \5642 , \5643 );
and \mul_6_18_g42436/U$2 ( \5645 , \5600 , \5644 );
nor \mul_6_18_g42505/U$1 ( \5646 , \5580 , \5599 );
nor \mul_6_18_g42436/U$1 ( \5647 , \5645 , \5646 );
not \mul_6_18_g42306/U$3 ( \5648 , \5647 );
xor \mul_6_18_g42559/U$1 ( \5649 , \5425 , \5436 );
xor \mul_6_18_g42559/U$1_r1 ( \5650 , \5649 , \5447 );
not \mul_6_18_g42306/U$4 ( \5651 , \5650 );
and \mul_6_18_g42306/U$2 ( \5652 , \5648 , \5651 );
and \mul_6_18_g42306/U$5 ( \5653 , \5647 , \5650 );
nor \mul_6_18_g42306/U$1 ( \5654 , \5652 , \5653 );
not \mul_6_18_g42214/U$3 ( \5655 , \5654 );
not \mul_6_18_g42680/U$3 ( \5656 , \5557 );
not \mul_6_18_g42948/U$1 ( \5657 , \5568 );
not \mul_6_18_g42680/U$4 ( \5658 , \5657 );
or \mul_6_18_g42680/U$2 ( \5659 , \5656 , \5658 );
nand \mul_6_18_g42680/U$1 ( \5660 , \5659 , \5579 );
or \mul_6_18_g45205/U$1 ( \5661 , \5657 , \5557 );
nand \mul_6_18_g42594/U$1 ( \5662 , \5660 , \5661 );
not \mul_6_18_g43370/U$3 ( \5663 , \5613 );
not \mul_6_18_g43370/U$4 ( \5664 , \2222 );
or \mul_6_18_g43370/U$2 ( \5665 , \5663 , \5664 );
nand \mul_6_18_g43612/U$1 ( \5666 , \5420 , \2934 );
nand \mul_6_18_g43370/U$1 ( \5667 , \5665 , \5666 );
not \mul_6_18_g42689/U$3 ( \5668 , \5667 );
not \mul_6_18_g43309/U$3 ( \5669 , \5639 );
not \mul_6_18_g43309/U$4 ( \5670 , \2274 );
or \mul_6_18_g43309/U$2 ( \5671 , \5669 , \5670 );
nand \mul_6_18_g43483/U$1 ( \5672 , \3449 , \5442 );
nand \mul_6_18_g43309/U$1 ( \5673 , \5671 , \5672 );
not \mul_6_18_g42689/U$4 ( \5674 , \5673 );
or \mul_6_18_g42689/U$2 ( \5675 , \5668 , \5674 );
or \mul_6_18_g42751/U$2 ( \5676 , \5673 , \5667 );
not \mul_6_18_g44099/U$3 ( \5677 , \2056 );
not \mul_6_18_g44099/U$4 ( \5678 , \2718 );
or \mul_6_18_g44099/U$2 ( \5679 , \5677 , \5678 );
nand \mul_6_18_g44379/U$1 ( \5680 , \2714 , \3360 );
nand \mul_6_18_g44099/U$1 ( \5681 , \5679 , \5680 );
not \mul_6_18_g43270/U$3 ( \5682 , \5681 );
not \mul_6_18_g43270/U$4 ( \5683 , \2729 );
or \mul_6_18_g43270/U$2 ( \5684 , \5682 , \5683 );
nand \mul_6_18_g43622/U$1 ( \5685 , \2733 , \5522 );
nand \mul_6_18_g43270/U$1 ( \5686 , \5684 , \5685 );
nand \mul_6_18_g42751/U$1 ( \5687 , \5676 , \5686 );
nand \mul_6_18_g42689/U$1 ( \5688 , \5675 , \5687 );
xor \mul_6_18_g42333/U$1 ( \5689 , \5662 , \5688 );
xor \mul_6_18_g42480/U$1 ( \5690 , \5527 , \5537 );
xor \mul_6_18_g42480/U$1_r1 ( \5691 , \5690 , \5542 );
xor \mul_6_18_g42333/U$1_r1 ( \5692 , \5689 , \5691 );
not \mul_6_18_g42214/U$4 ( \5693 , \5692 );
and \mul_6_18_g42214/U$2 ( \5694 , \5655 , \5693 );
and \mul_6_18_g42214/U$5 ( \5695 , \5692 , \5654 );
nor \mul_6_18_g42214/U$1 ( \5696 , \5694 , \5695 );
xor \mul_6_18_g42737/U$1 ( \5697 , \5667 , \5673 );
xnor \mul_6_18_g42737/U$1_r1 ( \5698 , \5697 , \5686 );
not \mul_6_18_g42644/U$1 ( \5699 , \5698 );
not \mul_6_18_g42242/U$3 ( \5700 , \5699 );
and \mul_6_18_g44134/U$2 ( \5701 , \2058 , \2972 );
not \mul_6_18_g44134/U$4 ( \5702 , \2058 );
and \mul_6_18_g44134/U$3 ( \5703 , \5702 , \2718 );
nor \mul_6_18_g44134/U$1 ( \5704 , \5701 , \5703 );
not \mul_6_18_g43273/U$3 ( \5705 , \5704 );
not \mul_6_18_g43273/U$4 ( \5706 , \2965 );
or \mul_6_18_g43273/U$2 ( \5707 , \5705 , \5706 );
nand \mul_6_18_g43631/U$1 ( \5708 , \3326 , \5681 );
nand \mul_6_18_g43273/U$1 ( \5709 , \5707 , \5708 );
not \mul_6_18_g42465/U$3 ( \5710 , \5709 );
not \mul_6_18_g42818/U$3 ( \5711 , \5598 );
not \mul_6_18_g42945/U$1 ( \5712 , \5590 );
not \mul_6_18_g42818/U$4 ( \5713 , \5712 );
or \mul_6_18_g42818/U$2 ( \5714 , \5711 , \5713 );
and \mul_6_18_g43670/U$2 ( \5715 , \2252 , \5592 );
nor \mul_6_18_g43670/U$1 ( \5716 , \5715 , \5597 );
not \mul_6_18_g42833/U$2 ( \5717 , \5716 );
nand \mul_6_18_g42833/U$1 ( \5718 , \5717 , \5590 );
nand \mul_6_18_g42818/U$1 ( \5719 , \5714 , \5718 );
not \mul_6_18_g42465/U$4 ( \5720 , \5719 );
or \mul_6_18_g42465/U$2 ( \5721 , \5710 , \5720 );
or \g45688/U$1 ( \5722 , \5719 , \5709 );
nand \mul_6_18_g43663/U$1 ( \5723 , \4327 , \2058 );
not \mul_6_18_g42681/U$3 ( \5724 , \5723 );
not \mul_6_18_g44033/U$3 ( \5725 , \2006 );
not \mul_6_18_g44033/U$4 ( \5726 , \2423 );
or \mul_6_18_g44033/U$2 ( \5727 , \5725 , \5726 );
nand \mul_6_18_g44350/U$1 ( \5728 , \2848 , \2795 );
nand \mul_6_18_g44033/U$1 ( \5729 , \5727 , \5728 );
not \mul_6_18_g42951/U$3 ( \5730 , \5729 );
not \mul_6_18_g42951/U$4 ( \5731 , \4014 );
or \mul_6_18_g42951/U$2 ( \5732 , \5730 , \5731 );
nand \mul_6_18_g43042/U$1 ( \5733 , \2434 , \5585 );
nand \mul_6_18_g42951/U$1 ( \5734 , \5732 , \5733 );
not \mul_6_18_g42950/U$1 ( \5735 , \5734 );
not \mul_6_18_g42681/U$4 ( \5736 , \5735 );
or \mul_6_18_g42681/U$2 ( \5737 , \5724 , \5736 );
not \mul_6_18_g44063/U$3 ( \5738 , \2168 );
not \mul_6_18_g44063/U$4 ( \5739 , \3186 );
or \mul_6_18_g44063/U$2 ( \5740 , \5738 , \5739 );
nand \mul_6_18_g44377/U$1 ( \5741 , \2626 , \3154 );
nand \mul_6_18_g44063/U$1 ( \5742 , \5740 , \5741 );
not \mul_6_18_g42981/U$3 ( \5743 , \5742 );
not \mul_6_18_g42981/U$4 ( \5744 , \2907 );
or \mul_6_18_g42981/U$2 ( \5745 , \5743 , \5744 );
nand \mul_6_18_g43043/U$1 ( \5746 , \2842 , \5620 );
nand \mul_6_18_g42981/U$1 ( \5747 , \5745 , \5746 );
nand \mul_6_18_g42681/U$1 ( \5748 , \5737 , \5747 );
not \mul_6_18_g42835/U$2 ( \5749 , \5723 );
nand \mul_6_18_g42835/U$1 ( \5750 , \5749 , \5734 );
nand \mul_6_18_g42593/U$1 ( \5751 , \5748 , \5750 );
nand \mul_6_18_g42516/U$1 ( \5752 , \5722 , \5751 );
nand \mul_6_18_g42465/U$1 ( \5753 , \5721 , \5752 );
not \mul_6_18_g42242/U$4 ( \5754 , \5753 );
or \mul_6_18_g42242/U$2 ( \5755 , \5700 , \5754 );
xor \mul_6_18_g42401/U$1 ( \5756 , \5599 , \5644 );
not \mul_6_18_g42564/U$1 ( \5757 , \5580 );
xnor \mul_6_18_g42401/U$1_r1 ( \5758 , \5756 , \5757 );
not \mul_6_18_g42388/U$2 ( \5759 , \5753 );
nand \mul_6_18_g42388/U$1 ( \5760 , \5759 , \5698 );
nand \mul_6_18_g42289/U$1 ( \5761 , \5758 , \5760 );
nand \mul_6_18_g42242/U$1 ( \5762 , \5755 , \5761 );
not \mul_6_18_g42234/U$1 ( \5763 , \5762 );
nand \mul_6_18_g42148/U$1 ( \5764 , \5696 , \5763 );
not \mul_6_18_g42382/U$3 ( \5765 , \5698 );
not \mul_6_18_g42382/U$4 ( \5766 , \5753 );
or \mul_6_18_g42382/U$2 ( \5767 , \5765 , \5766 );
or \mul_6_18_g42382/U$5 ( \5768 , \5753 , \5698 );
nand \mul_6_18_g42382/U$1 ( \5769 , \5767 , \5768 );
not \mul_6_18_g42361/U$1 ( \5770 , \5758 );
and \mul_6_18_g42270/U$2 ( \5771 , \5769 , \5770 );
not \mul_6_18_g42270/U$4 ( \5772 , \5769 );
and \mul_6_18_g42270/U$3 ( \5773 , \5772 , \5758 );
nor \mul_6_18_g42270/U$1 ( \5774 , \5771 , \5773 );
and \g45690/U$2 ( \5775 , \5605 , \2934 );
and \g45763/U$2 ( \5776 , \3422 , \1998 );
not \g45763/U$4 ( \5777 , \3422 );
and \g45763/U$3 ( \5778 , \5777 , \2489 );
or \g45763/U$1 ( \5779 , \5776 , \5778 );
and \g45690/U$3 ( \5780 , \2223 , \5779 );
nor \g45690/U$1 ( \5781 , \5775 , \5780 );
not \mul_6_18_g43386/U$1 ( \5782 , \5781 );
not \mul_6_18_g42601/U$3 ( \5783 , \5782 );
not \mul_6_18_g44088/U$3 ( \5784 , \2056 );
not \mul_6_18_g44088/U$4 ( \5785 , \2277 );
or \mul_6_18_g44088/U$2 ( \5786 , \5784 , \5785 );
nand \mul_6_18_g44381/U$1 ( \5787 , \2256 , \3360 );
nand \mul_6_18_g44088/U$1 ( \5788 , \5786 , \5787 );
not \mul_6_18_g43310/U$3 ( \5789 , \5788 );
not \mul_6_18_g43310/U$4 ( \5790 , \2274 );
or \mul_6_18_g43310/U$2 ( \5791 , \5789 , \5790 );
nand \mul_6_18_g43557/U$1 ( \5792 , \5631 , \3449 );
nand \mul_6_18_g43310/U$1 ( \5793 , \5791 , \5792 );
not \mul_6_18_g42601/U$4 ( \5794 , \5793 );
or \mul_6_18_g42601/U$2 ( \5795 , \5783 , \5794 );
not \mul_6_18_g44032/U$3 ( \5796 , \2179 );
not \mul_6_18_g44032/U$4 ( \5797 , \5141 );
or \mul_6_18_g44032/U$2 ( \5798 , \5796 , \5797 );
nand \mul_6_18_g44355/U$1 ( \5799 , \5561 , \2185 );
nand \mul_6_18_g44032/U$1 ( \5800 , \5798 , \5799 );
and \mul_6_18_g45222/U$2 ( \5801 , \4014 , \5800 );
and \mul_6_18_g45222/U$3 ( \5802 , \2434 , \5729 );
nor \mul_6_18_g45222/U$1 ( \5803 , \5801 , \5802 );
not \mul_6_18_g42952/U$1 ( \5804 , \5803 );
not \mul_6_18_g43725/U$3 ( \5805 , \2116 );
not \fopt45606/U$1 ( \5806 , \2263 );
not \mul_6_18_g43725/U$4 ( \5807 , \5806 );
or \mul_6_18_g43725/U$2 ( \5808 , \5805 , \5807 );
nand \mul_6_18_g43725/U$1 ( \5809 , \5808 , \2606 );
nand \mul_6_18_g44172/U$1 ( \5810 , \2263 , \2058 );
nand \mul_6_18_g43668/U$1 ( \5811 , \5809 , \2252 , \5810 );
not \mul_6_18_g43667/U$1 ( \5812 , \5811 );
nand \mul_6_18_g42846/U$1 ( \5813 , \5804 , \5812 );
not \mul_6_18_g45199/U$2 ( \5814 , \5813 );
not \mul_6_18_g42903/U$2 ( \5815 , \5793 );
nand \mul_6_18_g42903/U$1 ( \5816 , \5815 , \5781 );
nand \mul_6_18_g45199/U$1 ( \5817 , \5814 , \5816 );
nand \mul_6_18_g42601/U$1 ( \5818 , \5795 , \5817 );
not \g45787/U$3 ( \5819 , \5818 );
xor \mul_6_18_g42563/U$1 ( \5820 , \5615 , \5625 );
xor \mul_6_18_g42563/U$1_r1 ( \5821 , \5820 , \5641 );
not \g45787/U$4 ( \5822 , \5821 );
and \g45787/U$2 ( \5823 , \5819 , \5822 );
xor \mul_6_18_g42491/U$1 ( \5824 , \5709 , \5719 );
xnor \mul_6_18_g42491/U$1_r1 ( \5825 , \5824 , \5751 );
nor \g45787/U$1 ( \5826 , \5823 , \5825 );
and \mul_6_18_g42447/U$2 ( \5827 , \5821 , \5818 );
nor \g45786/U$1 ( \5828 , \5826 , \5827 );
nand \mul_6_18_g42186/U$1 ( \5829 , \5774 , \5828 );
and \mul_6_18_g42123/U$1 ( \5830 , \5764 , \5829 );
not \mul_6_18_g42021/U$3 ( \5831 , \5830 );
not \mul_6_18_g43381/U$3 ( \5832 , \2223 );
not \mul_6_18_g44020/U$3 ( \5833 , \2006 );
not \mul_6_18_g44020/U$4 ( \5834 , \5416 );
or \mul_6_18_g44020/U$2 ( \5835 , \5833 , \5834 );
nand \mul_6_18_g44345/U$1 ( \5836 , \2226 , \2795 );
nand \mul_6_18_g44020/U$1 ( \5837 , \5835 , \5836 );
not \mul_6_18_g43381/U$4 ( \5838 , \5837 );
or \mul_6_18_g43381/U$2 ( \5839 , \5832 , \5838 );
not \mul_6_18_g44002/U$3 ( \5840 , \2463 );
not \mul_6_18_g44002/U$4 ( \5841 , \3422 );
or \mul_6_18_g44002/U$2 ( \5842 , \5840 , \5841 );
nand \mul_6_18_g44322/U$1 ( \5843 , \2216 , \2468 );
nand \mul_6_18_g44002/U$1 ( \5844 , \5842 , \5843 );
nand \mul_6_18_g43525/U$1 ( \5845 , \5844 , \2934 );
nand \mul_6_18_g43381/U$1 ( \5846 , \5839 , \5845 );
not \mul_6_18_g42672/U$2 ( \5847 , \5846 );
not \mul_6_18_g44055/U$3 ( \5848 , \2144 );
not \mul_6_18_g44055/U$4 ( \5849 , \4008 );
or \mul_6_18_g44055/U$2 ( \5850 , \5848 , \5849 );
nand \mul_6_18_g44369/U$1 ( \5851 , \2418 , \2145 );
nand \mul_6_18_g44055/U$1 ( \5852 , \5850 , \5851 );
not \mul_6_18_g42928/U$3 ( \5853 , \5852 );
not \mul_6_18_g42928/U$4 ( \5854 , \4014 );
or \mul_6_18_g42928/U$2 ( \5855 , \5853 , \5854 );
not \mul_6_18_g44054/U$3 ( \5856 , \2168 );
not \mul_6_18_g44054/U$4 ( \5857 , \2423 );
or \mul_6_18_g44054/U$2 ( \5858 , \5856 , \5857 );
nand \mul_6_18_g44375/U$1 ( \5859 , \5561 , \3154 );
nand \mul_6_18_g44054/U$1 ( \5860 , \5858 , \5859 );
nand \mul_6_18_g43049/U$1 ( \5861 , \2434 , \5860 );
nand \mul_6_18_g42928/U$1 ( \5862 , \5855 , \5861 );
not \mul_6_18_g43732/U$3 ( \5863 , \2116 );
not \mul_6_18_g43732/U$4 ( \5864 , \1506 );
or \mul_6_18_g43732/U$2 ( \5865 , \5863 , \5864 );
nand \mul_6_18_g43732/U$1 ( \5866 , \5865 , \2848 );
nand \mul_6_18_g44189/U$1 ( \5867 , \1507 , \2058 );
and \mul_6_18_g43686/U$1 ( \5868 , \5866 , \2626 , \5867 );
nand \mul_6_18_g42847/U$1 ( \5869 , \5862 , \5868 );
nand \mul_6_18_g42672/U$1 ( \5870 , \5847 , \5869 );
not \mul_6_18_g42463/U$3 ( \5871 , \5870 );
not \mul_6_18_g43666/U$2 ( \5872 , \2284 );
nand \mul_6_18_g43666/U$1 ( \5873 , \5872 , \2058 );
not \mul_6_18_g42957/U$3 ( \5874 , \5860 );
not \mul_6_18_g42957/U$4 ( \5875 , \2586 );
or \mul_6_18_g42957/U$2 ( \5876 , \5874 , \5875 );
nand \mul_6_18_g43038/U$1 ( \5877 , \2434 , \5800 );
nand \mul_6_18_g42957/U$1 ( \5878 , \5876 , \5877 );
xor \mul_6_18_g42700/U$1 ( \5879 , \5873 , \5878 );
not \mul_6_18_g44080/U$3 ( \5880 , \2056 );
not \mul_6_18_g44080/U$4 ( \5881 , \2909 );
or \mul_6_18_g44080/U$2 ( \5882 , \5880 , \5881 );
nand \mul_6_18_g44385/U$1 ( \5883 , \2606 , \3360 );
nand \mul_6_18_g44080/U$1 ( \5884 , \5882 , \5883 );
not \mul_6_18_g42995/U$3 ( \5885 , \5884 );
not \mul_6_18_g42995/U$4 ( \5886 , \2907 );
or \mul_6_18_g42995/U$2 ( \5887 , \5885 , \5886 );
not \mul_6_18_g44062/U$3 ( \5888 , \2144 );
not \mul_6_18_g44062/U$4 ( \5889 , \2629 );
or \mul_6_18_g44062/U$2 ( \5890 , \5888 , \5889 );
nand \mul_6_18_g44378/U$1 ( \5891 , \2626 , \2145 );
nand \mul_6_18_g44062/U$1 ( \5892 , \5890 , \5891 );
nand \mul_6_18_g43047/U$1 ( \5893 , \2623 , \5892 );
nand \mul_6_18_g42995/U$1 ( \5894 , \5887 , \5893 );
xnor \mul_6_18_g42700/U$1_r1 ( \5895 , \5879 , \5894 );
not \mul_6_18_g42463/U$4 ( \5896 , \5895 );
or \mul_6_18_g42463/U$2 ( \5897 , \5871 , \5896 );
not \mul_6_18_g45198/U$2 ( \5898 , \5869 );
nand \mul_6_18_g45198/U$1 ( \5899 , \5898 , \5846 );
nand \mul_6_18_g42463/U$1 ( \5900 , \5897 , \5899 );
not \mul_6_18_g42819/U$3 ( \5901 , \5812 );
not \mul_6_18_g42819/U$4 ( \5902 , \5803 );
or \mul_6_18_g42819/U$2 ( \5903 , \5901 , \5902 );
nand \mul_6_18_g42834/U$1 ( \5904 , \5804 , \5811 );
nand \mul_6_18_g42819/U$1 ( \5905 , \5903 , \5904 );
not \mul_6_18_g42524/U$3 ( \5906 , \5905 );
not \mul_6_18_g42831/U$2 ( \5907 , \5894 );
nand \mul_6_18_g42831/U$1 ( \5908 , \5907 , \5873 );
and \mul_6_18_g45143/U$2 ( \5909 , \5908 , \5878 );
not \mul_6_18_g45146/U$2 ( \5910 , \5894 );
nor \mul_6_18_g45146/U$1 ( \5911 , \5910 , \5873 );
nor \mul_6_18_g45143/U$1 ( \5912 , \5909 , \5911 );
not \mul_6_18_g42524/U$4 ( \5913 , \5912 );
or \mul_6_18_g42524/U$2 ( \5914 , \5906 , \5913 );
or \mul_6_18_g42524/U$5 ( \5915 , \5912 , \5905 );
nand \mul_6_18_g42524/U$1 ( \5916 , \5914 , \5915 );
not \mul_6_18_g42441/U$3 ( \5917 , \5916 );
and \mul_6_18_g43383/U$2 ( \5918 , \2222 , \5844 );
and \mul_6_18_g43383/U$3 ( \5919 , \5779 , \2245 );
nor \mul_6_18_g43383/U$1 ( \5920 , \5918 , \5919 );
not \mul_6_18_g42994/U$3 ( \5921 , \5892 );
not \mul_6_18_g42994/U$4 ( \5922 , \3013 );
or \mul_6_18_g42994/U$2 ( \5923 , \5921 , \5922 );
nand \mul_6_18_g43046/U$1 ( \5924 , \2623 , \5742 );
nand \mul_6_18_g42994/U$1 ( \5925 , \5923 , \5924 );
not \mul_6_18_g42993/U$1 ( \5926 , \5925 );
xor \mul_6_18_g42566/U$1 ( \5927 , \5920 , \5926 );
not \mul_6_18_g44145/U$3 ( \5928 , \2058 );
not \mul_6_18_g44948/U$1 ( \5929 , \2280 );
not \mul_6_18_g44145/U$4 ( \5930 , \5929 );
or \mul_6_18_g44145/U$2 ( \5931 , \5928 , \5930 );
nand \mul_6_18_g44397/U$1 ( \5932 , \2256 , \2116 );
nand \mul_6_18_g44145/U$1 ( \5933 , \5931 , \5932 );
and \mul_6_18_g43311/U$2 ( \5934 , \2274 , \5933 );
and \mul_6_18_g43311/U$3 ( \5935 , \3232 , \5788 );
nor \mul_6_18_g43311/U$1 ( \5936 , \5934 , \5935 );
xor \mul_6_18_g42566/U$1_r1 ( \5937 , \5927 , \5936 );
not \mul_6_18_g42441/U$4 ( \5938 , \5937 );
or \mul_6_18_g42441/U$2 ( \5939 , \5917 , \5938 );
or \mul_6_18_g42441/U$5 ( \5940 , \5916 , \5937 );
nand \mul_6_18_g42441/U$1 ( \5941 , \5939 , \5940 );
xor \mul_6_18_g42107/U$4 ( \5942 , \5900 , \5941 );
not \mul_6_18_g42920/U$3 ( \5943 , \4265 );
and \mul_6_18_g44153/U$2 ( \5944 , \2116 , \2418 );
not \mul_6_18_g44153/U$4 ( \5945 , \2116 );
and \mul_6_18_g44153/U$3 ( \5946 , \5945 , \4008 );
nor \mul_6_18_g44153/U$1 ( \5947 , \5944 , \5946 );
not \mul_6_18_g42920/U$4 ( \5948 , \5947 );
and \mul_6_18_g42920/U$2 ( \5949 , \5943 , \5948 );
not \mul_6_18_g44070/U$3 ( \5950 , \2056 );
not \mul_6_18_g44070/U$4 ( \5951 , \2423 );
or \mul_6_18_g44070/U$2 ( \5952 , \5950 , \5951 );
nand \mul_6_18_g44384/U$1 ( \5953 , \2418 , \3360 );
nand \mul_6_18_g44070/U$1 ( \5954 , \5952 , \5953 );
and \mul_6_18_g42920/U$5 ( \5955 , \5954 , \2434 );
nor \mul_6_18_g42920/U$1 ( \5956 , \5949 , \5955 );
not \mul_6_18_g42821/U$3 ( \5957 , \5956 );
not \mul_6_18_g43733/U$3 ( \5958 , \2116 );
not \mul_6_18_g43733/U$4 ( \5959 , \2429 );
or \mul_6_18_g43733/U$2 ( \5960 , \5958 , \5959 );
nand \mul_6_18_g43733/U$1 ( \5961 , \5960 , \2236 );
nand \mul_6_18_g44190/U$1 ( \5962 , \1518 , \2058 );
and \mul_6_18_g43684/U$1 ( \5963 , \5961 , \2848 , \5962 );
not \mul_6_18_g42821/U$4 ( \5964 , \5963 );
and \mul_6_18_g42821/U$2 ( \5965 , \5957 , \5964 );
and \mul_6_18_g42821/U$5 ( \5966 , \5956 , \5963 );
nor \mul_6_18_g42821/U$1 ( \5967 , \5965 , \5966 );
not \mul_6_18_g44051/U$3 ( \5968 , \2168 );
not \mul_6_18_g44051/U$4 ( \5969 , \2929 );
or \mul_6_18_g44051/U$2 ( \5970 , \5968 , \5969 );
nand \mul_6_18_g44367/U$1 ( \5971 , \2236 , \3154 );
nand \mul_6_18_g44051/U$1 ( \5972 , \5970 , \5971 );
and \mul_6_18_g45240/U$2 ( \5973 , \5972 , \2934 );
not \mul_6_18_g44049/U$3 ( \5974 , \2144 );
not \mul_6_18_g44049/U$4 ( \5975 , \3422 );
or \mul_6_18_g44049/U$2 ( \5976 , \5974 , \5975 );
nand \mul_6_18_g44371/U$1 ( \5977 , \2236 , \2145 );
nand \mul_6_18_g44049/U$1 ( \5978 , \5976 , \5977 );
and \mul_6_18_g45240/U$3 ( \5979 , \2223 , \5978 );
nor \mul_6_18_g45240/U$1 ( \5980 , \5973 , \5979 );
nand \mul_6_18_g42663/U$1 ( \5981 , \5967 , \5980 );
not \g45742/U$3 ( \5982 , \5981 );
not \mul_6_18_g43391/U$3 ( \5983 , \3430 );
not \mul_6_18_g44066/U$3 ( \5984 , \2056 );
not \mul_6_18_g44066/U$4 ( \5985 , \3211 );
or \mul_6_18_g44066/U$2 ( \5986 , \5984 , \5985 );
nand \mul_6_18_g44382/U$1 ( \5987 , \2236 , \3360 );
nand \mul_6_18_g44066/U$1 ( \5988 , \5986 , \5987 );
not \mul_6_18_g43391/U$4 ( \5989 , \5988 );
or \mul_6_18_g43391/U$2 ( \5990 , \5983 , \5989 );
and \mul_6_18_g44156/U$2 ( \5991 , \2058 , \2236 );
not \mul_6_18_g44156/U$4 ( \5992 , \2058 );
and \mul_6_18_g44156/U$3 ( \5993 , \5992 , \3211 );
nor \mul_6_18_g44156/U$1 ( \5994 , \5991 , \5993 );
nand \mul_6_18_g43642/U$1 ( \5995 , \5994 , \2222 );
nand \mul_6_18_g43391/U$1 ( \5996 , \5990 , \5995 );
nand \mul_6_18_g44271/U$1 ( \5997 , \2244 , \2058 );
and \mul_6_18_g45147/U$1 ( \5998 , \5997 , \2226 );
nand \mul_6_18_g43051/U$1 ( \5999 , \5996 , \5998 );
nand \mul_6_18_g43055/U$1 ( \6000 , \2434 , \2058 );
not \mul_6_18_g42907/U$2 ( \6001 , \6000 );
buf \mul_6_18_g44873/U$1 ( \6002 , \2243 );
not \mul_6_18_g44872/U$1 ( \6003 , \6002 );
not \mul_6_18_g43376/U$3 ( \6004 , \6003 );
not \mul_6_18_g43376/U$4 ( \6005 , \5978 );
or \mul_6_18_g43376/U$2 ( \6006 , \6004 , \6005 );
nand \mul_6_18_g43482/U$1 ( \6007 , \5988 , \2222 );
nand \mul_6_18_g43376/U$1 ( \6008 , \6006 , \6007 );
nor \mul_6_18_g42907/U$1 ( \6009 , \6001 , \6008 );
or \mul_6_18_g42753/U$2 ( \6010 , \5999 , \6009 );
not \mul_6_18_g42906/U$2 ( \6011 , \6000 );
nand \mul_6_18_g42906/U$1 ( \6012 , \6011 , \6008 );
nand \mul_6_18_g42753/U$1 ( \6013 , \6010 , \6012 );
not \g45742/U$4 ( \6014 , \6013 );
or \g45742/U$2 ( \6015 , \5982 , \6014 );
not \mul_6_18_g42783/U$1 ( \6016 , \5967 );
not \mul_6_18_g43377/U$1 ( \6017 , \5980 );
nand \mul_6_18_g42669/U$1 ( \6018 , \6016 , \6017 );
nand \g45742/U$1 ( \6019 , \6015 , \6018 );
not \mul_6_18_g45232/U$2 ( \6020 , \5963 );
nor \mul_6_18_g45232/U$1 ( \6021 , \6020 , \5956 );
not \mul_6_18_g42538/U$2 ( \6022 , \6021 );
nand \mul_6_18_g43054/U$1 ( \6023 , \2622 , \2058 );
not \mul_6_18_g42959/U$3 ( \6024 , \5954 );
not \mul_6_18_g42959/U$4 ( \6025 , \4264 );
or \mul_6_18_g42959/U$2 ( \6026 , \6024 , \6025 );
nand \mul_6_18_g43045/U$1 ( \6027 , \5852 , \2434 );
nand \mul_6_18_g42959/U$1 ( \6028 , \6026 , \6027 );
xor \mul_6_18_g42699/U$1 ( \6029 , \6023 , \6028 );
not \mul_6_18_g43390/U$3 ( \6030 , \2222 );
not \mul_6_18_g43390/U$4 ( \6031 , \5972 );
or \mul_6_18_g43390/U$2 ( \6032 , \6030 , \6031 );
not \mul_6_18_g44022/U$3 ( \6033 , \2179 );
not \mul_6_18_g44022/U$4 ( \6034 , \3422 );
or \mul_6_18_g44022/U$2 ( \6035 , \6033 , \6034 );
nand \mul_6_18_g44346/U$1 ( \6036 , \3215 , \2185 );
nand \mul_6_18_g44022/U$1 ( \6037 , \6035 , \6036 );
nand \mul_6_18_g43640/U$1 ( \6038 , \6037 , \6003 );
nand \mul_6_18_g43390/U$1 ( \6039 , \6032 , \6038 );
not \mul_6_18_g43389/U$1 ( \6040 , \6039 );
xnor \mul_6_18_g42699/U$1_r1 ( \6041 , \6029 , \6040 );
nand \mul_6_18_g42538/U$1 ( \6042 , \6022 , \6041 );
nand \mul_6_18_g42432/U$1 ( \6043 , \6019 , \6042 );
not \mul_6_18_g45192/U$2 ( \6044 , \6041 );
nand \mul_6_18_g45192/U$1 ( \6045 , \6044 , \6021 );
nand \mul_6_18_g42396/U$1 ( \6046 , \6043 , \6045 );
not \mul_6_18_g42859/U$3 ( \6047 , \6023 );
not \mul_6_18_g42859/U$4 ( \6048 , \6040 );
or \mul_6_18_g42859/U$2 ( \6049 , \6047 , \6048 );
nand \mul_6_18_g42859/U$1 ( \6050 , \6049 , \6028 );
not \mul_6_18_g45209/U$2 ( \6051 , \6023 );
nand \mul_6_18_g45209/U$1 ( \6052 , \6051 , \6039 );
nand \mul_6_18_g42799/U$1 ( \6053 , \6050 , \6052 );
not \mul_6_18_g42508/U$2 ( \6054 , \6053 );
not \mul_6_18_g44392/U$1 ( \6055 , \2222 );
not \mul_6_18_g43385/U$3 ( \6056 , \6055 );
not \mul_6_18_g44021/U$1 ( \6057 , \6037 );
not \mul_6_18_g43385/U$4 ( \6058 , \6057 );
and \mul_6_18_g43385/U$2 ( \6059 , \6056 , \6058 );
and \mul_6_18_g43385/U$5 ( \6060 , \5837 , \2934 );
nor \mul_6_18_g43385/U$1 ( \6061 , \6059 , \6060 );
not \mul_6_18_g42997/U$3 ( \6062 , \2602 );
and \mul_6_18_g44149/U$2 ( \6063 , \2116 , \2606 );
not \mul_6_18_g44149/U$4 ( \6064 , \2116 );
and \mul_6_18_g44149/U$3 ( \6065 , \6064 , \2834 );
nor \mul_6_18_g44149/U$1 ( \6066 , \6063 , \6065 );
not \mul_6_18_g42997/U$4 ( \6067 , \6066 );
and \mul_6_18_g42997/U$2 ( \6068 , \6062 , \6067 );
and \mul_6_18_g42997/U$5 ( \6069 , \2842 , \5884 );
nor \mul_6_18_g42997/U$1 ( \6070 , \6068 , \6069 );
xor \mul_6_18_g42767/U$1 ( \6071 , \6061 , \6070 );
not \mul_6_18_g42658/U$3 ( \6072 , \6071 );
not \mul_6_18_g42927/U$1 ( \6073 , \5862 );
not \mul_6_18_g42820/U$3 ( \6074 , \6073 );
not \mul_6_18_g42820/U$4 ( \6075 , \5868 );
and \mul_6_18_g42820/U$2 ( \6076 , \6074 , \6075 );
and \mul_6_18_g42820/U$5 ( \6077 , \6073 , \5868 );
nor \mul_6_18_g42820/U$1 ( \6078 , \6076 , \6077 );
not \mul_6_18_g42658/U$4 ( \6079 , \6078 );
and \mul_6_18_g42658/U$2 ( \6080 , \6072 , \6079 );
and \mul_6_18_g42658/U$5 ( \6081 , \6078 , \6071 );
nor \mul_6_18_g42658/U$1 ( \6082 , \6080 , \6081 );
nand \mul_6_18_g42508/U$1 ( \6083 , \6054 , \6082 );
nand \mul_6_18_g42318/U$1 ( \6084 , \6046 , \6083 );
not \mul_6_18_g45188/U$2 ( \6085 , \6082 );
nand \mul_6_18_g45188/U$1 ( \6086 , \6085 , \6053 );
nand \mul_6_18_g42291/U$1 ( \6087 , \6084 , \6086 );
buf \mul_6_18_g42764/U$1 ( \6088 , \6078 );
and \mul_6_18_g42767/U$2 ( \6089 , \6061 , \6070 );
or \mul_6_18_g42603/U$2 ( \6090 , \6088 , \6089 );
or \mul_6_18_g45208/U$1 ( \6091 , \6070 , \6061 );
nand \mul_6_18_g42603/U$1 ( \6092 , \6090 , \6091 );
not \mul_6_18_g42390/U$2 ( \6093 , \6092 );
not \mul_6_18_g42467/U$3 ( \6094 , \5895 );
not \mul_6_18_g42613/U$3 ( \6095 , \5869 );
not \mul_6_18_g42613/U$4 ( \6096 , \5846 );
and \mul_6_18_g42613/U$2 ( \6097 , \6095 , \6096 );
and \mul_6_18_g42613/U$5 ( \6098 , \5869 , \5846 );
nor \mul_6_18_g42613/U$1 ( \6099 , \6097 , \6098 );
not \mul_6_18_g42467/U$4 ( \6100 , \6099 );
and \mul_6_18_g42467/U$2 ( \6101 , \6094 , \6100 );
and \mul_6_18_g42467/U$5 ( \6102 , \5895 , \6099 );
nor \mul_6_18_g42467/U$1 ( \6103 , \6101 , \6102 );
nand \mul_6_18_g42390/U$1 ( \6104 , \6093 , \6103 );
nand \mul_6_18_g42218/U$1 ( \6105 , \6087 , \6104 );
not \mul_6_18_g45180/U$2 ( \6106 , \6103 );
nand \mul_6_18_g45180/U$1 ( \6107 , \6106 , \6092 );
nand \mul_6_18_g42190/U$1 ( \6108 , \6105 , \6107 );
and \mul_6_18_g42107/U$3 ( \6109 , \5942 , \6108 );
and \mul_6_18_g42107/U$5 ( \6110 , \5900 , \5941 );
or \mul_6_18_g42107/U$2 ( \6111 , \6109 , \6110 );
not \mul_6_18_g42387/U$3 ( \6112 , \5825 );
xor \mul_6_18_g42447/U$1 ( \6113 , \5821 , \5818 );
not \mul_6_18_g42387/U$4 ( \6114 , \6113 );
and \mul_6_18_g42387/U$2 ( \6115 , \6112 , \6114 );
and \mul_6_18_g42387/U$5 ( \6116 , \5825 , \6113 );
nor \mul_6_18_g42387/U$1 ( \6117 , \6115 , \6116 );
xor \mul_6_18_g42566/U$4 ( \6118 , \5920 , \5926 );
and \mul_6_18_g42566/U$3 ( \6119 , \6118 , \5936 );
and \mul_6_18_g42566/U$5 ( \6120 , \5920 , \5926 );
or \mul_6_18_g42566/U$2 ( \6121 , \6119 , \6120 );
xor \mul_6_18_g42614/U$1 ( \6122 , \5723 , \5735 );
xnor \mul_6_18_g42614/U$1_r1 ( \6123 , \6122 , \5747 );
xor \mul_6_18_g42364/U$4 ( \6124 , \6121 , \6123 );
xor \mul_6_18_g42618/U$1 ( \6125 , \5781 , \5793 );
xnor \mul_6_18_g42618/U$1_r1 ( \6126 , \6125 , \5813 );
and \mul_6_18_g42364/U$3 ( \6127 , \6124 , \6126 );
and \mul_6_18_g42364/U$5 ( \6128 , \6121 , \6123 );
or \mul_6_18_g42364/U$2 ( \6129 , \6127 , \6128 );
nand \mul_6_18_g42281/U$1 ( \6130 , \6117 , \6129 );
xor \mul_6_18_g42364/U$1 ( \6131 , \6121 , \6123 );
xor \mul_6_18_g42364/U$1_r1 ( \6132 , \6131 , \6126 );
not \mul_6_18_g45187/U$2 ( \6133 , \5937 );
nand \mul_6_18_g45187/U$1 ( \6134 , \6133 , \5905 );
not \mul_6_18_g42769/U$1 ( \6135 , \5905 );
not \mul_6_18_g42459/U$3 ( \6136 , \6135 );
not \mul_6_18_g42459/U$4 ( \6137 , \5937 );
or \mul_6_18_g42459/U$2 ( \6138 , \6136 , \6137 );
not \mul_6_18_g42645/U$1 ( \6139 , \5912 );
nand \mul_6_18_g42459/U$1 ( \6140 , \6138 , \6139 );
and \mul_6_18_g42437/U$1 ( \6141 , \6134 , \6140 );
nand \mul_6_18_g42311/U$1 ( \6142 , \6132 , \6141 );
nand \mul_6_18_g42077/U$1 ( \6143 , \6111 , \6130 , \6142 );
nor \mul_6_18_g42317/U$1 ( \6144 , \6141 , \6132 );
and \mul_6_18_g42223/U$2 ( \6145 , \6130 , \6144 );
nor \mul_6_18_g42280/U$1 ( \6146 , \6117 , \6129 );
nor \mul_6_18_g42223/U$1 ( \6147 , \6145 , \6146 );
nand \mul_6_18_g42062/U$1 ( \6148 , \6143 , \6147 );
not \mul_6_18_g42021/U$4 ( \6149 , \6148 );
or \mul_6_18_g42021/U$2 ( \6150 , \5831 , \6149 );
nor \mul_6_18_g42184/U$1 ( \6151 , \5774 , \5828 );
and \mul_6_18_g42097/U$2 ( \6152 , \5764 , \6151 );
nor \mul_6_18_g42146/U$1 ( \6153 , \5696 , \5763 );
nor \mul_6_18_g42097/U$1 ( \6154 , \6152 , \6153 );
nand \mul_6_18_g42021/U$1 ( \6155 , \6150 , \6154 );
not \mul_6_18_g42213/U$3 ( \6156 , \5507 );
not \mul_6_18_g42328/U$1 ( \6157 , \5509 );
not \mul_6_18_g42266/U$3 ( \6158 , \6157 );
not \mul_6_18_g42330/U$1 ( \6159 , \5550 );
not \mul_6_18_g42266/U$4 ( \6160 , \6159 );
or \mul_6_18_g42266/U$2 ( \6161 , \6158 , \6160 );
nand \mul_6_18_g42273/U$1 ( \6162 , \5550 , \5509 );
nand \mul_6_18_g42266/U$1 ( \6163 , \6161 , \6162 );
not \mul_6_18_g42213/U$4 ( \6164 , \6163 );
or \mul_6_18_g42213/U$2 ( \6165 , \6156 , \6164 );
or \mul_6_18_g42213/U$5 ( \6166 , \6163 , \5507 );
nand \mul_6_18_g42213/U$1 ( \6167 , \6165 , \6166 );
not \mul_6_18_g42474/U$3 ( \6168 , \5450 );
not \mul_6_18_g42612/U$3 ( \6169 , \5469 );
not \mul_6_18_g42612/U$4 ( \6170 , \5479 );
and \mul_6_18_g42612/U$2 ( \6171 , \6169 , \6170 );
and \mul_6_18_g42612/U$5 ( \6172 , \5469 , \5479 );
nor \mul_6_18_g42612/U$1 ( \6173 , \6171 , \6172 );
not \mul_6_18_g42474/U$4 ( \6174 , \6173 );
or \mul_6_18_g42474/U$2 ( \6175 , \6168 , \6174 );
or \mul_6_18_g42474/U$5 ( \6176 , \6173 , \5450 );
nand \mul_6_18_g42474/U$1 ( \6177 , \6175 , \6176 );
xor \mul_6_18_g42333/U$4 ( \6178 , \5662 , \5688 );
and \mul_6_18_g42333/U$3 ( \6179 , \6178 , \5691 );
and \mul_6_18_g42333/U$5 ( \6180 , \5662 , \5688 );
or \mul_6_18_g42333/U$2 ( \6181 , \6179 , \6180 );
xor \mul_6_18_g42178/U$4 ( \6182 , \6177 , \6181 );
not \mul_6_18_g42488/U$3 ( \6183 , \5512 );
not \mul_6_18_g42488/U$4 ( \6184 , \5547 );
or \mul_6_18_g42488/U$2 ( \6185 , \6183 , \6184 );
nand \mul_6_18_g42496/U$1 ( \6186 , \5515 , \5548 );
nand \mul_6_18_g42488/U$1 ( \6187 , \6185 , \6186 );
xor \g45683/U$1 ( \6188 , \6187 , \5545 );
and \mul_6_18_g42178/U$3 ( \6189 , \6182 , \6188 );
and \mul_6_18_g42178/U$5 ( \6190 , \6177 , \6181 );
or \mul_6_18_g42178/U$2 ( \6191 , \6189 , \6190 );
nor \mul_6_18_g42145/U$1 ( \6192 , \6167 , \6191 );
xor \mul_6_18_g42178/U$1 ( \6193 , \6177 , \6181 );
xor \mul_6_18_g42178/U$1_r1 ( \6194 , \6193 , \6188 );
not \mul_6_18_g42314/U$2 ( \6195 , \5650 );
nand \mul_6_18_g42314/U$1 ( \6196 , \6195 , \5647 );
not \mul_6_18_g42191/U$3 ( \6197 , \6196 );
not \mul_6_18_g42191/U$4 ( \6198 , \5692 );
or \mul_6_18_g42191/U$2 ( \6199 , \6197 , \6198 );
not \mul_6_18_g45170/U$2 ( \6200 , \5647 );
nand \mul_6_18_g45170/U$1 ( \6201 , \6200 , \5650 );
nand \mul_6_18_g42191/U$1 ( \6202 , \6199 , \6201 );
nor \mul_6_18_g42142/U$1 ( \6203 , \6194 , \6202 );
nor \mul_6_18_g42122/U$1 ( \6204 , \6192 , \6203 );
and \mul_6_18_g42003/U$1 ( \6205 , \6155 , \6204 );
not \mul_6_18_g41969/U$4 ( \6206 , \6205 );
or \mul_6_18_g41969/U$2 ( \6207 , \5556 , \6206 );
nand \mul_6_18_g42140/U$1 ( \6208 , \6167 , \6191 );
nand \mul_6_18_g42150/U$1 ( \6209 , \6194 , \6202 );
nand \mul_6_18_g42124/U$1 ( \6210 , \6208 , \6209 );
not \mul_6_18_g42144/U$1 ( \6211 , \6192 );
and \mul_6_18_g42063/U$1 ( \6212 , \6210 , \5554 , \6211 );
not \mul_6_18_g42131/U$1 ( \6213 , \5505 );
not \mul_6_18_g42176/U$1 ( \6214 , \5553 );
nand \mul_6_18_g42093/U$1 ( \6215 , \6213 , \6214 );
nand \mul_6_18_g42059/U$1 ( \6216 , \5397 , \5494 );
nand \mul_6_18_g42040/U$1 ( \6217 , \6215 , \6216 );
or \mul_6_18_g42001/U$2 ( \6218 , \6212 , \6217 );
nand \mul_6_18_g42001/U$1 ( \6219 , \6218 , \5496 );
nand \mul_6_18_g41969/U$1 ( \6220 , \6207 , \6219 );
not \mul_6_18_g41851/U$3 ( \6221 , \6220 );
xor \mul_6_18_g42206/U$1 ( \6222 , \4846 , \4928 );
xor \mul_6_18_g42206/U$1_r1 ( \6223 , \6222 , \4931 );
xor \mul_6_18_g42728/U$1 ( \6224 , \4857 , \4868 );
xor \mul_6_18_g42728/U$1_r1 ( \6225 , \6224 , \4879 );
not \mul_6_18_g42726/U$1 ( \6226 , \6225 );
not \mul_6_18_g42514/U$3 ( \6227 , \6226 );
not \mul_6_18_g43910/U$3 ( \6228 , \2101 );
not \mul_6_18_g43910/U$4 ( \6229 , \3422 );
or \mul_6_18_g43910/U$2 ( \6230 , \6228 , \6229 );
nand \mul_6_18_g44236/U$1 ( \6231 , \2216 , \2670 );
nand \mul_6_18_g43910/U$1 ( \6232 , \6230 , \6231 );
not \mul_6_18_g43364/U$3 ( \6233 , \6232 );
not \mul_6_18_g43364/U$4 ( \6234 , \4076 );
or \mul_6_18_g43364/U$2 ( \6235 , \6233 , \6234 );
nand \mul_6_18_g43497/U$1 ( \6236 , \4852 , \2934 );
nand \mul_6_18_g43364/U$1 ( \6237 , \6235 , \6236 );
not \mul_6_18_g44012/U$3 ( \6238 , \2112 );
not \mul_6_18_g44012/U$4 ( \6239 , \2718 );
or \mul_6_18_g44012/U$2 ( \6240 , \6238 , \6239 );
nand \mul_6_18_g44299/U$1 ( \6241 , \2972 , \2824 );
nand \mul_6_18_g44012/U$1 ( \6242 , \6240 , \6241 );
not \mul_6_18_g43253/U$3 ( \6243 , \6242 );
not \mul_6_18_g43253/U$4 ( \6244 , \2965 );
or \mul_6_18_g43253/U$2 ( \6245 , \6243 , \6244 );
nand \mul_6_18_g43520/U$1 ( \6246 , \4863 , \4327 );
nand \mul_6_18_g43253/U$1 ( \6247 , \6245 , \6246 );
xor \mul_6_18_g42628/U$4 ( \6248 , \6237 , \6247 );
not \mul_6_18_g44058/U$3 ( \6249 , \1998 );
not \mul_6_18_g44058/U$4 ( \6250 , \2364 );
or \mul_6_18_g44058/U$2 ( \6251 , \6249 , \6250 );
nand \mul_6_18_g44337/U$1 ( \6252 , \5165 , \2489 );
nand \mul_6_18_g44058/U$1 ( \6253 , \6251 , \6252 );
not \mul_6_18_g43219/U$3 ( \6254 , \6253 );
not \mul_6_18_g43219/U$4 ( \6255 , \2399 );
or \mul_6_18_g43219/U$2 ( \6256 , \6254 , \6255 );
not \mul_6_18_g44023/U$3 ( \6257 , \2812 );
not \mul_6_18_g44023/U$4 ( \6258 , \2367 );
or \mul_6_18_g44023/U$2 ( \6259 , \6257 , \6258 );
nand \mul_6_18_g44306/U$1 ( \6260 , \5165 , \2811 );
nand \mul_6_18_g44023/U$1 ( \6261 , \6259 , \6260 );
nand \mul_6_18_g43506/U$1 ( \6262 , \2403 , \6261 );
nand \mul_6_18_g43219/U$1 ( \6263 , \6256 , \6262 );
and \mul_6_18_g42628/U$3 ( \6264 , \6248 , \6263 );
and \mul_6_18_g42628/U$5 ( \6265 , \6237 , \6247 );
or \mul_6_18_g42628/U$2 ( \6266 , \6264 , \6265 );
not \mul_6_18_g42626/U$1 ( \6267 , \6266 );
not \mul_6_18_g42514/U$4 ( \6268 , \6267 );
or \mul_6_18_g42514/U$2 ( \6269 , \6227 , \6268 );
xor \mul_6_18_g45217/U$1 ( \6270 , \4898 , \4888 );
xnor \mul_6_18_g45217/U$1_r1 ( \6271 , \6270 , \4909 );
not \mul_6_18_g42649/U$1 ( \6272 , \6271 );
nand \mul_6_18_g42514/U$1 ( \6273 , \6269 , \6272 );
nand \mul_6_18_g42534/U$1 ( \6274 , \6266 , \6225 );
nand \mul_6_18_g42470/U$1 ( \6275 , \6273 , \6274 );
not \mul_6_18_g42409/U$1 ( \6276 , \6275 );
not \mul_6_18_g42151/U$3 ( \6277 , \6276 );
and \mul_6_18_g44069/U$2 ( \6278 , \2058 , \3257 );
not \mul_6_18_g44069/U$4 ( \6279 , \2058 );
and \mul_6_18_g44069/U$3 ( \6280 , \6279 , \2816 );
nor \mul_6_18_g44069/U$1 ( \6281 , \6278 , \6280 );
not \mul_6_18_g43120/U$3 ( \6282 , \6281 );
not \mul_6_18_g43120/U$4 ( \6283 , \2510 );
or \mul_6_18_g43120/U$2 ( \6284 , \6282 , \6283 );
nand \mul_6_18_g43532/U$1 ( \6285 , \2514 , \4771 );
nand \mul_6_18_g43120/U$1 ( \6286 , \6284 , \6285 );
not \mul_6_18_g43931/U$3 ( \6287 , \2113 );
not \mul_6_18_g43931/U$4 ( \6288 , \2614 );
or \mul_6_18_g43931/U$2 ( \6289 , \6287 , \6288 );
nand \mul_6_18_g44239/U$1 ( \6290 , \2418 , \3899 );
nand \mul_6_18_g43931/U$1 ( \6291 , \6289 , \6290 );
not \mul_6_18_g42932/U$3 ( \6292 , \6291 );
not \mul_6_18_g42932/U$4 ( \6293 , \4264 );
or \mul_6_18_g42932/U$2 ( \6294 , \6292 , \6293 );
nand \mul_6_18_g43021/U$1 ( \6295 , \2434 , \4792 );
nand \mul_6_18_g42932/U$1 ( \6296 , \6294 , \6295 );
not \mul_6_18_g42597/U$3 ( \6297 , \6296 );
nand \mul_6_18_g43652/U$1 ( \6298 , \2514 , \2058 );
not \mul_6_18_g43651/U$1 ( \6299 , \6298 );
not \mul_6_18_g42597/U$4 ( \6300 , \6299 );
or \mul_6_18_g42597/U$2 ( \6301 , \6297 , \6300 );
or \mul_6_18_g42678/U$2 ( \6302 , \6299 , \6296 );
not \mul_6_18_g43955/U$3 ( \6303 , \2092 );
not \mul_6_18_g43955/U$4 ( \6304 , \2909 );
or \mul_6_18_g43955/U$2 ( \6305 , \6303 , \6304 );
nand \mul_6_18_g44266/U$1 ( \6306 , \2606 , \2754 );
nand \mul_6_18_g43955/U$1 ( \6307 , \6305 , \6306 );
not \mul_6_18_g42975/U$3 ( \6308 , \6307 );
not \mul_6_18_g42975/U$4 ( \6309 , \4002 );
or \mul_6_18_g42975/U$2 ( \6310 , \6308 , \6309 );
nand \mul_6_18_g43020/U$1 ( \6311 , \4005 , \4893 );
nand \mul_6_18_g42975/U$1 ( \6312 , \6310 , \6311 );
nand \mul_6_18_g42678/U$1 ( \6313 , \6302 , \6312 );
nand \mul_6_18_g42597/U$1 ( \6314 , \6301 , \6313 );
xor \mul_6_18_g42385/U$1 ( \6315 , \6286 , \6314 );
not \mul_6_18_g44114/U$3 ( \6316 , \2168 );
not \mul_6_18_g44114/U$4 ( \6317 , \3237 );
or \mul_6_18_g44114/U$2 ( \6318 , \6316 , \6317 );
nand \mul_6_18_g44365/U$1 ( \6319 , \2307 , \3154 );
nand \mul_6_18_g44114/U$1 ( \6320 , \6318 , \6319 );
not \mul_6_18_g43159/U$3 ( \6321 , \6320 );
not \mul_6_18_g43159/U$4 ( \6322 , \2302 );
or \mul_6_18_g43159/U$2 ( \6323 , \6321 , \6322 );
nand \mul_6_18_g43633/U$1 ( \6324 , \4904 , \2317 );
nand \mul_6_18_g43159/U$1 ( \6325 , \6323 , \6324 );
not \mul_6_18_g43982/U$3 ( \6326 , \2111 );
not \mul_6_18_g43982/U$4 ( \6327 , \5929 );
or \mul_6_18_g43982/U$2 ( \6328 , \6326 , \6327 );
nand \mul_6_18_g44278/U$1 ( \6329 , \2252 , \2779 );
nand \mul_6_18_g43982/U$1 ( \6330 , \6328 , \6329 );
not \mul_6_18_g43289/U$3 ( \6331 , \6330 );
not \mul_6_18_g43289/U$4 ( \6332 , \2938 );
or \mul_6_18_g43289/U$2 ( \6333 , \6331 , \6332 );
nand \mul_6_18_g43488/U$1 ( \6334 , \4883 , \3449 );
nand \mul_6_18_g43289/U$1 ( \6335 , \6333 , \6334 );
or \mul_6_18_g42857/U$2 ( \6336 , \6325 , \6335 );
not \mul_6_18_g44135/U$3 ( \6337 , \2056 );
not \mul_6_18_g44135/U$4 ( \6338 , \3920 );
or \mul_6_18_g44135/U$2 ( \6339 , \6337 , \6338 );
nand \mul_6_18_g44386/U$1 ( \6340 , \3330 , \3360 );
nand \mul_6_18_g44135/U$1 ( \6341 , \6339 , \6340 );
not \mul_6_18_g43133/U$3 ( \6342 , \6341 );
not \mul_6_18_g43133/U$4 ( \6343 , \2771 );
or \mul_6_18_g43133/U$2 ( \6344 , \6342 , \6343 );
nand \mul_6_18_g43625/U$1 ( \6345 , \2783 , \4874 );
nand \mul_6_18_g43133/U$1 ( \6346 , \6344 , \6345 );
nand \mul_6_18_g42857/U$1 ( \6347 , \6336 , \6346 );
nand \mul_6_18_g42891/U$1 ( \6348 , \6325 , \6335 );
nand \mul_6_18_g42807/U$1 ( \6349 , \6347 , \6348 );
xnor \mul_6_18_g42385/U$1_r1 ( \6350 , \6315 , \6349 );
not \mul_6_18_g43226/U$3 ( \6351 , \6261 );
not \mul_6_18_g43226/U$4 ( \6352 , \2399 );
or \mul_6_18_g43226/U$2 ( \6353 , \6351 , \6352 );
nand \mul_6_18_g43451/U$1 ( \6354 , \2403 , \4693 );
nand \mul_6_18_g43226/U$1 ( \6355 , \6353 , \6354 );
not \mul_6_18_g44068/U$3 ( \6356 , \2463 );
not \mul_6_18_g44068/U$4 ( \6357 , \2645 );
or \mul_6_18_g44068/U$2 ( \6358 , \6356 , \6357 );
nand \mul_6_18_g44335/U$1 ( \6359 , \3380 , \2468 );
nand \mul_6_18_g44068/U$1 ( \6360 , \6358 , \6359 );
and \mul_6_18_g43180/U$2 ( \6361 , \2349 , \6360 );
and \mul_6_18_g43180/U$3 ( \6362 , \2358 , \4782 );
nor \mul_6_18_g43180/U$1 ( \6363 , \6361 , \6362 );
not \mul_6_18_g43179/U$1 ( \6364 , \6363 );
xor \mul_6_18_g45200/U$1 ( \6365 , \6355 , \6364 );
and \mul_6_18_g43681/U$2 ( \6366 , \4798 , \2765 );
nor \mul_6_18_g43681/U$1 ( \6367 , \6366 , \4804 );
not \mul_6_18_g42814/U$3 ( \6368 , \6367 );
not \mul_6_18_g42922/U$1 ( \6369 , \4797 );
not \mul_6_18_g42814/U$4 ( \6370 , \6369 );
or \mul_6_18_g42814/U$2 ( \6371 , \6368 , \6370 );
or \mul_6_18_g42814/U$5 ( \6372 , \6369 , \4805 );
nand \mul_6_18_g42814/U$1 ( \6373 , \6371 , \6372 );
xnor \mul_6_18_g45200/U$1_r1 ( \6374 , \6365 , \6373 );
nand \mul_6_18_g42277/U$1 ( \6375 , \6350 , \6374 );
not \mul_6_18_g44086/U$3 ( \6376 , \2006 );
not \mul_6_18_g44086/U$4 ( \6377 , \2645 );
or \mul_6_18_g44086/U$2 ( \6378 , \6376 , \6377 );
nand \mul_6_18_g44344/U$1 ( \6379 , \3380 , \2795 );
nand \mul_6_18_g44086/U$1 ( \6380 , \6378 , \6379 );
not \mul_6_18_g43192/U$3 ( \6381 , \6380 );
not \mul_6_18_g43192/U$4 ( \6382 , \2349 );
or \mul_6_18_g43192/U$2 ( \6383 , \6381 , \6382 );
nand \mul_6_18_g43507/U$1 ( \6384 , \2359 , \6360 );
nand \mul_6_18_g43192/U$1 ( \6385 , \6383 , \6384 );
not \mul_6_18_g43929/U$3 ( \6386 , \2640 );
not \mul_6_18_g43929/U$4 ( \6387 , \2423 );
or \mul_6_18_g43929/U$2 ( \6388 , \6386 , \6387 );
nand \mul_6_18_g44253/U$1 ( \6389 , \5561 , \2639 );
nand \mul_6_18_g43929/U$1 ( \6390 , \6388 , \6389 );
not \mul_6_18_g42931/U$3 ( \6391 , \6390 );
not \mul_6_18_g42931/U$4 ( \6392 , \2586 );
or \mul_6_18_g42931/U$2 ( \6393 , \6391 , \6392 );
nand \mul_6_18_g43018/U$1 ( \6394 , \2434 , \6291 );
nand \mul_6_18_g42931/U$1 ( \6395 , \6393 , \6394 );
not \mul_6_18_g45144/U$2 ( \6396 , \6395 );
not \mul_6_18_g43721/U$3 ( \6397 , \2116 );
not \mul_6_18_g44750/U$1 ( \6398 , \1229 );
not \mul_6_18_g43721/U$4 ( \6399 , \6398 );
or \mul_6_18_g43721/U$2 ( \6400 , \6397 , \6399 );
nand \mul_6_18_g43721/U$1 ( \6401 , \6400 , \2311 );
not \mul_6_18_g45272/U$2 ( \6402 , \6398 );
nand \mul_6_18_g45272/U$1 ( \6403 , \6402 , \2058 );
nand \mul_6_18_g43679/U$1 ( \6404 , \6401 , \2761 , \6403 );
nor \mul_6_18_g45144/U$1 ( \6405 , \6396 , \6404 );
xor \mul_6_18_g42444/U$4 ( \6406 , \6385 , \6405 );
not \mul_6_18_g42619/U$3 ( \6407 , \6312 );
not \mul_6_18_g42812/U$3 ( \6408 , \6296 );
not \mul_6_18_g42812/U$4 ( \6409 , \6298 );
and \mul_6_18_g42812/U$2 ( \6410 , \6408 , \6409 );
and \mul_6_18_g42812/U$5 ( \6411 , \6296 , \6298 );
nor \mul_6_18_g42812/U$1 ( \6412 , \6410 , \6411 );
not \mul_6_18_g42619/U$4 ( \6413 , \6412 );
or \mul_6_18_g42619/U$2 ( \6414 , \6407 , \6413 );
or \mul_6_18_g42619/U$5 ( \6415 , \6412 , \6312 );
nand \mul_6_18_g42619/U$1 ( \6416 , \6414 , \6415 );
and \mul_6_18_g42444/U$3 ( \6417 , \6406 , \6416 );
and \mul_6_18_g42444/U$5 ( \6418 , \6385 , \6405 );
or \mul_6_18_g42444/U$2 ( \6419 , \6417 , \6418 );
and \mul_6_18_g42226/U$2 ( \6420 , \6375 , \6419 );
nor \mul_6_18_g42276/U$1 ( \6421 , \6350 , \6374 );
nor \mul_6_18_g42226/U$1 ( \6422 , \6420 , \6421 );
not \mul_6_18_g42151/U$4 ( \6423 , \6422 );
or \mul_6_18_g42151/U$2 ( \6424 , \6277 , \6423 );
xor \mul_6_18_g42711/U$1 ( \6425 , \4687 , \4698 );
xor \mul_6_18_g42711/U$1_r1 ( \6426 , \6425 , \4710 );
not \mul_6_18_g43225/U$1 ( \6427 , \6355 );
not \mul_6_18_g43224/U$1 ( \6428 , \6427 );
not \mul_6_18_g42602/U$3 ( \6429 , \6428 );
not \mul_6_18_g42602/U$4 ( \6430 , \6364 );
or \mul_6_18_g42602/U$2 ( \6431 , \6429 , \6430 );
not \mul_6_18_g42683/U$3 ( \6432 , \6427 );
not \mul_6_18_g42683/U$4 ( \6433 , \6363 );
or \mul_6_18_g42683/U$2 ( \6434 , \6432 , \6433 );
nand \mul_6_18_g42683/U$1 ( \6435 , \6434 , \6373 );
nand \mul_6_18_g42602/U$1 ( \6436 , \6431 , \6435 );
xor \mul_6_18_g45196/U$1 ( \6437 , \6426 , \6436 );
xor \mul_6_18_g45215/U$1 ( \6438 , \4733 , \4723 );
xnor \mul_6_18_g45215/U$1_r1 ( \6439 , \6438 , \4743 );
xnor \mul_6_18_g45196/U$1_r1 ( \6440 , \6437 , \6439 );
nand \mul_6_18_g42151/U$1 ( \6441 , \6424 , \6440 );
not \mul_6_18_g45173/U$2 ( \6442 , \6276 );
not \mul_6_18_g42198/U$1 ( \6443 , \6422 );
nand \mul_6_18_g45173/U$1 ( \6444 , \6442 , \6443 );
nand \mul_6_18_g42130/U$1 ( \6445 , \6441 , \6444 );
xor \g45358/U$1 ( \6446 , \6223 , \6445 );
xor \g45813/U$1 ( \6447 , \4806 , \4787 );
xor \g45813/U$1_r1 ( \6448 , \6447 , \4777 );
not \mul_6_18_g42482/U$1 ( \6449 , \6448 );
not \mul_6_18_g42246/U$3 ( \6450 , \6449 );
not \mul_6_18_g42484/U$3 ( \6451 , \4912 );
not \mul_6_18_g42484/U$4 ( \6452 , \4924 );
or \mul_6_18_g42484/U$2 ( \6453 , \6451 , \6452 );
or \mul_6_18_g42484/U$5 ( \6454 , \4912 , \4924 );
nand \mul_6_18_g42484/U$1 ( \6455 , \6453 , \6454 );
not \mul_6_18_g42727/U$1 ( \6456 , \4882 );
and \mul_6_18_g42427/U$2 ( \6457 , \6455 , \6456 );
not \mul_6_18_g42427/U$4 ( \6458 , \6455 );
and \mul_6_18_g42427/U$3 ( \6459 , \6458 , \4882 );
nor \mul_6_18_g42427/U$1 ( \6460 , \6457 , \6459 );
not \mul_6_18_g42375/U$1 ( \6461 , \6460 );
not \mul_6_18_g42246/U$4 ( \6462 , \6461 );
or \mul_6_18_g42246/U$2 ( \6463 , \6450 , \6462 );
not \mul_6_18_g42284/U$3 ( \6464 , \6448 );
not \mul_6_18_g42284/U$4 ( \6465 , \6460 );
or \mul_6_18_g42284/U$2 ( \6466 , \6464 , \6465 );
not \mul_6_18_g43119/U$1 ( \6467 , \6286 );
not \mul_6_18_g43118/U$1 ( \6468 , \6467 );
not \mul_6_18_g42349/U$3 ( \6469 , \6468 );
not \mul_6_18_g42554/U$1 ( \6470 , \6314 );
not \mul_6_18_g42553/U$1 ( \6471 , \6470 );
not \mul_6_18_g42349/U$4 ( \6472 , \6471 );
or \mul_6_18_g42349/U$2 ( \6473 , \6469 , \6472 );
not \mul_6_18_g42393/U$3 ( \6474 , \6467 );
not \mul_6_18_g42393/U$4 ( \6475 , \6470 );
or \mul_6_18_g42393/U$2 ( \6476 , \6474 , \6475 );
nand \mul_6_18_g42393/U$1 ( \6477 , \6476 , \6349 );
nand \mul_6_18_g42349/U$1 ( \6478 , \6473 , \6477 );
nand \mul_6_18_g42284/U$1 ( \6479 , \6466 , \6478 );
nand \mul_6_18_g42246/U$1 ( \6480 , \6463 , \6479 );
not \mul_6_18_g42138/U$3 ( \6481 , \6480 );
xor \mul_6_18_g42261/U$1 ( \6482 , \4757 , \4766 );
xor \mul_6_18_g42261/U$1_r1 ( \6483 , \6482 , \4809 );
not \mul_6_18_g42208/U$3 ( \6484 , \6483 );
not \mul_6_18_g42710/U$1 ( \6485 , \6426 );
not \mul_6_18_g42434/U$3 ( \6486 , \6485 );
not \mul_6_18_g42434/U$4 ( \6487 , \6439 );
or \mul_6_18_g42434/U$2 ( \6488 , \6486 , \6487 );
nand \mul_6_18_g42434/U$1 ( \6489 , \6488 , \6436 );
not \mul_6_18_g45178/U$2 ( \6490 , \6489 );
nor \mul_6_18_g42590/U$1 ( \6491 , \6439 , \6485 );
nor \mul_6_18_g45178/U$1 ( \6492 , \6490 , \6491 );
not \mul_6_18_g42208/U$4 ( \6493 , \6492 );
and \mul_6_18_g42208/U$2 ( \6494 , \6484 , \6493 );
and \mul_6_18_g42208/U$5 ( \6495 , \6483 , \6492 );
nor \mul_6_18_g42208/U$1 ( \6496 , \6494 , \6495 );
not \mul_6_18_g42138/U$4 ( \6497 , \6496 );
and \mul_6_18_g42138/U$2 ( \6498 , \6481 , \6497 );
and \mul_6_18_g42138/U$5 ( \6499 , \6480 , \6496 );
nor \mul_6_18_g42138/U$1 ( \6500 , \6498 , \6499 );
and \g45357/U$2 ( \6501 , \6446 , \6500 );
not \g45357/U$4 ( \6502 , \6446 );
not \mul_6_18_g42103/U$1 ( \6503 , \6500 );
and \g45357/U$3 ( \6504 , \6502 , \6503 );
nor \g45357/U$1 ( \6505 , \6501 , \6504 );
not \mul_6_18_g42264/U$3 ( \6506 , \6449 );
not \mul_6_18_g42339/U$1 ( \6507 , \6478 );
not \mul_6_18_g42264/U$4 ( \6508 , \6507 );
or \mul_6_18_g42264/U$2 ( \6509 , \6506 , \6508 );
nand \mul_6_18_g42275/U$1 ( \6510 , \6478 , \6448 );
nand \mul_6_18_g42264/U$1 ( \6511 , \6509 , \6510 );
and \mul_6_18_g42210/U$2 ( \6512 , \6511 , \6460 );
not \mul_6_18_g42210/U$4 ( \6513 , \6511 );
and \mul_6_18_g42210/U$3 ( \6514 , \6513 , \6461 );
nor \mul_6_18_g42210/U$1 ( \6515 , \6512 , \6514 );
not \mul_6_18_g44113/U$3 ( \6516 , \2144 );
not \mul_6_18_g44113/U$4 ( \6517 , \3237 );
or \mul_6_18_g44113/U$2 ( \6518 , \6516 , \6517 );
nand \mul_6_18_g44364/U$1 ( \6519 , \2307 , \2145 );
nand \mul_6_18_g44113/U$1 ( \6520 , \6518 , \6519 );
not \mul_6_18_g43161/U$3 ( \6521 , \6520 );
not \mul_6_18_g43161/U$4 ( \6522 , \4049 );
or \mul_6_18_g43161/U$2 ( \6523 , \6521 , \6522 );
nand \mul_6_18_g43505/U$1 ( \6524 , \2317 , \6320 );
nand \mul_6_18_g43161/U$1 ( \6525 , \6523 , \6524 );
not \g45790/U$3 ( \6526 , \6525 );
not \mul_6_18_g43956/U$3 ( \6527 , \2107 );
not \mul_6_18_g43956/U$4 ( \6528 , \3186 );
or \mul_6_18_g43956/U$2 ( \6529 , \6527 , \6528 );
nand \mul_6_18_g44268/U$1 ( \6530 , \2606 , \5229 );
nand \mul_6_18_g43956/U$1 ( \6531 , \6529 , \6530 );
not \mul_6_18_g42973/U$3 ( \6532 , \6531 );
not \mul_6_18_g42973/U$4 ( \6533 , \4002 );
or \mul_6_18_g42973/U$2 ( \6534 , \6532 , \6533 );
nand \mul_6_18_g43019/U$1 ( \6535 , \4005 , \6307 );
nand \mul_6_18_g42973/U$1 ( \6536 , \6534 , \6535 );
not \g45790/U$4 ( \6537 , \6536 );
or \g45790/U$2 ( \6538 , \6526 , \6537 );
not \mul_6_18_g42972/U$1 ( \6539 , \6536 );
not \g45791/U$3 ( \6540 , \6539 );
not \mul_6_18_fopt45130/U$1 ( \6541 , \6525 );
not \g45791/U$4 ( \6542 , \6541 );
or \g45791/U$2 ( \6543 , \6540 , \6542 );
and \g45520/U$2 ( \6544 , \2251 , \2094 );
not \g45520/U$4 ( \6545 , \2251 );
and \g45520/U$3 ( \6546 , \6545 , \2500 );
or \g45520/U$1 ( \6547 , \6544 , \6546 );
not \mul_6_18_g43293/U$3 ( \6548 , \6547 );
not \mul_6_18_g43293/U$4 ( \6549 , \2938 );
or \mul_6_18_g43293/U$2 ( \6550 , \6548 , \6549 );
nand \mul_6_18_g43601/U$1 ( \6551 , \3232 , \6330 );
nand \mul_6_18_g43293/U$1 ( \6552 , \6550 , \6551 );
nand \g45791/U$1 ( \6553 , \6543 , \6552 );
nand \g45790/U$1 ( \6554 , \6538 , \6553 );
xnor \mul_6_18_g45563/U$1 ( \6555 , \2225 , \1970 );
not \mul_6_18_g43908/U$1 ( \6556 , \6555 );
not \mul_6_18_g43365/U$3 ( \6557 , \6556 );
not \mul_6_18_g43365/U$4 ( \6558 , \2222 );
or \mul_6_18_g43365/U$2 ( \6559 , \6557 , \6558 );
nand \mul_6_18_g43604/U$1 ( \6560 , \6232 , \3430 );
nand \mul_6_18_g43365/U$1 ( \6561 , \6559 , \6560 );
not \mul_6_18_g44013/U$3 ( \6562 , \2810 );
not \mul_6_18_g44013/U$4 ( \6563 , \2718 );
or \mul_6_18_g44013/U$2 ( \6564 , \6562 , \6563 );
nand \mul_6_18_g44305/U$1 ( \6565 , \2714 , \2811 );
nand \mul_6_18_g44013/U$1 ( \6566 , \6564 , \6565 );
not \mul_6_18_g43256/U$3 ( \6567 , \6566 );
not \mul_6_18_g43256/U$4 ( \6568 , \2965 );
or \mul_6_18_g43256/U$2 ( \6569 , \6567 , \6568 );
nand \mul_6_18_g43502/U$1 ( \6570 , \6242 , \2733 );
nand \mul_6_18_g43256/U$1 ( \6571 , \6569 , \6570 );
xor \mul_6_18_g42732/U$4 ( \6572 , \6561 , \6571 );
and \mul_6_18_g44089/U$2 ( \6573 , \2116 , \3331 );
not \mul_6_18_g44089/U$4 ( \6574 , \2116 );
and \mul_6_18_g44089/U$3 ( \6575 , \6574 , \3330 );
nor \mul_6_18_g44089/U$1 ( \6576 , \6573 , \6575 );
not \mul_6_18_g43134/U$3 ( \6577 , \6576 );
not \mul_6_18_g43134/U$4 ( \6578 , \2771 );
or \mul_6_18_g43134/U$2 ( \6579 , \6577 , \6578 );
nand \mul_6_18_g43503/U$1 ( \6580 , \6341 , \2783 );
nand \mul_6_18_g43134/U$1 ( \6581 , \6579 , \6580 );
and \mul_6_18_g42732/U$3 ( \6582 , \6572 , \6581 );
and \mul_6_18_g42732/U$5 ( \6583 , \6561 , \6571 );
or \mul_6_18_g42732/U$2 ( \6584 , \6582 , \6583 );
xor \mul_6_18_g42325/U$4 ( \6585 , \6554 , \6584 );
not \mul_6_18_g44059/U$3 ( \6586 , \2463 );
not \mul_6_18_g44059/U$4 ( \6587 , \2367 );
or \mul_6_18_g44059/U$2 ( \6588 , \6586 , \6587 );
nand \mul_6_18_g44326/U$1 ( \6589 , \5165 , \2468 );
nand \mul_6_18_g44059/U$1 ( \6590 , \6588 , \6589 );
not \mul_6_18_g43220/U$3 ( \6591 , \6590 );
not \mul_6_18_g43220/U$4 ( \6592 , \2399 );
or \mul_6_18_g43220/U$2 ( \6593 , \6591 , \6592 );
nand \mul_6_18_g43565/U$1 ( \6594 , \2403 , \6253 );
nand \mul_6_18_g43220/U$1 ( \6595 , \6593 , \6594 );
not \mul_6_18_g44087/U$3 ( \6596 , \2179 );
not \mul_6_18_g44087/U$4 ( \6597 , \2330 );
or \mul_6_18_g44087/U$2 ( \6598 , \6596 , \6597 );
nand \mul_6_18_g44354/U$1 ( \6599 , \2329 , \2185 );
nand \mul_6_18_g44087/U$1 ( \6600 , \6598 , \6599 );
not \mul_6_18_g43199/U$3 ( \6601 , \6600 );
not \mul_6_18_g43199/U$4 ( \6602 , \2349 );
or \mul_6_18_g43199/U$2 ( \6603 , \6601 , \6602 );
nand \mul_6_18_g43500/U$1 ( \6604 , \2359 , \6380 );
nand \mul_6_18_g43199/U$1 ( \6605 , \6603 , \6604 );
xor \mul_6_18_g42483/U$4 ( \6606 , \6595 , \6605 );
not \mul_6_18_g42815/U$3 ( \6607 , \6404 );
not \mul_6_18_g42815/U$4 ( \6608 , \6395 );
or \mul_6_18_g42815/U$2 ( \6609 , \6607 , \6608 );
or \mul_6_18_g42815/U$5 ( \6610 , \6404 , \6395 );
nand \mul_6_18_g42815/U$1 ( \6611 , \6609 , \6610 );
and \mul_6_18_g42483/U$3 ( \6612 , \6606 , \6611 );
and \mul_6_18_g42483/U$5 ( \6613 , \6595 , \6605 );
or \mul_6_18_g42483/U$2 ( \6614 , \6612 , \6613 );
and \mul_6_18_g42325/U$3 ( \6615 , \6585 , \6614 );
and \mul_6_18_g42325/U$5 ( \6616 , \6554 , \6584 );
or \mul_6_18_g42325/U$2 ( \6617 , \6615 , \6616 );
not \mul_6_18_g42324/U$1 ( \6618 , \6617 );
not \mul_6_18_g42189/U$3 ( \6619 , \6618 );
xor \mul_6_18_g45139/U$1 ( \6620 , \6266 , \6225 );
xor \mul_6_18_g45139/U$1_r1 ( \6621 , \6620 , \6271 );
not \mul_6_18_g42189/U$4 ( \6622 , \6621 );
or \mul_6_18_g42189/U$2 ( \6623 , \6619 , \6622 );
xor \mul_6_18_g42628/U$1 ( \6624 , \6237 , \6247 );
xor \mul_6_18_g42628/U$1_r1 ( \6625 , \6624 , \6263 );
not \mul_6_18_g45190/U$2 ( \6626 , \6625 );
xor \g45454/U$1 ( \6627 , \6325 , \6346 );
xor \g45454/U$1_r1 ( \6628 , \6627 , \6335 );
not \mul_6_18_g42709/U$1 ( \6629 , \6628 );
nand \mul_6_18_g45190/U$1 ( \6630 , \6626 , \6629 );
not \mul_6_18_g42292/U$3 ( \6631 , \6630 );
nor \mul_6_18_g43655/U$1 ( \6632 , \2782 , \2116 );
not \g45798/U$3 ( \6633 , \2434 );
not \g45798/U$4 ( \6634 , \6390 );
or \g45798/U$2 ( \6635 , \6633 , \6634 );
not \g45799/U$2 ( \6636 , \2447 );
nand \g45799/U$1 ( \6637 , \6636 , \5310 );
nand \g45798/U$1 ( \6638 , \6635 , \6637 );
xor \mul_6_18_g42584/U$4 ( \6639 , \6632 , \6638 );
not \g45749/U$3 ( \6640 , \2842 );
not \g45749/U$4 ( \6641 , \6531 );
or \g45749/U$2 ( \6642 , \6640 , \6641 );
not \mul_6_18_g43976/U$1 ( \6643 , \5043 );
or \g45749/U$5 ( \6644 , \6643 , \5046 );
nand \g45749/U$1 ( \6645 , \6642 , \6644 );
and \mul_6_18_g42584/U$3 ( \6646 , \6639 , \6645 );
and \mul_6_18_g42584/U$5 ( \6647 , \6632 , \6638 );
or \mul_6_18_g42584/U$2 ( \6648 , \6646 , \6647 );
not \mul_6_18_g43187/U$3 ( \6649 , \4120 );
not \mul_6_18_g43187/U$4 ( \6650 , \5288 );
or \mul_6_18_g43187/U$2 ( \6651 , \6649 , \6650 );
nand \mul_6_18_g43534/U$1 ( \6652 , \2358 , \6600 );
nand \mul_6_18_g43187/U$1 ( \6653 , \6651 , \6652 );
buf \mul_6_18_g43186/U$1 ( \6654 , \6653 );
not \mul_6_18_g43218/U$3 ( \6655 , \4996 );
not \mul_6_18_g43218/U$4 ( \6656 , \2400 );
or \mul_6_18_g43218/U$2 ( \6657 , \6655 , \6656 );
nand \mul_6_18_g43493/U$1 ( \6658 , \2403 , \6590 );
nand \mul_6_18_g43218/U$1 ( \6659 , \6657 , \6658 );
or \mul_6_18_g42855/U$2 ( \6660 , \6654 , \6659 );
not \mul_6_18_g43252/U$3 ( \6661 , \5015 );
not \mul_6_18_g43252/U$4 ( \6662 , \2729 );
or \mul_6_18_g43252/U$2 ( \6663 , \6661 , \6662 );
nand \mul_6_18_g43495/U$1 ( \6664 , \4327 , \6566 );
nand \mul_6_18_g43252/U$1 ( \6665 , \6663 , \6664 );
nand \mul_6_18_g42855/U$1 ( \6666 , \6660 , \6665 );
nand \mul_6_18_g42887/U$1 ( \6667 , \6654 , \6659 );
nand \mul_6_18_g42805/U$1 ( \6668 , \6666 , \6667 );
xor \mul_6_18_g42377/U$4 ( \6669 , \6648 , \6668 );
not \mul_6_18_g43362/U$3 ( \6670 , \6555 );
not \mul_6_18_g43362/U$4 ( \6671 , \6002 );
and \mul_6_18_g43362/U$2 ( \6672 , \6670 , \6671 );
and \mul_6_18_g43362/U$5 ( \6673 , \5035 , \2222 );
nor \mul_6_18_g43362/U$1 ( \6674 , \6672 , \6673 );
not \mul_6_18_g42744/U$3 ( \6675 , \6674 );
not \mul_6_18_g43155/U$3 ( \6676 , \5065 );
not \mul_6_18_g43155/U$4 ( \6677 , \4049 );
or \mul_6_18_g43155/U$2 ( \6678 , \6676 , \6677 );
nand \mul_6_18_g43489/U$1 ( \6679 , \4287 , \6520 );
nand \mul_6_18_g43155/U$1 ( \6680 , \6678 , \6679 );
not \mul_6_18_g43153/U$1 ( \6681 , \6680 );
not \mul_6_18_g42744/U$4 ( \6682 , \6681 );
or \mul_6_18_g42744/U$2 ( \6683 , \6675 , \6682 );
not \mul_6_18_g43285/U$3 ( \6684 , \4979 );
not \mul_6_18_g43285/U$4 ( \6685 , \2274 );
or \mul_6_18_g43285/U$2 ( \6686 , \6684 , \6685 );
nand \mul_6_18_g43491/U$1 ( \6687 , \3232 , \6547 );
nand \mul_6_18_g43285/U$1 ( \6688 , \6686 , \6687 );
nand \mul_6_18_g42744/U$1 ( \6689 , \6683 , \6688 );
not \mul_6_18_g45225/U$2 ( \6690 , \6674 );
nand \mul_6_18_g45225/U$1 ( \6691 , \6690 , \6680 );
nand \mul_6_18_g42687/U$1 ( \6692 , \6689 , \6691 );
and \mul_6_18_g42377/U$3 ( \6693 , \6669 , \6692 );
and \mul_6_18_g42377/U$5 ( \6694 , \6648 , \6668 );
or \mul_6_18_g42377/U$2 ( \6695 , \6693 , \6694 );
not \mul_6_18_g42292/U$4 ( \6696 , \6695 );
or \mul_6_18_g42292/U$2 ( \6697 , \6631 , \6696 );
nand \mul_6_18_g42540/U$1 ( \6698 , \6625 , \6628 );
nand \mul_6_18_g42292/U$1 ( \6699 , \6697 , \6698 );
nand \mul_6_18_g42189/U$1 ( \6700 , \6623 , \6699 );
not \mul_6_18_g42407/U$1 ( \6701 , \6621 );
nand \mul_6_18_g42282/U$1 ( \6702 , \6701 , \6617 );
and \mul_6_18_g42170/U$1 ( \6703 , \6700 , \6702 );
xor \mul_6_18_g42005/U$4 ( \6704 , \6515 , \6703 );
xor \mul_6_18_g42162/U$1 ( \6705 , \6275 , \6440 );
xnor \mul_6_18_g42162/U$1_r1 ( \6706 , \6705 , \6443 );
and \mul_6_18_g42005/U$3 ( \6707 , \6704 , \6706 );
and \mul_6_18_g42005/U$5 ( \6708 , \6515 , \6703 );
or \mul_6_18_g42005/U$2 ( \6709 , \6707 , \6708 );
nand \mul_6_18_g41976/U$1 ( \6710 , \6505 , \6709 );
xor \mul_6_18_g42005/U$1 ( \6711 , \6515 , \6703 );
xor \mul_6_18_g42005/U$1_r1 ( \6712 , \6711 , \6706 );
not \mul_6_18_g42263/U$3 ( \6713 , \6618 );
not \mul_6_18_g42263/U$4 ( \6714 , \6701 );
or \mul_6_18_g42263/U$2 ( \6715 , \6713 , \6714 );
nand \mul_6_18_g42274/U$1 ( \6716 , \6621 , \6617 );
nand \mul_6_18_g42263/U$1 ( \6717 , \6715 , \6716 );
and \mul_6_18_g45137/U$2 ( \6718 , \6717 , \6699 );
not \mul_6_18_g45137/U$4 ( \6719 , \6717 );
not \mul_6_18_g42248/U$1 ( \6720 , \6699 );
and \mul_6_18_g45137/U$3 ( \6721 , \6719 , \6720 );
nor \mul_6_18_g45137/U$1 ( \6722 , \6718 , \6721 );
xor \mul_6_18_g42444/U$1 ( \6723 , \6385 , \6405 );
xor \mul_6_18_g42444/U$1_r1 ( \6724 , \6723 , \6416 );
xor \mul_6_18_g42325/U$1 ( \6725 , \6554 , \6584 );
xor \mul_6_18_g42325/U$1_r1 ( \6726 , \6725 , \6614 );
xor \mul_6_18_g42159/U$4 ( \6727 , \6724 , \6726 );
xor \mul_6_18_g42732/U$1 ( \6728 , \6561 , \6571 );
xor \mul_6_18_g42732/U$1_r1 ( \6729 , \6728 , \6581 );
not \mul_6_18_g42824/U$3 ( \6730 , \6525 );
not \mul_6_18_g42824/U$4 ( \6731 , \6539 );
or \mul_6_18_g42824/U$2 ( \6732 , \6730 , \6731 );
nand \mul_6_18_g42828/U$1 ( \6733 , \6541 , \6536 );
nand \mul_6_18_g42824/U$1 ( \6734 , \6732 , \6733 );
xor \mul_6_18_g45220/U$1 ( \6735 , \6734 , \6552 );
xor \mul_6_18_g42301/U$4 ( \6736 , \6729 , \6735 );
xor \mul_6_18_g42483/U$1 ( \6737 , \6595 , \6605 );
xor \mul_6_18_g42483/U$1_r1 ( \6738 , \6737 , \6611 );
and \mul_6_18_g42301/U$3 ( \6739 , \6736 , \6738 );
and \mul_6_18_g42301/U$5 ( \6740 , \6729 , \6735 );
or \mul_6_18_g42301/U$2 ( \6741 , \6739 , \6740 );
and \mul_6_18_g42159/U$3 ( \6742 , \6727 , \6741 );
and \mul_6_18_g42159/U$5 ( \6743 , \6724 , \6726 );
or \mul_6_18_g42159/U$2 ( \6744 , \6742 , \6743 );
xor \g45735/U$1 ( \6745 , \6374 , \6419 );
buf \mul_6_18_g42338/U$1 ( \6746 , \6350 );
xor \g45735/U$1_r1 ( \6747 , \6745 , \6746 );
or \mul_6_18_g45158/U$1 ( \6748 , \6744 , \6747 );
and \mul_6_18_g42041/U$2 ( \6749 , \6722 , \6748 );
and \mul_6_18_g42082/U$2 ( \6750 , \6747 , \6744 );
nor \mul_6_18_g42041/U$1 ( \6751 , \6749 , \6750 );
nand \mul_6_18_g41974/U$1 ( \6752 , \6712 , \6751 );
and \mul_6_18_g41958/U$1 ( \6753 , \6710 , \6752 );
xor \mul_6_18_g41953/U$1 ( \6754 , \4828 , \4939 );
xor \mul_6_18_g41953/U$1_r1 ( \6755 , \6754 , \4942 );
not \mul_6_18_g41951/U$1 ( \6756 , \6755 );
not \mul_6_18_g42139/U$3 ( \6757 , \4934 );
and \g45364/U$2 ( \6758 , \4834 , \4831 );
not \g45364/U$4 ( \6759 , \4834 );
and \g45364/U$3 ( \6760 , \6759 , \4830 );
nor \g45364/U$1 ( \6761 , \6758 , \6760 );
not \mul_6_18_g42139/U$4 ( \6762 , \6761 );
and \mul_6_18_g42139/U$2 ( \6763 , \6757 , \6762 );
and \mul_6_18_g42139/U$5 ( \6764 , \4934 , \6761 );
nor \mul_6_18_g42139/U$1 ( \6765 , \6763 , \6764 );
not \mul_6_18_fopt45122/U$1 ( \6766 , \6765 );
xor \mul_6_18_g42163/U$1 ( \6767 , \4812 , \4752 );
xor \mul_6_18_g42163/U$1_r1 ( \6768 , \6767 , \4754 );
or \mul_6_18_g42019/U$2 ( \6769 , \6766 , \6768 );
not \mul_6_18_g45163/U$2 ( \6770 , \6483 );
nand \mul_6_18_g45163/U$1 ( \6771 , \6770 , \6492 );
not \mul_6_18_g42129/U$3 ( \6772 , \6771 );
not \mul_6_18_g42129/U$4 ( \6773 , \6480 );
or \mul_6_18_g42129/U$2 ( \6774 , \6772 , \6773 );
not \mul_6_18_g45164/U$2 ( \6775 , \6492 );
nand \mul_6_18_g45164/U$1 ( \6776 , \6775 , \6483 );
nand \mul_6_18_g42129/U$1 ( \6777 , \6774 , \6776 );
nand \mul_6_18_g42019/U$1 ( \6778 , \6769 , \6777 );
not \mul_6_18_g42135/U$1 ( \6779 , \6768 );
not \mul_6_18_g42076/U$2 ( \6780 , \6779 );
nand \mul_6_18_g42076/U$1 ( \6781 , \6780 , \6766 );
nand \mul_6_18_g42004/U$1 ( \6782 , \6778 , \6781 );
not \mul_6_18_g41992/U$1 ( \6783 , \6782 );
nand \mul_6_18_g41918/U$1 ( \6784 , \6756 , \6783 );
not \mul_6_18_g42241/U$3 ( \6785 , \5281 );
not \mul_6_18_g42241/U$4 ( \6786 , \5340 );
or \mul_6_18_g42241/U$2 ( \6787 , \6785 , \6786 );
or \mul_6_18_g42287/U$2 ( \6788 , \5340 , \5281 );
nand \mul_6_18_g42287/U$1 ( \6789 , \6788 , \5395 );
nand \mul_6_18_g42241/U$1 ( \6790 , \6787 , \6789 );
not \mul_6_18_g42099/U$3 ( \6791 , \6790 );
xor \mul_6_18_g42872/U$1 ( \6792 , \6665 , \6653 );
not \mul_6_18_g43217/U$1 ( \6793 , \6659 );
and \mul_6_18_g42791/U$2 ( \6794 , \6792 , \6793 );
not \mul_6_18_g42791/U$4 ( \6795 , \6792 );
and \mul_6_18_g42791/U$3 ( \6796 , \6795 , \6659 );
nor \mul_6_18_g42791/U$1 ( \6797 , \6794 , \6796 );
not \mul_6_18_g42707/U$1 ( \6798 , \6797 );
not \mul_6_18_g42586/U$3 ( \6799 , \6798 );
not \g45792/U$3 ( \6800 , \5021 );
not \g45792/U$4 ( \6801 , \4981 );
or \g45792/U$2 ( \6802 , \6800 , \6801 );
not \g45793/U$3 ( \6803 , \4982 );
not \g45793/U$4 ( \6804 , \5018 );
or \g45793/U$2 ( \6805 , \6803 , \6804 );
nand \g45793/U$1 ( \6806 , \6805 , \4998 );
nand \g45792/U$1 ( \6807 , \6802 , \6806 );
not \mul_6_18_g42706/U$1 ( \6808 , \6807 );
not \mul_6_18_g42586/U$4 ( \6809 , \6808 );
or \mul_6_18_g42586/U$2 ( \6810 , \6799 , \6809 );
nand \mul_6_18_g42591/U$1 ( \6811 , \6797 , \6807 );
nand \mul_6_18_g42586/U$1 ( \6812 , \6810 , \6811 );
xor \mul_6_18_g45218/U$1 ( \6813 , \6674 , \6680 );
xor \mul_6_18_g45218/U$1_r1 ( \6814 , \6813 , \6688 );
buf \mul_6_18_g42653/U$1 ( \6815 , \6814 );
not \mul_6_18_g42652/U$1 ( \6816 , \6815 );
and \mul_6_18_g42489/U$2 ( \6817 , \6812 , \6816 );
not \mul_6_18_g42489/U$4 ( \6818 , \6812 );
and \mul_6_18_g42489/U$3 ( \6819 , \6818 , \6815 );
nor \mul_6_18_g42489/U$1 ( \6820 , \6817 , \6819 );
not \mul_6_18_g42099/U$4 ( \6821 , \6820 );
or \mul_6_18_g42099/U$2 ( \6822 , \6791 , \6821 );
or \g45843/U$2 ( \6823 , \6820 , \6790 );
xor \mul_6_18_g42446/U$4 ( \6824 , \5290 , \5313 );
and \mul_6_18_g42446/U$3 ( \6825 , \6824 , \5339 );
and \mul_6_18_g42446/U$5 ( \6826 , \5290 , \5313 );
or \mul_6_18_g42446/U$2 ( \6827 , \6825 , \6826 );
nand \mul_6_18_g42536/U$1 ( \6828 , \5023 , \5107 );
and \mul_6_18_g42471/U$2 ( \6829 , \6828 , \5068 );
nor \mul_6_18_g42535/U$1 ( \6830 , \5023 , \5107 );
nor \mul_6_18_g42471/U$1 ( \6831 , \6829 , \6830 );
not \mul_6_18_g42356/U$1 ( \6832 , \6831 );
xor \g45677/U$1 ( \6833 , \6827 , \6832 );
and \mul_6_18_g42771/U$2 ( \6834 , \5297 , \5312 );
xor \mul_6_18_g42550/U$4 ( \6835 , \5037 , \5052 );
and \mul_6_18_g42550/U$3 ( \6836 , \6835 , \5067 );
and \mul_6_18_g42550/U$5 ( \6837 , \5037 , \5052 );
or \mul_6_18_g42550/U$2 ( \6838 , \6836 , \6837 );
xor \mul_6_18_g42323/U$1 ( \6839 , \6834 , \6838 );
xor \mul_6_18_g42584/U$1 ( \6840 , \6632 , \6638 );
xor \mul_6_18_g42584/U$1_r1 ( \6841 , \6840 , \6645 );
xor \mul_6_18_g42323/U$1_r1 ( \6842 , \6839 , \6841 );
xor \g45677/U$1_r1 ( \6843 , \6833 , \6842 );
nand \g45843/U$1 ( \6844 , \6823 , \6843 );
nand \mul_6_18_g42099/U$1 ( \6845 , \6822 , \6844 );
not \g45671/U$2 ( \6846 , \6845 );
xor \mul_6_18_g42301/U$1 ( \6847 , \6729 , \6735 );
xor \mul_6_18_g42301/U$1_r1 ( \6848 , \6847 , \6738 );
not \mul_6_18_g42247/U$3 ( \6849 , \6827 );
not \mul_6_18_g42247/U$4 ( \6850 , \6832 );
or \mul_6_18_g42247/U$2 ( \6851 , \6849 , \6850 );
not \mul_6_18_g45179/U$2 ( \6852 , \6827 );
nand \mul_6_18_g45179/U$1 ( \6853 , \6852 , \6831 );
nand \mul_6_18_g42286/U$1 ( \6854 , \6842 , \6853 );
nand \mul_6_18_g42247/U$1 ( \6855 , \6851 , \6854 );
and \mul_6_18_g45157/U$2 ( \6856 , \6848 , \6855 );
not \mul_6_18_g45157/U$4 ( \6857 , \6848 );
not \mul_6_18_g42175/U$1 ( \6858 , \6855 );
and \mul_6_18_g45157/U$3 ( \6859 , \6857 , \6858 );
nor \mul_6_18_g45157/U$1 ( \6860 , \6856 , \6859 );
xor \mul_6_18_g42323/U$4 ( \6861 , \6834 , \6838 );
and \mul_6_18_g42323/U$3 ( \6862 , \6861 , \6841 );
and \mul_6_18_g42323/U$5 ( \6863 , \6834 , \6838 );
or \mul_6_18_g42323/U$2 ( \6864 , \6862 , \6863 );
not \mul_6_18_g42513/U$3 ( \6865 , \6814 );
not \mul_6_18_g42513/U$4 ( \6866 , \6808 );
or \mul_6_18_g42513/U$2 ( \6867 , \6865 , \6866 );
nand \mul_6_18_g42513/U$1 ( \6868 , \6867 , \6798 );
not \mul_6_18_g45193/U$2 ( \6869 , \6814 );
nand \mul_6_18_g45193/U$1 ( \6870 , \6869 , \6807 );
nand \mul_6_18_g42469/U$1 ( \6871 , \6868 , \6870 );
xor \mul_6_18_g42158/U$1 ( \6872 , \6864 , \6871 );
xor \mul_6_18_g42377/U$1 ( \6873 , \6648 , \6668 );
xor \mul_6_18_g42377/U$1_r1 ( \6874 , \6873 , \6692 );
xor \mul_6_18_g42158/U$1_r1 ( \6875 , \6872 , \6874 );
not \mul_6_18_g42157/U$1 ( \6876 , \6875 );
and \mul_6_18_g42088/U$2 ( \6877 , \6860 , \6876 );
not \mul_6_18_g42088/U$4 ( \6878 , \6860 );
and \mul_6_18_g42088/U$3 ( \6879 , \6878 , \6875 );
nor \mul_6_18_g42088/U$1 ( \6880 , \6877 , \6879 );
nand \g45671/U$1 ( \6881 , \6846 , \6880 );
xor \mul_6_18_g42112/U$1 ( \6882 , \6820 , \6790 );
xnor \mul_6_18_g42112/U$1_r1 ( \6883 , \6882 , \6843 );
xor \mul_6_18_g42085/U$4 ( \6884 , \5111 , \5274 );
and \mul_6_18_g42085/U$3 ( \6885 , \6884 , \5396 );
and \mul_6_18_g42085/U$5 ( \6886 , \5111 , \5274 );
or \mul_6_18_g42085/U$2 ( \6887 , \6885 , \6886 );
not \mul_6_18_g42084/U$1 ( \6888 , \6887 );
nand \mul_6_18_g42054/U$1 ( \6889 , \6883 , \6888 );
and \mul_6_18_g42018/U$1 ( \6890 , \6881 , \6889 );
xor \mul_6_18_g42082/U$1 ( \6891 , \6747 , \6744 );
and \mul_6_18_g42051/U$2 ( \6892 , \6891 , \6722 );
not \mul_6_18_g42051/U$4 ( \6893 , \6891 );
and \mul_6_18_g2/U$2 ( \6894 , \6717 , \6699 );
not \mul_6_18_g2/U$4 ( \6895 , \6717 );
and \mul_6_18_g2/U$3 ( \6896 , \6895 , \6720 );
or \mul_6_18_g2/U$1 ( \6897 , \6894 , \6896 );
and \mul_6_18_g42051/U$3 ( \6898 , \6893 , \6897 );
nor \mul_6_18_g42051/U$1 ( \6899 , \6892 , \6898 );
not \mul_6_18_g42028/U$1 ( \6900 , \6899 );
and \mul_6_18_g42525/U$2 ( \6901 , \6625 , \6628 );
not \mul_6_18_g42525/U$4 ( \6902 , \6625 );
and \mul_6_18_g42525/U$3 ( \6903 , \6902 , \6629 );
nor \mul_6_18_g42525/U$1 ( \6904 , \6901 , \6903 );
xor \g45393/U$1 ( \6905 , \6695 , \6904 );
xor \mul_6_18_g42158/U$4 ( \6906 , \6864 , \6871 );
and \mul_6_18_g42158/U$3 ( \6907 , \6906 , \6874 );
and \mul_6_18_g42158/U$5 ( \6908 , \6864 , \6871 );
or \mul_6_18_g42158/U$2 ( \6909 , \6907 , \6908 );
xor \mul_6_18_g42044/U$4 ( \6910 , \6905 , \6909 );
xor \mul_6_18_g42159/U$1 ( \6911 , \6724 , \6726 );
xor \mul_6_18_g42159/U$1_r1 ( \6912 , \6911 , \6741 );
and \mul_6_18_g42044/U$3 ( \6913 , \6910 , \6912 );
and \mul_6_18_g42044/U$5 ( \6914 , \6905 , \6909 );
or \mul_6_18_g42044/U$2 ( \6915 , \6913 , \6914 );
not \mul_6_18_g42043/U$1 ( \6916 , \6915 );
nand \mul_6_18_g41999/U$1 ( \6917 , \6900 , \6916 );
xor \mul_6_18_g42044/U$1 ( \6918 , \6905 , \6909 );
xor \mul_6_18_g42044/U$1_r1 ( \6919 , \6918 , \6912 );
not \mul_6_18_g42017/U$2 ( \6920 , \6919 );
not \g45730/U$3 ( \6921 , \6875 );
not \g45730/U$4 ( \6922 , \6848 );
or \g45730/U$2 ( \6923 , \6921 , \6922 );
or \mul_6_18_g42096/U$2 ( \6924 , \6875 , \6848 );
nand \mul_6_18_g42096/U$1 ( \6925 , \6924 , \6855 );
nand \g45730/U$1 ( \6926 , \6923 , \6925 );
not \mul_6_18_g42067/U$1 ( \6927 , \6926 );
nand \mul_6_18_g42017/U$1 ( \6928 , \6920 , \6927 );
and \mul_6_18_g41967/U$1 ( \6929 , \6890 , \6917 , \6928 );
not \mul_6_18_g42071/U$3 ( \6930 , \6779 );
not \mul_6_18_fopt45123/U$1 ( \6931 , \6765 );
not \mul_6_18_g42071/U$4 ( \6932 , \6931 );
or \mul_6_18_g42071/U$2 ( \6933 , \6930 , \6932 );
nand \mul_6_18_g42075/U$1 ( \6934 , \6765 , \6768 );
nand \mul_6_18_g42071/U$1 ( \6935 , \6933 , \6934 );
not \mul_6_18_g42104/U$1 ( \6936 , \6777 );
and \mul_6_18_g42007/U$2 ( \6937 , \6935 , \6936 );
not \mul_6_18_g42007/U$4 ( \6938 , \6935 );
and \mul_6_18_g42007/U$3 ( \6939 , \6938 , \6777 );
nor \mul_6_18_g42007/U$1 ( \6940 , \6937 , \6939 );
not \mul_6_18_g42205/U$1 ( \6941 , \6223 );
not \mul_6_18_g42060/U$3 ( \6942 , \6941 );
not \mul_6_18_g42060/U$4 ( \6943 , \6500 );
or \mul_6_18_g42060/U$2 ( \6944 , \6942 , \6943 );
nand \mul_6_18_g42060/U$1 ( \6945 , \6944 , \6445 );
nand \mul_6_18_g42074/U$1 ( \6946 , \6503 , \6223 );
and \mul_6_18_g42042/U$1 ( \6947 , \6945 , \6946 );
nand \mul_6_18_g41966/U$1 ( \6948 , \6940 , \6947 );
and \mul_6_18_g41888/U$1 ( \6949 , \6753 , \6784 , \6929 , \6948 );
not \mul_6_18_g41851/U$4 ( \6950 , \6949 );
or \mul_6_18_g41851/U$2 ( \6951 , \6221 , \6950 );
nand \mul_6_18_g42000/U$1 ( \6952 , \6899 , \6915 );
nand \mul_6_18_g45140/U$1 ( \6953 , \6919 , \6926 );
and \mul_6_18_g41977/U$1 ( \6954 , \6952 , \6953 );
not \mul_6_18_g42066/U$1 ( \6955 , \6880 );
nand \mul_6_18_g42035/U$1 ( \6956 , \6955 , \6845 );
not \mul_6_18_g42086/U$1 ( \6957 , \6883 );
nand \mul_6_18_g42052/U$1 ( \6958 , \6957 , \6887 );
nand \mul_6_18_g42015/U$1 ( \6959 , \6956 , \6958 );
buf \mul_6_18_fopt45053/U$1 ( \6960 , \6881 );
nand \mul_6_18_g41982/U$1 ( \6961 , \6959 , \6928 , \6960 );
nand \mul_6_18_g41968/U$1 ( \6962 , \6954 , \6961 );
not \mul_6_18_g41998/U$1 ( \6963 , \6917 );
not \mul_6_18_g41996/U$1 ( \6964 , \6963 );
and \mul_6_18_g41927/U$1 ( \6965 , \6753 , \6962 , \6964 );
nor \mul_6_18_g41962/U$1 ( \6966 , \6940 , \6947 );
nor \mul_6_18_g41979/U$1 ( \6967 , \6505 , \6709 );
nor \mul_6_18_g41938/U$1 ( \6968 , \6966 , \6967 );
nor \mul_6_18_g41981/U$1 ( \6969 , \6712 , \6751 );
nand \mul_6_18_g41963/U$1 ( \6970 , \6710 , \6969 );
nand \mul_6_18_g41921/U$1 ( \6971 , \6755 , \6782 );
nand \mul_6_18_g41887/U$1 ( \6972 , \6968 , \6970 , \6971 );
or \mul_6_18_g41853/U$2 ( \6973 , \6965 , \6972 );
not \g45729/U$3 ( \6974 , \6784 );
not \g45729/U$4 ( \6975 , \6948 );
or \g45729/U$2 ( \6976 , \6974 , \6975 );
nand \g45729/U$1 ( \6977 , \6976 , \6971 );
nand \mul_6_18_g41853/U$1 ( \6978 , \6973 , \6977 );
nand \mul_6_18_g41851/U$1 ( \6979 , \6951 , \6978 );
not \mul_6_18_g41922/U$2 ( \6980 , \4822 );
not \mul_6_18_g41952/U$1 ( \6981 , \4945 );
nand \mul_6_18_g41922/U$1 ( \6982 , \6980 , \6981 );
nand \mul_6_18_g41875/U$1 ( \6983 , \6982 , \4957 );
nor \mul_6_18_g41863/U$1 ( \6984 , \4671 , \6983 );
and \mul_6_18_g41854/U$1 ( \6985 , \6984 , \4423 );
nand \mul_6_18_g41848/U$1 ( \6986 , \6979 , \6985 );
nand \mul_6_18_g41842/U$1 ( \6987 , \4968 , \6986 );
not \mul_6_18_g41837/U$4 ( \6988 , \6987 );
or \mul_6_18_g41837/U$2 ( \6989 , \4200 , \6988 );
not \mul_6_18_g41872/U$1 ( \6990 , \3761 );
not \mul_6_18_g41936/U$1 ( \6991 , \3985 );
not \mul_6_18_g41989/U$1 ( \6992 , \3987 );
not \mul_6_18_g41947/U$1 ( \6993 , \4196 );
nand \mul_6_18_g41924/U$1 ( \6994 , \6992 , \6993 );
or \mul_6_18_g41882/U$2 ( \6995 , \6991 , \6994 );
not \mul_6_18_g45151/U$2 ( \6996 , \3984 );
buf \mul_6_18_fopt/U$1 ( \6997 , \3763 );
nand \mul_6_18_g45151/U$1 ( \6998 , \6996 , \6997 );
nand \mul_6_18_g41882/U$1 ( \6999 , \6995 , \6998 );
and \mul_6_18_g41856/U$2 ( \7000 , \6990 , \6999 );
and \mul_6_18_g41876/U$1 ( \7001 , \3702 , \3760 );
nor \mul_6_18_g41856/U$1 ( \7002 , \7000 , \7001 );
nand \mul_6_18_g41837/U$1 ( \7003 , \6989 , \7002 );
xor \mul_6_18_g41910/U$4 ( \7004 , \3094 , \3504 );
and \mul_6_18_g41910/U$3 ( \7005 , \7004 , \3701 );
and \mul_6_18_g41910/U$5 ( \7006 , \3094 , \3504 );
or \mul_6_18_g41910/U$2 ( \7007 , \7005 , \7006 );
xor \mul_6_18_g42068/U$4 ( \7008 , \2459 , \2867 );
and \mul_6_18_g42068/U$3 ( \7009 , \7008 , \3093 );
and \mul_6_18_g42068/U$5 ( \7010 , \2459 , \2867 );
or \mul_6_18_g42068/U$2 ( \7011 , \7009 , \7010 );
xor \mul_6_18_g42202/U$4 ( \7012 , \2921 , \3003 );
and \mul_6_18_g42202/U$3 ( \7013 , \7012 , \3092 );
and \mul_6_18_g42202/U$5 ( \7014 , \2921 , \3003 );
or \mul_6_18_g42202/U$2 ( \7015 , \7013 , \7014 );
not \mul_6_18_g42154/U$3 ( \7016 , \7015 );
or \mul_6_18_g42886/U$1 ( \7017 , \2361 , \2408 );
and \mul_6_18_g42604/U$2 ( \7018 , \2457 , \7017 );
and \mul_6_18_g42885/U$1 ( \7019 , \2361 , \2408 );
nor \mul_6_18_g42604/U$1 ( \7020 , \7018 , \7019 );
xor \mul_6_18_g42715/U$4 ( \7021 , \3587 , \3596 );
and \mul_6_18_g42715/U$3 ( \7022 , \7021 , \3607 );
and \mul_6_18_g42715/U$5 ( \7023 , \3587 , \3596 );
or \mul_6_18_g42715/U$2 ( \7024 , \7022 , \7023 );
xnor \g45411/U$1 ( \7025 , \7020 , \7024 );
not \mul_6_18_g42425/U$1 ( \7026 , \7025 );
not \mul_6_18_g42321/U$3 ( \7027 , \7026 );
not \mul_6_18_g43001/U$3 ( \7028 , \2447 );
not \mul_6_18_g43753/U$1 ( \7029 , \2894 );
not \mul_6_18_g43001/U$4 ( \7030 , \7029 );
and \mul_6_18_g43001/U$2 ( \7031 , \7028 , \7030 );
and \mul_6_18_g43752/U$2 ( \7032 , \1807 , \2424 );
not \mul_6_18_g43752/U$4 ( \7033 , \1807 );
and \mul_6_18_g43752/U$3 ( \7034 , \7033 , \2423 );
nor \mul_6_18_g43752/U$1 ( \7035 , \7032 , \7034 );
and \mul_6_18_g43001/U$5 ( \7036 , \2434 , \7035 );
nor \mul_6_18_g43001/U$1 ( \7037 , \7031 , \7036 );
not \mul_6_18_g42801/U$3 ( \7038 , \7037 );
not \mul_6_18_g43071/U$3 ( \7039 , \3594 );
not \mul_6_18_g43071/U$4 ( \7040 , \2202 );
or \mul_6_18_g43071/U$2 ( \7041 , \7039 , \7040 );
and \mul_6_18_g44122/U$2 ( \7042 , \1998 , \2181 );
not \mul_6_18_g44122/U$4 ( \7043 , \1998 );
and \mul_6_18_g44122/U$3 ( \7044 , \7043 , \2182 );
nor \mul_6_18_g44122/U$1 ( \7045 , \7042 , \7044 );
nand \mul_6_18_g43494/U$1 ( \7046 , \7045 , \2210 );
nand \mul_6_18_g43071/U$1 ( \7047 , \7041 , \7046 );
not \mul_6_18_g42801/U$4 ( \7048 , \7047 );
or \mul_6_18_g42801/U$2 ( \7049 , \7038 , \7048 );
or \mul_6_18_g42801/U$5 ( \7050 , \7047 , \7037 );
nand \mul_6_18_g42801/U$1 ( \7051 , \7049 , \7050 );
not \g45797/U$3 ( \7052 , \3573 );
not \g45797/U$4 ( \7053 , \2692 );
or \g45797/U$2 ( \7054 , \7052 , \7053 );
and \mul_6_18_g45247/U$2 ( \7055 , \2694 , \2779 );
not \mul_6_18_g45247/U$4 ( \7056 , \2694 );
and \mul_6_18_g45247/U$3 ( \7057 , \7056 , \2111 );
nor \mul_6_18_g45247/U$1 ( \7058 , \7055 , \7057 );
nand \mul_6_18_g43435/U$1 ( \7059 , \2701 , \7058 );
nand \g45797/U$1 ( \7060 , \7054 , \7059 );
not \fopt45574/U$1 ( \7061 , \5426 );
not \mul_6_18_g42971/U$3 ( \7062 , \7061 );
not \mul_6_18_g42971/U$4 ( \7063 , \2917 );
and \mul_6_18_g42971/U$2 ( \7064 , \7062 , \7063 );
and \mul_6_18_g43756/U$2 ( \7065 , \1784 , \2606 );
not \mul_6_18_g43756/U$4 ( \7066 , \1784 );
and \mul_6_18_g43756/U$3 ( \7067 , \7066 , \2607 );
nor \mul_6_18_g43756/U$1 ( \7068 , \7065 , \7067 );
and \mul_6_18_g42971/U$5 ( \7069 , \2842 , \7068 );
nor \mul_6_18_g42971/U$1 ( \7070 , \7064 , \7069 );
xor \g45796/U$1 ( \7071 , \7060 , \7070 );
xor \g45871/U$1 ( \7072 , \7051 , \7071 );
not \mul_6_18_g43132/U$3 ( \7073 , \3564 );
not \mul_6_18_g43132/U$4 ( \7074 , \2773 );
or \mul_6_18_g43132/U$2 ( \7075 , \7073 , \7074 );
or \mul_6_18_g43981/U$2 ( \7076 , \2765 , \2312 );
or \mul_6_18_g43981/U$3 ( \7077 , \2762 , \2305 );
nand \mul_6_18_g43981/U$1 ( \7078 , \7076 , \7077 );
nand \mul_6_18_g43429/U$1 ( \7079 , \2784 , \7078 );
nand \mul_6_18_g43132/U$1 ( \7080 , \7075 , \7079 );
or \mul_6_18_g43906/U$2 ( \7081 , \2335 , \2369 );
or \mul_6_18_g43906/U$3 ( \7082 , \2336 , \2110 );
nand \mul_6_18_g43906/U$1 ( \7083 , \7081 , \7082 );
and \g45802/U$2 ( \7084 , \2359 , \7083 );
not \g45803/U$2 ( \7085 , \2349 );
nor \g45803/U$1 ( \7086 , \7085 , \2356 );
nor \g45802/U$1 ( \7087 , \7084 , \7086 );
xor \g45768/U$1 ( \7088 , \7080 , \7087 );
not \mul_6_18_g45228/U$2 ( \7089 , \2938 );
nor \mul_6_18_g45228/U$1 ( \7090 , \7089 , \2282 );
and \mul_6_18_g43859/U$2 ( \7091 , \2251 , \2098 );
and \mul_6_18_g43859/U$3 ( \7092 , \2256 , \2582 );
nor \mul_6_18_g43859/U$1 ( \7093 , \7091 , \7092 );
nor \mul_6_18_g43479/U$1 ( \7094 , \7093 , \2284 );
nor \mul_6_18_g43281/U$1 ( \7095 , \7090 , \7094 );
not \mul_6_18_g42867/U$3 ( \7096 , \7095 );
not \mul_6_18_fopt45089/U$1 ( \7097 , \2323 );
not \mul_6_18_g43152/U$3 ( \7098 , \7097 );
not \mul_6_18_g43152/U$4 ( \7099 , \2303 );
or \mul_6_18_g43152/U$2 ( \7100 , \7098 , \7099 );
or \mul_6_18_g43943/U$2 ( \7101 , \2307 , \2670 );
or \mul_6_18_g43943/U$3 ( \7102 , \2308 , \2101 );
nand \mul_6_18_g43943/U$1 ( \7103 , \7101 , \7102 );
nand \mul_6_18_g43638/U$1 ( \7104 , \2318 , \7103 );
nand \mul_6_18_g43152/U$1 ( \7105 , \7100 , \7104 );
not \mul_6_18_g42867/U$4 ( \7106 , \7105 );
or \mul_6_18_g42867/U$2 ( \7107 , \7096 , \7106 );
or \mul_6_18_g42867/U$5 ( \7108 , \7105 , \7095 );
nand \mul_6_18_g42867/U$1 ( \7109 , \7107 , \7108 );
xor \g45768/U$1_r1 ( \7110 , \7088 , \7109 );
xnor \g45871/U$1_r1 ( \7111 , \7072 , \7110 );
not \mul_6_18_g42545/U$1 ( \7112 , \7111 );
not \mul_6_18_g42321/U$4 ( \7113 , \7112 );
or \mul_6_18_g42321/U$2 ( \7114 , \7027 , \7113 );
nand \mul_6_18_g42346/U$1 ( \7115 , \7111 , \7025 );
nand \mul_6_18_g42321/U$1 ( \7116 , \7114 , \7115 );
xor \mul_6_18_g42704/U$4 ( \7117 , \3557 , \3566 );
and \mul_6_18_g42704/U$3 ( \7118 , \7117 , \3575 );
and \mul_6_18_g42704/U$5 ( \7119 , \3557 , \3566 );
or \mul_6_18_g42704/U$2 ( \7120 , \7118 , \7119 );
not \mul_6_18_g44038/U$1 ( \7121 , \2875 );
not \mul_6_18_g43063/U$3 ( \7122 , \7121 );
not \mul_6_18_g43063/U$4 ( \7123 , \2162 );
or \mul_6_18_g43063/U$2 ( \7124 , \7122 , \7123 );
and \mul_6_18_g44037/U$2 ( \7125 , \2006 , \2536 );
not \mul_6_18_g44037/U$4 ( \7126 , \2006 );
and \mul_6_18_g44037/U$3 ( \7127 , \7126 , \2159 );
nor \mul_6_18_g44037/U$1 ( \7128 , \7125 , \7127 );
nand \mul_6_18_g43542/U$1 ( \7129 , \7128 , \2155 );
nand \mul_6_18_g43063/U$1 ( \7130 , \7124 , \7129 );
and \mul_6_18_g43945/U$2 ( \7131 , \2117 , \2168 );
and \mul_6_18_g43945/U$3 ( \7132 , \2414 , \3154 );
nor \mul_6_18_g43945/U$1 ( \7133 , \7131 , \7132 );
not \mul_6_18_g43060/U$3 ( \7134 , \7133 );
not \mul_6_18_g43863/U$1 ( \7135 , \2129 );
not \mul_6_18_g43060/U$4 ( \7136 , \7135 );
and \mul_6_18_g43060/U$2 ( \7137 , \7134 , \7136 );
and \mul_6_18_g43060/U$5 ( \7138 , \2879 , \2886 );
nor \mul_6_18_g43060/U$1 ( \7139 , \7137 , \7138 );
xnor \g45554/U$1 ( \7140 , \7130 , \7139 );
not \mul_6_18_g43708/U$1 ( \7141 , \2511 );
or \mul_6_18_g43112/U$2 ( \7142 , \7141 , \3604 );
not \mul_6_18_g43819/U$1 ( \7143 , \2515 );
and \mul_6_18_g44035/U$2 ( \7144 , \2497 , \2092 );
and \mul_6_18_g44035/U$3 ( \7145 , \2496 , \2754 );
nor \mul_6_18_g44035/U$1 ( \7146 , \7144 , \7145 );
or \mul_6_18_g43112/U$3 ( \7147 , \7143 , \7146 );
nand \mul_6_18_g43112/U$1 ( \7148 , \7142 , \7147 );
not \mul_6_18_g43111/U$1 ( \7149 , \7148 );
and \mul_6_18_g42759/U$2 ( \7150 , \7140 , \7149 );
not \mul_6_18_g42759/U$4 ( \7151 , \7140 );
and \mul_6_18_g42759/U$3 ( \7152 , \7151 , \7148 );
nor \mul_6_18_g42759/U$1 ( \7153 , \7150 , \7152 );
xnor \g45433/U$1 ( \7154 , \7120 , \7153 );
xor \mul_6_18_g42450/U$4 ( \7155 , \2877 , \2888 );
and \mul_6_18_g42450/U$3 ( \7156 , \7155 , \2920 );
and \mul_6_18_g42450/U$5 ( \7157 , \2877 , \2888 );
or \mul_6_18_g42450/U$2 ( \7158 , \7156 , \7157 );
not \mul_6_18_g42449/U$1 ( \7159 , \7158 );
and \mul_6_18_g42353/U$2 ( \7160 , \7154 , \7159 );
not \mul_6_18_g42353/U$4 ( \7161 , \7154 );
and \mul_6_18_g42353/U$3 ( \7162 , \7161 , \7158 );
nor \mul_6_18_g42353/U$1 ( \7163 , \7160 , \7162 );
xor \mul_6_18_g45169/U$1 ( \7164 , \7116 , \7163 );
not \mul_6_18_g42154/U$4 ( \7165 , \7164 );
and \mul_6_18_g42154/U$2 ( \7166 , \7016 , \7165 );
and \mul_6_18_g42154/U$5 ( \7167 , \7015 , \7164 );
nor \mul_6_18_g42154/U$1 ( \7168 , \7166 , \7167 );
not \mul_6_18_g42153/U$1 ( \7169 , \7168 );
and \mul_6_18_g42025/U$2 ( \7170 , \7011 , \7169 );
not \mul_6_18_g42025/U$4 ( \7171 , \7011 );
and \mul_6_18_g42025/U$3 ( \7172 , \7171 , \7168 );
nor \mul_6_18_g42025/U$1 ( \7173 , \7170 , \7172 );
xor \mul_6_18_g42203/U$4 ( \7174 , \3542 , \3546 );
and \mul_6_18_g42203/U$3 ( \7175 , \7174 , \3609 );
and \mul_6_18_g42203/U$5 ( \7176 , \3542 , \3546 );
or \mul_6_18_g42203/U$2 ( \7177 , \7175 , \7176 );
or \mul_6_18_g43255/U$2 ( \7178 , \3079 , \3555 );
and \mul_6_18_g43877/U$2 ( \7179 , \2969 , \2099 );
and \mul_6_18_g43877/U$3 ( \7180 , \3083 , \2257 );
nor \mul_6_18_g43877/U$1 ( \7181 , \7179 , \7180 );
or \mul_6_18_g43255/U$3 ( \7182 , \3086 , \7181 );
nand \mul_6_18_g43255/U$1 ( \7183 , \7178 , \7182 );
not \mul_6_18_g42871/U$3 ( \7184 , \7183 );
and \mul_6_18_g43221/U$2 ( \7185 , \2400 , \2406 );
and \g45701/U$2 ( \7186 , \2364 , \2568 );
not \g45701/U$4 ( \7187 , \2364 );
and \g45701/U$3 ( \7188 , \7187 , \2105 );
nor \g45701/U$1 ( \7189 , \7186 , \7188 );
and \mul_6_18_g43221/U$3 ( \7190 , \2403 , \7189 );
nor \mul_6_18_g43221/U$1 ( \7191 , \7185 , \7190 );
not \mul_6_18_g42871/U$4 ( \7192 , \7191 );
or \mul_6_18_g42871/U$2 ( \7193 , \7184 , \7192 );
or \mul_6_18_g42871/U$5 ( \7194 , \7191 , \7183 );
nand \mul_6_18_g42871/U$1 ( \7195 , \7193 , \7194 );
not \mul_6_18_g44137/U$1 ( \7196 , \3583 );
not \mul_6_18_g43702/U$1 ( \7197 , \2482 );
or \mul_6_18_g43075/U$2 ( \7198 , \7196 , \7197 );
not \mul_6_18_g43834/U$1 ( \7199 , \2485 );
and \mul_6_18_g45276/U$2 ( \7200 , \2195 , \2112 );
not \mul_6_18_g45276/U$4 ( \7201 , \2195 );
and \mul_6_18_g45276/U$3 ( \7202 , \7201 , \2824 );
nor \mul_6_18_g45276/U$1 ( \7203 , \7200 , \7202 );
or \mul_6_18_g43075/U$3 ( \7204 , \7199 , \7203 );
nand \mul_6_18_g43075/U$1 ( \7205 , \7198 , \7204 );
nand \mul_6_18_g44168/U$1 ( \7206 , \875 , \2058 );
not \mul_6_18_g43718/U$3 ( \7207 , \2116 );
not \mul_6_18_g43718/U$4 ( \7208 , \2902 );
or \mul_6_18_g43718/U$2 ( \7209 , \7207 , \7208 );
nand \mul_6_18_g43718/U$1 ( \7210 , \7209 , \2414 );
nand \g45753/U$1 ( \7211 , \7206 , \840 , \7210 );
not \mul_6_18_g43417/U$3 ( \7212 , \2240 );
not \mul_6_18_g43417/U$4 ( \7213 , \2223 );
or \mul_6_18_g43417/U$2 ( \7214 , \7212 , \7213 );
not \mul_6_18_g43745/U$3 ( \7215 , \2236 );
not \mul_6_18_g44973/U$1 ( \7216 , \2115 );
not \mul_6_18_g43745/U$4 ( \7217 , \7216 );
or \mul_6_18_g43745/U$2 ( \7218 , \7215 , \7217 );
or \mul_6_18_g43745/U$5 ( \7219 , \2226 , \7216 );
nand \mul_6_18_g43745/U$1 ( \7220 , \7218 , \7219 );
nand \mul_6_18_g43653/U$1 ( \7221 , \7220 , \2245 );
nand \mul_6_18_g43417/U$1 ( \7222 , \7214 , \7221 );
xor \g45769/U$1 ( \7223 , \7211 , \7222 );
and \mul_6_18_g43826/U$2 ( \7224 , \2058 , \840 );
not \mul_6_18_g43826/U$4 ( \7225 , \2058 );
not \mul_6_18_g44715/U$1 ( \7226 , \840 );
and \mul_6_18_g43826/U$3 ( \7227 , \7225 , \7226 );
nor \mul_6_18_g43826/U$1 ( \7228 , \7224 , \7227 );
and \mul_6_18_g43932/U$2 ( \7229 , \875 , \840 );
not \mul_6_18_g43932/U$4 ( \7230 , \875 );
and \mul_6_18_g43932/U$3 ( \7231 , \7230 , \7226 );
nor \mul_6_18_g43932/U$1 ( \7232 , \7229 , \7231 );
nand \mul_6_18_g43486/U$1 ( \7233 , \7228 , \7232 );
or \mul_6_18_g43056/U$2 ( \7234 , \2904 , \7233 );
and \mul_6_18_g43862/U$2 ( \7235 , \2056 , \840 );
not \mul_6_18_g43862/U$4 ( \7236 , \2056 );
and \mul_6_18_g43862/U$3 ( \7237 , \7236 , \7226 );
nor \mul_6_18_g43862/U$1 ( \7238 , \7235 , \7237 );
nand \mul_6_18_g43600/U$1 ( \7239 , \2904 , \7238 );
nand \mul_6_18_g43056/U$1 ( \7240 , \7234 , \7239 );
xnor \g45769/U$1_r1 ( \7241 , \7223 , \7240 );
xnor \g45452/U$1 ( \7242 , \7205 , \7241 );
xor \g45613/U$1 ( \7243 , \7195 , \7242 );
xor \mul_6_18_g42650/U$4 ( \7244 , \2248 , \2287 );
and \mul_6_18_g42650/U$3 ( \7245 , \7244 , \2325 );
and \mul_6_18_g42650/U$5 ( \7246 , \2248 , \2287 );
or \mul_6_18_g42650/U$2 ( \7247 , \7245 , \7246 );
xor \mul_6_18_g42583/U$4 ( \7248 , \2899 , \2905 );
and \mul_6_18_g42583/U$3 ( \7249 , \7248 , \2919 );
and \mul_6_18_g42583/U$5 ( \7250 , \2899 , \2905 );
or \mul_6_18_g42583/U$2 ( \7251 , \7249 , \7250 );
xor \mul_6_18_g45189/U$1 ( \7252 , \7247 , \7251 );
xor \g45613/U$1_r1 ( \7253 , \7243 , \7252 );
not \mul_6_18_g42294/U$3 ( \7254 , \7253 );
xor \mul_6_18_g42374/U$4 ( \7255 , \3551 , \3576 );
and \mul_6_18_g42374/U$3 ( \7256 , \7255 , \3608 );
and \mul_6_18_g42374/U$5 ( \7257 , \3551 , \3576 );
or \mul_6_18_g42374/U$2 ( \7258 , \7256 , \7257 );
not \mul_6_18_g42294/U$4 ( \7259 , \7258 );
and \mul_6_18_g42294/U$2 ( \7260 , \7254 , \7259 );
and \mul_6_18_g42294/U$5 ( \7261 , \7258 , \7253 );
nor \mul_6_18_g42294/U$1 ( \7262 , \7260 , \7261 );
xor \g45731/U$1 ( \7263 , \7177 , \7262 );
xor \mul_6_18_g42373/U$4 ( \7264 , \2215 , \2326 );
and \mul_6_18_g42373/U$3 ( \7265 , \7264 , \2458 );
and \mul_6_18_g42373/U$5 ( \7266 , \2215 , \2326 );
or \mul_6_18_g42373/U$2 ( \7267 , \7265 , \7266 );
xor \mul_6_18_g42372/U$4 ( \7268 , \3028 , \3061 );
and \mul_6_18_g42372/U$3 ( \7269 , \7268 , \3091 );
and \mul_6_18_g42372/U$5 ( \7270 , \3028 , \3061 );
or \mul_6_18_g42372/U$2 ( \7271 , \7269 , \7270 );
xnor \mul_6_18_g45172/U$1 ( \7272 , \7267 , \7271 );
xor \g45731/U$1_r1 ( \7273 , \7263 , \7272 );
and \mul_6_18_g41987/U$2 ( \7274 , \7173 , \7273 );
not \mul_6_18_g41987/U$4 ( \7275 , \7173 );
not \mul_6_18_g42155/U$1 ( \7276 , \7273 );
and \mul_6_18_g41987/U$3 ( \7277 , \7275 , \7276 );
nor \mul_6_18_g41987/U$1 ( \7278 , \7274 , \7277 );
xor \mul_6_18_g42027/U$4 ( \7279 , \3509 , \3610 );
and \mul_6_18_g42027/U$3 ( \7280 , \7279 , \3700 );
and \mul_6_18_g42027/U$5 ( \7281 , \3509 , \3610 );
or \mul_6_18_g42027/U$2 ( \7282 , \7280 , \7281 );
not \mul_6_18_g42026/U$1 ( \7283 , \7282 );
and \mul_6_18_g41945/U$2 ( \7284 , \7278 , \7283 );
not \mul_6_18_g41945/U$4 ( \7285 , \7278 );
and \mul_6_18_g41945/U$3 ( \7286 , \7285 , \7282 );
nor \mul_6_18_g41945/U$1 ( \7287 , \7284 , \7286 );
not \mul_6_18_g41944/U$1 ( \7288 , \7287 );
and \mul_6_18_g41866/U$2 ( \7289 , \7007 , \7288 );
not \mul_6_18_g41866/U$4 ( \7290 , \7007 );
and \mul_6_18_g41866/U$3 ( \7291 , \7290 , \7287 );
nor \mul_6_18_g41866/U$1 ( \7292 , \7289 , \7291 );
and \mul_6_18_g41832/U$2 ( \7293 , \7003 , \7292 );
not \mul_6_18_g41832/U$4 ( \7294 , \7003 );
not \mul_6_18_g41865/U$1 ( \7295 , \7292 );
and \mul_6_18_g41832/U$3 ( \7296 , \7294 , \7295 );
nor \mul_6_18_g41832/U$1 ( \7297 , \7293 , \7296 );
not \mul_6_18_g41903/U$1 ( \7298 , \4198 );
not \mul_6_18_g41835/U$3 ( \7299 , \7298 );
not \mul_6_18_g41835/U$4 ( \7300 , \6987 );
or \mul_6_18_g41835/U$2 ( \7301 , \7299 , \7300 );
not \mul_6_18_g41881/U$1 ( \7302 , \6999 );
nand \mul_6_18_g41835/U$1 ( \7303 , \7301 , \7302 );
not \mul_6_18_g41861/U$2 ( \7304 , \7001 );
nand \mul_6_18_g41861/U$1 ( \7305 , \7304 , \6990 );
not \mul_6_18_g41860/U$1 ( \7306 , \7305 );
and \mul_6_18_g41833/U$2 ( \7307 , \7303 , \7306 );
not \mul_6_18_g41833/U$4 ( \7308 , \7303 );
and \mul_6_18_g41833/U$3 ( \7309 , \7308 , \7305 );
nor \mul_6_18_g41833/U$1 ( \7310 , \7307 , \7309 );
buf \mul_6_18_g41919/U$1 ( \7311 , \4197 );
not \mul_6_18_g41836/U$3 ( \7312 , \7311 );
not \mul_6_18_g41836/U$4 ( \7313 , \6987 );
or \mul_6_18_g41836/U$2 ( \7314 , \7312 , \7313 );
buf \mul_6_18_g41923/U$1 ( \7315 , \6994 );
nand \mul_6_18_g41836/U$1 ( \7316 , \7314 , \7315 );
not \mul_6_18_g45149/U$2 ( \7317 , \6991 );
nand \mul_6_18_g45149/U$1 ( \7318 , \7317 , \6998 );
not \mul_6_18_g41911/U$1 ( \7319 , \7318 );
and \mul_6_18_g41834/U$2 ( \7320 , \7316 , \7319 );
not \mul_6_18_g41834/U$4 ( \7321 , \7316 );
and \mul_6_18_g41834/U$3 ( \7322 , \7321 , \7318 );
nor \mul_6_18_g41834/U$1 ( \7323 , \7320 , \7322 );
buf \fopt/U$1 ( \7324 , \6987 );
nand \mul_6_18_g41890/U$1 ( \7325 , \7315 , \7311 );
not \mul_6_18_g41889/U$1 ( \7326 , \7325 );
and \mul_6_18_g41838/U$2 ( \7327 , \7324 , \7326 );
not \mul_6_18_g41838/U$4 ( \7328 , \7324 );
and \mul_6_18_g41838/U$3 ( \7329 , \7328 , \7325 );
nor \mul_6_18_g41838/U$1 ( \7330 , \7327 , \7329 );
not \mul_6_18_g41845/U$3 ( \7331 , \6984 );
not \mul_6_18_g41845/U$4 ( \7332 , \6979 );
or \mul_6_18_g41845/U$2 ( \7333 , \7331 , \7332 );
nand \mul_6_18_g41845/U$1 ( \7334 , \7333 , \4962 );
nand \mul_6_18_g41892/U$1 ( \7335 , \4423 , \4965 );
not \mul_6_18_g41891/U$1 ( \7336 , \7335 );
and \mul_6_18_g41839/U$2 ( \7337 , \7334 , \7336 );
not \mul_6_18_g41839/U$4 ( \7338 , \7334 );
and \mul_6_18_g41839/U$3 ( \7339 , \7338 , \7335 );
nor \mul_6_18_g41839/U$1 ( \7340 , \7337 , \7339 );
not \mul_6_18_g41874/U$1 ( \7341 , \6983 );
not \mul_6_18_g41843/U$3 ( \7342 , \7341 );
not \mul_6_18_g41843/U$4 ( \7343 , \6979 );
or \mul_6_18_g41843/U$2 ( \7344 , \7342 , \7343 );
nand \mul_6_18_g41843/U$1 ( \7345 , \7344 , \4958 );
not \mul_6_18_g45148/U$2 ( \7346 , \4671 );
nand \mul_6_18_g45148/U$1 ( \7347 , \7346 , \4960 );
not \mul_6_18_g41867/U$1 ( \7348 , \7347 );
and \mul_6_18_g41840/U$2 ( \7349 , \7345 , \7348 );
not \mul_6_18_g41840/U$4 ( \7350 , \7345 );
and \mul_6_18_g41840/U$3 ( \7351 , \7350 , \7347 );
nor \mul_6_18_g41840/U$1 ( \7352 , \7349 , \7351 );
buf \mul_6_18_fopt45086/U$1 ( \7353 , \6982 );
not \mul_6_18_g41844/U$3 ( \7354 , \7353 );
not \mul_6_18_g41844/U$4 ( \7355 , \6979 );
or \mul_6_18_g41844/U$2 ( \7356 , \7354 , \7355 );
buf \mul_6_18_g41914/U$1 ( \7357 , \4946 );
nand \mul_6_18_g41844/U$1 ( \7358 , \7356 , \7357 );
nand \mul_6_18_g41870/U$1 ( \7359 , \4953 , \4957 );
not \mul_6_18_g41869/U$1 ( \7360 , \7359 );
and \mul_6_18_g41841/U$2 ( \7361 , \7358 , \7360 );
not \mul_6_18_g41841/U$4 ( \7362 , \7358 );
and \mul_6_18_g41841/U$3 ( \7363 , \7362 , \7359 );
nor \mul_6_18_g41841/U$1 ( \7364 , \7361 , \7363 );
buf \fopt45636/U$1 ( \7365 , \6979 );
nand \mul_6_18_g41894/U$1 ( \7366 , \7353 , \7357 );
not \mul_6_18_g41893/U$1 ( \7367 , \7366 );
and \mul_6_18_g41846/U$2 ( \7368 , \7365 , \7367 );
not \mul_6_18_g41846/U$4 ( \7369 , \7365 );
and \mul_6_18_g41846/U$3 ( \7370 , \7369 , \7366 );
nor \mul_6_18_g41846/U$1 ( \7371 , \7368 , \7370 );
not \mul_6_18_g41886/U$3 ( \7372 , \6753 );
not \mul_6_18_g41925/U$3 ( \7373 , \6929 );
not \mul_6_18_g41925/U$4 ( \7374 , \6220 );
or \mul_6_18_g41925/U$2 ( \7375 , \7373 , \7374 );
not \g45356/U$2 ( \7376 , \6963 );
nand \g45356/U$1 ( \7377 , \7376 , \6962 );
nand \mul_6_18_g41925/U$1 ( \7378 , \7375 , \7377 );
not \mul_6_18_g41886/U$4 ( \7379 , \7378 );
or \mul_6_18_g41886/U$2 ( \7380 , \7372 , \7379 );
not \mul_6_18_g41978/U$1 ( \7381 , \6967 );
and \mul_6_18_g41932/U$1 ( \7382 , \6970 , \7381 );
nand \mul_6_18_g41886/U$1 ( \7383 , \7380 , \7382 );
buf \mul_6_18_g41965/U$1 ( \7384 , \6948 );
and \mul_6_18_g41855/U$2 ( \7385 , \7383 , \7384 );
buf \mul_6_18_g41961/U$1 ( \7386 , \6966 );
nor \mul_6_18_g41855/U$1 ( \7387 , \7385 , \7386 );
nand \mul_6_18_g41896/U$1 ( \7388 , \6784 , \6971 );
and \mul_6_18_g41849/U$2 ( \7389 , \7387 , \7388 );
not \mul_6_18_g41849/U$4 ( \7390 , \7387 );
not \mul_6_18_g41895/U$1 ( \7391 , \7388 );
and \mul_6_18_g41849/U$3 ( \7392 , \7390 , \7391 );
nor \mul_6_18_g41849/U$1 ( \7393 , \7389 , \7392 );
not \mul_6_18_g45150/U$2 ( \7394 , \7386 );
nand \mul_6_18_g45150/U$1 ( \7395 , \7394 , \7384 );
not \mul_6_18_g41933/U$1 ( \7396 , \7395 );
and \mul_6_18_g41857/U$2 ( \7397 , \7383 , \7396 );
not \mul_6_18_g41857/U$4 ( \7398 , \7383 );
and \mul_6_18_g41857/U$3 ( \7399 , \7398 , \7395 );
nor \mul_6_18_g41857/U$1 ( \7400 , \7397 , \7399 );
not \mul_6_18_g41877/U$3 ( \7401 , \6752 );
not \mul_6_18_g41877/U$4 ( \7402 , \7378 );
or \mul_6_18_g41877/U$2 ( \7403 , \7401 , \7402 );
not \mul_6_18_g41980/U$1 ( \7404 , \6969 );
nand \mul_6_18_g41877/U$1 ( \7405 , \7403 , \7404 );
nand \mul_6_18_g41956/U$1 ( \7406 , \6710 , \7381 );
not \mul_6_18_g41955/U$1 ( \7407 , \7406 );
and \mul_6_18_g41858/U$2 ( \7408 , \7405 , \7407 );
not \mul_6_18_g41858/U$4 ( \7409 , \7405 );
and \mul_6_18_g41858/U$3 ( \7410 , \7409 , \7406 );
nor \mul_6_18_g41858/U$1 ( \7411 , \7408 , \7410 );
not \mul_6_18_g41972/U$2 ( \7412 , \6952 );
nor \mul_6_18_g41972/U$1 ( \7413 , \7412 , \6963 );
buf \mul_6_18_g42016/U$1 ( \7414 , \6928 );
not \mul_6_18_g41879/U$3 ( \7415 , \7414 );
not \mul_6_18_g41928/U$3 ( \7416 , \6890 );
not \mul_6_18_g41928/U$4 ( \7417 , \6220 );
or \mul_6_18_g41928/U$2 ( \7418 , \7416 , \7417 );
nand \mul_6_18_g41993/U$1 ( \7419 , \6959 , \6960 );
nand \mul_6_18_g41928/U$1 ( \7420 , \7418 , \7419 );
not \mul_6_18_g41879/U$4 ( \7421 , \7420 );
or \mul_6_18_g41879/U$2 ( \7422 , \7415 , \7421 );
buf \mul_6_18_g42013/U$1 ( \7423 , \6953 );
nand \mul_6_18_g41879/U$1 ( \7424 , \7422 , \7423 );
and \mul_6_18_g41859/U$2 ( \7425 , \7413 , \7424 );
not \mul_6_18_g41859/U$4 ( \7426 , \7413 );
not \mul_6_18_g41878/U$1 ( \7427 , \7424 );
and \mul_6_18_g41859/U$3 ( \7428 , \7426 , \7427 );
nor \mul_6_18_g41859/U$1 ( \7429 , \7425 , \7428 );
nand \mul_6_18_g41957/U$1 ( \7430 , \7404 , \6752 );
not \mul_6_18_g41883/U$3 ( \7431 , \7430 );
not \mul_6_18_g41883/U$4 ( \7432 , \7378 );
or \mul_6_18_g41883/U$2 ( \7433 , \7431 , \7432 );
or \mul_6_18_g41883/U$5 ( \7434 , \7430 , \7378 );
nand \mul_6_18_g41883/U$1 ( \7435 , \7433 , \7434 );
nand \mul_6_18_g41995/U$1 ( \7436 , \7423 , \7414 );
not \mul_6_18_g41994/U$1 ( \7437 , \7436 );
and \mul_6_18_g41884/U$2 ( \7438 , \7420 , \7437 );
not \mul_6_18_g41884/U$4 ( \7439 , \7420 );
and \mul_6_18_g41884/U$3 ( \7440 , \7439 , \7436 );
nor \mul_6_18_g41884/U$1 ( \7441 , \7438 , \7440 );
not \mul_6_18_g41926/U$3 ( \7442 , \6889 );
not \mul_6_18_g41926/U$4 ( \7443 , \6220 );
or \mul_6_18_g41926/U$2 ( \7444 , \7442 , \7443 );
buf \mul_6_18_fopt45083/U$1 ( \7445 , \6958 );
nand \mul_6_18_g41926/U$1 ( \7446 , \7444 , \7445 );
nand \mul_6_18_g42009/U$1 ( \7447 , \6956 , \6960 );
not \mul_6_18_g42008/U$1 ( \7448 , \7447 );
and \mul_6_18_g41885/U$2 ( \7449 , \7446 , \7448 );
not \mul_6_18_g41885/U$4 ( \7450 , \7446 );
and \mul_6_18_g41885/U$3 ( \7451 , \7450 , \7447 );
nor \mul_6_18_g41885/U$1 ( \7452 , \7449 , \7451 );
not \mul_6_18_g41940/U$3 ( \7453 , \5554 );
not \mul_6_18_g45152/U$2 ( \7454 , \6205 );
nand \mul_6_18_g42090/U$1 ( \7455 , \6210 , \6211 );
nand \mul_6_18_g45152/U$1 ( \7456 , \7454 , \7455 );
not \mul_6_18_g41940/U$4 ( \7457 , \7456 );
or \mul_6_18_g41940/U$2 ( \7458 , \7453 , \7457 );
nand \mul_6_18_g41940/U$1 ( \7459 , \7458 , \6215 );
nand \mul_6_18_g42032/U$1 ( \7460 , \6216 , \5496 );
not \mul_6_18_g42031/U$1 ( \7461 , \7460 );
and \mul_6_18_g41909/U$2 ( \7462 , \7459 , \7461 );
not \mul_6_18_g41909/U$4 ( \7463 , \7459 );
and \mul_6_18_g41909/U$3 ( \7464 , \7463 , \7460 );
nor \mul_6_18_g41909/U$1 ( \7465 , \7462 , \7464 );
nand \mul_6_18_g42033/U$1 ( \7466 , \7445 , \6889 );
not \mul_6_18_g41929/U$3 ( \7467 , \7466 );
not \mul_6_18_g41929/U$4 ( \7468 , \6220 );
or \mul_6_18_g41929/U$2 ( \7469 , \7467 , \7468 );
or \mul_6_18_g41929/U$5 ( \7470 , \7466 , \6220 );
nand \mul_6_18_g41929/U$1 ( \7471 , \7469 , \7470 );
nand \mul_6_18_g42073/U$1 ( \7472 , \5554 , \6215 );
not \mul_6_18_g42072/U$1 ( \7473 , \7472 );
and \mul_6_18_g41942/U$2 ( \7474 , \7456 , \7473 );
not \mul_6_18_g41942/U$4 ( \7475 , \7456 );
and \mul_6_18_g41942/U$3 ( \7476 , \7475 , \7472 );
nor \mul_6_18_g41942/U$1 ( \7477 , \7474 , \7476 );
not \mul_6_18_g42141/U$1 ( \7478 , \6203 );
not \mul_6_18_g41983/U$3 ( \7479 , \7478 );
buf \mul_6_18_g42020/U$1 ( \7480 , \6155 );
not \mul_6_18_g41983/U$4 ( \7481 , \7480 );
or \mul_6_18_g41983/U$2 ( \7482 , \7479 , \7481 );
buf \mul_6_18_g42149/U$1 ( \7483 , \6209 );
nand \mul_6_18_g41983/U$1 ( \7484 , \7482 , \7483 );
nand \mul_6_18_g42115/U$1 ( \7485 , \6208 , \6211 );
not \mul_6_18_g42114/U$1 ( \7486 , \7485 );
and \mul_6_18_g41943/U$2 ( \7487 , \7484 , \7486 );
not \mul_6_18_g41943/U$4 ( \7488 , \7484 );
and \mul_6_18_g41943/U$3 ( \7489 , \7488 , \7485 );
nor \mul_6_18_g41943/U$1 ( \7490 , \7487 , \7489 );
nand \mul_6_18_g42117/U$1 ( \7491 , \7483 , \7478 );
not \mul_6_18_g42116/U$1 ( \7492 , \7491 );
and \mul_6_18_g41985/U$2 ( \7493 , \7480 , \7492 );
not \mul_6_18_g41985/U$4 ( \7494 , \7480 );
and \mul_6_18_g41985/U$3 ( \7495 , \7494 , \7491 );
nor \mul_6_18_g41985/U$1 ( \7496 , \7493 , \7495 );
not \mul_6_18_g42022/U$3 ( \7497 , \5829 );
buf \mul_6_18_g42061/U$1 ( \7498 , \6148 );
not \mul_6_18_g42022/U$4 ( \7499 , \7498 );
or \mul_6_18_g42022/U$2 ( \7500 , \7497 , \7499 );
not \mul_6_18_g42183/U$1 ( \7501 , \6151 );
nand \mul_6_18_g42022/U$1 ( \7502 , \7500 , \7501 );
not \mul_6_18_g42119/U$2 ( \7503 , \6153 );
nand \mul_6_18_g42119/U$1 ( \7504 , \7503 , \5764 );
not \mul_6_18_g42118/U$1 ( \7505 , \7504 );
and \mul_6_18_g41986/U$2 ( \7506 , \7502 , \7505 );
not \mul_6_18_g41986/U$4 ( \7507 , \7502 );
and \mul_6_18_g41986/U$3 ( \7508 , \7507 , \7504 );
nor \mul_6_18_g41986/U$1 ( \7509 , \7506 , \7508 );
buf \mul_6_18_g42106/U$1 ( \7510 , \6111 );
and \mul_6_18_g42064/U$2 ( \7511 , \7510 , \6142 );
nor \mul_6_18_g42064/U$1 ( \7512 , \7511 , \6144 );
xor \mul_6_18_g42107/U$1 ( \7513 , \5900 , \5941 );
xor \mul_6_18_g42107/U$1_r1 ( \7514 , \7513 , \6108 );
nand \mul_6_18_g42166/U$1 ( \7515 , \7501 , \5829 );
not \mul_6_18_g42240/U$2 ( \7516 , \6146 );
nand \mul_6_18_g42240/U$1 ( \7517 , \7516 , \6130 );
nand \mul_6_18_g42342/U$1 ( \7518 , \6107 , \6104 );
nand \mul_6_18_g42510/U$1 ( \7519 , \6045 , \6042 );
and \mul_6_18_g42588/U$1 ( \7520 , \6018 , \5981 );
not \mul_6_18_g42838/U$2 ( \7521 , \6009 );
nand \mul_6_18_g42838/U$1 ( \7522 , \7521 , \6012 );
or \mul_6_18_g42915/U$2 ( \7523 , \5996 , \5998 );
nand \mul_6_18_g42915/U$1 ( \7524 , \7523 , \5999 );
not \mul_6_18_g42914/U$1 ( \7525 , \7524 );
not \mul_6_18_g44270/U$1 ( \7526 , \5997 );
not \mul_6_18_g45166/U$2 ( \7527 , \6144 );
nand \mul_6_18_g45166/U$1 ( \7528 , \7527 , \6142 );
xnor \mul_6_18_g45154/U$1 ( \7529 , \7510 , \7528 );
xor \mul_6_18_g45160/U$1 ( \7530 , \7512 , \7517 );
xnor \mul_6_18_g45161/U$1 ( \7531 , \6087 , \7518 );
and \mul_6_18_g45182/U$1 ( \7532 , \6086 , \6083 );
xor \mul_6_18_g45171/U$1 ( \7533 , \7532 , \6046 );
xnor \mul_6_18_g45181/U$1 ( \7534 , \7519 , \6019 );
xor \mul_6_18_g45195/U$1 ( \7535 , \7520 , \6013 );
xor \mul_6_18_g45204/U$1 ( \7536 , \7522 , \5999 );
not \mul_6_18_g45296/U$2 ( \7537 , \7515 );
xor \mul_6_18_g45296/U$1 ( \7538 , \7498 , \7537 );
endmodule

