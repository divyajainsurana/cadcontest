//
// Conformal-LEC Version 19.20-d255 (16-Apr-2020)
//
module top(\a[15] ,\a[14] ,\a[13] ,\a[12] ,\a[11] ,\a[10] ,\a[9] ,\a[8] ,\a[7] ,
        \a[6] ,\a[5] ,\a[4] ,\a[3] ,\a[2] ,\a[1] ,\a[0] ,\b[15] ,\b[14] ,\b[13] ,
        \b[12] ,\b[11] ,\b[10] ,\b[9] ,\b[8] ,\b[7] ,\b[6] ,\b[5] ,\b[4] ,\b[3] ,
        \b[2] ,\b[1] ,\b[0] ,\c[15] ,\c[14] ,\c[13] ,\c[12] ,\c[11] ,\c[10] ,\c[9] ,
        \c[8] ,\c[7] ,\c[6] ,\c[5] ,\c[4] ,\c[3] ,\c[2] ,\c[1] ,\c[0] ,\d[15] ,
        \d[14] ,\d[13] ,\d[12] ,\d[11] ,\d[10] ,\d[9] ,\d[8] ,\d[7] ,\d[6] ,\d[5] ,
        \d[4] ,\d[3] ,\d[2] ,\d[1] ,\d[0] ,\o[31] ,\o[30] ,\o[29] ,\o[28] ,\o[27] ,
        \o[26] ,\o[25] ,\o[24] ,\o[23] ,\o[22] ,\o[21] ,\o[20] ,\o[19] ,\o[18] ,\o[17] ,
        \o[16] ,\o[15] ,\o[14] ,\o[13] ,\o[12] ,\o[11] ,\o[10] ,\o[9] ,\o[8] ,\o[7] ,
        \o[6] ,\o[5] ,\o[4] ,\o[3] ,\o[2] ,\o[1] ,\o[0] );
input \a[15] ,\a[14] ,\a[13] ,\a[12] ,\a[11] ,\a[10] ,\a[9] ,\a[8] ,\a[7] ,
        \a[6] ,\a[5] ,\a[4] ,\a[3] ,\a[2] ,\a[1] ,\a[0] ,\b[15] ,\b[14] ,\b[13] ,
        \b[12] ,\b[11] ,\b[10] ,\b[9] ,\b[8] ,\b[7] ,\b[6] ,\b[5] ,\b[4] ,\b[3] ,
        \b[2] ,\b[1] ,\b[0] ,\c[15] ,\c[14] ,\c[13] ,\c[12] ,\c[11] ,\c[10] ,\c[9] ,
        \c[8] ,\c[7] ,\c[6] ,\c[5] ,\c[4] ,\c[3] ,\c[2] ,\c[1] ,\c[0] ,\d[15] ,
        \d[14] ,\d[13] ,\d[12] ,\d[11] ,\d[10] ,\d[9] ,\d[8] ,\d[7] ,\d[6] ,\d[5] ,
        \d[4] ,\d[3] ,\d[2] ,\d[1] ,\d[0] ;
output \o[31] ,\o[30] ,\o[29] ,\o[28] ,\o[27] ,\o[26] ,\o[25] ,\o[24] ,\o[23] ,
        \o[22] ,\o[21] ,\o[20] ,\o[19] ,\o[18] ,\o[17] ,\o[16] ,\o[15] ,\o[14] ,\o[13] ,
        \o[12] ,\o[11] ,\o[10] ,\o[9] ,\o[8] ,\o[7] ,\o[6] ,\o[5] ,\o[4] ,\o[3] ,
        \o[2] ,\o[1] ,\o[0] ;

wire \97_ZERO , \98_ONE , \99 , \100 , \101 , \102 , \103 , \104 , \105 ,
         \106 , \107 , \108 , \109 , \110 , \111 , \112 , \113 , \114 , \115 ,
         \116 , \117 , \118 , \119 , \120 , \121 , \122 , \123 , \124 , \125 ,
         \126 , \127 , \128 , \129 , \130 , \131 , \132 , \133 , \134 , \135 ,
         \136 , \137 , \138 , \139 , \140 , \141 , \142 , \143 , \144 , \145 ,
         \146 , \147 , \148 , \149 , \150 , \151 , \152 , \153 , \154 , \155 ,
         \156 , \157 , \158 , \159 , \160 , \161 , \162 , \163 , \164 , \165 ,
         \166 , \167 , \168 , \169 , \170 , \171 , \172 , \173 , \174 , \175 ,
         \176 , \177 , \178 , \179 , \180 , \181 , \182 , \183 , \184 , \185 ,
         \186 , \187 , \188 , \189 , \190 , \191 , \192 , \193 , \194 , \195 ,
         \196 , \197 , \198 , \199 , \200 , \201 , \202 , \203 , \204 , \205 ,
         \206 , \207 , \208 , \209 , \210 , \211 , \212 , \213 , \214 , \215 ,
         \216 , \217 , \218 , \219 , \220 , \221 , \222 , \223 , \224 , \225 ,
         \226 , \227 , \228 , \229 , \230 , \231 , \232 , \233 , \234 , \235 ,
         \236 , \237 , \238 , \239 , \240 , \241 , \242 , \243 , \244 , \245 ,
         \246 , \247 , \248 , \249 , \250 , \251 , \252 , \253 , \254 , \255 ,
         \256 , \257 , \258 , \259 , \260 , \261 , \262 , \263 , \264 , \265 ,
         \266 , \267 , \268 , \269 , \270 , \271 , \272 , \273 , \274 , \275 ,
         \276 , \277 , \278 , \279 , \280 , \281 , \282 , \283 , \284 , \285 ,
         \286 , \287 , \288 , \289 , \290 , \291 , \292 , \293 , \294 , \295 ,
         \296 , \297 , \298 , \299 , \300 , \301 , \302 , \303 , \304 , \305 ,
         \306 , \307 , \308 , \309 , \310 , \311 , \312 , \313 , \314 , \315 ,
         \316 , \317 , \318 , \319 , \320 , \321 , \322 , \323 , \324 , \325 ,
         \326 , \327 , \328 , \329 , \330 , \331 , \332 , \333 , \334 , \335 ,
         \336 , \337 , \338 , \339 , \340 , \341 , \342 , \343 , \344 , \345 ,
         \346 , \347 , \348 , \349 , \350 , \351 , \352 , \353 , \354 , \355 ,
         \356 , \357 , \358 , \359 , \360 , \361 , \362 , \363 , \364 , \365 ,
         \366 , \367 , \368 , \369 , \370 , \371 , \372 , \373 , \374 , \375 ,
         \376 , \377 , \378 , \379 , \380 , \381 , \382 , \383 , \384 , \385 ,
         \386 , \387 , \388 , \389 , \390 , \391 , \392 , \393 , \394 , \395 ,
         \396 , \397 , \398 , \399 , \400 , \401 , \402 , \403 , \404 , \405 ,
         \406 , \407 , \408 , \409 , \410 , \411 , \412 , \413 , \414 , \415 ,
         \416 , \417 , \418 , \419 , \420 , \421 , \422 , \423 , \424 , \425 ,
         \426 , \427 , \428 , \429 , \430 , \431 , \432 , \433 , \434 , \435 ,
         \436 , \437 , \438 , \439 , \440 , \441 , \442 , \443 , \444 , \445 ,
         \446 , \447 , \448 , \449 , \450 , \451 , \452 , \453 , \454 , \455 ,
         \456 , \457 , \458 , \459 , \460 , \461 , \462 , \463 , \464 , \465 ,
         \466 , \467 , \468 , \469 , \470 , \471 , \472 , \473 , \474 , \475 ,
         \476 , \477 , \478 , \479 , \480 , \481 , \482 , \483 , \484 , \485 ,
         \486 , \487 , \488 , \489 , \490 , \491 , \492 , \493 , \494 , \495 ,
         \496 , \497 , \498 , \499 , \500 , \501 , \502 , \503 , \504 , \505 ,
         \506 , \507 , \508 , \509 , \510 , \511 , \512 , \513 , \514 , \515 ,
         \516 , \517 , \518 , \519 , \520 , \521 , \522 , \523 , \524 , \525 ,
         \526 , \527 , \528 , \529 , \530 , \531 , \532 , \533 , \534 , \535 ,
         \536 , \537 , \538 , \539 , \540 , \541 , \542 , \543 , \544 , \545 ,
         \546 , \547 , \548 , \549 , \550 , \551 , \552 , \553 , \554 , \555 ,
         \556 , \557 , \558 , \559 , \560 , \561 , \562 , \563 , \564 , \565 ,
         \566 , \567 , \568 , \569 , \570 , \571 , \572 , \573 , \574 , \575 ,
         \576 , \577 , \578 , \579 , \580 , \581 , \582 , \583 , \584 , \585 ,
         \586 , \587 , \588 , \589 , \590 , \591 , \592 , \593 , \594 , \595 ,
         \596 , \597 , \598 , \599 , \600 , \601 , \602 , \603 , \604 , \605 ,
         \606 , \607 , \608 , \609 , \610 , \611 , \612 , \613 , \614 , \615 ,
         \616 , \617 , \618 , \619 , \620 , \621 , \622 , \623 , \624 , \625 ,
         \626 , \627 , \628 , \629 , \630 , \631 , \632 , \633 , \634 , \635 ,
         \636 , \637 , \638 , \639 , \640 , \641 , \642 , \643 , \644 , \645 ,
         \646 , \647 , \648 , \649 , \650 , \651 , \652 , \653 , \654 , \655 ,
         \656 , \657 , \658 , \659 , \660 , \661 , \662 , \663 , \664 , \665 ,
         \666 , \667 , \668 , \669 , \670 , \671 , \672 , \673 , \674 , \675 ,
         \676 , \677 , \678 , \679 , \680 , \681 , \682 , \683 , \684 , \685 ,
         \686 , \687 , \688 , \689 , \690 , \691 , \692 , \693 , \694 , \695 ,
         \696 , \697 , \698 , \699 , \700 , \701 , \702 , \703 , \704 , \705 ,
         \706 , \707 , \708 , \709 , \710 , \711 , \712 , \713 , \714 , \715 ,
         \716 , \717 , \718 , \719 , \720 , \721 , \722 , \723 , \724 , \725 ,
         \726 , \727 , \728 , \729 , \730 , \731 , \732 , \733 , \734 , \735 ,
         \736 , \737 , \738 , \739 , \740 , \741 , \742 , \743 , \744 , \745 ,
         \746 , \747 , \748 , \749 , \750 , \751 , \752 , \753 , \754 , \755 ,
         \756 , \757 , \758 , \759 , \760 , \761 , \762 , \763 , \764 , \765 ,
         \766 , \767 , \768 , \769 , \770 , \771 , \772 , \773 , \774 , \775 ,
         \776 , \777 , \778 , \779 , \780 , \781 , \782 , \783 , \784 , \785 ,
         \786 , \787 , \788 , \789 , \790 , \791 , \792 , \793 , \794 , \795 ,
         \796 , \797 , \798 , \799 , \800 , \801 , \802 , \803 , \804 , \805 ,
         \806 , \807 , \808 , \809 , \810 , \811 , \812 , \813 , \814 , \815 ,
         \816 , \817 , \818 , \819 , \820 , \821 , \822 , \823 , \824 , \825 ,
         \826 , \827 , \828 , \829 , \830 , \831 , \832 , \833 , \834 , \835 ,
         \836 , \837 , \838 , \839 , \840 , \841 , \842 , \843 , \844 , \845 ,
         \846 , \847 , \848 , \849 , \850 , \851 , \852 , \853 , \854 , \855 ,
         \856 , \857 , \858 , \859 , \860 , \861 , \862 , \863 , \864 , \865 ,
         \866 , \867 , \868 , \869 , \870 , \871 , \872 , \873 , \874 , \875 ,
         \876 , \877 , \878 , \879 , \880 , \881 , \882 , \883 , \884 , \885 ,
         \886 , \887 , \888 , \889 , \890 , \891 , \892 , \893 , \894 , \895 ,
         \896 , \897 , \898 , \899 , \900 , \901 , \902 , \903 , \904 , \905 ,
         \906 , \907 , \908 , \909 , \910 , \911 , \912 , \913 , \914 , \915 ,
         \916 , \917 , \918 , \919 , \920 , \921 , \922 , \923 , \924 , \925 ,
         \926 , \927 , \928 , \929 , \930 , \931 , \932 , \933 , \934 , \935 ,
         \936 , \937 , \938 , \939 , \940 , \941 , \942 , \943 , \944 , \945 ,
         \946 , \947 , \948 , \949 , \950 , \951 , \952 , \953 , \954 , \955 ,
         \956 , \957 , \958 , \959 , \960 , \961 , \962 , \963 , \964 , \965 ,
         \966 , \967 , \968 , \969 , \970 , \971 , \972 , \973 , \974 , \975 ,
         \976 , \977 , \978 , \979 , \980 , \981 , \982 , \983 , \984 , \985 ,
         \986 , \987 , \988 , \989 , \990 , \991 , \992 , \993 , \994 , \995 ,
         \996 , \997 , \998 , \999 , \1000 , \1001 , \1002 , \1003 , \1004 , \1005 ,
         \1006 , \1007 , \1008 , \1009 , \1010 , \1011 , \1012 , \1013 , \1014 , \1015 ,
         \1016 , \1017 , \1018 , \1019 , \1020 , \1021 , \1022 , \1023 , \1024 , \1025 ,
         \1026 , \1027 , \1028 , \1029 , \1030 , \1031 , \1032 , \1033 , \1034 , \1035 ,
         \1036 , \1037 , \1038 , \1039 , \1040 , \1041 , \1042 , \1043 , \1044 , \1045 ,
         \1046 , \1047 , \1048 , \1049 , \1050 , \1051 , \1052 , \1053 , \1054 , \1055 ,
         \1056 , \1057 , \1058 , \1059 , \1060 , \1061 , \1062 , \1063 , \1064 , \1065 ,
         \1066 , \1067 , \1068 , \1069 , \1070 , \1071 , \1072 , \1073 , \1074 , \1075 ,
         \1076 , \1077 , \1078 , \1079 , \1080 , \1081 , \1082 , \1083 , \1084 , \1085 ,
         \1086 , \1087 , \1088 , \1089 , \1090 , \1091 , \1092 , \1093 , \1094 , \1095 ,
         \1096 , \1097 , \1098 , \1099 , \1100 , \1101 , \1102 , \1103 , \1104 , \1105 ,
         \1106 , \1107 , \1108 , \1109 , \1110 , \1111 , \1112 , \1113 , \1114 , \1115 ,
         \1116 , \1117 , \1118 , \1119 , \1120 , \1121 , \1122 , \1123 , \1124 , \1125 ,
         \1126 , \1127 , \1128 , \1129 , \1130 , \1131 , \1132 , \1133 , \1134 , \1135 ,
         \1136 , \1137 , \1138 , \1139 , \1140 , \1141 , \1142 , \1143 , \1144 , \1145 ,
         \1146 , \1147 , \1148 , \1149 , \1150 , \1151 , \1152 , \1153 , \1154 , \1155 ,
         \1156 , \1157 , \1158 , \1159 , \1160 , \1161 , \1162 , \1163 , \1164 , \1165 ,
         \1166 , \1167 , \1168 , \1169 , \1170 , \1171 , \1172 , \1173 , \1174 , \1175 ,
         \1176 , \1177 , \1178 , \1179 , \1180 , \1181 , \1182 , \1183 , \1184 , \1185 ,
         \1186 , \1187 , \1188 , \1189 , \1190 , \1191 , \1192 , \1193 , \1194 , \1195 ,
         \1196 , \1197 , \1198 , \1199 , \1200 , \1201 , \1202 , \1203 , \1204 , \1205 ,
         \1206 , \1207 , \1208 , \1209 , \1210 , \1211 , \1212 , \1213 , \1214 , \1215 ,
         \1216 , \1217 , \1218 , \1219 , \1220 , \1221 , \1222 , \1223 , \1224 , \1225 ,
         \1226 , \1227 , \1228 , \1229 , \1230 , \1231 , \1232 , \1233 , \1234 , \1235 ,
         \1236 , \1237 , \1238 , \1239 , \1240 , \1241 , \1242 , \1243 , \1244 , \1245 ,
         \1246 , \1247 , \1248 , \1249 , \1250 , \1251 , \1252 , \1253 , \1254 , \1255 ,
         \1256 , \1257 , \1258 , \1259 , \1260 , \1261 , \1262 , \1263 , \1264 , \1265 ,
         \1266 , \1267 , \1268 , \1269 , \1270 , \1271 , \1272 , \1273 , \1274 , \1275 ,
         \1276 , \1277 , \1278 , \1279 , \1280 , \1281 , \1282 , \1283 , \1284 , \1285 ,
         \1286 , \1287 , \1288 , \1289 , \1290 , \1291 , \1292 , \1293 , \1294 , \1295 ,
         \1296 , \1297 , \1298 , \1299 , \1300 , \1301 , \1302 , \1303 , \1304 , \1305 ,
         \1306 , \1307 , \1308 , \1309 , \1310 , \1311 , \1312 , \1313 , \1314 , \1315 ,
         \1316 , \1317 , \1318 , \1319 , \1320 , \1321 , \1322 , \1323 , \1324 , \1325 ,
         \1326 , \1327 , \1328 , \1329 , \1330 , \1331 , \1332 , \1333 , \1334 , \1335 ,
         \1336 , \1337 , \1338 , \1339 , \1340 , \1341 , \1342 , \1343 , \1344 , \1345 ,
         \1346 , \1347 , \1348 , \1349 , \1350 , \1351 , \1352 , \1353 , \1354 , \1355 ,
         \1356 , \1357 , \1358 , \1359 , \1360 , \1361 , \1362 , \1363 , \1364 , \1365 ,
         \1366 , \1367 , \1368 , \1369 , \1370 , \1371 , \1372 , \1373 , \1374 , \1375 ,
         \1376 , \1377 , \1378 , \1379 , \1380 , \1381 , \1382 , \1383 , \1384 , \1385 ,
         \1386 , \1387 , \1388 , \1389 , \1390 , \1391 , \1392 , \1393 , \1394 , \1395 ,
         \1396 , \1397 , \1398 , \1399 , \1400 , \1401 , \1402 , \1403 , \1404 , \1405 ,
         \1406 , \1407 , \1408 , \1409 , \1410 , \1411 , \1412 , \1413 , \1414 , \1415 ,
         \1416 , \1417 , \1418 , \1419 , \1420 , \1421 , \1422 , \1423 , \1424 , \1425 ,
         \1426 , \1427 , \1428 , \1429 , \1430 , \1431 , \1432 , \1433 , \1434 , \1435 ,
         \1436 , \1437 , \1438 , \1439 , \1440 , \1441 , \1442 , \1443 , \1444 , \1445 ,
         \1446 , \1447 , \1448 , \1449 , \1450 , \1451 , \1452 , \1453 , \1454 , \1455 ,
         \1456 , \1457 , \1458 , \1459 , \1460 , \1461 , \1462 , \1463 , \1464 , \1465 ,
         \1466 , \1467 , \1468 , \1469 , \1470 , \1471 , \1472 , \1473 , \1474 , \1475 ,
         \1476 , \1477 , \1478 , \1479 , \1480 , \1481 , \1482 , \1483 , \1484 , \1485 ,
         \1486 , \1487 , \1488 , \1489 , \1490 , \1491 , \1492 , \1493 , \1494 , \1495 ,
         \1496 , \1497 , \1498 , \1499 , \1500 , \1501 , \1502 , \1503 , \1504 , \1505 ,
         \1506 , \1507 , \1508 , \1509 , \1510 , \1511 , \1512 , \1513 , \1514 , \1515 ,
         \1516 , \1517 , \1518 , \1519 , \1520 , \1521 , \1522 , \1523 , \1524 , \1525 ,
         \1526 , \1527 , \1528 , \1529 , \1530 , \1531 , \1532 , \1533 , \1534 , \1535 ,
         \1536 , \1537 , \1538 , \1539 , \1540 , \1541 , \1542 , \1543 , \1544 , \1545 ,
         \1546 , \1547 , \1548 , \1549 , \1550 , \1551 , \1552 , \1553 , \1554 , \1555 ,
         \1556 , \1557 , \1558 , \1559 , \1560 , \1561 , \1562 , \1563 , \1564 , \1565 ,
         \1566 , \1567 , \1568 , \1569 , \1570 , \1571 , \1572 , \1573 , \1574 , \1575 ,
         \1576 , \1577 , \1578 , \1579 , \1580 , \1581 , \1582 , \1583 , \1584 , \1585 ,
         \1586 , \1587 , \1588 , \1589 , \1590 , \1591 , \1592 , \1593 , \1594 , \1595 ,
         \1596 , \1597 , \1598 , \1599 , \1600 , \1601 , \1602 , \1603 , \1604 , \1605 ,
         \1606 , \1607 , \1608 , \1609 , \1610 , \1611 , \1612 , \1613 , \1614 , \1615 ,
         \1616 , \1617 , \1618 , \1619 , \1620 , \1621 , \1622 , \1623 , \1624 , \1625 ,
         \1626 , \1627 , \1628 , \1629 , \1630 , \1631 , \1632 , \1633 , \1634 , \1635 ,
         \1636 , \1637 , \1638 , \1639 , \1640 , \1641 , \1642 , \1643 , \1644 , \1645 ,
         \1646 , \1647 , \1648 , \1649 , \1650 , \1651 , \1652 , \1653 , \1654 , \1655 ,
         \1656 , \1657 , \1658 , \1659 , \1660 , \1661 , \1662 , \1663 , \1664 , \1665 ,
         \1666 , \1667 , \1668 , \1669 , \1670 , \1671 , \1672 , \1673 , \1674 , \1675 ,
         \1676 , \1677 , \1678 , \1679 , \1680 , \1681 , \1682 , \1683 , \1684 , \1685 ,
         \1686 , \1687 , \1688 , \1689 , \1690 , \1691 , \1692 , \1693 , \1694 , \1695 ,
         \1696 , \1697 , \1698 , \1699 , \1700 , \1701 , \1702 , \1703 , \1704 , \1705 ,
         \1706 , \1707 , \1708 , \1709 , \1710 , \1711 , \1712 , \1713 , \1714 , \1715 ,
         \1716 , \1717 , \1718 , \1719 , \1720 , \1721 , \1722 , \1723 , \1724 , \1725 ,
         \1726 , \1727 , \1728 , \1729 , \1730 , \1731 , \1732 , \1733 , \1734 , \1735 ,
         \1736 , \1737 , \1738 , \1739 , \1740 , \1741 , \1742 , \1743 , \1744 , \1745 ,
         \1746 , \1747 , \1748 , \1749 , \1750 , \1751 , \1752 , \1753 , \1754 , \1755 ,
         \1756 , \1757 , \1758 , \1759 , \1760 , \1761 , \1762 , \1763 , \1764 , \1765 ,
         \1766 , \1767 , \1768 , \1769 , \1770 , \1771 , \1772 , \1773 , \1774 , \1775 ,
         \1776 , \1777 , \1778 , \1779 , \1780 , \1781 , \1782 , \1783 , \1784 , \1785 ,
         \1786 , \1787 , \1788 , \1789 , \1790 , \1791 , \1792 , \1793 , \1794 , \1795 ,
         \1796 , \1797 , \1798 , \1799 , \1800 , \1801 , \1802 , \1803 , \1804 , \1805 ,
         \1806 , \1807 , \1808 , \1809 , \1810 , \1811 , \1812 , \1813 , \1814 , \1815 ,
         \1816 , \1817 , \1818 , \1819 , \1820 , \1821 , \1822 , \1823 , \1824 , \1825 ,
         \1826 , \1827 , \1828 , \1829 , \1830 , \1831 , \1832 , \1833 , \1834 , \1835 ,
         \1836 , \1837 , \1838 , \1839 , \1840 , \1841 , \1842 , \1843 , \1844 , \1845 ,
         \1846 , \1847 , \1848 , \1849 , \1850 , \1851 , \1852 , \1853 , \1854 , \1855 ,
         \1856 , \1857 , \1858 , \1859 , \1860 , \1861 , \1862 , \1863 , \1864 , \1865 ,
         \1866 , \1867 , \1868 , \1869 , \1870 , \1871 , \1872 , \1873 , \1874 , \1875 ,
         \1876 , \1877 , \1878 , \1879 , \1880 , \1881 , \1882 , \1883 , \1884 , \1885 ,
         \1886 , \1887 , \1888 , \1889 , \1890 , \1891 , \1892 , \1893 , \1894 , \1895 ,
         \1896 , \1897 , \1898 , \1899 , \1900 , \1901 , \1902 , \1903 , \1904 , \1905 ,
         \1906 , \1907 , \1908 , \1909 , \1910 , \1911 , \1912 , \1913 , \1914 , \1915 ,
         \1916 , \1917 , \1918 , \1919 , \1920 , \1921 , \1922 , \1923 , \1924 , \1925 ,
         \1926 , \1927 , \1928 , \1929 , \1930 , \1931 , \1932 , \1933 , \1934 , \1935 ,
         \1936 , \1937 , \1938 , \1939 , \1940 , \1941 , \1942 , \1943 , \1944 , \1945 ,
         \1946 , \1947 , \1948 , \1949 , \1950 , \1951 , \1952 , \1953 , \1954 , \1955 ,
         \1956 , \1957 , \1958 , \1959 , \1960 , \1961 , \1962 , \1963 , \1964 , \1965 ,
         \1966 , \1967 , \1968 , \1969 , \1970 , \1971 , \1972 , \1973 , \1974 , \1975 ,
         \1976 , \1977 , \1978 , \1979 , \1980 , \1981 , \1982 , \1983 , \1984 , \1985 ,
         \1986 , \1987 , \1988 , \1989 , \1990 , \1991 , \1992 , \1993 , \1994 , \1995 ,
         \1996 , \1997 , \1998 , \1999 , \2000 , \2001 , \2002 , \2003 , \2004 , \2005 ,
         \2006 , \2007 , \2008 , \2009 , \2010 , \2011 , \2012 , \2013 , \2014 , \2015 ,
         \2016 , \2017 , \2018 , \2019 , \2020 , \2021 , \2022 , \2023 , \2024 , \2025 ,
         \2026 , \2027 , \2028 , \2029 , \2030 , \2031 , \2032 , \2033 , \2034 , \2035 ,
         \2036 , \2037 , \2038 , \2039 , \2040 , \2041 , \2042 , \2043 , \2044 , \2045 ,
         \2046 , \2047 , \2048 , \2049 , \2050 , \2051 , \2052 , \2053 , \2054 , \2055 ,
         \2056 , \2057 , \2058 , \2059 , \2060 , \2061 , \2062 , \2063 , \2064 , \2065 ,
         \2066 , \2067 , \2068 , \2069 , \2070 , \2071 , \2072 , \2073 , \2074 , \2075 ,
         \2076 , \2077 , \2078 , \2079 , \2080 , \2081 , \2082 , \2083 , \2084 , \2085 ,
         \2086 , \2087 , \2088 , \2089 , \2090 , \2091 , \2092 , \2093 , \2094 , \2095 ,
         \2096 , \2097 , \2098 , \2099 , \2100 , \2101 , \2102 , \2103 , \2104 , \2105 ,
         \2106 , \2107 , \2108 , \2109 , \2110 , \2111 , \2112 , \2113 , \2114 , \2115 ,
         \2116 , \2117 , \2118 , \2119 , \2120 , \2121 , \2122 , \2123 , \2124 , \2125 ,
         \2126 , \2127 , \2128 , \2129 , \2130 , \2131 , \2132 , \2133 , \2134 , \2135 ,
         \2136 , \2137 , \2138 , \2139 , \2140 , \2141 , \2142 , \2143 , \2144 , \2145 ,
         \2146 , \2147 , \2148 , \2149 , \2150 , \2151 , \2152 , \2153 , \2154 , \2155 ,
         \2156 , \2157 , \2158 , \2159 , \2160 , \2161 , \2162 , \2163 , \2164 , \2165 ,
         \2166 , \2167 , \2168 , \2169 , \2170 , \2171 , \2172 , \2173 , \2174 , \2175 ,
         \2176 , \2177 , \2178 , \2179 , \2180 , \2181 , \2182 , \2183 , \2184 , \2185 ,
         \2186 , \2187 , \2188 , \2189 , \2190 , \2191 , \2192 , \2193 , \2194 , \2195 ,
         \2196 , \2197 , \2198 , \2199 , \2200 , \2201 , \2202 , \2203 , \2204 , \2205 ,
         \2206 , \2207 , \2208 , \2209 , \2210 , \2211 , \2212 , \2213 , \2214 , \2215 ,
         \2216 , \2217 , \2218 , \2219 , \2220 , \2221 , \2222 , \2223 , \2224 , \2225 ,
         \2226 , \2227 , \2228 , \2229 , \2230 , \2231 , \2232 , \2233 , \2234 , \2235 ,
         \2236 , \2237 , \2238 , \2239 , \2240 , \2241 , \2242 , \2243 , \2244 , \2245 ,
         \2246 , \2247 , \2248 , \2249 , \2250 , \2251 , \2252 , \2253 , \2254 , \2255 ,
         \2256 , \2257 , \2258 , \2259 , \2260 , \2261 , \2262 , \2263 , \2264 , \2265 ,
         \2266 , \2267 , \2268 , \2269 , \2270 , \2271 , \2272 , \2273 , \2274 , \2275 ,
         \2276 , \2277 , \2278 , \2279 , \2280 , \2281 , \2282 , \2283 , \2284 , \2285 ,
         \2286 , \2287 , \2288 , \2289 , \2290 , \2291 , \2292 , \2293 , \2294 , \2295 ,
         \2296 , \2297 , \2298 , \2299 , \2300 , \2301 , \2302 , \2303 , \2304 , \2305 ,
         \2306 , \2307 , \2308 , \2309 , \2310 , \2311 , \2312 , \2313 , \2314 , \2315 ,
         \2316 , \2317 , \2318 , \2319 , \2320 , \2321 , \2322 , \2323 , \2324 , \2325 ,
         \2326 , \2327 , \2328 , \2329 , \2330 , \2331 , \2332 , \2333 , \2334 , \2335 ,
         \2336 , \2337 , \2338 , \2339 , \2340 , \2341 , \2342 , \2343 , \2344 , \2345 ,
         \2346 , \2347 , \2348 , \2349 , \2350 , \2351 , \2352 , \2353 , \2354 , \2355 ,
         \2356 , \2357 , \2358 , \2359 , \2360 , \2361 , \2362 , \2363 , \2364 , \2365 ,
         \2366 , \2367 , \2368 , \2369 , \2370 , \2371 , \2372 , \2373 , \2374 , \2375 ,
         \2376 , \2377 , \2378 , \2379 , \2380 , \2381 , \2382 , \2383 , \2384 , \2385 ,
         \2386 , \2387 , \2388 , \2389 , \2390 , \2391 , \2392 , \2393 , \2394 , \2395 ,
         \2396 , \2397 , \2398 , \2399 , \2400 , \2401 , \2402 , \2403 , \2404 , \2405 ,
         \2406 , \2407 , \2408 , \2409 , \2410 , \2411 , \2412 , \2413 , \2414 , \2415 ,
         \2416 , \2417 , \2418 , \2419 , \2420 , \2421 , \2422 , \2423 , \2424 , \2425 ,
         \2426 , \2427 , \2428 , \2429 , \2430 , \2431 , \2432 , \2433 , \2434 , \2435 ,
         \2436 , \2437 , \2438 , \2439 , \2440 , \2441 , \2442 , \2443 , \2444 , \2445 ,
         \2446 , \2447 , \2448 , \2449 , \2450 , \2451 , \2452 , \2453 , \2454 , \2455 ,
         \2456 , \2457 , \2458 , \2459 , \2460 , \2461 , \2462 , \2463 , \2464 , \2465 ,
         \2466 , \2467 , \2468 , \2469 , \2470 , \2471 , \2472 , \2473 , \2474 , \2475 ,
         \2476 , \2477 , \2478 , \2479 , \2480 , \2481 , \2482 , \2483 , \2484 , \2485 ,
         \2486 , \2487 , \2488 , \2489 , \2490 , \2491 , \2492 , \2493 , \2494 , \2495 ,
         \2496 , \2497 , \2498 , \2499 , \2500 , \2501 , \2502 , \2503 , \2504 , \2505 ,
         \2506 , \2507 , \2508 , \2509 , \2510 , \2511 , \2512 , \2513 , \2514 , \2515 ,
         \2516 , \2517 , \2518 , \2519 , \2520 , \2521 , \2522 , \2523 , \2524 , \2525 ,
         \2526 , \2527 , \2528 , \2529 , \2530 , \2531 , \2532 , \2533 , \2534 , \2535 ,
         \2536 , \2537 , \2538 , \2539 , \2540 , \2541 , \2542 , \2543 , \2544 , \2545 ,
         \2546 , \2547 , \2548 , \2549 , \2550 , \2551 , \2552 , \2553 , \2554 , \2555 ,
         \2556 , \2557 , \2558 , \2559 , \2560 , \2561 , \2562 , \2563 , \2564 , \2565 ,
         \2566 , \2567 , \2568 , \2569 , \2570 , \2571 , \2572 , \2573 , \2574 , \2575 ,
         \2576 , \2577 , \2578 , \2579 , \2580 , \2581 , \2582 , \2583 , \2584 , \2585 ,
         \2586 , \2587 , \2588 , \2589 , \2590 , \2591 , \2592 , \2593 , \2594 , \2595 ,
         \2596 , \2597 , \2598 , \2599 , \2600 , \2601 , \2602 , \2603 , \2604 , \2605 ,
         \2606 , \2607 , \2608 , \2609 , \2610 , \2611 , \2612 , \2613 , \2614 , \2615 ,
         \2616 , \2617 , \2618 , \2619 , \2620 , \2621 , \2622 , \2623 , \2624 , \2625 ,
         \2626 , \2627 , \2628 , \2629 , \2630 , \2631 , \2632 , \2633 , \2634 , \2635 ,
         \2636 , \2637 , \2638 , \2639 , \2640 , \2641 , \2642 , \2643 , \2644 , \2645 ,
         \2646 , \2647 , \2648 , \2649 , \2650 , \2651 , \2652 , \2653 , \2654 , \2655 ,
         \2656 , \2657 , \2658 , \2659 , \2660 , \2661 , \2662 , \2663 , \2664 , \2665 ,
         \2666 , \2667 , \2668 , \2669 , \2670 , \2671 , \2672 , \2673 , \2674 , \2675 ,
         \2676 , \2677 , \2678 , \2679 , \2680 , \2681 , \2682 , \2683 , \2684 , \2685 ,
         \2686 , \2687 , \2688 , \2689 , \2690 , \2691 , \2692 , \2693 , \2694 , \2695 ,
         \2696 , \2697 , \2698 , \2699 , \2700 , \2701 , \2702 , \2703 , \2704 , \2705 ,
         \2706 , \2707 , \2708 , \2709 , \2710 , \2711 , \2712 , \2713 , \2714 , \2715 ,
         \2716 , \2717 , \2718 , \2719 , \2720 , \2721 , \2722 , \2723 , \2724 , \2725 ,
         \2726 , \2727 , \2728 , \2729 , \2730 , \2731 , \2732 , \2733 , \2734 , \2735 ,
         \2736 , \2737 , \2738 , \2739 , \2740 , \2741 , \2742 , \2743 , \2744 , \2745 ,
         \2746 , \2747 , \2748 , \2749 , \2750 , \2751 , \2752 , \2753 , \2754 , \2755 ,
         \2756 , \2757 , \2758 , \2759 , \2760 , \2761 , \2762 , \2763 , \2764 , \2765 ,
         \2766 , \2767 , \2768 , \2769 , \2770 , \2771 , \2772 , \2773 , \2774 , \2775 ,
         \2776 , \2777 , \2778 , \2779 , \2780 , \2781 , \2782 , \2783 , \2784 , \2785 ,
         \2786 , \2787 , \2788 , \2789 , \2790 , \2791 , \2792 , \2793 , \2794 , \2795 ,
         \2796 , \2797 , \2798 , \2799 , \2800 , \2801 , \2802 , \2803 , \2804 , \2805 ,
         \2806 , \2807 , \2808 , \2809 , \2810 , \2811 , \2812 , \2813 , \2814 , \2815 ,
         \2816 , \2817 , \2818 , \2819 , \2820 , \2821 , \2822 , \2823 , \2824 , \2825 ,
         \2826 , \2827 , \2828 , \2829 , \2830 , \2831 , \2832 , \2833 , \2834 , \2835 ,
         \2836 , \2837 , \2838 , \2839 , \2840 , \2841 , \2842 , \2843 , \2844 , \2845 ,
         \2846 , \2847 , \2848 , \2849 , \2850 , \2851 , \2852 , \2853 , \2854 , \2855 ,
         \2856 , \2857 , \2858 , \2859 , \2860 , \2861 , \2862 , \2863 , \2864 , \2865 ,
         \2866 , \2867 , \2868 , \2869 , \2870 , \2871 , \2872 , \2873 , \2874 , \2875 ,
         \2876 , \2877 , \2878 , \2879 , \2880 , \2881 , \2882 , \2883 , \2884 , \2885 ,
         \2886 , \2887 , \2888 , \2889 , \2890 , \2891 , \2892 , \2893 , \2894 , \2895 ,
         \2896 , \2897 , \2898 , \2899 , \2900 , \2901 , \2902 , \2903 , \2904 , \2905 ,
         \2906 , \2907 , \2908 , \2909 , \2910 , \2911 , \2912 , \2913 , \2914 , \2915 ,
         \2916 , \2917 , \2918 , \2919 , \2920 , \2921 , \2922 , \2923 , \2924 , \2925 ,
         \2926 , \2927 , \2928 , \2929 , \2930 , \2931 , \2932 , \2933 , \2934 , \2935 ,
         \2936 , \2937 , \2938 , \2939 , \2940 , \2941 , \2942 , \2943 , \2944 , \2945 ,
         \2946 , \2947 , \2948 , \2949 , \2950 , \2951 , \2952 , \2953 , \2954 , \2955 ,
         \2956 , \2957 , \2958 , \2959 , \2960 , \2961 , \2962 , \2963 , \2964 , \2965 ,
         \2966 , \2967 , \2968 , \2969 , \2970 , \2971 , \2972 , \2973 , \2974 , \2975 ,
         \2976 , \2977 , \2978 , \2979 , \2980 , \2981 , \2982 , \2983 , \2984 , \2985 ,
         \2986 , \2987 , \2988 , \2989 , \2990 , \2991 , \2992 , \2993 , \2994 , \2995 ,
         \2996 , \2997 , \2998 , \2999 , \3000 , \3001 , \3002 , \3003 , \3004 , \3005 ,
         \3006 , \3007 , \3008 , \3009 , \3010 , \3011 , \3012 , \3013 , \3014 , \3015 ,
         \3016 , \3017 , \3018 , \3019 , \3020 , \3021 , \3022 , \3023 , \3024 , \3025 ,
         \3026 , \3027 , \3028 , \3029 , \3030 , \3031 , \3032 , \3033 , \3034 , \3035 ,
         \3036 , \3037 , \3038 , \3039 , \3040 , \3041 , \3042 , \3043 , \3044 , \3045 ,
         \3046 , \3047 , \3048 , \3049 , \3050 , \3051 , \3052 , \3053 , \3054 , \3055 ,
         \3056 , \3057 , \3058 , \3059 , \3060 , \3061 , \3062 , \3063 , \3064 , \3065 ,
         \3066 , \3067 , \3068 , \3069 , \3070 , \3071 , \3072 , \3073 , \3074 , \3075 ,
         \3076 , \3077 , \3078 , \3079 , \3080 , \3081 , \3082 , \3083 , \3084 , \3085 ,
         \3086 , \3087 , \3088 , \3089 , \3090 , \3091 , \3092 , \3093 , \3094 , \3095 ,
         \3096 , \3097 , \3098 , \3099 , \3100 , \3101 , \3102 , \3103 , \3104 , \3105 ,
         \3106 , \3107 , \3108 , \3109 , \3110 , \3111 , \3112 , \3113 , \3114 , \3115 ,
         \3116 , \3117 , \3118 , \3119 , \3120 , \3121 , \3122 , \3123 , \3124 , \3125 ,
         \3126 , \3127 , \3128 , \3129 , \3130 , \3131 , \3132 , \3133 , \3134 , \3135 ,
         \3136 , \3137 , \3138 , \3139 , \3140 , \3141 , \3142 , \3143 , \3144 , \3145 ,
         \3146 , \3147 , \3148 , \3149 , \3150 , \3151 , \3152 , \3153 , \3154 , \3155 ,
         \3156 , \3157 , \3158 , \3159 , \3160 , \3161 , \3162 , \3163 , \3164 , \3165 ,
         \3166 , \3167 , \3168 , \3169 , \3170 , \3171 , \3172 , \3173 , \3174 , \3175 ,
         \3176 , \3177 , \3178 , \3179 , \3180 , \3181 , \3182 , \3183 , \3184 , \3185 ,
         \3186 , \3187 , \3188 , \3189 , \3190 , \3191 , \3192 , \3193 , \3194 , \3195 ,
         \3196 , \3197 , \3198 , \3199 , \3200 , \3201 , \3202 , \3203 , \3204 , \3205 ,
         \3206 , \3207 , \3208 , \3209 , \3210 , \3211 , \3212 , \3213 , \3214 , \3215 ,
         \3216 , \3217 , \3218 , \3219 , \3220 , \3221 , \3222 , \3223 , \3224 , \3225 ,
         \3226 , \3227 , \3228 , \3229 , \3230 , \3231 , \3232 , \3233 , \3234 , \3235 ,
         \3236 , \3237 , \3238 , \3239 , \3240 , \3241 , \3242 , \3243 , \3244 , \3245 ,
         \3246 , \3247 , \3248 , \3249 , \3250 , \3251 , \3252 , \3253 , \3254 , \3255 ,
         \3256 , \3257 , \3258 , \3259 , \3260 , \3261 , \3262 , \3263 , \3264 , \3265 ,
         \3266 , \3267 , \3268 , \3269 , \3270 , \3271 , \3272 , \3273 , \3274 , \3275 ,
         \3276 , \3277 , \3278 , \3279 , \3280 , \3281 , \3282 , \3283 , \3284 , \3285 ,
         \3286 , \3287 , \3288 , \3289 , \3290 , \3291 , \3292 , \3293 , \3294 , \3295 ,
         \3296 , \3297 , \3298 , \3299 , \3300 , \3301 , \3302 , \3303 , \3304 , \3305 ,
         \3306 , \3307 , \3308 , \3309 , \3310 , \3311 , \3312 , \3313 , \3314 , \3315 ,
         \3316 , \3317 , \3318 , \3319 , \3320 , \3321 , \3322 , \3323 , \3324 , \3325 ,
         \3326 , \3327 , \3328 , \3329 , \3330 , \3331 , \3332 , \3333 , \3334 , \3335 ,
         \3336 , \3337 , \3338 , \3339 , \3340 , \3341 , \3342 , \3343 , \3344 , \3345 ,
         \3346 , \3347 , \3348 , \3349 , \3350 , \3351 , \3352 , \3353 , \3354 , \3355 ,
         \3356 , \3357 , \3358 , \3359 , \3360 , \3361 , \3362 , \3363 , \3364 , \3365 ,
         \3366 , \3367 , \3368 , \3369 , \3370 , \3371 , \3372 , \3373 , \3374 , \3375 ,
         \3376 , \3377 , \3378 , \3379 , \3380 , \3381 , \3382 , \3383 , \3384 , \3385 ,
         \3386 , \3387 , \3388 , \3389 , \3390 , \3391 , \3392 , \3393 , \3394 , \3395 ,
         \3396 , \3397 , \3398 , \3399 , \3400 , \3401 , \3402 , \3403 , \3404 , \3405 ,
         \3406 , \3407 , \3408 , \3409 , \3410 , \3411 , \3412 , \3413 , \3414 , \3415 ,
         \3416 , \3417 , \3418 , \3419 , \3420 , \3421 , \3422 , \3423 , \3424 , \3425 ,
         \3426 , \3427 , \3428 , \3429 , \3430 , \3431 , \3432 , \3433 , \3434 , \3435 ,
         \3436 , \3437 , \3438 , \3439 , \3440 , \3441 , \3442 , \3443 , \3444 , \3445 ,
         \3446 , \3447 , \3448 , \3449 , \3450 , \3451 , \3452 , \3453 , \3454 , \3455 ,
         \3456 , \3457 , \3458 , \3459 , \3460 , \3461 , \3462 , \3463 , \3464 , \3465 ,
         \3466 , \3467 , \3468 , \3469 , \3470 , \3471 , \3472 , \3473 , \3474 , \3475 ,
         \3476 , \3477 , \3478 , \3479 , \3480 , \3481 , \3482 , \3483 , \3484 , \3485 ,
         \3486 , \3487 , \3488 , \3489 , \3490 , \3491 , \3492 , \3493 , \3494 , \3495 ,
         \3496 , \3497 , \3498 , \3499 , \3500 , \3501 , \3502 , \3503 , \3504 , \3505 ,
         \3506 , \3507 , \3508 , \3509 , \3510 , \3511 , \3512 , \3513 , \3514 , \3515 ,
         \3516 , \3517 , \3518 , \3519 , \3520 , \3521 , \3522 , \3523 , \3524 , \3525 ,
         \3526 , \3527 , \3528 , \3529 , \3530 , \3531 , \3532 , \3533 , \3534 , \3535 ,
         \3536 , \3537 , \3538 , \3539 , \3540 , \3541 , \3542 , \3543 , \3544 , \3545 ,
         \3546 , \3547 , \3548 , \3549 , \3550 , \3551 , \3552 , \3553 , \3554 , \3555 ,
         \3556 , \3557 , \3558 , \3559 , \3560 , \3561 , \3562 , \3563 , \3564 , \3565 ,
         \3566 , \3567 , \3568 , \3569 , \3570 , \3571 , \3572 , \3573 , \3574 , \3575 ,
         \3576 , \3577 , \3578 , \3579 , \3580 , \3581 , \3582 , \3583 , \3584 , \3585 ,
         \3586 , \3587 , \3588 , \3589 , \3590 , \3591 , \3592 , \3593 , \3594 , \3595 ,
         \3596 , \3597 , \3598 , \3599 , \3600 , \3601 , \3602 , \3603 , \3604 , \3605 ,
         \3606 , \3607 , \3608 , \3609 , \3610 , \3611 , \3612 , \3613 , \3614 , \3615 ,
         \3616 , \3617 , \3618 , \3619 , \3620 , \3621 , \3622 , \3623 , \3624 , \3625 ,
         \3626 , \3627 , \3628 , \3629 , \3630 , \3631 , \3632 , \3633 , \3634 , \3635 ,
         \3636 , \3637 , \3638 , \3639 , \3640 , \3641 , \3642 , \3643 , \3644 , \3645 ,
         \3646 , \3647 , \3648 , \3649 , \3650 , \3651 , \3652 , \3653 , \3654 , \3655 ,
         \3656 , \3657 , \3658 , \3659 , \3660 , \3661 , \3662 , \3663 , \3664 , \3665 ,
         \3666 , \3667 , \3668 , \3669 , \3670 , \3671 , \3672 , \3673 , \3674 , \3675 ,
         \3676 , \3677 , \3678 , \3679 , \3680 , \3681 , \3682 , \3683 , \3684 , \3685 ,
         \3686 , \3687 , \3688 , \3689 , \3690 , \3691 , \3692 , \3693 , \3694 , \3695 ,
         \3696 , \3697 , \3698 , \3699 , \3700 , \3701 , \3702 , \3703 , \3704 , \3705 ,
         \3706 , \3707 , \3708 , \3709 , \3710 , \3711 , \3712 , \3713 , \3714 , \3715 ,
         \3716 , \3717 , \3718 , \3719 , \3720 , \3721 , \3722 , \3723 , \3724 , \3725 ,
         \3726 , \3727 , \3728 , \3729 , \3730 , \3731 , \3732 , \3733 , \3734 , \3735 ,
         \3736 , \3737 , \3738 , \3739 , \3740 , \3741 , \3742 , \3743 , \3744 , \3745 ,
         \3746 , \3747 , \3748 , \3749 , \3750 , \3751 , \3752 , \3753 , \3754 , \3755 ,
         \3756 , \3757 , \3758 , \3759 , \3760 , \3761 , \3762 , \3763 , \3764 , \3765 ,
         \3766 , \3767 , \3768 , \3769 , \3770 , \3771 , \3772 , \3773 , \3774 , \3775 ,
         \3776 , \3777 , \3778 , \3779 , \3780 , \3781 , \3782 , \3783 , \3784 , \3785 ,
         \3786 , \3787 , \3788 , \3789 , \3790 , \3791 , \3792 , \3793 , \3794 , \3795 ,
         \3796 , \3797 , \3798 , \3799 , \3800 , \3801 , \3802 , \3803 , \3804 , \3805 ,
         \3806 , \3807 , \3808 , \3809 , \3810 , \3811 , \3812 , \3813 , \3814 , \3815 ,
         \3816 , \3817 , \3818 , \3819 , \3820 , \3821 , \3822 , \3823 , \3824 , \3825 ,
         \3826 , \3827 , \3828 , \3829 , \3830 , \3831 , \3832 , \3833 , \3834 , \3835 ,
         \3836 , \3837 , \3838 , \3839 , \3840 , \3841 , \3842 , \3843 , \3844 , \3845 ,
         \3846 , \3847 , \3848 , \3849 , \3850 , \3851 , \3852 , \3853 , \3854 , \3855 ,
         \3856 , \3857 , \3858 , \3859 , \3860 , \3861 , \3862 , \3863 , \3864 , \3865 ,
         \3866 , \3867 , \3868 , \3869 , \3870 , \3871 , \3872 , \3873 , \3874 , \3875 ,
         \3876 , \3877 , \3878 , \3879 , \3880 , \3881 , \3882 , \3883 , \3884 , \3885 ,
         \3886 , \3887 , \3888 , \3889 , \3890 , \3891 , \3892 , \3893 , \3894 , \3895 ,
         \3896 , \3897 , \3898 , \3899 , \3900 , \3901 , \3902 , \3903 , \3904 , \3905 ,
         \3906 , \3907 , \3908 , \3909 , \3910 , \3911 , \3912 , \3913 , \3914 , \3915 ,
         \3916 , \3917 , \3918 , \3919 , \3920 , \3921 , \3922 , \3923 , \3924 , \3925 ,
         \3926 , \3927 , \3928 , \3929 , \3930 , \3931 , \3932 , \3933 , \3934 , \3935 ,
         \3936 , \3937 , \3938 , \3939 , \3940 , \3941 , \3942 , \3943 , \3944 , \3945 ,
         \3946 , \3947 , \3948 , \3949 , \3950 , \3951 , \3952 , \3953 , \3954 , \3955 ,
         \3956 , \3957 , \3958 , \3959 , \3960 , \3961 , \3962 , \3963 , \3964 , \3965 ,
         \3966 , \3967 , \3968 , \3969 , \3970 , \3971 , \3972 , \3973 , \3974 , \3975 ,
         \3976 , \3977 , \3978 , \3979 , \3980 , \3981 , \3982 , \3983 , \3984 , \3985 ,
         \3986 , \3987 , \3988 , \3989 , \3990 , \3991 , \3992 , \3993 , \3994 , \3995 ,
         \3996 , \3997 , \3998 , \3999 , \4000 , \4001 , \4002 , \4003 , \4004 , \4005 ,
         \4006 , \4007 , \4008 , \4009 , \4010 , \4011 , \4012 , \4013 , \4014 , \4015 ,
         \4016 , \4017 , \4018 , \4019 , \4020 , \4021 , \4022 , \4023 , \4024 , \4025 ,
         \4026 , \4027 , \4028 , \4029 , \4030 , \4031 , \4032 , \4033 , \4034 , \4035 ,
         \4036 , \4037 , \4038 , \4039 , \4040 , \4041 , \4042 , \4043 , \4044 , \4045 ,
         \4046 , \4047 , \4048 , \4049 , \4050 , \4051 , \4052 , \4053 , \4054 , \4055 ,
         \4056 , \4057 , \4058 , \4059 , \4060 , \4061 , \4062 , \4063 , \4064 , \4065 ,
         \4066 , \4067 , \4068 , \4069 , \4070 , \4071 , \4072 , \4073 , \4074 , \4075 ,
         \4076 , \4077 , \4078 , \4079 , \4080 , \4081 , \4082 , \4083 , \4084 , \4085 ,
         \4086 , \4087 , \4088 , \4089 , \4090 , \4091 , \4092 , \4093 , \4094 , \4095 ,
         \4096 , \4097 , \4098 , \4099 , \4100 , \4101 , \4102 , \4103 , \4104 , \4105 ,
         \4106 , \4107 , \4108 , \4109 , \4110 , \4111 , \4112 , \4113 , \4114 , \4115 ,
         \4116 , \4117 , \4118 , \4119 , \4120 , \4121 , \4122 , \4123 , \4124 , \4125 ,
         \4126 , \4127 , \4128 , \4129 , \4130 , \4131 , \4132 , \4133 , \4134 , \4135 ,
         \4136 , \4137 , \4138 , \4139 , \4140 , \4141 , \4142 , \4143 , \4144 , \4145 ,
         \4146 , \4147 , \4148 , \4149 , \4150 , \4151 , \4152 , \4153 , \4154 , \4155 ,
         \4156 , \4157 , \4158 , \4159 , \4160 , \4161 , \4162 , \4163 , \4164 , \4165 ,
         \4166 , \4167 , \4168 , \4169 , \4170 , \4171 , \4172 , \4173 , \4174 , \4175 ,
         \4176 , \4177 , \4178 , \4179 , \4180 , \4181 , \4182 , \4183 , \4184 , \4185 ,
         \4186 , \4187 , \4188 , \4189 , \4190 , \4191 , \4192 , \4193 , \4194 , \4195 ,
         \4196 , \4197 , \4198 , \4199 , \4200 , \4201 , \4202 , \4203 , \4204 , \4205 ,
         \4206 , \4207 , \4208 , \4209 , \4210 , \4211 , \4212 , \4213 , \4214 , \4215 ,
         \4216 , \4217 , \4218 , \4219 , \4220 , \4221 , \4222 , \4223 , \4224 , \4225 ,
         \4226 , \4227 , \4228 , \4229 , \4230 , \4231 , \4232 , \4233 , \4234 , \4235 ,
         \4236 , \4237 , \4238 , \4239 , \4240 , \4241 , \4242 , \4243 , \4244 , \4245 ,
         \4246 , \4247 , \4248 , \4249 , \4250 , \4251 , \4252 , \4253 , \4254 , \4255 ,
         \4256 , \4257 , \4258 , \4259 , \4260 , \4261 , \4262 , \4263 , \4264 , \4265 ,
         \4266 , \4267 , \4268 , \4269 , \4270 , \4271 , \4272 , \4273 , \4274 , \4275 ,
         \4276 , \4277 , \4278 , \4279 , \4280 , \4281 , \4282 , \4283 , \4284 , \4285 ,
         \4286 , \4287 , \4288 , \4289 , \4290 , \4291 , \4292 , \4293 , \4294 , \4295 ,
         \4296 , \4297 , \4298 , \4299 , \4300 , \4301 , \4302 , \4303 , \4304 , \4305 ,
         \4306 , \4307 , \4308 , \4309 , \4310 , \4311 , \4312 , \4313 , \4314 , \4315 ,
         \4316 , \4317 , \4318 , \4319 , \4320 , \4321 , \4322 , \4323 , \4324 , \4325 ,
         \4326 , \4327 , \4328 , \4329 , \4330 , \4331 , \4332 , \4333 , \4334 , \4335 ,
         \4336 , \4337 , \4338 , \4339 , \4340 , \4341 , \4342 , \4343 , \4344 , \4345 ,
         \4346 , \4347 , \4348 , \4349 , \4350 , \4351 , \4352 , \4353 , \4354 , \4355 ,
         \4356 , \4357 , \4358 , \4359 , \4360 , \4361 , \4362 , \4363 , \4364 , \4365 ,
         \4366 , \4367 , \4368 , \4369 , \4370 , \4371 , \4372 , \4373 , \4374 , \4375 ,
         \4376 , \4377 , \4378 , \4379 , \4380 , \4381 , \4382 , \4383 , \4384 , \4385 ,
         \4386 , \4387 , \4388 , \4389 , \4390 , \4391 , \4392 , \4393 , \4394 , \4395 ,
         \4396 , \4397 , \4398 , \4399 , \4400 , \4401 , \4402 , \4403 , \4404 , \4405 ,
         \4406 , \4407 , \4408 , \4409 , \4410 , \4411 , \4412 , \4413 , \4414 , \4415 ,
         \4416 , \4417 , \4418 , \4419 , \4420 , \4421 , \4422 , \4423 , \4424 , \4425 ,
         \4426 , \4427 , \4428 , \4429 , \4430 , \4431 , \4432 , \4433 , \4434 , \4435 ,
         \4436 , \4437 , \4438 , \4439 , \4440 , \4441 , \4442 , \4443 , \4444 , \4445 ,
         \4446 , \4447 , \4448 , \4449 , \4450 , \4451 , \4452 , \4453 , \4454 , \4455 ,
         \4456 , \4457 , \4458 , \4459 , \4460 , \4461 , \4462 , \4463 , \4464 , \4465 ,
         \4466 , \4467 , \4468 , \4469 , \4470 , \4471 , \4472 , \4473 , \4474 , \4475 ,
         \4476 , \4477 , \4478 , \4479 , \4480 , \4481 , \4482 , \4483 , \4484 , \4485 ,
         \4486 , \4487 , \4488 , \4489 , \4490 , \4491 , \4492 , \4493 , \4494 , \4495 ,
         \4496 , \4497 , \4498 , \4499 , \4500 , \4501 , \4502 , \4503 , \4504 , \4505 ,
         \4506 , \4507 , \4508 , \4509 , \4510 , \4511 , \4512 , \4513 , \4514 , \4515 ,
         \4516 , \4517 , \4518 , \4519 , \4520 , \4521 , \4522 , \4523 , \4524 , \4525 ,
         \4526 , \4527 , \4528 , \4529 , \4530 , \4531 , \4532 , \4533 , \4534 , \4535 ,
         \4536 , \4537 , \4538 , \4539 , \4540 , \4541 , \4542 , \4543 , \4544 , \4545 ,
         \4546 , \4547 , \4548 , \4549 , \4550 , \4551 , \4552 , \4553 , \4554 , \4555 ,
         \4556 , \4557 , \4558 , \4559 , \4560 , \4561 , \4562 , \4563 , \4564 , \4565 ,
         \4566 , \4567 , \4568 , \4569 , \4570 , \4571 , \4572 , \4573 , \4574 , \4575 ,
         \4576 , \4577 , \4578 , \4579 , \4580 , \4581 , \4582 , \4583 , \4584 , \4585 ,
         \4586 , \4587 , \4588 , \4589 , \4590 , \4591 , \4592 , \4593 , \4594 , \4595 ,
         \4596 , \4597 , \4598 , \4599 , \4600 , \4601 , \4602 , \4603 , \4604 , \4605 ,
         \4606 , \4607 , \4608 , \4609 , \4610 , \4611 , \4612 , \4613 , \4614 , \4615 ,
         \4616 , \4617 , \4618 , \4619 , \4620 , \4621 , \4622 , \4623 , \4624 , \4625 ,
         \4626 , \4627 , \4628 , \4629 , \4630 , \4631 , \4632 , \4633 , \4634 , \4635 ,
         \4636 , \4637 , \4638 , \4639 , \4640 , \4641 , \4642 , \4643 , \4644 , \4645 ,
         \4646 , \4647 , \4648 , \4649 , \4650 , \4651 , \4652 , \4653 , \4654 , \4655 ,
         \4656 , \4657 , \4658 , \4659 , \4660 , \4661 , \4662 , \4663 , \4664 , \4665 ,
         \4666 , \4667 , \4668 , \4669 , \4670 , \4671 , \4672 , \4673 , \4674 , \4675 ,
         \4676 , \4677 , \4678 , \4679 , \4680 , \4681 , \4682 , \4683 , \4684 , \4685 ,
         \4686 , \4687 , \4688 , \4689 , \4690 , \4691 , \4692 , \4693 , \4694 , \4695 ,
         \4696 , \4697 , \4698 , \4699 , \4700 , \4701 , \4702 , \4703 , \4704 , \4705 ,
         \4706 , \4707 , \4708 , \4709 , \4710 , \4711 , \4712 , \4713 , \4714 , \4715 ,
         \4716 , \4717 , \4718 , \4719 , \4720 , \4721 , \4722 , \4723 , \4724 , \4725 ,
         \4726 , \4727 , \4728 , \4729 , \4730 , \4731 , \4732 , \4733 , \4734 , \4735 ,
         \4736 , \4737 , \4738 , \4739 , \4740 , \4741 , \4742 , \4743 , \4744 , \4745 ,
         \4746 , \4747 , \4748 , \4749 , \4750 , \4751 , \4752 , \4753 , \4754 , \4755 ,
         \4756 , \4757 , \4758 , \4759 , \4760 , \4761 , \4762 , \4763 , \4764 , \4765 ,
         \4766 , \4767 , \4768 , \4769 , \4770 , \4771 , \4772 , \4773 , \4774 , \4775 ,
         \4776 , \4777 , \4778 , \4779 , \4780 , \4781 , \4782 , \4783 , \4784 , \4785 ,
         \4786 , \4787 , \4788 , \4789 , \4790 , \4791 , \4792 , \4793 , \4794 , \4795 ,
         \4796 , \4797 , \4798 , \4799 , \4800 , \4801 , \4802 , \4803 , \4804 , \4805 ,
         \4806 , \4807 , \4808 , \4809 , \4810 , \4811 , \4812 , \4813 , \4814 , \4815 ,
         \4816 , \4817 , \4818 , \4819 , \4820 , \4821 , \4822 , \4823 , \4824 , \4825 ,
         \4826 , \4827 , \4828 , \4829 , \4830 , \4831 , \4832 , \4833 , \4834 , \4835 ,
         \4836 , \4837 , \4838 , \4839 , \4840 , \4841 , \4842 , \4843 , \4844 , \4845 ,
         \4846 , \4847 , \4848 , \4849 , \4850 , \4851 , \4852 , \4853 , \4854 , \4855 ,
         \4856 , \4857 , \4858 , \4859 , \4860 , \4861 , \4862 , \4863 , \4864 , \4865 ,
         \4866 , \4867 , \4868 , \4869 , \4870 , \4871 , \4872 , \4873 , \4874 , \4875 ,
         \4876 , \4877 , \4878 , \4879 , \4880 , \4881 , \4882 , \4883 , \4884 , \4885 ,
         \4886 , \4887 , \4888 , \4889 , \4890 , \4891 , \4892 , \4893 , \4894 , \4895 ,
         \4896 , \4897 , \4898 , \4899 , \4900 , \4901 , \4902 , \4903 , \4904 , \4905 ,
         \4906 , \4907 , \4908 , \4909 , \4910 , \4911 , \4912 , \4913 , \4914 , \4915 ,
         \4916 , \4917 , \4918 , \4919 , \4920 , \4921 , \4922 , \4923 , \4924 , \4925 ,
         \4926 , \4927 , \4928 , \4929 , \4930 , \4931 , \4932 , \4933 , \4934 , \4935 ,
         \4936 , \4937 , \4938 , \4939 , \4940 , \4941 , \4942 , \4943 , \4944 , \4945 ,
         \4946 , \4947 , \4948 , \4949 , \4950 , \4951 , \4952 , \4953 , \4954 , \4955 ,
         \4956 , \4957 , \4958 , \4959 , \4960 , \4961 , \4962 , \4963 , \4964 , \4965 ,
         \4966 , \4967 , \4968 , \4969 , \4970 , \4971 , \4972 , \4973 , \4974 , \4975 ,
         \4976 , \4977 , \4978 , \4979 , \4980 , \4981 , \4982 , \4983 , \4984 , \4985 ,
         \4986 , \4987 , \4988 , \4989 , \4990 , \4991 , \4992 , \4993 , \4994 , \4995 ,
         \4996 , \4997 , \4998 , \4999 , \5000 , \5001 , \5002 , \5003 , \5004 , \5005 ,
         \5006 , \5007 , \5008 , \5009 , \5010 , \5011 , \5012 , \5013 , \5014 , \5015 ,
         \5016 , \5017 , \5018 , \5019 , \5020 , \5021 , \5022 , \5023 , \5024 , \5025 ,
         \5026 , \5027 , \5028 , \5029 , \5030 , \5031 , \5032 , \5033 , \5034 , \5035 ,
         \5036 , \5037 , \5038 , \5039 , \5040 , \5041 , \5042 , \5043 , \5044 , \5045 ,
         \5046 , \5047 , \5048 , \5049 , \5050 , \5051 , \5052 , \5053 , \5054 , \5055 ,
         \5056 , \5057 , \5058 , \5059 , \5060 , \5061 , \5062 , \5063 , \5064 , \5065 ,
         \5066 , \5067 , \5068 , \5069 , \5070 , \5071 , \5072 , \5073 , \5074 , \5075 ,
         \5076 , \5077 , \5078 , \5079 , \5080 , \5081 , \5082 , \5083 , \5084 , \5085 ,
         \5086 , \5087 , \5088 , \5089 , \5090 , \5091 , \5092 , \5093 , \5094 , \5095 ,
         \5096 , \5097 , \5098 , \5099 , \5100 , \5101 , \5102 , \5103 , \5104 , \5105 ,
         \5106 , \5107 , \5108 , \5109 , \5110 , \5111 , \5112 , \5113 , \5114 , \5115 ,
         \5116 , \5117 , \5118 , \5119 , \5120 , \5121 , \5122 , \5123 , \5124 , \5125 ,
         \5126 , \5127 , \5128 , \5129 , \5130 , \5131 , \5132 , \5133 , \5134 , \5135 ,
         \5136 , \5137 , \5138 , \5139 , \5140 , \5141 , \5142 , \5143 , \5144 , \5145 ,
         \5146 , \5147 , \5148 , \5149 , \5150 , \5151 , \5152 , \5153 , \5154 , \5155 ,
         \5156 , \5157 , \5158 , \5159 , \5160 , \5161 , \5162 , \5163 , \5164 , \5165 ,
         \5166 , \5167 , \5168 , \5169 , \5170 , \5171 , \5172 , \5173 , \5174 , \5175 ,
         \5176 , \5177 , \5178 , \5179 , \5180 , \5181 , \5182 , \5183 , \5184 , \5185 ,
         \5186 , \5187 , \5188 , \5189 , \5190 , \5191 , \5192 , \5193 , \5194 , \5195 ,
         \5196 , \5197 , \5198 , \5199 , \5200 , \5201 , \5202 , \5203 , \5204 , \5205 ,
         \5206 , \5207 , \5208 , \5209 , \5210 , \5211 , \5212 , \5213 , \5214 , \5215 ,
         \5216 , \5217 , \5218 , \5219 , \5220 , \5221 , \5222 , \5223 , \5224 , \5225 ,
         \5226 , \5227 , \5228 , \5229 , \5230 , \5231 , \5232 , \5233 , \5234 , \5235 ,
         \5236 , \5237 , \5238 , \5239 , \5240 , \5241 , \5242 , \5243 , \5244 , \5245 ,
         \5246 , \5247 , \5248 , \5249 , \5250 , \5251 , \5252 , \5253 , \5254 , \5255 ,
         \5256 , \5257 , \5258 , \5259 , \5260 , \5261 , \5262 , \5263 , \5264 , \5265 ,
         \5266 , \5267 , \5268 , \5269 , \5270 , \5271 , \5272 , \5273 , \5274 , \5275 ,
         \5276 , \5277 , \5278 , \5279 , \5280 , \5281 , \5282 , \5283 , \5284 , \5285 ,
         \5286 , \5287 , \5288 , \5289 , \5290 , \5291 , \5292 , \5293 , \5294 , \5295 ,
         \5296 , \5297 , \5298 , \5299 , \5300 , \5301 , \5302 , \5303 , \5304 , \5305 ,
         \5306 , \5307 , \5308 , \5309 , \5310 , \5311 , \5312 , \5313 , \5314 , \5315 ,
         \5316 , \5317 , \5318 , \5319 , \5320 , \5321 , \5322 , \5323 , \5324 , \5325 ,
         \5326 , \5327 , \5328 , \5329 , \5330 , \5331 , \5332 , \5333 , \5334 , \5335 ,
         \5336 , \5337 , \5338 , \5339 , \5340 , \5341 , \5342 , \5343 , \5344 , \5345 ,
         \5346 , \5347 , \5348 , \5349 , \5350 , \5351 , \5352 , \5353 , \5354 , \5355 ,
         \5356 , \5357 , \5358 , \5359 , \5360 , \5361 , \5362 , \5363 , \5364 , \5365 ,
         \5366 , \5367 , \5368 , \5369 , \5370 , \5371 , \5372 , \5373 , \5374 , \5375 ,
         \5376 , \5377 , \5378 , \5379 , \5380 , \5381 , \5382 , \5383 , \5384 , \5385 ,
         \5386 , \5387 , \5388 , \5389 , \5390 , \5391 , \5392 , \5393 , \5394 , \5395 ,
         \5396 , \5397 , \5398 , \5399 , \5400 , \5401 , \5402 , \5403 , \5404 , \5405 ,
         \5406 , \5407 , \5408 , \5409 , \5410 , \5411 , \5412 , \5413 , \5414 , \5415 ,
         \5416 , \5417 , \5418 , \5419 , \5420 , \5421 , \5422 , \5423 , \5424 , \5425 ,
         \5426 , \5427 , \5428 , \5429 , \5430 , \5431 , \5432 , \5433 , \5434 , \5435 ,
         \5436 , \5437 , \5438 , \5439 , \5440 , \5441 , \5442 , \5443 , \5444 , \5445 ,
         \5446 , \5447 , \5448 , \5449 , \5450 , \5451 , \5452 , \5453 , \5454 , \5455 ,
         \5456 , \5457 , \5458 , \5459 , \5460 , \5461 , \5462 , \5463 , \5464 , \5465 ,
         \5466 , \5467 , \5468 , \5469 , \5470 , \5471 , \5472 , \5473 , \5474 , \5475 ,
         \5476 , \5477 , \5478 , \5479 , \5480 , \5481 , \5482 , \5483 , \5484 , \5485 ,
         \5486 , \5487 , \5488 , \5489 , \5490 , \5491 , \5492 , \5493 , \5494 , \5495 ,
         \5496 , \5497 , \5498 , \5499 , \5500 , \5501 , \5502 , \5503 , \5504 , \5505 ,
         \5506 , \5507 , \5508 , \5509 , \5510 , \5511 , \5512 , \5513 , \5514 , \5515 ,
         \5516 , \5517 , \5518 , \5519 , \5520 , \5521 , \5522 , \5523 , \5524 , \5525 ,
         \5526 , \5527 , \5528 , \5529 , \5530 , \5531 , \5532 , \5533 , \5534 , \5535 ,
         \5536 , \5537 , \5538 , \5539 , \5540 , \5541 , \5542 , \5543 , \5544 , \5545 ,
         \5546 , \5547 , \5548 , \5549 , \5550 , \5551 , \5552 , \5553 , \5554 , \5555 ,
         \5556 , \5557 , \5558 , \5559 , \5560 , \5561 , \5562 , \5563 , \5564 , \5565 ,
         \5566 , \5567 , \5568 , \5569 , \5570 , \5571 , \5572 , \5573 , \5574 , \5575 ,
         \5576 , \5577 , \5578 , \5579 , \5580 , \5581 , \5582 , \5583 , \5584 , \5585 ,
         \5586 , \5587 , \5588 , \5589 , \5590 , \5591 , \5592 , \5593 , \5594 , \5595 ,
         \5596 , \5597 , \5598 , \5599 , \5600 , \5601 , \5602 , \5603 , \5604 , \5605 ,
         \5606 , \5607 , \5608 , \5609 , \5610 , \5611 , \5612 , \5613 , \5614 , \5615 ,
         \5616 , \5617 , \5618 , \5619 , \5620 , \5621 , \5622 , \5623 , \5624 , \5625 ,
         \5626 , \5627 , \5628 , \5629 , \5630 , \5631 , \5632 , \5633 , \5634 , \5635 ,
         \5636 , \5637 , \5638 , \5639 , \5640 , \5641 , \5642 , \5643 , \5644 , \5645 ,
         \5646 , \5647 , \5648 , \5649 , \5650 , \5651 , \5652 , \5653 , \5654 , \5655 ,
         \5656 , \5657 , \5658 , \5659 , \5660 , \5661 , \5662 , \5663 , \5664 , \5665 ,
         \5666 , \5667 , \5668 , \5669 , \5670 , \5671 , \5672 , \5673 , \5674 , \5675 ,
         \5676 , \5677 , \5678 , \5679 , \5680 , \5681 , \5682 , \5683 , \5684 , \5685 ,
         \5686 , \5687 , \5688 , \5689 , \5690 , \5691 , \5692 , \5693 , \5694 , \5695 ,
         \5696 , \5697 , \5698 , \5699 , \5700 , \5701 , \5702 , \5703 , \5704 , \5705 ,
         \5706 , \5707 , \5708 , \5709 , \5710 , \5711 , \5712 , \5713 , \5714 , \5715 ,
         \5716 , \5717 , \5718 , \5719 , \5720 , \5721 , \5722 , \5723 , \5724 , \5725 ,
         \5726 , \5727 , \5728 , \5729 , \5730 , \5731 , \5732 , \5733 , \5734 , \5735 ,
         \5736 , \5737 , \5738 , \5739 , \5740 , \5741 , \5742 , \5743 , \5744 , \5745 ,
         \5746 , \5747 , \5748 , \5749 , \5750 , \5751 , \5752 , \5753 , \5754 , \5755 ,
         \5756 , \5757 , \5758 , \5759 , \5760 , \5761 , \5762 , \5763 , \5764 , \5765 ,
         \5766 , \5767 , \5768 , \5769 , \5770 , \5771 , \5772 , \5773 , \5774 , \5775 ,
         \5776 , \5777 , \5778 , \5779 , \5780 , \5781 , \5782 , \5783 , \5784 , \5785 ,
         \5786 , \5787 , \5788 , \5789 , \5790 , \5791 , \5792 , \5793 , \5794 , \5795 ,
         \5796 , \5797 , \5798 , \5799 , \5800 , \5801 , \5802 , \5803 , \5804 , \5805 ,
         \5806 , \5807 , \5808 , \5809 , \5810 , \5811 , \5812 , \5813 , \5814 , \5815 ,
         \5816 , \5817 , \5818 , \5819 , \5820 , \5821 , \5822 , \5823 , \5824 , \5825 ,
         \5826 , \5827 , \5828 , \5829 , \5830 , \5831 , \5832 , \5833 , \5834 , \5835 ,
         \5836 , \5837 , \5838 , \5839 , \5840 , \5841 , \5842 , \5843 , \5844 , \5845 ,
         \5846 , \5847 , \5848 , \5849 , \5850 , \5851 , \5852 , \5853 , \5854 , \5855 ,
         \5856 , \5857 , \5858 , \5859 , \5860 , \5861 , \5862 , \5863 , \5864 , \5865 ,
         \5866 , \5867 , \5868 , \5869 , \5870 , \5871 , \5872 , \5873 , \5874 , \5875 ,
         \5876 , \5877 , \5878 , \5879 , \5880 , \5881 , \5882 , \5883 , \5884 , \5885 ,
         \5886 , \5887 , \5888 , \5889 , \5890 , \5891 , \5892 , \5893 , \5894 , \5895 ,
         \5896 , \5897 , \5898 , \5899 , \5900 , \5901 , \5902 , \5903 , \5904 , \5905 ,
         \5906 , \5907 , \5908 , \5909 , \5910 , \5911 , \5912 , \5913 , \5914 , \5915 ,
         \5916 , \5917 , \5918 , \5919 , \5920 , \5921 , \5922 , \5923 , \5924 , \5925 ,
         \5926 , \5927 , \5928 , \5929 , \5930 , \5931 , \5932 , \5933 , \5934 , \5935 ,
         \5936 , \5937 , \5938 , \5939 , \5940 , \5941 , \5942 , \5943 , \5944 , \5945 ,
         \5946 , \5947 , \5948 , \5949 , \5950 , \5951 , \5952 , \5953 , \5954 , \5955 ,
         \5956 , \5957 , \5958 , \5959 , \5960 , \5961 , \5962 , \5963 , \5964 , \5965 ,
         \5966 , \5967 , \5968 , \5969 , \5970 , \5971 , \5972 , \5973 , \5974 , \5975 ,
         \5976 , \5977 , \5978 , \5979 , \5980 , \5981 , \5982 , \5983 , \5984 , \5985 ,
         \5986 , \5987 , \5988 , \5989 , \5990 , \5991 , \5992 , \5993 , \5994 , \5995 ,
         \5996 , \5997 , \5998 , \5999 , \6000 , \6001 , \6002 , \6003 , \6004 , \6005 ,
         \6006 , \6007 , \6008 , \6009 , \6010 , \6011 , \6012 , \6013 , \6014 , \6015 ,
         \6016 , \6017 , \6018 , \6019 , \6020 , \6021 , \6022 , \6023 , \6024 , \6025 ,
         \6026 , \6027 , \6028 , \6029 , \6030 , \6031 , \6032 , \6033 , \6034 , \6035 ,
         \6036 , \6037 , \6038 , \6039 , \6040 , \6041 , \6042 , \6043 , \6044 , \6045 ,
         \6046 , \6047 , \6048 , \6049 , \6050 , \6051 , \6052 , \6053 , \6054 , \6055 ,
         \6056 , \6057 , \6058 , \6059 , \6060 , \6061 , \6062 , \6063 , \6064 , \6065 ,
         \6066 , \6067 , \6068 , \6069 , \6070 , \6071 , \6072 , \6073 , \6074 , \6075 ,
         \6076 , \6077 , \6078 , \6079 , \6080 , \6081 , \6082 , \6083 , \6084 , \6085 ,
         \6086 , \6087 , \6088 , \6089 , \6090 , \6091 , \6092 , \6093 , \6094 , \6095 ,
         \6096 , \6097 , \6098 , \6099 , \6100 , \6101 , \6102 , \6103 , \6104 , \6105 ,
         \6106 , \6107 , \6108 , \6109 , \6110 , \6111 , \6112 , \6113 , \6114 , \6115 ,
         \6116 , \6117 , \6118 , \6119 , \6120 , \6121 , \6122 , \6123 , \6124 , \6125 ,
         \6126 , \6127 , \6128 , \6129 , \6130 , \6131 , \6132 , \6133 , \6134 , \6135 ,
         \6136 , \6137 , \6138 , \6139 , \6140 , \6141 , \6142 , \6143 , \6144 , \6145 ,
         \6146 , \6147 , \6148 , \6149 , \6150 , \6151 , \6152 , \6153 , \6154 , \6155 ,
         \6156 , \6157 , \6158 , \6159 , \6160 , \6161 , \6162 , \6163 , \6164 , \6165 ,
         \6166 , \6167 , \6168 , \6169 , \6170 , \6171 , \6172 , \6173 , \6174 , \6175 ,
         \6176 , \6177 , \6178 , \6179 , \6180 , \6181 , \6182 , \6183 , \6184 , \6185 ,
         \6186 , \6187 , \6188 , \6189 , \6190 , \6191 , \6192 , \6193 , \6194 , \6195 ,
         \6196 , \6197 , \6198 , \6199 , \6200 , \6201 , \6202 , \6203 , \6204 , \6205 ,
         \6206 , \6207 , \6208 , \6209 , \6210 , \6211 , \6212 , \6213 , \6214 , \6215 ,
         \6216 , \6217 , \6218 , \6219 , \6220 , \6221 , \6222 , \6223 , \6224 , \6225 ,
         \6226 , \6227 , \6228 , \6229 , \6230 , \6231 , \6232 , \6233 , \6234 , \6235 ,
         \6236 , \6237 , \6238 , \6239 , \6240 , \6241 , \6242 , \6243 , \6244 , \6245 ,
         \6246 , \6247 , \6248 , \6249 , \6250 , \6251 , \6252 , \6253 , \6254 , \6255 ,
         \6256 , \6257 , \6258 , \6259 , \6260 , \6261 , \6262 , \6263 , \6264 , \6265 ,
         \6266 , \6267 , \6268 , \6269 , \6270 , \6271 , \6272 , \6273 , \6274 , \6275 ,
         \6276 , \6277 , \6278 , \6279 , \6280 , \6281 , \6282 , \6283 , \6284 , \6285 ,
         \6286 , \6287 , \6288 , \6289 , \6290 , \6291 , \6292 , \6293 , \6294 , \6295 ,
         \6296 , \6297 , \6298 , \6299 , \6300 , \6301 , \6302 , \6303 , \6304 , \6305 ,
         \6306 , \6307 , \6308 , \6309 , \6310 , \6311 , \6312 , \6313 , \6314 , \6315 ,
         \6316 , \6317 , \6318 , \6319 , \6320 , \6321 , \6322 , \6323 , \6324 , \6325 ,
         \6326 , \6327 , \6328 , \6329 , \6330 , \6331 , \6332 , \6333 , \6334 , \6335 ,
         \6336 , \6337 , \6338 , \6339 , \6340 , \6341 , \6342 , \6343 , \6344 , \6345 ,
         \6346 , \6347 , \6348 , \6349 , \6350 , \6351 , \6352 , \6353 , \6354 , \6355 ,
         \6356 , \6357 , \6358 , \6359 , \6360 , \6361 , \6362 , \6363 , \6364 , \6365 ,
         \6366 , \6367 , \6368 , \6369 , \6370 , \6371 , \6372 , \6373 , \6374 , \6375 ,
         \6376 , \6377 , \6378 , \6379 , \6380 , \6381 , \6382 , \6383 , \6384 , \6385 ,
         \6386 , \6387 , \6388 , \6389 , \6390 , \6391 , \6392 , \6393 , \6394 , \6395 ,
         \6396 , \6397 , \6398 , \6399 , \6400 , \6401 , \6402 , \6403 , \6404 , \6405 ,
         \6406 , \6407 , \6408 , \6409 , \6410 , \6411 , \6412 , \6413 , \6414 , \6415 ,
         \6416 , \6417 , \6418 , \6419 , \6420 , \6421 , \6422 , \6423 , \6424 , \6425 ,
         \6426 , \6427 , \6428 , \6429 , \6430 , \6431 , \6432 , \6433 , \6434 , \6435 ,
         \6436 , \6437 , \6438 , \6439 , \6440 , \6441 , \6442 , \6443 , \6444 , \6445 ,
         \6446 , \6447 , \6448 , \6449 , \6450 , \6451 , \6452 , \6453 , \6454 , \6455 ,
         \6456 , \6457 , \6458 , \6459 , \6460 , \6461 , \6462 , \6463 , \6464 , \6465 ,
         \6466 , \6467 , \6468 , \6469 , \6470 , \6471 , \6472 , \6473 , \6474 , \6475 ,
         \6476 , \6477 , \6478 , \6479 , \6480 , \6481 , \6482 , \6483 , \6484 , \6485 ,
         \6486 , \6487 , \6488 , \6489 , \6490 , \6491 , \6492 , \6493 , \6494 , \6495 ,
         \6496 , \6497 , \6498 , \6499 , \6500 , \6501 , \6502 , \6503 , \6504 , \6505 ,
         \6506 , \6507 , \6508 , \6509 , \6510 , \6511 , \6512 , \6513 , \6514 , \6515 ,
         \6516 , \6517 , \6518 , \6519 , \6520 , \6521 , \6522 , \6523 , \6524 , \6525 ,
         \6526 , \6527 , \6528 , \6529 , \6530 , \6531 , \6532 , \6533 , \6534 , \6535 ,
         \6536 , \6537 , \6538 , \6539 , \6540 , \6541 , \6542 , \6543 , \6544 , \6545 ,
         \6546 , \6547 , \6548 , \6549 , \6550 , \6551 , \6552 , \6553 , \6554 , \6555 ,
         \6556 , \6557 , \6558 , \6559 , \6560 , \6561 , \6562 , \6563 , \6564 , \6565 ,
         \6566 , \6567 , \6568 , \6569 , \6570 , \6571 , \6572 , \6573 , \6574 , \6575 ,
         \6576 , \6577 , \6578 , \6579 , \6580 , \6581 , \6582 , \6583 , \6584 , \6585 ,
         \6586 , \6587 , \6588 , \6589 , \6590 , \6591 , \6592 , \6593 , \6594 , \6595 ,
         \6596 , \6597 , \6598 , \6599 , \6600 , \6601 , \6602 , \6603 , \6604 , \6605 ,
         \6606 , \6607 , \6608 , \6609 , \6610 , \6611 , \6612 , \6613 , \6614 , \6615 ,
         \6616 , \6617 , \6618 , \6619 , \6620 , \6621 , \6622 , \6623 , \6624 , \6625 ,
         \6626 , \6627 , \6628 , \6629 , \6630 , \6631 , \6632 , \6633 , \6634 , \6635 ,
         \6636 , \6637 , \6638 , \6639 , \6640 , \6641 , \6642 , \6643 , \6644 , \6645 ,
         \6646 , \6647 , \6648 , \6649 , \6650 , \6651 , \6652 , \6653 , \6654 , \6655 ,
         \6656 , \6657 , \6658 , \6659 , \6660 , \6661 , \6662 , \6663 , \6664 , \6665 ,
         \6666 , \6667 , \6668 , \6669 , \6670 , \6671 , \6672 , \6673 , \6674 , \6675 ,
         \6676 , \6677 , \6678 , \6679 , \6680 , \6681 , \6682 , \6683 , \6684 , \6685 ,
         \6686 , \6687 , \6688 , \6689 , \6690 , \6691 , \6692 , \6693 , \6694 , \6695 ,
         \6696 , \6697 , \6698 , \6699 , \6700 , \6701 , \6702 , \6703 , \6704 , \6705 ,
         \6706 , \6707 , \6708 , \6709 , \6710 , \6711 , \6712 , \6713 , \6714 , \6715 ,
         \6716 , \6717 , \6718 , \6719 , \6720 , \6721 , \6722 , \6723 , \6724 , \6725 ,
         \6726 , \6727 , \6728 , \6729 , \6730 , \6731 , \6732 , \6733 , \6734 , \6735 ,
         \6736 , \6737 , \6738 , \6739 , \6740 , \6741 , \6742 , \6743 , \6744 , \6745 ,
         \6746 , \6747 , \6748 , \6749 , \6750 , \6751 , \6752 , \6753 , \6754 , \6755 ,
         \6756 , \6757 , \6758 , \6759 , \6760 , \6761 , \6762 , \6763 , \6764 , \6765 ,
         \6766 , \6767 , \6768 , \6769 , \6770 , \6771 , \6772 , \6773 , \6774 , \6775 ,
         \6776 , \6777 , \6778 , \6779 , \6780 , \6781 , \6782 , \6783 , \6784 , \6785 ,
         \6786 , \6787 , \6788 , \6789 , \6790 , \6791 , \6792 , \6793 , \6794 , \6795 ,
         \6796 , \6797 , \6798 , \6799 , \6800 , \6801 , \6802 , \6803 , \6804 , \6805 ,
         \6806 , \6807 , \6808 , \6809 , \6810 , \6811 , \6812 , \6813 , \6814 , \6815 ,
         \6816 , \6817 , \6818 , \6819 , \6820 , \6821 , \6822 , \6823 , \6824 , \6825 ,
         \6826 , \6827 , \6828 , \6829 , \6830 , \6831 , \6832 , \6833 , \6834 , \6835 ,
         \6836 , \6837 , \6838 , \6839 , \6840 , \6841 , \6842 , \6843 , \6844 , \6845 ,
         \6846 , \6847 , \6848 , \6849 , \6850 , \6851 , \6852 , \6853 , \6854 , \6855 ,
         \6856 , \6857 , \6858 , \6859 , \6860 , \6861 , \6862 , \6863 , \6864 , \6865 ,
         \6866 , \6867 , \6868 , \6869 , \6870 , \6871 , \6872 , \6873 , \6874 , \6875 ,
         \6876 , \6877 , \6878 , \6879 , \6880 , \6881 , \6882 , \6883 , \6884 , \6885 ,
         \6886 , \6887 , \6888 , \6889 , \6890 , \6891 , \6892 , \6893 , \6894 , \6895 ,
         \6896 , \6897 , \6898 , \6899 , \6900 , \6901 , \6902 , \6903 , \6904 , \6905 ,
         \6906 , \6907 , \6908 , \6909 , \6910 , \6911 , \6912 , \6913 , \6914 , \6915 ,
         \6916 , \6917 , \6918 , \6919 , \6920 , \6921 , \6922 , \6923 , \6924 , \6925 ,
         \6926 , \6927 , \6928 , \6929 , \6930 , \6931 , \6932 , \6933 , \6934 , \6935 ,
         \6936 , \6937 , \6938 , \6939 , \6940 , \6941 , \6942 , \6943 , \6944 , \6945 ,
         \6946 , \6947 , \6948 , \6949 , \6950 , \6951 , \6952 , \6953 , \6954 , \6955 ,
         \6956 , \6957 , \6958 , \6959 , \6960 , \6961 , \6962 , \6963 , \6964 , \6965 ,
         \6966 , \6967 , \6968 , \6969 , \6970 , \6971 , \6972 , \6973 , \6974 , \6975 ,
         \6976 , \6977 , \6978 , \6979 , \6980 , \6981 , \6982 , \6983 , \6984 , \6985 ,
         \6986 , \6987 , \6988 , \6989 , \6990 , \6991 , \6992 , \6993 , \6994 , \6995 ,
         \6996 , \6997 , \6998 , \6999 , \7000 , \7001 , \7002 , \7003 , \7004 , \7005 ,
         \7006 , \7007 , \7008 , \7009 , \7010 , \7011 , \7012 , \7013 , \7014 , \7015 ,
         \7016 , \7017 , \7018 , \7019 , \7020 , \7021 , \7022 , \7023 , \7024 , \7025 ,
         \7026 , \7027 , \7028 , \7029 , \7030 , \7031 , \7032 , \7033 , \7034 , \7035 ,
         \7036 , \7037 , \7038 , \7039 , \7040 , \7041 , \7042 , \7043 , \7044 , \7045 ,
         \7046 , \7047 , \7048 , \7049 , \7050 , \7051 , \7052 , \7053 , \7054 , \7055 ,
         \7056 , \7057 , \7058 , \7059 , \7060 , \7061 , \7062 , \7063 , \7064 , \7065 ,
         \7066 , \7067 , \7068 , \7069 , \7070 , \7071 , \7072 , \7073 , \7074 , \7075 ,
         \7076 , \7077 , \7078 , \7079 , \7080 , \7081 , \7082 , \7083 , \7084 , \7085 ,
         \7086 , \7087 , \7088 , \7089 , \7090 , \7091 , \7092 , \7093 , \7094 , \7095 ,
         \7096 , \7097 , \7098 , \7099 , \7100 , \7101 , \7102 , \7103 , \7104 , \7105 ,
         \7106 , \7107 , \7108 , \7109 , \7110 , \7111 , \7112 , \7113 , \7114 , \7115 ,
         \7116 , \7117 , \7118 , \7119 , \7120 , \7121 , \7122 , \7123 , \7124 , \7125 ,
         \7126 , \7127 , \7128 , \7129 , \7130 , \7131 , \7132 , \7133 , \7134 , \7135 ,
         \7136 , \7137 , \7138 , \7139 , \7140 , \7141 , \7142 , \7143 , \7144 , \7145 ,
         \7146 , \7147 , \7148 , \7149 , \7150 , \7151 , \7152 , \7153 , \7154 , \7155 ,
         \7156 , \7157 , \7158 , \7159 , \7160 , \7161 , \7162 , \7163 , \7164 , \7165 ,
         \7166 , \7167 , \7168 , \7169 , \7170 , \7171 , \7172 , \7173 , \7174 , \7175 ,
         \7176 , \7177 , \7178 , \7179 , \7180 , \7181 , \7182 , \7183 , \7184 , \7185 ,
         \7186 , \7187 , \7188 , \7189 , \7190 , \7191 , \7192 , \7193 , \7194 , \7195 ,
         \7196 , \7197 , \7198 , \7199 , \7200 , \7201 , \7202 , \7203 , \7204 , \7205 ,
         \7206 , \7207 , \7208 , \7209 , \7210 , \7211 , \7212 , \7213 , \7214 , \7215 ,
         \7216 ;
buf \U$labaj739 ( \o[31] , \6967 );
buf \U$labaj740 ( \o[30] , \7061 );
buf \U$labaj741 ( \o[29] , \6979 );
buf \U$labaj742 ( \o[28] , \6991 );
buf \U$labaj743 ( \o[27] , \7007 );
buf \U$labaj744 ( \o[26] , \7020 );
buf \U$labaj745 ( \o[25] , \7030 );
buf \U$labaj746 ( \o[24] , \7216 );
buf \U$labaj747 ( \o[23] , \7046 );
buf \U$labaj748 ( \o[22] , \7206 );
buf \U$labaj749 ( \o[21] , \7072 );
buf \U$labaj750 ( \o[20] , \7078 );
buf \U$labaj751 ( \o[19] , \7095 );
buf \U$labaj752 ( \o[18] , \7102 );
buf \U$labaj753 ( \o[17] , \7112 );
buf \U$labaj754 ( \o[16] , \7118 );
buf \U$labaj755 ( \o[15] , \7132 );
buf \U$labaj756 ( \o[14] , \7138 );
buf \U$labaj757 ( \o[13] , \7147 );
buf \U$labaj758 ( \o[12] , \7154 );
buf \U$labaj759 ( \o[11] , \7171 );
buf \U$labaj760 ( \o[10] , \7178 );
buf \U$labaj761 ( \o[9] , \7188 );
buf \U$labaj762 ( \o[8] , \7194 );
buf \U$labaj763 ( \o[7] , \7215 );
buf \U$labaj764 ( \o[6] , \7207 );
buf \U$labaj765 ( \o[5] , \7210 );
buf \U$labaj766 ( \o[4] , \7211 );
buf \U$labaj767 ( \o[3] , \7212 );
buf \U$labaj768 ( \o[2] , \7213 );
buf \U$labaj769 ( \o[1] , \7203 );
buf \U$labaj770 ( \o[0] , \7204 );
not \g35732/U$3 ( \99 , \a[7] );
not \g35732/U$4 ( \100 , \d[7] );
and \g35732/U$2 ( \101 , \99 , \100 );
xor \mul_6_11_g13942/U$1 ( \102 , \a[0] , \b[9] );
not \mul_6_11_g13735/U$3 ( \103 , \102 );
xor \mul_6_11_g35491/U$1 ( \104 , \b[8] , \b[7] );
xnor \mul_6_11_g13984/U$1 ( \105 , \b[9] , \b[8] );
nor \mul_6_11_g13868/U$1 ( \106 , \104 , \105 );
not \mul_6_11_g13735/U$4 ( \107 , \106 );
or \mul_6_11_g13735/U$2 ( \108 , \103 , \107 );
xor \mul_6_11_g13947/U$1 ( \109 , \a[1] , \b[9] );
nand \mul_6_11_g13812/U$1 ( \110 , \104 , \109 );
nand \mul_6_11_g13735/U$1 ( \111 , \108 , \110 );
or \mul_6_11_g13875/U$2 ( \112 , \a[0] , \b[8] );
nand \mul_6_11_g13875/U$1 ( \113 , \112 , \b[7] );
nand \mul_6_11_g13956/U$1 ( \114 , \a[0] , \b[8] );
and \mul_6_11_g13982/U$1 ( \115 , \113 , \114 , \b[9] );
xor \mul_6_11_g14016/U$1 ( \116 , \a[4] , \b[5] );
xor \mul_6_11_g13976/U$1 ( \117 , \b[5] , \b[4] );
nand \mul_6_11_g13826/U$1 ( \118 , \116 , \117 );
xor \mul_6_11_g35494/U$1 ( \119 , \b[4] , \b[3] );
or \g35917/U$2 ( \120 , \118 , \119 );
xor \mul_6_11_g13974/U$1 ( \121 , \b[4] , \b[3] );
xor \mul_6_11_g13922/U$1 ( \122 , \a[5] , \b[5] );
nand \mul_6_11_g13802/U$1 ( \123 , \121 , \122 );
nand \g35917/U$1 ( \124 , \120 , \123 );
xor \mul_6_11_g13686/U$1 ( \125 , \115 , \124 );
xor \g35624/U$1 ( \126 , \111 , \125 );
nand \mul_6_11_g13840/U$1 ( \127 , \104 , \a[0] );
not \mul_6_11_g35696/U$1 ( \128 , \127 );
xor \mul_6_11_g13887/U$1 ( \129 , \a[7] , \b[1] );
not \mul_6_11_g13776/U$3 ( \130 , \129 );
not \mul_6_11_g35730/U$2 ( \131 , \b[0] );
nand \mul_6_11_g35730/U$1 ( \132 , \131 , \b[1] );
not \mul_6_11_g13969/U$1 ( \133 , \132 );
not \mul_6_11_g13776/U$4 ( \134 , \133 );
or \mul_6_11_g13776/U$2 ( \135 , \130 , \134 );
xor \g35753/U$1 ( \136 , \b[1] , \a[8] );
nand \mul_6_11_g13843/U$1 ( \137 , \136 , \b[0] );
nand \mul_6_11_g13776/U$1 ( \138 , \135 , \137 );
or \g35850/U$1 ( \139 , \128 , \138 );
not \mul_6_11_g13704/U$3 ( \140 , \139 );
xor \mul_6_11_g35953/U$1 ( \141 , \a[5] , \b[3] );
not \mul_6_11_g13754/U$3 ( \142 , \141 );
xnor \mul_6_11_g35613/U$1 ( \143 , \b[3] , \b[2] );
xor \mul_6_11_g35773/U$1 ( \144 , \b[2] , \b[1] );
nor \mul_6_11_g13821/U$1 ( \145 , \143 , \144 );
not \mul_6_11_g13820/U$1 ( \146 , \145 );
not \mul_6_11_g13818/U$1 ( \147 , \146 );
not \mul_6_11_g13754/U$4 ( \148 , \147 );
or \mul_6_11_g13754/U$2 ( \149 , \142 , \148 );
xor \mul_6_11_g13977/U$1 ( \150 , \b[2] , \b[1] );
xor \mul_6_11_g13896/U$1 ( \151 , \a[6] , \b[3] );
nand \mul_6_11_g13806/U$1 ( \152 , \150 , \151 );
nand \mul_6_11_g13754/U$1 ( \153 , \149 , \152 );
not \mul_6_11_g13704/U$4 ( \154 , \153 );
or \mul_6_11_g13704/U$2 ( \155 , \140 , \154 );
nand \mul_6_11_g13718/U$1 ( \156 , \138 , \128 );
nand \mul_6_11_g13704/U$1 ( \157 , \155 , \156 );
xnor \g35624/U$1_r1 ( \158 , \126 , \157 );
not \mul_6_11_g13579/U$3 ( \159 , \158 );
xor \mul_6_11_g35748/U$1 ( \160 , \a[9] , \b[1] );
and \mul_6_11_g14014/U$2 ( \161 , \160 , \b[0] );
not \g35729/U$2 ( \162 , \b[1] );
nor \g35729/U$1 ( \163 , \162 , \b[0] );
and \mul_6_11_g14014/U$3 ( \164 , \163 , \136 );
nor \mul_6_11_g14014/U$1 ( \165 , \161 , \164 );
not \mul_6_11_g13756/U$3 ( \166 , \151 );
not \mul_6_11_g13756/U$4 ( \167 , \145 );
or \mul_6_11_g13756/U$2 ( \168 , \166 , \167 );
xor \mul_6_11_g13903/U$1 ( \169 , \a[7] , \b[3] );
nand \mul_6_11_g13823/U$1 ( \170 , \150 , \169 );
nand \mul_6_11_g13756/U$1 ( \171 , \168 , \170 );
xor \mul_6_11_g13677/U$1 ( \172 , \165 , \171 );
xor \mul_6_11_g13937/U$1 ( \173 , \a[2] , \b[7] );
not \mul_6_11_g13747/U$3 ( \174 , \173 );
xor \mul_6_11_g35751/U$1 ( \175 , \b[7] , \b[6] );
not \mul_6_11_g13832/U$2 ( \176 , \175 );
xor \mul_6_11_g13975/U$1 ( \177 , \b[6] , \b[5] );
nor \mul_6_11_g13832/U$1 ( \178 , \176 , \177 );
not \mul_6_11_g13747/U$4 ( \179 , \178 );
or \mul_6_11_g13747/U$2 ( \180 , \174 , \179 );
xor \mul_6_11_g13938/U$1 ( \181 , \a[3] , \b[7] );
nand \mul_6_11_g13815/U$1 ( \182 , \177 , \181 );
nand \mul_6_11_g13747/U$1 ( \183 , \180 , \182 );
not \mul_6_11_g13746/U$1 ( \184 , \183 );
xnor \mul_6_11_g13677/U$1_r1 ( \185 , \172 , \184 );
buf \fopt35776/U$1 ( \186 , \185 );
not \mul_6_11_g13579/U$4 ( \187 , \186 );
or \mul_6_11_g13579/U$2 ( \188 , \159 , \187 );
xor \mul_6_11_g35715/U$1 ( \189 , \a[1] , \b[7] );
not \mul_6_11_g13744/U$3 ( \190 , \189 );
not \mul_6_11_g13744/U$4 ( \191 , \178 );
or \mul_6_11_g13744/U$2 ( \192 , \190 , \191 );
nand \mul_6_11_g13799/U$1 ( \193 , \173 , \177 );
nand \mul_6_11_g13744/U$1 ( \194 , \192 , \193 );
xor \mul_6_11_g35954/U$1 ( \195 , \a[3] , \b[5] );
not \mul_6_11_g13738/U$3 ( \196 , \195 );
not \mul_6_11_g13904/U$1 ( \197 , \117 );
nor \mul_6_11_g13811/U$1 ( \198 , \197 , \121 );
not \mul_6_11_g13738/U$4 ( \199 , \198 );
or \mul_6_11_g13738/U$2 ( \200 , \196 , \199 );
nand \mul_6_11_g13801/U$1 ( \201 , \121 , \116 );
nand \mul_6_11_g13738/U$1 ( \202 , \200 , \201 );
xor \mul_6_11_g13641/U$4 ( \203 , \194 , \202 );
or \mul_6_11_g13876/U$2 ( \204 , \a[0] , \b[6] );
nand \mul_6_11_g13876/U$1 ( \205 , \204 , \b[5] );
nand \mul_6_11_g13955/U$1 ( \206 , \a[0] , \b[6] );
and \mul_6_11_g13981/U$1 ( \207 , \205 , \206 , \b[7] );
not \mul_6_11_g13726/U$3 ( \208 , \141 );
not \mul_6_11_g13726/U$4 ( \209 , \150 );
or \mul_6_11_g13726/U$2 ( \210 , \208 , \209 );
not \mul_6_11_g14013/U$2 ( \211 , \144 );
xnor \mul_6_11_g13986/U$1 ( \212 , \a[4] , \b[3] );
nor \mul_6_11_g13807/U$1 ( \213 , \212 , \143 );
nand \mul_6_11_g14013/U$1 ( \214 , \211 , \213 );
nand \mul_6_11_g13726/U$1 ( \215 , \210 , \214 );
and \mul_6_11_g13691/U$2 ( \216 , \207 , \215 );
and \mul_6_11_g13641/U$3 ( \217 , \203 , \216 );
and \mul_6_11_g13641/U$5 ( \218 , \194 , \202 );
or \mul_6_11_g13641/U$2 ( \219 , \217 , \218 );
buf \fopt35789/U$1 ( \220 , \219 );
nand \mul_6_11_g13579/U$1 ( \221 , \188 , \220 );
not \mul_6_11_g13585/U$2 ( \222 , \186 );
not \mul_6_11_g13606/U$1 ( \223 , \158 );
nand \mul_6_11_g13585/U$1 ( \224 , \222 , \223 );
nand \mul_6_11_g13571/U$1 ( \225 , \221 , \224 );
not \mul_6_11_g13531/U$2 ( \226 , \225 );
not \mul_6_11_g13731/U$3 ( \227 , \109 );
nor \mul_6_11_g13867/U$1 ( \228 , \104 , \105 );
not \mul_6_11_g13731/U$4 ( \229 , \228 );
or \mul_6_11_g13731/U$2 ( \230 , \227 , \229 );
xor \mul_6_11_g13943/U$1 ( \231 , \a[2] , \b[9] );
nand \mul_6_11_g13793/U$1 ( \232 , \104 , \231 );
nand \mul_6_11_g13731/U$1 ( \233 , \230 , \232 );
not \mul_6_11_g13748/U$3 ( \234 , \181 );
not \mul_6_11_g13748/U$4 ( \235 , \178 );
or \mul_6_11_g13748/U$2 ( \236 , \234 , \235 );
xor \mul_6_11_g13926/U$1 ( \237 , \a[4] , \b[7] );
nand \mul_6_11_g13827/U$1 ( \238 , \177 , \237 );
nand \mul_6_11_g13748/U$1 ( \239 , \236 , \238 );
xor \mul_6_11_g13655/U$1 ( \240 , \233 , \239 );
not \mul_6_11_g13760/U$3 ( \241 , \169 );
not \mul_6_11_g13819/U$1 ( \242 , \146 );
not \mul_6_11_g13760/U$4 ( \243 , \242 );
or \mul_6_11_g13760/U$2 ( \244 , \241 , \243 );
xor \mul_6_11_g13895/U$1 ( \245 , \a[8] , \b[3] );
nand \mul_6_11_g13856/U$1 ( \246 , \150 , \245 );
nand \mul_6_11_g13760/U$1 ( \247 , \244 , \246 );
xor \mul_6_11_g13655/U$1_r1 ( \248 , \240 , \247 );
not \mul_6_11_g13615/U$3 ( \249 , \111 );
not \mul_6_11_g13615/U$4 ( \250 , \125 );
or \mul_6_11_g13615/U$2 ( \251 , \249 , \250 );
or \g35915/U$2 ( \252 , \125 , \111 );
nand \g35915/U$1 ( \253 , \252 , \157 );
nand \mul_6_11_g13615/U$1 ( \254 , \251 , \253 );
xor \mul_6_11_g13555/U$1 ( \255 , \248 , \254 );
and \mul_6_11_g13686/U$2 ( \256 , \115 , \124 );
xor \mul_6_11_g13916/U$1 ( \257 , \b[10] , \b[9] );
and \mul_6_11_g13805/U$1 ( \258 , \257 , \a[0] );
not \mul_6_11_g13767/U$3 ( \259 , \160 );
not \mul_6_11_g13767/U$4 ( \260 , \163 );
or \mul_6_11_g13767/U$2 ( \261 , \259 , \260 );
xor \mul_6_11_g13894/U$1 ( \262 , \a[10] , \b[1] );
nand \mul_6_11_g13842/U$1 ( \263 , \b[0] , \262 );
nand \mul_6_11_g13767/U$1 ( \264 , \261 , \263 );
xor \mul_6_11_g13662/U$1 ( \265 , \258 , \264 );
not \mul_6_11_g13739/U$3 ( \266 , \122 );
nor \mul_6_11_g13810/U$1 ( \267 , \119 , \197 );
not \mul_6_11_g13739/U$4 ( \268 , \267 );
or \mul_6_11_g13739/U$2 ( \269 , \266 , \268 );
xor \mul_6_11_g13907/U$1 ( \270 , \a[6] , \b[5] );
nand \mul_6_11_g13808/U$1 ( \271 , \121 , \270 );
nand \mul_6_11_g13739/U$1 ( \272 , \269 , \271 );
xor \mul_6_11_g13662/U$1_r1 ( \273 , \265 , \272 );
xor \mul_6_11_g13592/U$1 ( \274 , \256 , \273 );
not \mul_6_11_g13693/U$3 ( \275 , \165 );
not \mul_6_11_g13693/U$4 ( \276 , \184 );
or \mul_6_11_g13693/U$2 ( \277 , \275 , \276 );
nand \mul_6_11_g13693/U$1 ( \278 , \277 , \171 );
not \g35845/U$2 ( \279 , \165 );
nand \g35845/U$1 ( \280 , \279 , \183 );
nand \mul_6_11_g13692/U$1 ( \281 , \278 , \280 );
xor \mul_6_11_g13592/U$1_r1 ( \282 , \274 , \281 );
xnor \mul_6_11_g13555/U$1_r1 ( \283 , \255 , \282 );
nand \mul_6_11_g13531/U$1 ( \284 , \226 , \283 );
not \mul_6_11_g13520/U$3 ( \285 , \284 );
not \mul_6_11_g13617/U$3 ( \286 , \219 );
not \mul_6_11_g13617/U$4 ( \287 , \185 );
and \mul_6_11_g13617/U$2 ( \288 , \286 , \287 );
and \mul_6_11_g13617/U$5 ( \289 , \219 , \185 );
nor \mul_6_11_g13617/U$1 ( \290 , \288 , \289 );
and \mul_6_11_g13580/U$2 ( \291 , \290 , \158 );
not \mul_6_11_g13580/U$4 ( \292 , \290 );
and \mul_6_11_g13580/U$3 ( \293 , \292 , \223 );
nor \mul_6_11_g13580/U$1 ( \294 , \291 , \293 );
not \mul_6_11_g13559/U$1 ( \295 , \294 );
not \mul_6_11_g13967/U$1 ( \296 , \132 );
not \mul_6_11_g13780/U$3 ( \297 , \296 );
xor \mul_6_11_g13890/U$1 ( \298 , \a[6] , \b[1] );
not \mul_6_11_g13780/U$4 ( \299 , \298 );
or \mul_6_11_g13780/U$2 ( \300 , \297 , \299 );
nand \mul_6_11_g13814/U$1 ( \301 , \129 , \b[0] );
nand \mul_6_11_g13780/U$1 ( \302 , \300 , \301 );
xor \mul_6_11_g13946/U$1 ( \303 , \a[0] , \b[7] );
nand \mul_6_11_g13817/U$1 ( \304 , \303 , \175 );
or \mul_6_11_g13727/U$2 ( \305 , \304 , \177 );
nand \mul_6_11_g13816/U$1 ( \306 , \189 , \177 );
nand \mul_6_11_g13727/U$1 ( \307 , \305 , \306 );
xor \mul_6_11_g13644/U$4 ( \308 , \302 , \307 );
xor \mul_6_11_g13933/U$1 ( \309 , \a[2] , \b[5] );
not \mul_6_11_g13740/U$3 ( \310 , \309 );
not \mul_6_11_g13740/U$4 ( \311 , \267 );
or \mul_6_11_g13740/U$2 ( \312 , \310 , \311 );
nand \mul_6_11_g13813/U$1 ( \313 , \121 , \195 );
nand \mul_6_11_g13740/U$1 ( \314 , \312 , \313 );
and \mul_6_11_g13644/U$3 ( \315 , \308 , \314 );
and \mul_6_11_g13644/U$5 ( \316 , \302 , \307 );
or \mul_6_11_g13644/U$2 ( \317 , \315 , \316 );
xor \mul_6_11_g13641/U$1 ( \318 , \194 , \202 );
xor \mul_6_11_g13641/U$1_r1 ( \319 , \318 , \216 );
xor \g35770/U$4 ( \320 , \317 , \319 );
xor \g35695/U$1 ( \321 , \127 , \138 );
xnor \g35695/U$1_r1 ( \322 , \321 , \153 );
buf \fopt35790/U$1 ( \323 , \322 );
and \g35770/U$3 ( \324 , \320 , \323 );
and \g35770/U$5 ( \325 , \317 , \319 );
or \g35770/U$2 ( \326 , \324 , \325 );
not \fopt35587/U$1 ( \327 , \326 );
nand \mul_6_11_g13551/U$1 ( \328 , \295 , \327 );
xor \mul_6_11_g35955/U$1 ( \329 , \a[5] , \b[1] );
not \mul_6_11_g13789/U$3 ( \330 , \329 );
not \mul_6_11_g13789/U$4 ( \331 , \133 );
or \mul_6_11_g13789/U$2 ( \332 , \330 , \331 );
nand \mul_6_11_g13803/U$1 ( \333 , \298 , \b[0] );
nand \mul_6_11_g13789/U$1 ( \334 , \332 , \333 );
not \mul_6_11_g13788/U$1 ( \335 , \334 );
not \mul_6_11_g13648/U$3 ( \336 , \335 );
or \mul_6_11_g13877/U$2 ( \337 , \a[0] , \b[4] );
nand \mul_6_11_g13877/U$1 ( \338 , \337 , \b[3] );
nand \mul_6_11_g13954/U$1 ( \339 , \a[0] , \b[4] );
nand \mul_6_11_g13860/U$1 ( \340 , \338 , \339 , \b[5] );
not \mul_6_11_g14012/U$2 ( \341 , \340 );
xor \mul_6_11_g35979/U$1 ( \342 , \a[2] , \b[3] );
xor \g35977/U$1 ( \343 , \b[3] , \b[2] );
nand \g35611/U$1 ( \344 , \342 , \343 );
or \mul_6_11_g13730/U$2 ( \345 , \344 , \150 );
xor \g35486/U$1 ( \346 , \b[3] , \a[3] );
nand \mul_6_11_g35702/U$1 ( \347 , \346 , \150 );
nand \mul_6_11_g13730/U$1 ( \348 , \345 , \347 );
nand \mul_6_11_g14012/U$1 ( \349 , \341 , \348 );
not \mul_6_11_g13709/U$1 ( \350 , \349 );
not \mul_6_11_g13648/U$4 ( \351 , \350 );
or \mul_6_11_g13648/U$2 ( \352 , \336 , \351 );
or \mul_6_11_g13648/U$5 ( \353 , \350 , \335 );
nand \mul_6_11_g13648/U$1 ( \354 , \352 , \353 );
not \mul_6_11_g13645/U$1 ( \355 , \354 );
not \mul_6_11_g13619/U$3 ( \356 , \355 );
nand \mul_6_11_g35754/U$1 ( \357 , \177 , \a[0] );
not \mul_6_11_g13847/U$1 ( \358 , \357 );
xor \mul_6_11_g13941/U$1 ( \359 , \a[1] , \b[5] );
nand \mul_6_11_g13825/U$1 ( \360 , \359 , \117 );
or \mul_6_11_g13729/U$2 ( \361 , \360 , \119 );
nand \mul_6_11_g13822/U$1 ( \362 , \309 , \119 );
nand \mul_6_11_g13729/U$1 ( \363 , \361 , \362 );
xor \mul_6_11_g13672/U$1 ( \364 , \358 , \363 );
not \mul_6_11_g13757/U$3 ( \365 , \346 );
not \mul_6_11_g13757/U$4 ( \366 , \147 );
or \mul_6_11_g13757/U$2 ( \367 , \365 , \366 );
not \mul_6_11_g13824/U$2 ( \368 , \212 );
nand \mul_6_11_g13824/U$1 ( \369 , \368 , \150 );
nand \mul_6_11_g13757/U$1 ( \370 , \367 , \369 );
xnor \mul_6_11_g13672/U$1_r1 ( \371 , \364 , \370 );
not \mul_6_11_g13660/U$1 ( \372 , \371 );
not \mul_6_11_g13619/U$4 ( \373 , \372 );
or \mul_6_11_g13619/U$2 ( \374 , \356 , \373 );
nand \mul_6_11_g13622/U$1 ( \375 , \354 , \371 );
nand \mul_6_11_g13619/U$1 ( \376 , \374 , \375 );
not \mul_6_11_g13603/U$1 ( \377 , \376 );
not \mul_6_11_g13697/U$3 ( \378 , \348 );
not \mul_6_11_g13697/U$4 ( \379 , \340 );
and \mul_6_11_g13697/U$2 ( \380 , \378 , \379 );
and \mul_6_11_g13697/U$5 ( \381 , \348 , \340 );
nor \mul_6_11_g13697/U$1 ( \382 , \380 , \381 );
not \mul_6_11_g13687/U$1 ( \383 , \382 );
xor \g35483/U$1 ( \384 , \b[1] , \a[4] );
not \mul_6_11_g13785/U$3 ( \385 , \384 );
not \mul_6_11_g13785/U$4 ( \386 , \133 );
or \mul_6_11_g13785/U$2 ( \387 , \385 , \386 );
nand \mul_6_11_g13829/U$1 ( \388 , \329 , \b[0] );
nand \mul_6_11_g13785/U$1 ( \389 , \387 , \388 );
or \mul_6_11_g13647/U$2 ( \390 , \383 , \389 );
xor \mul_6_11_g13948/U$1 ( \391 , \a[0] , \b[5] );
not \mul_6_11_g13743/U$3 ( \392 , \391 );
not \mul_6_11_g13743/U$4 ( \393 , \198 );
or \mul_6_11_g13743/U$2 ( \394 , \392 , \393 );
nand \mul_6_11_g13795/U$1 ( \395 , \121 , \359 );
nand \mul_6_11_g13743/U$1 ( \396 , \394 , \395 );
nand \mul_6_11_g13647/U$1 ( \397 , \390 , \396 );
not \mul_6_11_g13784/U$1 ( \398 , \389 );
not \mul_6_11_g13666/U$2 ( \399 , \398 );
nand \mul_6_11_g13666/U$1 ( \400 , \399 , \383 );
nand \mul_6_11_g13635/U$1 ( \401 , \397 , \400 );
not \fopt35591/U$1 ( \402 , \401 );
nand \mul_6_11_g13584/U$1 ( \403 , \377 , \402 );
not \mul_6_11_g13583/U$1 ( \404 , \403 );
xor \mul_6_11_g13691/U$1 ( \405 , \207 , \215 );
xor \mul_6_11_g13644/U$1 ( \406 , \302 , \307 );
xor \mul_6_11_g13644/U$1_r1 ( \407 , \406 , \314 );
xor \mul_6_11_g13598/U$1 ( \408 , \405 , \407 );
not \mul_6_11_g13707/U$2 ( \409 , \363 );
nand \mul_6_11_g13707/U$1 ( \410 , \409 , \357 );
not \mul_6_11_g13682/U$3 ( \411 , \410 );
not \mul_6_11_g13682/U$4 ( \412 , \370 );
or \mul_6_11_g13682/U$2 ( \413 , \411 , \412 );
nand \mul_6_11_g13705/U$1 ( \414 , \363 , \358 );
nand \mul_6_11_g13682/U$1 ( \415 , \413 , \414 );
xor \mul_6_11_g13598/U$1_r1 ( \416 , \408 , \415 );
nand \mul_6_11_g13668/U$1 ( \417 , \349 , \335 );
not \mul_6_11_g13616/U$3 ( \418 , \417 );
not \mul_6_11_g13616/U$4 ( \419 , \372 );
or \mul_6_11_g13616/U$2 ( \420 , \418 , \419 );
nand \mul_6_11_g13667/U$1 ( \421 , \350 , \334 );
nand \mul_6_11_g13616/U$1 ( \422 , \420 , \421 );
nand \mul_6_11_g13575/U$1 ( \423 , \416 , \422 );
and \mul_6_11_g13558/U$2 ( \424 , \404 , \423 );
nor \mul_6_11_g13577/U$1 ( \425 , \416 , \422 );
nor \mul_6_11_g13558/U$1 ( \426 , \424 , \425 );
not \mul_6_11_g13792/U$3 ( \427 , \163 );
xor \g35978/U$1 ( \428 , \b[1] , \a[3] );
not \mul_6_11_g13792/U$4 ( \429 , \428 );
or \mul_6_11_g13792/U$2 ( \430 , \427 , \429 );
nand \mul_6_11_g13828/U$1 ( \431 , \384 , \b[0] );
nand \mul_6_11_g13792/U$1 ( \432 , \430 , \431 );
not \mul_6_11_g13719/U$2 ( \433 , \432 );
nand \mul_6_11_g13978/U$1 ( \434 , \121 , \a[0] );
nand \mul_6_11_g13719/U$1 ( \435 , \433 , \434 );
not \mul_6_11_g13669/U$3 ( \436 , \435 );
xor \mul_6_11_g13936/U$1 ( \437 , \a[1] , \b[3] );
not \mul_6_11_g13758/U$3 ( \438 , \437 );
not \mul_6_11_g13758/U$4 ( \439 , \242 );
or \mul_6_11_g13758/U$2 ( \440 , \438 , \439 );
nand \mul_6_11_g13804/U$1 ( \441 , \150 , \342 );
nand \mul_6_11_g13758/U$1 ( \442 , \440 , \441 );
not \mul_6_11_g13669/U$4 ( \443 , \442 );
or \mul_6_11_g13669/U$2 ( \444 , \436 , \443 );
not \mul_6_11_g14010/U$2 ( \445 , \434 );
nand \mul_6_11_g14010/U$1 ( \446 , \445 , \432 );
nand \mul_6_11_g13669/U$1 ( \447 , \444 , \446 );
not \g35609/U$2 ( \448 , \447 );
not \mul_6_11_g13698/U$3 ( \449 , \398 );
not \mul_6_11_g13698/U$4 ( \450 , \396 );
or \mul_6_11_g13698/U$2 ( \451 , \449 , \450 );
or \mul_6_11_g13698/U$5 ( \452 , \396 , \398 );
nand \mul_6_11_g13698/U$1 ( \453 , \451 , \452 );
and \mul_6_11_g13650/U$2 ( \454 , \453 , \382 );
not \mul_6_11_g13650/U$4 ( \455 , \453 );
and \mul_6_11_g13650/U$3 ( \456 , \455 , \383 );
nor \mul_6_11_g13650/U$1 ( \457 , \454 , \456 );
nand \g35609/U$1 ( \458 , \448 , \457 );
not \g35608/U$3 ( \459 , \458 );
nand \mul_6_11_g13958/U$1 ( \460 , \a[0] , \b[2] );
and \mul_6_11_g13983/U$1 ( \461 , \460 , \b[3] );
or \mul_6_11_g13878/U$2 ( \462 , \a[0] , \b[2] );
nand \mul_6_11_g13878/U$1 ( \463 , \462 , \b[1] );
nand \mul_6_11_g13858/U$1 ( \464 , \461 , \463 );
not \mul_6_11_g14011/U$2 ( \465 , \464 );
xor \mul_6_11_g13928/U$1 ( \466 , \a[2] , \b[1] );
not \mul_6_11_g13778/U$3 ( \467 , \466 );
not \mul_6_11_g13778/U$4 ( \468 , \163 );
or \mul_6_11_g13778/U$2 ( \469 , \467 , \468 );
nand \mul_6_11_g13794/U$1 ( \470 , \428 , \b[0] );
nand \mul_6_11_g13778/U$1 ( \471 , \469 , \470 );
nand \mul_6_11_g14011/U$1 ( \472 , \465 , \471 );
not \mul_6_11_g13610/U$3 ( \473 , \472 );
not \mul_6_11_g13712/U$3 ( \474 , \432 );
not \mul_6_11_g13712/U$4 ( \475 , \434 );
and \mul_6_11_g13712/U$2 ( \476 , \474 , \475 );
and \mul_6_11_g13712/U$5 ( \477 , \432 , \434 );
nor \mul_6_11_g13712/U$1 ( \478 , \476 , \477 );
not \mul_6_11_g13673/U$3 ( \479 , \478 );
not \mul_6_11_g13673/U$4 ( \480 , \442 );
and \mul_6_11_g13673/U$2 ( \481 , \479 , \480 );
and \mul_6_11_g13673/U$5 ( \482 , \442 , \478 );
nor \mul_6_11_g13673/U$1 ( \483 , \481 , \482 );
not \mul_6_11_g13610/U$4 ( \484 , \483 );
or \mul_6_11_g13610/U$2 ( \485 , \473 , \484 );
xor \g35487/U$1 ( \486 , \b[3] , \a[0] );
not \mul_6_11_g13753/U$3 ( \487 , \486 );
not \mul_6_11_g13753/U$4 ( \488 , \242 );
or \mul_6_11_g13753/U$2 ( \489 , \487 , \488 );
nand \mul_6_11_g13796/U$1 ( \490 , \150 , \437 );
nand \mul_6_11_g13753/U$1 ( \491 , \489 , \490 );
not \mul_6_11_g14006/U$2 ( \492 , \491 );
not \mul_6_11_g13713/U$3 ( \493 , \471 );
not \mul_6_11_g13713/U$4 ( \494 , \464 );
and \mul_6_11_g13713/U$2 ( \495 , \493 , \494 );
and \mul_6_11_g13713/U$5 ( \496 , \471 , \464 );
nor \mul_6_11_g13713/U$1 ( \497 , \495 , \496 );
nand \mul_6_11_g14006/U$1 ( \498 , \492 , \497 );
xor \mul_6_11_g13935/U$1 ( \499 , \a[1] , \b[1] );
not \mul_6_11_g13779/U$3 ( \500 , \499 );
not \mul_6_11_g13779/U$4 ( \501 , \133 );
or \mul_6_11_g13779/U$2 ( \502 , \500 , \501 );
nand \mul_6_11_g13798/U$1 ( \503 , \466 , \b[0] );
nand \mul_6_11_g13779/U$1 ( \504 , \502 , \503 );
and \mul_6_11_g13980/U$1 ( \505 , \144 , \a[0] );
nor \mul_6_11_g13721/U$1 ( \506 , \504 , \505 );
nand \mul_6_11_g13959/U$1 ( \507 , \a[0] , \b[0] );
nand \mul_6_11_g13882/U$1 ( \508 , \507 , \b[1] );
nor \mul_6_11_g13841/U$1 ( \509 , \508 , \a[0] );
not \mul_6_11_g13809/U$2 ( \510 , \499 );
nand \mul_6_11_g13809/U$1 ( \511 , \510 , \b[0] );
nand \mul_6_11_g13766/U$1 ( \512 , \509 , \511 );
or \mul_6_11_g13694/U$2 ( \513 , \506 , \512 );
nand \mul_6_11_g35965/U$1 ( \514 , \504 , \505 );
nand \mul_6_11_g13694/U$1 ( \515 , \513 , \514 );
nand \mul_6_11_g13646/U$1 ( \516 , \498 , \515 );
not \mul_6_11_g14005/U$2 ( \517 , \497 );
nand \mul_6_11_g14005/U$1 ( \518 , \517 , \491 );
nand \mul_6_11_g13634/U$1 ( \519 , \516 , \518 );
nand \mul_6_11_g13610/U$1 ( \520 , \485 , \519 );
not \fopt35791/U$1 ( \521 , \483 );
not \mul_6_11_g13703/U$1 ( \522 , \472 );
nand \mul_6_11_g13633/U$1 ( \523 , \521 , \522 );
nand \mul_6_11_g13600/U$1 ( \524 , \520 , \523 );
not \g35608/U$4 ( \525 , \524 );
or \g35608/U$2 ( \526 , \459 , \525 );
not \mul_6_11_g13997/U$2 ( \527 , \457 );
nand \mul_6_11_g13997/U$1 ( \528 , \527 , \447 );
nand \g35608/U$1 ( \529 , \526 , \528 );
not \mul_6_11_g13546/U$2 ( \530 , \529 );
nand \mul_6_11_g13587/U$1 ( \531 , \376 , \401 );
nand \mul_6_11_g13546/U$1 ( \532 , \530 , \423 , \531 );
xor \mul_6_11_g13590/U$1 ( \533 , \317 , \322 );
xnor \mul_6_11_g13590/U$1_r1 ( \534 , \533 , \319 );
xor \mul_6_11_g13598/U$4 ( \535 , \405 , \407 );
and \mul_6_11_g13598/U$3 ( \536 , \535 , \415 );
and \mul_6_11_g13598/U$5 ( \537 , \405 , \407 );
or \mul_6_11_g13598/U$2 ( \538 , \536 , \537 );
not \mul_6_11_g35630/U$1 ( \539 , \538 );
nand \mul_6_11_g35716/U$1 ( \540 , \534 , \539 );
and \mul_6_11_g13526/U$1 ( \541 , \328 , \426 , \532 , \540 );
not \mul_6_11_g13520/U$4 ( \542 , \541 );
or \mul_6_11_g13520/U$2 ( \543 , \285 , \542 );
not \mul_6_11_g13561/U$1 ( \544 , \225 );
nand \mul_6_11_g13532/U$1 ( \545 , \283 , \544 );
not \g35626/U$3 ( \546 , \326 );
not \g35626/U$4 ( \547 , \294 );
or \g35626/U$2 ( \548 , \546 , \547 );
not \g35627/U$2 ( \549 , \534 );
nand \g35627/U$1 ( \550 , \549 , \538 );
nand \g35626/U$1 ( \551 , \548 , \550 );
or \mul_6_11_g13990/U$1 ( \552 , \294 , \326 );
and \mul_6_11_g13522/U$2 ( \553 , \545 , \551 , \552 );
nor \mul_6_11_g13534/U$1 ( \554 , \283 , \544 );
nor \mul_6_11_g13522/U$1 ( \555 , \553 , \554 );
nand \mul_6_11_g13520/U$1 ( \556 , \543 , \555 );
not \mul_6_11_g13737/U$3 ( \557 , \231 );
not \mul_6_11_g13737/U$4 ( \558 , \106 );
or \mul_6_11_g13737/U$2 ( \559 , \557 , \558 );
xor \mul_6_11_g13944/U$1 ( \560 , \a[3] , \b[9] );
nand \mul_6_11_g13835/U$1 ( \561 , \104 , \560 );
nand \mul_6_11_g13737/U$1 ( \562 , \559 , \561 );
not \mul_6_11_g13736/U$1 ( \563 , \562 );
not \mul_6_11_g13759/U$3 ( \564 , \245 );
not \mul_6_11_g13759/U$4 ( \565 , \242 );
or \mul_6_11_g13759/U$2 ( \566 , \564 , \565 );
not \mul_6_11_g13953/U$2 ( \567 , \b[3] );
nand \mul_6_11_g13953/U$1 ( \568 , \567 , \a[9] );
not \mul_6_11_g13855/U$3 ( \569 , \568 );
not \mul_6_11_g13952/U$2 ( \570 , \a[9] );
nand \mul_6_11_g13952/U$1 ( \571 , \570 , \b[3] );
not \mul_6_11_g13855/U$4 ( \572 , \571 );
or \mul_6_11_g13855/U$2 ( \573 , \569 , \572 );
nand \mul_6_11_g13855/U$1 ( \574 , \573 , \150 );
nand \mul_6_11_g13759/U$1 ( \575 , \566 , \574 );
xor \g35949/U$1 ( \576 , \563 , \575 );
xor \mul_6_11_g13939/U$1 ( \577 , \b[11] , \b[10] );
xor \mul_6_11_g13915/U$1 ( \578 , \a[0] , \b[11] );
nand \mul_6_11_g13834/U$1 ( \579 , \577 , \578 );
or \mul_6_11_g13724/U$2 ( \580 , \579 , \257 );
xor \mul_6_11_g13932/U$1 ( \581 , \a[1] , \b[11] );
nand \mul_6_11_g13797/U$1 ( \582 , \257 , \581 );
nand \mul_6_11_g13724/U$1 ( \583 , \580 , \582 );
or \mul_6_11_g13874/U$2 ( \584 , \a[0] , \b[10] );
nand \mul_6_11_g13874/U$1 ( \585 , \584 , \b[9] );
nand \mul_6_11_g13957/U$1 ( \586 , \a[0] , \b[10] );
nand \mul_6_11_g13866/U$1 ( \587 , \585 , \586 , \b[11] );
not \mul_6_11_g13865/U$1 ( \588 , \587 );
and \mul_6_11_g13696/U$2 ( \589 , \583 , \588 );
not \mul_6_11_g13696/U$4 ( \590 , \583 );
and \mul_6_11_g13696/U$3 ( \591 , \590 , \587 );
nor \mul_6_11_g13696/U$1 ( \592 , \589 , \591 );
not \mul_6_11_g13772/U$3 ( \593 , \262 );
not \mul_6_11_g13772/U$4 ( \594 , \133 );
or \mul_6_11_g13772/U$2 ( \595 , \593 , \594 );
xor \mul_6_11_g13886/U$1 ( \596 , \a[11] , \b[1] );
nand \mul_6_11_g13844/U$1 ( \597 , \596 , \b[0] );
nand \mul_6_11_g13772/U$1 ( \598 , \595 , \597 );
xnor \mul_6_11_g14008/U$1 ( \599 , \592 , \598 );
xnor \g35949/U$1_r1 ( \600 , \576 , \599 );
not \mul_6_11_g13750/U$3 ( \601 , \237 );
not \mul_6_11_g13750/U$4 ( \602 , \178 );
or \mul_6_11_g13750/U$2 ( \603 , \601 , \602 );
xor \mul_6_11_g13925/U$1 ( \604 , \a[5] , \b[7] );
nand \mul_6_11_g13800/U$1 ( \605 , \177 , \604 );
nand \mul_6_11_g13750/U$1 ( \606 , \603 , \605 );
not \mul_6_11_g13741/U$3 ( \607 , \270 );
not \mul_6_11_g13741/U$4 ( \608 , \198 );
or \mul_6_11_g13741/U$2 ( \609 , \607 , \608 );
xor \mul_6_11_g13911/U$1 ( \610 , \a[7] , \b[5] );
nand \mul_6_11_g13830/U$1 ( \611 , \121 , \610 );
nand \mul_6_11_g13741/U$1 ( \612 , \609 , \611 );
not \g36021/U$2 ( \613 , \612 );
xor \g36021/U$1 ( \614 , \606 , \613 );
and \g35948/U$2 ( \615 , \600 , \614 );
not \g35948/U$4 ( \616 , \600 );
not \mul_6_11_g13699/U$1 ( \617 , \614 );
and \g35948/U$3 ( \618 , \616 , \617 );
nor \g35948/U$1 ( \619 , \615 , \618 );
xor \mul_6_11_g13655/U$4 ( \620 , \233 , \239 );
and \mul_6_11_g13655/U$3 ( \621 , \620 , \247 );
and \mul_6_11_g13655/U$5 ( \622 , \233 , \239 );
or \mul_6_11_g13655/U$2 ( \623 , \621 , \622 );
xor \mul_6_11_g13662/U$4 ( \624 , \258 , \264 );
and \mul_6_11_g13662/U$3 ( \625 , \624 , \272 );
and \mul_6_11_g13662/U$5 ( \626 , \258 , \264 );
or \mul_6_11_g13662/U$2 ( \627 , \625 , \626 );
xor \mul_6_11_g14001/U$1 ( \628 , \623 , \627 );
xor \g35947/U$1 ( \629 , \619 , \628 );
xor \mul_6_11_g13592/U$4 ( \630 , \256 , \273 );
and \mul_6_11_g13592/U$3 ( \631 , \630 , \281 );
and \mul_6_11_g13592/U$5 ( \632 , \256 , \273 );
or \mul_6_11_g13592/U$2 ( \633 , \631 , \632 );
xor \g35946/U$1 ( \634 , \629 , \633 );
buf \fopt35792/U$1 ( \635 , \248 );
or \mul_6_11_g14000/U$1 ( \636 , \254 , \635 );
not \mul_6_11_g13554/U$3 ( \637 , \636 );
not \mul_6_11_g13554/U$4 ( \638 , \282 );
or \mul_6_11_g13554/U$2 ( \639 , \637 , \638 );
nand \mul_6_11_g13588/U$1 ( \640 , \254 , \635 );
nand \mul_6_11_g13554/U$1 ( \641 , \639 , \640 );
xor \g35946/U$1_r1 ( \642 , \634 , \641 );
xor \mul_6_11_g35498/U$1 ( \643 , \556 , \642 );
buf \fopt35678/U$1 ( \644 , \643 );
not \fopt35676/U$1 ( \645 , \644 );
nor \g35732/U$1 ( \646 , \101 , \645 );
not \g5053/U$2 ( \647 , \b[7] );
not \g5113/U$1 ( \648 , \a[7] );
nand \g5053/U$1 ( \649 , \647 , \648 );
not \g4855/U$3 ( \650 , \649 );
not \mul_6_11_g13525/U$3 ( \651 , \540 );
or \g35844/U$1 ( \652 , \416 , \422 );
not \mul_6_11_g13544/U$3 ( \653 , \652 );
nand \mul_6_11_g13567/U$1 ( \654 , \423 , \531 );
not \mul_6_11_g13544/U$4 ( \655 , \654 );
or \mul_6_11_g13544/U$2 ( \656 , \653 , \655 );
nand \mul_6_11_g13553/U$1 ( \657 , \652 , \529 , \403 );
nand \mul_6_11_g13544/U$1 ( \658 , \656 , \657 );
not \mul_6_11_g13525/U$4 ( \659 , \658 );
or \mul_6_11_g13525/U$2 ( \660 , \651 , \659 );
nor \mul_6_11_g35629/U$1 ( \661 , \539 , \534 );
not \mul_6_11_g35628/U$1 ( \662 , \661 );
nand \mul_6_11_g13525/U$1 ( \663 , \660 , \662 );
and \mul_6_11_g2/U$1 ( \664 , \294 , \326 );
not \mul_6_11_g13542/U$2 ( \665 , \664 );
nand \mul_6_11_g13542/U$1 ( \666 , \665 , \552 );
not \mul_6_11_g13541/U$1 ( \667 , \666 );
and \mul_6_11_g13519/U$2 ( \668 , \663 , \667 );
not \mul_6_11_g13519/U$4 ( \669 , \663 );
and \mul_6_11_g13519/U$3 ( \670 , \669 , \666 );
nor \mul_6_11_g13519/U$1 ( \671 , \668 , \670 );
buf \g5124/U$1 ( \672 , \671 );
not \g4855/U$4 ( \673 , \672 );
or \g4855/U$2 ( \674 , \650 , \673 );
xor \mul_17_13_g35959/U$1 ( \675 , \b[6] , \c[1] );
not \mul_17_13_g20405/U$3 ( \676 , \675 );
not \mul_17_13_g20703/U$2 ( \677 , \c[0] );
nand \mul_17_13_g20703/U$1 ( \678 , \677 , \c[1] );
not \mul_17_13_g20691/U$1 ( \679 , \678 );
not \mul_17_13_g20405/U$4 ( \680 , \679 );
or \mul_17_13_g20405/U$2 ( \681 , \676 , \680 );
xor \mul_17_13_g20613/U$1 ( \682 , \b[7] , \c[1] );
nand \mul_17_13_g20461/U$1 ( \683 , \682 , \c[0] );
nand \mul_17_13_g20405/U$1 ( \684 , \681 , \683 );
not \mul_17_13_g20298/U$3 ( \685 , \684 );
or \mul_17_13_g20548/U$2 ( \686 , \b[0] , \c[6] );
nand \mul_17_13_g20548/U$1 ( \687 , \686 , \c[5] );
nand \mul_17_13_g20671/U$1 ( \688 , \b[0] , \c[6] );
nand \mul_17_13_g20527/U$1 ( \689 , \687 , \688 , \c[7] );
not \mul_17_13_g20298/U$4 ( \690 , \689 );
and \mul_17_13_g20298/U$2 ( \691 , \685 , \690 );
and \mul_17_13_g20298/U$5 ( \692 , \684 , \689 );
nor \mul_17_13_g20298/U$1 ( \693 , \691 , \692 );
xor \mul_17_13_g20636/U$1 ( \694 , \b[3] , \c[3] );
not \mul_17_13_g20388/U$3 ( \695 , \694 );
xor \mul_17_13_g20568/U$1 ( \696 , \c[3] , \c[2] );
not \mul_17_13_g20486/U$2 ( \697 , \696 );
xor \mul_17_13_g35707/U$1 ( \698 , \c[2] , \c[1] );
nor \mul_17_13_g20486/U$1 ( \699 , \697 , \698 );
not \mul_17_13_g20388/U$4 ( \700 , \699 );
or \mul_17_13_g20388/U$2 ( \701 , \695 , \700 );
buf \mul_17_13_g20559/U$1 ( \702 , \698 );
xor \mul_17_13_g20625/U$1 ( \703 , \b[4] , \c[3] );
nand \mul_17_13_g20459/U$1 ( \704 , \702 , \703 );
nand \mul_17_13_g20388/U$1 ( \705 , \701 , \704 );
not \mul_17_13_g20237/U$3 ( \706 , \705 );
xor \mul_17_13_g35957/U$1 ( \707 , \b[5] , \c[1] );
not \mul_17_13_g20413/U$3 ( \708 , \707 );
not \mul_17_13_g20413/U$4 ( \709 , \679 );
or \mul_17_13_g20413/U$2 ( \710 , \708 , \709 );
nand \mul_17_13_g20462/U$1 ( \711 , \675 , \c[0] );
nand \mul_17_13_g20413/U$1 ( \712 , \710 , \711 );
xor \mul_17_13_g35490/U$1 ( \713 , \c[6] , \c[5] );
buf \mul_17_13_g20582/U$1 ( \714 , \713 );
nand \mul_17_13_g20705/U$1 ( \715 , \714 , \b[0] );
not \mul_17_13_g20512/U$1 ( \716 , \715 );
or \mul_17_13_g20707/U$1 ( \717 , \712 , \716 );
not \mul_17_13_g20237/U$4 ( \718 , \717 );
or \mul_17_13_g20237/U$2 ( \719 , \706 , \718 );
nand \mul_17_13_g20305/U$1 ( \720 , \712 , \716 );
nand \mul_17_13_g20237/U$1 ( \721 , \719 , \720 );
xor \mul_17_13_g20159/U$1 ( \722 , \693 , \721 );
xor \mul_17_13_g20659/U$1 ( \723 , \b[0] , \c[7] );
not \mul_17_13_g20347/U$3 ( \724 , \723 );
xnor \mul_17_13_g20718/U$1 ( \725 , \c[7] , \c[6] );
nor \mul_17_13_g20444/U$1 ( \726 , \725 , \713 );
not \mul_17_13_g20347/U$4 ( \727 , \726 );
or \mul_17_13_g20347/U$2 ( \728 , \724 , \727 );
xor \mul_17_13_g20653/U$1 ( \729 , \b[1] , \c[7] );
nand \mul_17_13_g20490/U$1 ( \730 , \714 , \729 );
nand \mul_17_13_g20347/U$1 ( \731 , \728 , \730 );
xor \mul_17_13_g20640/U$1 ( \732 , \b[2] , \c[5] );
not \mul_17_13_g20372/U$3 ( \733 , \732 );
xor \mul_17_13_g35650/U$1 ( \734 , \c[4] , \c[3] );
xnor \mul_17_13_g20717/U$1 ( \735 , \c[5] , \c[4] );
nor \mul_17_13_g20704/U$1 ( \736 , \734 , \735 );
not \mul_17_13_g20372/U$4 ( \737 , \736 );
or \mul_17_13_g20372/U$2 ( \738 , \733 , \737 );
xor \g35708/U$1 ( \739 , \c[4] , \c[3] );
xor \mul_17_13_g20639/U$1 ( \740 , \b[3] , \c[5] );
nand \mul_17_13_g20478/U$1 ( \741 , \739 , \740 );
nand \mul_17_13_g20372/U$1 ( \742 , \738 , \741 );
xor \mul_17_13_g20205/U$1 ( \743 , \731 , \742 );
not \mul_17_13_g20391/U$3 ( \744 , \703 );
not \mul_17_13_g20756/U$2 ( \745 , \696 );
nor \mul_17_13_g20756/U$1 ( \746 , \745 , \698 );
not \mul_17_13_g20391/U$4 ( \747 , \746 );
or \mul_17_13_g20391/U$2 ( \748 , \744 , \747 );
xor \mul_17_13_g20624/U$1 ( \749 , \b[5] , \c[3] );
nand \mul_17_13_g20496/U$1 ( \750 , \702 , \749 );
nand \mul_17_13_g20391/U$1 ( \751 , \748 , \750 );
xor \mul_17_13_g20205/U$1_r1 ( \752 , \743 , \751 );
xnor \mul_17_13_g20159/U$1_r1 ( \753 , \722 , \752 );
xor \mul_17_13_g20623/U$1 ( \754 , \b[4] , \c[1] );
not \mul_17_13_g20408/U$3 ( \755 , \754 );
not \mul_17_13_g20408/U$4 ( \756 , \679 );
or \mul_17_13_g20408/U$2 ( \757 , \755 , \756 );
nand \mul_17_13_g20452/U$1 ( \758 , \707 , \c[0] );
nand \mul_17_13_g20408/U$1 ( \759 , \757 , \758 );
not \mul_17_13_g20752/U$2 ( \760 , \759 );
or \mul_17_13_g20549/U$2 ( \761 , \b[0] , \c[4] );
nand \mul_17_13_g20549/U$1 ( \762 , \761 , \c[3] );
nand \mul_17_13_g20667/U$1 ( \763 , \b[0] , \c[4] );
nand \mul_17_13_g20524/U$1 ( \764 , \762 , \763 , \c[5] );
nor \mul_17_13_g20752/U$1 ( \765 , \760 , \764 );
not \mul_17_13_g20741/U$2 ( \766 , \765 );
xor \mul_17_13_g20648/U$1 ( \767 , \b[1] , \c[5] );
not \mul_17_13_g20371/U$3 ( \768 , \767 );
not \mul_17_13_g20371/U$4 ( \769 , \736 );
or \mul_17_13_g20371/U$2 ( \770 , \768 , \769 );
nand \mul_17_13_g20475/U$1 ( \771 , \734 , \732 );
nand \mul_17_13_g20371/U$1 ( \772 , \770 , \771 );
not \mul_17_13_g20370/U$1 ( \773 , \772 );
nand \mul_17_13_g20741/U$1 ( \774 , \766 , \773 );
not \mul_17_13_g20185/U$3 ( \775 , \774 );
xor \g35922/U$1 ( \776 , \715 , \712 );
xnor \g35922/U$1_r1 ( \777 , \776 , \705 );
not \mul_17_13_g20185/U$4 ( \778 , \777 );
or \mul_17_13_g20185/U$2 ( \779 , \775 , \778 );
nand \mul_17_13_g20246/U$1 ( \780 , \772 , \765 );
nand \mul_17_13_g20185/U$1 ( \781 , \779 , \780 );
or \mul_17_13_g20732/U$1 ( \782 , \753 , \781 );
nand \mul_17_13_g20112/U$1 ( \783 , \753 , \781 );
nand \mul_17_13_g20729/U$1 ( \784 , \782 , \783 );
xor \mul_17_13_g20661/U$1 ( \785 , \b[0] , \c[5] );
not \mul_17_13_g20375/U$3 ( \786 , \785 );
not \mul_17_13_g20375/U$4 ( \787 , \736 );
or \mul_17_13_g20375/U$2 ( \788 , \786 , \787 );
nand \mul_17_13_g20434/U$1 ( \789 , \739 , \767 );
nand \mul_17_13_g20375/U$1 ( \790 , \788 , \789 );
not \mul_17_13_g20299/U$3 ( \791 , \759 );
not \mul_17_13_g20299/U$4 ( \792 , \764 );
and \mul_17_13_g20299/U$2 ( \793 , \791 , \792 );
and \mul_17_13_g20299/U$5 ( \794 , \759 , \764 );
nor \mul_17_13_g20299/U$1 ( \795 , \793 , \794 );
xor \mul_17_13_g20192/U$1 ( \796 , \790 , \795 );
xor \mul_17_13_g20637/U$1 ( \797 , \b[2] , \c[3] );
not \mul_17_13_g20392/U$3 ( \798 , \797 );
not \mul_17_13_g20392/U$4 ( \799 , \746 );
or \mul_17_13_g20392/U$2 ( \800 , \798 , \799 );
nand \mul_17_13_g20438/U$1 ( \801 , \702 , \694 );
nand \mul_17_13_g20392/U$1 ( \802 , \800 , \801 );
xor \mul_17_13_g20192/U$1_r1 ( \803 , \796 , \802 );
nand \mul_17_13_g20516/U$1 ( \804 , \739 , \b[0] );
and \g35471/U$2 ( \805 , \702 , \797 );
not \g35471/U$4 ( \806 , \702 );
xor \mul_17_13_g20644/U$1 ( \807 , \b[1] , \c[3] );
and \g35472/U$1 ( \808 , \696 , \807 );
and \g35471/U$3 ( \809 , \806 , \808 );
nor \g35471/U$1 ( \810 , \805 , \809 );
xor \mul_17_13_g20220/U$4 ( \811 , \804 , \810 );
xor \mul_17_13_g20634/U$1 ( \812 , \b[3] , \c[1] );
and \mul_17_13_g20416/U$2 ( \813 , \679 , \812 );
and \mul_17_13_g20710/U$1 ( \814 , \754 , \c[0] );
nor \mul_17_13_g20416/U$1 ( \815 , \813 , \814 );
and \mul_17_13_g20220/U$3 ( \816 , \811 , \815 );
and \mul_17_13_g20220/U$5 ( \817 , \804 , \810 );
or \mul_17_13_g20220/U$2 ( \818 , \816 , \817 );
nand \mul_17_13_g20148/U$1 ( \819 , \803 , \818 );
xor \mul_17_13_g20664/U$1 ( \820 , \b[0] , \c[3] );
not \mul_17_13_g20396/U$3 ( \821 , \820 );
not \mul_17_13_g20396/U$4 ( \822 , \746 );
or \mul_17_13_g20396/U$2 ( \823 , \821 , \822 );
nand \mul_17_13_g20491/U$1 ( \824 , \702 , \807 );
nand \mul_17_13_g20396/U$1 ( \825 , \823 , \824 );
not \mul_17_13_g20750/U$2 ( \826 , \825 );
xor \mul_17_13_g20633/U$1 ( \827 , \b[2] , \c[1] );
not \mul_17_13_g20410/U$3 ( \828 , \827 );
not \mul_17_13_g20410/U$4 ( \829 , \679 );
or \mul_17_13_g20410/U$2 ( \830 , \828 , \829 );
nand \mul_17_13_g20454/U$1 ( \831 , \812 , \c[0] );
nand \mul_17_13_g20410/U$1 ( \832 , \830 , \831 );
not \mul_17_13_g20300/U$3 ( \833 , \832 );
nand \mul_17_13_g20669/U$1 ( \834 , \b[0] , \c[2] );
or \mul_17_13_g20550/U$2 ( \835 , \b[0] , \c[2] );
nand \mul_17_13_g20550/U$1 ( \836 , \835 , \c[1] );
nand \g35912/U$1 ( \837 , \834 , \c[3] , \836 );
not \mul_17_13_g20300/U$4 ( \838 , \837 );
and \mul_17_13_g20300/U$2 ( \839 , \833 , \838 );
and \mul_17_13_g20300/U$5 ( \840 , \832 , \837 );
nor \mul_17_13_g20300/U$1 ( \841 , \839 , \840 );
nand \mul_17_13_g20750/U$1 ( \842 , \826 , \841 );
not \g35910/U$3 ( \843 , \842 );
xor \g35476/U$1 ( \844 , \c[1] , \b[1] );
not \mul_17_13_g20420/U$3 ( \845 , \844 );
not \mul_17_13_g20420/U$4 ( \846 , \679 );
or \mul_17_13_g20420/U$2 ( \847 , \845 , \846 );
nand \mul_17_13_g20476/U$1 ( \848 , \827 , \c[0] );
nand \mul_17_13_g20420/U$1 ( \849 , \847 , \848 );
and \mul_17_13_g20713/U$1 ( \850 , \702 , \b[0] );
nor \mul_17_13_g20309/U$1 ( \851 , \849 , \850 );
nand \mul_17_13_g20681/U$1 ( \852 , \b[0] , \c[0] );
nand \mul_17_13_g20543/U$1 ( \853 , \852 , \c[1] );
not \mul_17_13_g20755/U$2 ( \854 , \853 );
xor \mul_17_13_g20665/U$1 ( \855 , \b[0] , \c[1] );
not \mul_17_13_g20407/U$3 ( \856 , \855 );
not \mul_17_13_g20407/U$4 ( \857 , \679 );
or \mul_17_13_g20407/U$2 ( \858 , \856 , \857 );
nand \mul_17_13_g20477/U$1 ( \859 , \844 , \c[0] );
nand \mul_17_13_g20407/U$1 ( \860 , \858 , \859 );
nand \mul_17_13_g20755/U$1 ( \861 , \854 , \860 );
or \mul_17_13_g20235/U$2 ( \862 , \851 , \861 );
nand \mul_17_13_g20308/U$1 ( \863 , \849 , \850 );
nand \mul_17_13_g20235/U$1 ( \864 , \862 , \863 );
not \g35910/U$4 ( \865 , \864 );
or \g35910/U$2 ( \866 , \843 , \865 );
not \mul_17_13_g20742/U$2 ( \867 , \841 );
nand \mul_17_13_g20742/U$1 ( \868 , \867 , \825 );
nand \g35910/U$1 ( \869 , \866 , \868 );
not \mul_17_13_g20132/U$3 ( \870 , \869 );
xor \mul_17_13_g20220/U$1 ( \871 , \804 , \810 );
xor \mul_17_13_g20220/U$1_r1 ( \872 , \871 , \815 );
not \mul_17_13_g20751/U$2 ( \873 , \837 );
nand \mul_17_13_g20751/U$1 ( \874 , \873 , \832 );
nand \mul_17_13_g20198/U$1 ( \875 , \872 , \874 );
not \mul_17_13_g20132/U$4 ( \876 , \875 );
or \mul_17_13_g20132/U$2 ( \877 , \870 , \876 );
or \g35839/U$1 ( \878 , \872 , \874 );
nand \mul_17_13_g20132/U$1 ( \879 , \877 , \878 );
nand \mul_17_13_g20100/U$1 ( \880 , \819 , \879 );
not \mul_17_13_g20239/U$3 ( \881 , \765 );
not \mul_17_13_g20239/U$4 ( \882 , \773 );
and \mul_17_13_g20239/U$2 ( \883 , \881 , \882 );
and \mul_17_13_g20239/U$5 ( \884 , \765 , \773 );
nor \mul_17_13_g20239/U$1 ( \885 , \883 , \884 );
xnor \g35464/U$1 ( \886 , \777 , \885 );
not \mul_17_13_g20740/U$2 ( \887 , \795 );
nand \mul_17_13_g20740/U$1 ( \888 , \887 , \790 );
not \mul_17_13_g20374/U$1 ( \889 , \790 );
not \mul_17_13_g20200/U$3 ( \890 , \889 );
not \mul_17_13_g20200/U$4 ( \891 , \795 );
or \mul_17_13_g20200/U$2 ( \892 , \890 , \891 );
nand \mul_17_13_g20200/U$1 ( \893 , \892 , \802 );
nand \mul_17_13_g35706/U$1 ( \894 , \888 , \893 );
nor \mul_17_13_g20146/U$1 ( \895 , \886 , \894 );
nor \mul_17_13_g20087/U$1 ( \896 , \880 , \895 );
not \mul_17_13_g20172/U$1 ( \897 , \803 );
not \mul_17_13_g20219/U$1 ( \898 , \818 );
nand \mul_17_13_g20152/U$1 ( \899 , \897 , \898 );
or \mul_17_13_g20115/U$2 ( \900 , \895 , \899 );
nand \mul_17_13_g20150/U$1 ( \901 , \886 , \894 );
nand \mul_17_13_g20115/U$1 ( \902 , \900 , \901 );
nor \mul_17_13_g20078/U$1 ( \903 , \896 , \902 );
not \fopt35684/U$1 ( \904 , \903 );
xor \g35815/U$1 ( \905 , \784 , \904 );
not \g4878/U$3 ( \906 , \905 );
not \mul_6_11_g13545/U$3 ( \907 , \403 );
not \mul_6_11_g13545/U$4 ( \908 , \529 );
or \mul_6_11_g13545/U$2 ( \909 , \907 , \908 );
nand \mul_6_11_g13545/U$1 ( \910 , \909 , \531 );
not \mul_6_11_g13568/U$2 ( \911 , \425 );
nand \mul_6_11_g13568/U$1 ( \912 , \911 , \423 );
nor \mul_6_11_g13536/U$1 ( \913 , \910 , \912 );
not \mul_6_11_g13528/U$2 ( \914 , \913 );
nand \mul_6_11_g13535/U$1 ( \915 , \910 , \912 );
nand \mul_6_11_g13528/U$1 ( \916 , \914 , \915 );
not \fopt5205/U$1 ( \917 , \916 );
not \g4878/U$4 ( \918 , \917 );
and \g4878/U$2 ( \919 , \906 , \918 );
xor \g5024/U$1 ( \920 , \c[7] , \d[7] );
not \g4889/U$3 ( \921 , \920 );
not \g35360/U$2 ( \922 , \661 );
nand \g35360/U$1 ( \923 , \922 , \540 );
xor \g35703/U$1 ( \924 , \923 , \658 );
not \fopt5177/U$1 ( \925 , \924 );
not \g4889/U$4 ( \926 , \925 );
or \g4889/U$2 ( \927 , \921 , \926 );
xor \mul_16_12_g20591/U$1 ( \928 , \a[4] , \d[1] );
not \mul_16_12_g20389/U$3 ( \929 , \928 );
not \mul_16_12_g20670/U$2 ( \930 , \d[0] );
nand \mul_16_12_g20670/U$1 ( \931 , \930 , \d[1] );
not \mul_16_12_g20661/U$1 ( \932 , \931 );
not \mul_16_12_g20389/U$4 ( \933 , \932 );
or \mul_16_12_g20389/U$2 ( \934 , \929 , \933 );
xor \mul_16_12_g35958/U$1 ( \935 , \a[5] , \d[1] );
nand \mul_16_12_g20452/U$1 ( \936 , \935 , \d[0] );
nand \mul_16_12_g20389/U$1 ( \937 , \934 , \936 );
not \mul_16_12_g20721/U$2 ( \938 , \937 );
or \mul_16_12_g20523/U$2 ( \939 , \a[0] , \d[4] );
nand \mul_16_12_g20523/U$1 ( \940 , \939 , \d[3] );
nand \mul_16_12_g20643/U$1 ( \941 , \a[0] , \d[4] );
nand \mul_16_12_g20500/U$1 ( \942 , \940 , \941 , \d[5] );
nor \mul_16_12_g20721/U$1 ( \943 , \938 , \942 );
xor \mul_16_12_g20619/U$1 ( \944 , \a[1] , \d[5] );
not \mul_16_12_g20358/U$3 ( \945 , \944 );
xnor \mul_16_12_g20684/U$1 ( \946 , \d[5] , \d[4] );
xor \mul_16_12_g35496/U$1 ( \947 , \d[4] , \d[3] );
nor \mul_16_12_g20424/U$1 ( \948 , \946 , \947 );
not \mul_16_12_g20358/U$4 ( \949 , \948 );
or \mul_16_12_g20358/U$2 ( \950 , \945 , \949 );
buf \mul_16_12_g20548/U$1 ( \951 , \947 );
xor \mul_16_12_g20610/U$1 ( \952 , \a[2] , \d[5] );
nand \mul_16_12_g20440/U$1 ( \953 , \951 , \952 );
nand \mul_16_12_g20358/U$1 ( \954 , \950 , \953 );
not \mul_16_12_g20357/U$1 ( \955 , \954 );
xor \g35450/U$1 ( \956 , \943 , \955 );
xor \mul_16_12_g20667/U$1 ( \957 , \d[6] , \d[5] );
buf \mul_16_12_g20556/U$1 ( \958 , \957 );
and \mul_16_12_g20491/U$1 ( \959 , \958 , \a[0] );
not \mul_16_12_g20388/U$3 ( \960 , \935 );
not \mul_16_12_g20388/U$4 ( \961 , \932 );
or \mul_16_12_g20388/U$2 ( \962 , \960 , \961 );
xor \mul_16_12_g20584/U$1 ( \963 , \a[6] , \d[1] );
nand \mul_16_12_g20436/U$1 ( \964 , \963 , \d[0] );
nand \mul_16_12_g20388/U$1 ( \965 , \962 , \964 );
xor \mul_16_12_g20226/U$1 ( \966 , \959 , \965 );
xor \mul_16_12_g20606/U$1 ( \967 , \a[3] , \d[3] );
not \mul_16_12_g20368/U$3 ( \968 , \967 );
xor \mul_16_12_g35756/U$1 ( \969 , \d[2] , \d[1] );
not \mul_16_12_g20432/U$2 ( \970 , \969 );
xor \mul_16_12_g35759/U$1 ( \971 , \d[3] , \d[2] );
nand \mul_16_12_g20432/U$1 ( \972 , \970 , \971 );
not \fopt35583/U$1 ( \973 , \972 );
not \mul_16_12_g20368/U$4 ( \974 , \973 );
or \mul_16_12_g20368/U$2 ( \975 , \968 , \974 );
buf \mul_16_12_g20538/U$1 ( \976 , \969 );
xor \mul_16_12_g20594/U$1 ( \977 , \a[4] , \d[3] );
nand \mul_16_12_g20465/U$1 ( \978 , \976 , \977 );
nand \mul_16_12_g20368/U$1 ( \979 , \975 , \978 );
xor \mul_16_12_g20226/U$1_r1 ( \980 , \966 , \979 );
xnor \g35450/U$1_r1 ( \981 , \956 , \980 );
not \mul_16_12_g20151/U$1 ( \982 , \981 );
xor \mul_16_12_g20633/U$1 ( \983 , \a[0] , \d[5] );
not \mul_16_12_g20361/U$3 ( \984 , \983 );
not \mul_16_12_g20361/U$4 ( \985 , \948 );
or \mul_16_12_g20361/U$2 ( \986 , \984 , \985 );
nand \mul_16_12_g20406/U$1 ( \987 , \951 , \944 );
nand \mul_16_12_g20361/U$1 ( \988 , \986 , \987 );
not \mul_16_12_g20360/U$1 ( \989 , \988 );
not \mul_16_12_g20184/U$3 ( \990 , \989 );
not \mul_16_12_g20289/U$3 ( \991 , \937 );
not \mul_16_12_g20289/U$4 ( \992 , \942 );
and \mul_16_12_g20289/U$2 ( \993 , \991 , \992 );
and \mul_16_12_g20289/U$5 ( \994 , \937 , \942 );
nor \mul_16_12_g20289/U$1 ( \995 , \993 , \994 );
not \mul_16_12_g20184/U$4 ( \996 , \995 );
or \mul_16_12_g20184/U$2 ( \997 , \990 , \996 );
xor \mul_16_12_g20607/U$1 ( \998 , \a[2] , \d[3] );
not \mul_16_12_g20375/U$3 ( \999 , \998 );
not \mul_16_12_g20375/U$4 ( \1000 , \973 );
or \mul_16_12_g20375/U$2 ( \1001 , \999 , \1000 );
nand \mul_16_12_g20463/U$1 ( \1002 , \976 , \967 );
nand \mul_16_12_g20375/U$1 ( \1003 , \1001 , \1002 );
nand \mul_16_12_g20184/U$1 ( \1004 , \997 , \1003 );
or \mul_16_12_g20705/U$1 ( \1005 , \995 , \989 );
nand \mul_16_12_g20171/U$1 ( \1006 , \1004 , \1005 );
not \mul_16_12_g20158/U$1 ( \1007 , \1006 );
nand \mul_16_12_g20134/U$1 ( \1008 , \982 , \1007 );
not \mul_16_12_g20071/U$3 ( \1009 , \1008 );
xor \mul_16_12_g35966/U$1 ( \1010 , \988 , \995 );
xor \mul_16_12_g35966/U$1_r1 ( \1011 , \1010 , \1003 );
nand \mul_16_12_g20492/U$1 ( \1012 , \951 , \a[0] );
and \g35746/U$2 ( \1013 , \976 , \998 );
not \g35746/U$4 ( \1014 , \976 );
xor \mul_16_12_g20615/U$1 ( \1015 , \a[1] , \d[3] );
and \g35747/U$1 ( \1016 , \971 , \1015 );
and \g35746/U$3 ( \1017 , \1014 , \1016 );
nor \g35746/U$1 ( \1018 , \1013 , \1017 );
xor \mul_16_12_g20231/U$4 ( \1019 , \1012 , \1018 );
xor \mul_16_12_g35956/U$1 ( \1020 , \a[3] , \d[1] );
and \mul_16_12_g20393/U$2 ( \1021 , \932 , \1020 );
and \mul_16_12_g20676/U$1 ( \1022 , \928 , \d[0] );
nor \mul_16_12_g20393/U$1 ( \1023 , \1021 , \1022 );
and \mul_16_12_g20231/U$3 ( \1024 , \1019 , \1023 );
and \mul_16_12_g20231/U$5 ( \1025 , \1012 , \1018 );
or \mul_16_12_g20231/U$2 ( \1026 , \1024 , \1025 );
nand \mul_16_12_g20136/U$1 ( \1027 , \1011 , \1026 );
nand \mul_16_12_g20496/U$1 ( \1028 , \976 , \a[0] );
not \mul_16_12_g20719/U$2 ( \1029 , \1028 );
xor \mul_16_12_g20613/U$1 ( \1030 , \a[1] , \d[1] );
not \mul_16_12_g20397/U$3 ( \1031 , \1030 );
not \mul_16_12_g20397/U$4 ( \1032 , \932 );
or \mul_16_12_g20397/U$2 ( \1033 , \1031 , \1032 );
xor \mul_16_12_g20604/U$1 ( \1034 , \a[2] , \d[1] );
nand \mul_16_12_g20460/U$1 ( \1035 , \1034 , \d[0] );
nand \mul_16_12_g20397/U$1 ( \1036 , \1033 , \1035 );
nor \mul_16_12_g20719/U$1 ( \1037 , \1029 , \1036 );
xor \mul_16_12_g20637/U$1 ( \1038 , \a[0] , \d[1] );
not \mul_16_12_g20398/U$3 ( \1039 , \1038 );
not \mul_16_12_g20398/U$4 ( \1040 , \932 );
or \mul_16_12_g20398/U$2 ( \1041 , \1039 , \1040 );
nand \mul_16_12_g20469/U$1 ( \1042 , \1030 , \d[0] );
nand \mul_16_12_g20398/U$1 ( \1043 , \1041 , \1042 );
nand \mul_16_12_g20652/U$1 ( \1044 , \a[0] , \d[0] );
and \mul_16_12_g20517/U$1 ( \1045 , \1044 , \d[1] );
nand \mul_16_12_g20293/U$1 ( \1046 , \1043 , \1045 );
or \mul_16_12_g20242/U$2 ( \1047 , \1037 , \1046 );
not \mul_16_12_g20296/U$2 ( \1048 , \1028 );
nand \mul_16_12_g20296/U$1 ( \1049 , \1048 , \1036 );
nand \mul_16_12_g20242/U$1 ( \1050 , \1047 , \1049 );
not \mul_16_12_g20168/U$3 ( \1051 , \1050 );
not \mul_16_12_g20396/U$3 ( \1052 , \1034 );
not \mul_16_12_g20396/U$4 ( \1053 , \932 );
or \mul_16_12_g20396/U$2 ( \1054 , \1052 , \1053 );
nand \mul_16_12_g20407/U$1 ( \1055 , \d[0] , \1020 );
nand \mul_16_12_g20396/U$1 ( \1056 , \1054 , \1055 );
not \mul_16_12_g20290/U$3 ( \1057 , \1056 );
nand \mul_16_12_g20640/U$1 ( \1058 , \a[0] , \d[2] );
and \mul_16_12_g20681/U$1 ( \1059 , \1058 , \d[3] );
or \mul_16_12_g20524/U$2 ( \1060 , \a[0] , \d[2] );
nand \mul_16_12_g20524/U$1 ( \1061 , \1060 , \d[1] );
nand \mul_16_12_g20498/U$1 ( \1062 , \1059 , \1061 );
not \mul_16_12_g20290/U$4 ( \1063 , \1062 );
and \mul_16_12_g20290/U$2 ( \1064 , \1057 , \1063 );
and \mul_16_12_g20290/U$5 ( \1065 , \1056 , \1062 );
nor \mul_16_12_g20290/U$1 ( \1066 , \1064 , \1065 );
buf \fopt35582/U$1 ( \1067 , \973 );
xor \mul_16_12_g20636/U$1 ( \1068 , \a[0] , \d[3] );
nand \mul_16_12_g35657/U$1 ( \1069 , \1067 , \1068 );
nand \mul_16_12_g20448/U$1 ( \1070 , \976 , \1015 );
nand \mul_16_12_g20241/U$1 ( \1071 , \1066 , \1069 , \1070 );
not \mul_16_12_g20168/U$4 ( \1072 , \1071 );
or \mul_16_12_g20168/U$2 ( \1073 , \1051 , \1072 );
not \mul_16_12_g20704/U$2 ( \1074 , \1066 );
nand \mul_16_12_g20291/U$1 ( \1075 , \1069 , \1070 );
nand \mul_16_12_g20704/U$1 ( \1076 , \1074 , \1075 );
nand \mul_16_12_g20168/U$1 ( \1077 , \1073 , \1076 );
not \g35905/U$3 ( \1078 , \1077 );
xor \mul_16_12_g20231/U$1 ( \1079 , \1012 , \1018 );
xor \mul_16_12_g20231/U$1_r1 ( \1080 , \1079 , \1023 );
not \mul_16_12_g20720/U$2 ( \1081 , \1062 );
nand \mul_16_12_g20720/U$1 ( \1082 , \1081 , \1056 );
nand \mul_16_12_g20182/U$1 ( \1083 , \1080 , \1082 );
not \g35905/U$4 ( \1084 , \1083 );
or \g35905/U$2 ( \1085 , \1078 , \1084 );
not \mul_16_12_g20229/U$1 ( \1086 , \1080 );
not \mul_16_12_g20268/U$1 ( \1087 , \1082 );
nand \mul_16_12_g20180/U$1 ( \1088 , \1086 , \1087 );
nand \g35905/U$1 ( \1089 , \1085 , \1088 );
and \mul_16_12_g20097/U$1 ( \1090 , \1027 , \1089 );
not \mul_16_12_g20071/U$4 ( \1091 , \1090 );
or \mul_16_12_g20071/U$2 ( \1092 , \1009 , \1091 );
not \mul_16_12_g20157/U$1 ( \1093 , \1011 );
not \mul_16_12_g20230/U$1 ( \1094 , \1026 );
nand \mul_16_12_g20139/U$1 ( \1095 , \1093 , \1094 );
not \g35903/U$3 ( \1096 , \1095 );
nand \mul_16_12_g20141/U$1 ( \1097 , \981 , \1006 );
not \g35903/U$4 ( \1098 , \1097 );
or \g35903/U$2 ( \1099 , \1096 , \1098 );
nand \g35903/U$1 ( \1100 , \1099 , \1008 );
nand \mul_16_12_g20071/U$1 ( \1101 , \1092 , \1100 );
not \mul_16_12_g20048/U$3 ( \1102 , \1101 );
not \mul_16_12_g20387/U$3 ( \1103 , \963 );
not \mul_16_12_g20387/U$4 ( \1104 , \932 );
or \mul_16_12_g20387/U$2 ( \1105 , \1103 , \1104 );
xor \mul_16_12_g20583/U$1 ( \1106 , \a[7] , \d[1] );
nand \mul_16_12_g20422/U$1 ( \1107 , \1106 , \d[0] );
nand \mul_16_12_g20387/U$1 ( \1108 , \1105 , \1107 );
or \mul_16_12_g20522/U$2 ( \1109 , \a[0] , \d[6] );
nand \mul_16_12_g20522/U$1 ( \1110 , \1109 , \d[5] );
nand \mul_16_12_g20641/U$1 ( \1111 , \a[0] , \d[6] );
nand \mul_16_12_g20504/U$1 ( \1112 , \1110 , \1111 , \d[7] );
not \mul_16_12_g20503/U$1 ( \1113 , \1112 );
and \mul_16_12_g20288/U$2 ( \1114 , \1108 , \1113 );
not \mul_16_12_g20288/U$4 ( \1115 , \1108 );
and \mul_16_12_g20288/U$3 ( \1116 , \1115 , \1112 );
nor \mul_16_12_g20288/U$1 ( \1117 , \1114 , \1116 );
xor \mul_16_12_g20226/U$4 ( \1118 , \959 , \965 );
and \mul_16_12_g20226/U$3 ( \1119 , \1118 , \979 );
and \mul_16_12_g20226/U$5 ( \1120 , \959 , \965 );
or \mul_16_12_g20226/U$2 ( \1121 , \1119 , \1120 );
xor \mul_16_12_g20109/U$1 ( \1122 , \1117 , \1121 );
xor \mul_16_12_g20631/U$1 ( \1123 , \a[0] , \d[7] );
not \mul_16_12_g20329/U$3 ( \1124 , \1123 );
xor \mul_16_12_g35769/U$1 ( \1125 , \d[7] , \d[6] );
not \fopt35663/U$1 ( \1126 , \1125 );
nor \mul_16_12_g20409/U$1 ( \1127 , \957 , \1126 );
buf \fopt35575/U$1 ( \1128 , \1127 );
not \mul_16_12_g20329/U$4 ( \1129 , \1128 );
or \mul_16_12_g20329/U$2 ( \1130 , \1124 , \1129 );
xor \mul_16_12_g20624/U$1 ( \1131 , \a[1] , \d[7] );
nand \mul_16_12_g20468/U$1 ( \1132 , \958 , \1131 );
nand \mul_16_12_g20329/U$1 ( \1133 , \1130 , \1132 );
not \mul_16_12_g20353/U$3 ( \1134 , \952 );
nor \mul_16_12_g20425/U$1 ( \1135 , \946 , \947 );
not \mul_16_12_g20353/U$4 ( \1136 , \1135 );
or \mul_16_12_g20353/U$2 ( \1137 , \1134 , \1136 );
xor \mul_16_12_g20609/U$1 ( \1138 , \a[3] , \d[5] );
nand \mul_16_12_g20443/U$1 ( \1139 , \951 , \1138 );
nand \mul_16_12_g20353/U$1 ( \1140 , \1137 , \1139 );
xor \mul_16_12_g20202/U$1 ( \1141 , \1133 , \1140 );
not \mul_16_12_g20370/U$3 ( \1142 , \977 );
not \mul_16_12_g20370/U$4 ( \1143 , \1067 );
or \mul_16_12_g20370/U$2 ( \1144 , \1142 , \1143 );
xor \mul_16_12_g20593/U$1 ( \1145 , \a[5] , \d[3] );
nand \mul_16_12_g20441/U$1 ( \1146 , \976 , \1145 );
nand \mul_16_12_g20370/U$1 ( \1147 , \1144 , \1146 );
xor \mul_16_12_g20202/U$1_r1 ( \1148 , \1141 , \1147 );
xor \mul_16_12_g20109/U$1_r1 ( \1149 , \1122 , \1148 );
not \mul_16_12_g20706/U$2 ( \1150 , \943 );
nand \mul_16_12_g20706/U$1 ( \1151 , \1150 , \955 );
not \mul_16_12_g20170/U$3 ( \1152 , \1151 );
not \mul_16_12_g20170/U$4 ( \1153 , \980 );
or \mul_16_12_g20170/U$2 ( \1154 , \1152 , \1153 );
nand \mul_16_12_g20247/U$1 ( \1155 , \943 , \954 );
nand \mul_16_12_g20170/U$1 ( \1156 , \1154 , \1155 );
or \g35902/U$2 ( \1157 , \1149 , \1156 );
nand \mul_16_12_g20672/U$1 ( \1158 , \1149 , \1156 );
nand \g35902/U$1 ( \1159 , \1157 , \1158 );
not \mul_16_12_g20048/U$4 ( \1160 , \1159 );
or \mul_16_12_g20048/U$2 ( \1161 , \1102 , \1160 );
or \mul_16_12_g20048/U$5 ( \1162 , \1159 , \1101 );
nand \mul_16_12_g20048/U$1 ( \1163 , \1161 , \1162 );
and \mul_6_11_g13992/U$1 ( \1164 , \403 , \531 );
buf \mul_6_11_g13564/U$1 ( \1165 , \529 );
xor \mul_6_11_g13991/U$1 ( \1166 , \1164 , \1165 );
not \fopt35537/U$1 ( \1167 , \1166 );
not \fopt35538/U$1 ( \1168 , \1167 );
and \g4907/U$2 ( \1169 , \1163 , \1168 );
nor \add_15_12_g7242/U$1 ( \1170 , \b[2] , \d[2] );
nor \add_15_12_g7236/U$1 ( \1171 , \b[3] , \d[3] );
nor \add_15_12_g7218/U$1 ( \1172 , \1170 , \1171 );
not \add_15_12_g7167/U$3 ( \1173 , \1172 );
nand \add_15_12_g7275/U$1 ( \1174 , \b[0] , \d[0] );
not \add_15_12_g7200/U$1 ( \1175 , \1174 );
not \add_15_12_g7175/U$3 ( \1176 , \1175 );
or \add_15_12_g7276/U$1 ( \1177 , \b[1] , \d[1] );
not \add_15_12_g7175/U$4 ( \1178 , \1177 );
or \add_15_12_g7175/U$2 ( \1179 , \1176 , \1178 );
nand \add_15_12_g7262/U$1 ( \1180 , \b[1] , \d[1] );
nand \add_15_12_g7175/U$1 ( \1181 , \1179 , \1180 );
not \add_15_12_g7167/U$4 ( \1182 , \1181 );
or \add_15_12_g7167/U$2 ( \1183 , \1173 , \1182 );
nand \add_15_12_g7268/U$1 ( \1184 , \b[3] , \d[3] );
not \add_15_12_g7280/U$2 ( \1185 , \1184 );
nand \add_15_12_g7257/U$1 ( \1186 , \b[2] , \d[2] );
nor \add_15_12_g7210/U$1 ( \1187 , \1171 , \1186 );
nor \add_15_12_g7280/U$1 ( \1188 , \1185 , \1187 );
nand \add_15_12_g7167/U$1 ( \1189 , \1183 , \1188 );
nor \add_15_12_g7234/U$1 ( \1190 , \b[4] , \d[4] );
not \add_15_12_g7279/U$2 ( \1191 , \1190 );
or \add_15_12_g2/U$1 ( \1192 , \b[5] , \d[5] );
nand \add_15_12_g7279/U$1 ( \1193 , \1191 , \1192 );
nor \add_15_12_g7231/U$1 ( \1194 , \b[6] , \d[6] );
nor \add_15_12_g7189/U$1 ( \1195 , \1193 , \1194 );
nand \add_15_12_g7161/U$1 ( \1196 , \1189 , \1195 );
nand \add_15_12_g7245/U$1 ( \1197 , \b[4] , \d[4] );
not \add_15_12_g7244/U$1 ( \1198 , \1197 );
nand \add_15_12_g7203/U$1 ( \1199 , \1192 , \1198 );
nand \add_15_12_g7256/U$1 ( \1200 , \b[5] , \d[5] );
nand \add_15_12_g7188/U$1 ( \1201 , \1199 , \1200 );
not \add_15_12_g7229/U$1 ( \1202 , \1194 );
and \add_15_12_g7176/U$2 ( \1203 , \1201 , \1202 );
nand \add_15_12_g7239/U$1 ( \1204 , \b[6] , \d[6] );
not \add_15_12_g7238/U$1 ( \1205 , \1204 );
nor \add_15_12_g7176/U$1 ( \1206 , \1203 , \1205 );
nand \add_15_12_g7156/U$1 ( \1207 , \1196 , \1206 );
nor \add_15_12_g7261/U$1 ( \1208 , \b[7] , \d[7] );
not \add_15_12_g7260/U$1 ( \1209 , \1208 );
nand \add_15_12_g7272/U$1 ( \1210 , \b[7] , \d[7] );
nand \add_15_12_g7212/U$1 ( \1211 , \1209 , \1210 );
xnor \add_15_12_g7278/U$1 ( \1212 , \1207 , \1211 );
not \g4923/U$3 ( \1213 , \1212 );
not \mul_6_11_g35610/U$1 ( \1214 , \447 );
not \mul_6_11_g13601/U$3 ( \1215 , \1214 );
not \mul_6_11_g13601/U$4 ( \1216 , \457 );
or \mul_6_11_g13601/U$2 ( \1217 , \1215 , \1216 );
nand \mul_6_11_g13601/U$1 ( \1218 , \1217 , \528 );
buf \mul_6_11_g13594/U$1 ( \1219 , \524 );
xnor \g35816/U$1 ( \1220 , \1218 , \1219 );
not \g4923/U$4 ( \1221 , \1220 );
or \g4923/U$2 ( \1222 , \1213 , \1221 );
buf \fopt35585/U$1 ( \1223 , \519 );
not \mul_6_11_g13602/U$3 ( \1224 , \1223 );
not \mul_6_11_g13624/U$3 ( \1225 , \472 );
not \mul_6_11_g13624/U$4 ( \1226 , \483 );
or \mul_6_11_g13624/U$2 ( \1227 , \1225 , \1226 );
nand \mul_6_11_g13624/U$1 ( \1228 , \1227 , \523 );
not \mul_6_11_g13602/U$4 ( \1229 , \1228 );
or \mul_6_11_g13602/U$2 ( \1230 , \1224 , \1229 );
or \mul_6_11_g13995/U$1 ( \1231 , \1228 , \1223 );
nand \mul_6_11_g13602/U$1 ( \1232 , \1230 , \1231 );
nor \add_14_12_g7242/U$1 ( \1233 , \a[2] , \c[2] );
nor \add_14_12_g7236/U$1 ( \1234 , \a[3] , \c[3] );
nor \add_14_12_g7218/U$1 ( \1235 , \1233 , \1234 );
not \add_14_12_g7167/U$3 ( \1236 , \1235 );
nand \add_14_12_g7275/U$1 ( \1237 , \a[0] , \c[0] );
not \add_14_12_g7200/U$1 ( \1238 , \1237 );
not \add_14_12_g7175/U$3 ( \1239 , \1238 );
or \add_14_12_g7276/U$1 ( \1240 , \a[1] , \c[1] );
not \add_14_12_g7175/U$4 ( \1241 , \1240 );
or \add_14_12_g7175/U$2 ( \1242 , \1239 , \1241 );
nand \add_14_12_g7262/U$1 ( \1243 , \a[1] , \c[1] );
nand \add_14_12_g7175/U$1 ( \1244 , \1242 , \1243 );
not \add_14_12_g7167/U$4 ( \1245 , \1244 );
or \add_14_12_g7167/U$2 ( \1246 , \1236 , \1245 );
nand \add_14_12_g7268/U$1 ( \1247 , \a[3] , \c[3] );
not \add_14_12_g7280/U$2 ( \1248 , \1247 );
nand \add_14_12_g7257/U$1 ( \1249 , \a[2] , \c[2] );
nor \add_14_12_g7210/U$1 ( \1250 , \1234 , \1249 );
nor \add_14_12_g7280/U$1 ( \1251 , \1248 , \1250 );
nand \add_14_12_g7167/U$1 ( \1252 , \1246 , \1251 );
nor \add_14_12_g7234/U$1 ( \1253 , \a[4] , \c[4] );
not \add_14_12_g7279/U$2 ( \1254 , \1253 );
or \add_14_12_g2/U$1 ( \1255 , \a[5] , \c[5] );
nand \add_14_12_g7279/U$1 ( \1256 , \1254 , \1255 );
nor \add_14_12_g7231/U$1 ( \1257 , \a[6] , \c[6] );
nor \add_14_12_g7189/U$1 ( \1258 , \1256 , \1257 );
nand \add_14_12_g7161/U$1 ( \1259 , \1252 , \1258 );
nand \add_14_12_g7245/U$1 ( \1260 , \a[4] , \c[4] );
not \add_14_12_g7244/U$1 ( \1261 , \1260 );
nand \add_14_12_g7203/U$1 ( \1262 , \1255 , \1261 );
nand \add_14_12_g7256/U$1 ( \1263 , \a[5] , \c[5] );
nand \add_14_12_g7188/U$1 ( \1264 , \1262 , \1263 );
not \add_14_12_g7229/U$1 ( \1265 , \1257 );
and \add_14_12_g7176/U$2 ( \1266 , \1264 , \1265 );
nand \add_14_12_g7239/U$1 ( \1267 , \a[6] , \c[6] );
not \add_14_12_g7238/U$1 ( \1268 , \1267 );
nor \add_14_12_g7176/U$1 ( \1269 , \1266 , \1268 );
nand \add_14_12_g7156/U$1 ( \1270 , \1259 , \1269 );
nor \add_14_12_g7261/U$1 ( \1271 , \a[7] , \c[7] );
not \add_14_12_g7260/U$1 ( \1272 , \1271 );
nand \add_14_12_g7272/U$1 ( \1273 , \a[7] , \c[7] );
nand \add_14_12_g7212/U$1 ( \1274 , \1272 , \1273 );
xnor \add_14_12_g7278/U$1 ( \1275 , \1270 , \1274 );
and \g4943/U$2 ( \1276 , \1232 , \1275 );
not \g4968/U$3 ( \1277 , \d[7] );
nand \mul_6_11_g13665/U$1 ( \1278 , \518 , \498 );
buf \mul_6_11_g13675/U$1 ( \1279 , \515 );
xnor \mul_6_11_g14003/U$1 ( \1280 , \1278 , \1279 );
not \g5173/U$1 ( \1281 , \1280 );
not \g5167/U$1 ( \1282 , \1281 );
not \g4968/U$4 ( \1283 , \1282 );
or \g4968/U$2 ( \1284 , \1277 , \1283 );
not \mul_6_11_g13711/U$2 ( \1285 , \506 );
nand \mul_6_11_g13711/U$1 ( \1286 , \1285 , \514 );
xor \mul_6_11_g14007/U$1 ( \1287 , \1286 , \512 );
and \g5005/U$2 ( \1288 , \1287 , \c[7] );
not \mul_6_11_g13763/U$3 ( \1289 , \b[0] );
not \mul_6_11_g13763/U$4 ( \1290 , \499 );
or \mul_6_11_g13763/U$2 ( \1291 , \1289 , \1290 );
nand \mul_6_11_g13763/U$1 ( \1292 , \1291 , \508 );
and \mul_6_11_g13979/U$1 ( \1293 , \512 , \1292 );
and \g5060/U$1 ( \1294 , \1293 , \b[7] );
nor \g5005/U$1 ( \1295 , \1288 , \1294 );
nand \g4968/U$1 ( \1296 , \1284 , \1295 );
nor \g4943/U$1 ( \1297 , \1276 , \1296 );
nand \g4923/U$1 ( \1298 , \1222 , \1297 );
nor \g4907/U$1 ( \1299 , \1169 , \1298 );
nand \g4889/U$1 ( \1300 , \927 , \1299 );
nor \g4878/U$1 ( \1301 , \919 , \1300 );
nand \g4855/U$1 ( \1302 , \674 , \1301 );
not \g5238/U$2 ( \1303 , \1302 );
nand \mul_6_11_g13539/U$1 ( \1304 , \551 , \328 );
not \mul_6_11_g13988/U$2 ( \1305 , \1304 );
nor \mul_6_11_g13988/U$1 ( \1306 , \1305 , \541 );
not \mul_6_11_g13533/U$2 ( \1307 , \544 );
not \mul_6_11_g13548/U$1 ( \1308 , \283 );
nand \mul_6_11_g13533/U$1 ( \1309 , \1307 , \1308 );
nand \mul_6_11_g13524/U$1 ( \1310 , \1309 , \284 );
and \mul_6_11_g13518/U$2 ( \1311 , \1306 , \1310 );
not \mul_6_11_g13518/U$4 ( \1312 , \1306 );
not \mul_6_11_g13523/U$1 ( \1313 , \1310 );
and \mul_6_11_g13518/U$3 ( \1314 , \1312 , \1313 );
nor \mul_6_11_g13518/U$1 ( \1315 , \1311 , \1314 );
buf \fopt35669/U$1 ( \1316 , \1315 );
and \g5039/U$1 ( \1317 , \b[7] , \c[7] );
nand \g4988/U$1 ( \1318 , \1316 , \1317 );
not \g4860/U$2 ( \1319 , \1316 );
not \fopt5183/U$1 ( \1320 , \924 );
not \g35820/U$2 ( \1321 , \1320 );
not \g5251/U$2 ( \1322 , \1232 );
not \fopt35570/U$1 ( \1323 , \1287 );
not \g5114/U$1 ( \1324 , \1293 );
nand \g5097/U$1 ( \1325 , \1323 , \1324 );
nor \g4990/U$1 ( \1326 , \1280 , \1325 );
nand \g5251/U$1 ( \1327 , \1322 , \1326 );
nor \g4935/U$1 ( \1328 , \1220 , \1327 );
nand \g4929/U$1 ( \1329 , \1167 , \1328 );
nor \g4902/U$1 ( \1330 , \916 , \1329 );
nand \g35820/U$1 ( \1331 , \1321 , \1330 );
nor \g4866/U$1 ( \1332 , \1331 , \648 );
nand \g4860/U$1 ( \1333 , \1319 , \1332 );
nand \g5238/U$1 ( \1334 , \1303 , \1318 , \1333 );
nor \g35731/U$1 ( \1335 , \646 , \1334 );
not \g4807/U$1 ( \1336 , \1335 );
not \g4809/U$3 ( \1337 , \a[1] );
nor \g4867/U$1 ( \1338 , \1316 , \1331 );
not \g4809/U$4 ( \1339 , \1338 );
or \g4809/U$2 ( \1340 , \1337 , \1339 );
not \fopt35682/U$1 ( \1341 , \643 );
not \fopt35679/U$1 ( \1342 , \1341 );
or \g5087/U$1 ( \1343 , \a[1] , \d[1] );
and \g4824/U$2 ( \1344 , \1342 , \1343 );
and \g5045/U$1 ( \1345 , \b[1] , \c[1] );
not \g4842/U$3 ( \1346 , \1345 );
not \g4842/U$4 ( \1347 , \1316 );
or \g4842/U$2 ( \1348 , \1346 , \1347 );
or \g5042/U$1 ( \1349 , \a[1] , \b[1] );
not \g5120/U$1 ( \1350 , \671 );
not \g5117/U$1 ( \1351 , \1350 );
and \g4853/U$2 ( \1352 , \1349 , \1351 );
not \fopt35536/U$1 ( \1353 , \1167 );
or \mul_16_12_g20294/U$1 ( \1354 , \1043 , \1045 );
and \mul_16_12_g20286/U$1 ( \1355 , \1354 , \1046 );
and \g4901/U$2 ( \1356 , \1353 , \1355 );
not \add_15_12_g7182/U$3 ( \1357 , \1175 );
nand \add_15_12_g7201/U$1 ( \1358 , \1177 , \1180 );
not \add_15_12_g7182/U$4 ( \1359 , \1358 );
or \add_15_12_g7182/U$2 ( \1360 , \1357 , \1359 );
or \add_15_12_g7182/U$5 ( \1361 , \1358 , \1175 );
nand \add_15_12_g7182/U$1 ( \1362 , \1360 , \1361 );
not \g4920/U$3 ( \1363 , \1362 );
not \g4920/U$4 ( \1364 , \1220 );
or \g4920/U$2 ( \1365 , \1363 , \1364 );
not \add_14_12_g7182/U$3 ( \1366 , \1238 );
nand \add_14_12_g7201/U$1 ( \1367 , \1240 , \1243 );
not \add_14_12_g7182/U$4 ( \1368 , \1367 );
or \add_14_12_g7182/U$2 ( \1369 , \1366 , \1368 );
or \add_14_12_g7182/U$5 ( \1370 , \1367 , \1238 );
nand \add_14_12_g7182/U$1 ( \1371 , \1369 , \1370 );
and \g4939/U$2 ( \1372 , \1232 , \1371 );
not \g4962/U$3 ( \1373 , \d[1] );
not \g4962/U$4 ( \1374 , \1282 );
or \g4962/U$2 ( \1375 , \1373 , \1374 );
and \g4997/U$2 ( \1376 , \1287 , \c[1] );
and \g5040/U$1 ( \1377 , \1293 , \b[1] );
nor \g4997/U$1 ( \1378 , \1376 , \1377 );
nand \g4962/U$1 ( \1379 , \1375 , \1378 );
nor \g4939/U$1 ( \1380 , \1372 , \1379 );
nand \g4920/U$1 ( \1381 , \1365 , \1380 );
nor \g4901/U$1 ( \1382 , \1356 , \1381 );
not \fopt5178/U$1 ( \1383 , \924 );
xor \g5020/U$1 ( \1384 , \c[1] , \d[1] );
nand \g4956/U$1 ( \1385 , \1383 , \1384 );
not \mul_17_13_g20406/U$1 ( \1386 , \860 );
and \mul_17_13_g20295/U$2 ( \1387 , \1386 , \853 );
not \mul_17_13_g20301/U$1 ( \1388 , \861 );
nor \mul_17_13_g20295/U$1 ( \1389 , \1387 , \1388 );
nand \g5043/U$1 ( \1390 , \916 , \1389 );
nand \g4874/U$1 ( \1391 , \1382 , \1385 , \1390 );
nor \g4853/U$1 ( \1392 , \1352 , \1391 );
nand \g4842/U$1 ( \1393 , \1348 , \1392 );
nor \g4824/U$1 ( \1394 , \1344 , \1393 );
nand \g4809/U$1 ( \1395 , \1340 , \1394 );
not \g4833/U$3 ( \1396 , \a[4] );
nor \g4871/U$1 ( \1397 , \1316 , \1331 );
not \g4833/U$4 ( \1398 , \1397 );
or \g4833/U$2 ( \1399 , \1396 , \1398 );
and \g5074/U$1 ( \1400 , \b[4] , \c[4] );
and \g4844/U$2 ( \1401 , \1400 , \1316 );
or \g5084/U$1 ( \1402 , \a[4] , \b[4] );
not \g4857/U$3 ( \1403 , \1402 );
not \g4857/U$4 ( \1404 , \671 );
or \g4857/U$2 ( \1405 , \1403 , \1404 );
xor \g5030/U$1 ( \1406 , \c[4] , \d[4] );
nand \g4957/U$1 ( \1407 , \1383 , \1406 );
nand \mul_17_13_g20734/U$1 ( \1408 , \875 , \878 );
xnor \g35357/U$1 ( \1409 , \869 , \1408 );
nand \g35356/U$1 ( \1410 , \1409 , \916 );
nand \mul_16_12_g20163/U$1 ( \1411 , \1088 , \1083 );
xnor \mul_16_12_g20145/U$1 ( \1412 , \1411 , \1077 );
and \g4913/U$2 ( \1413 , \1168 , \1412 );
nor \add_15_12_g7224/U$1 ( \1414 , \1198 , \1190 );
not \add_15_12_g7158/U$3 ( \1415 , \1414 );
not \add_15_12_g7166/U$1 ( \1416 , \1189 );
not \add_15_12_g7158/U$4 ( \1417 , \1416 );
or \add_15_12_g7158/U$2 ( \1418 , \1415 , \1417 );
or \add_15_12_g7158/U$5 ( \1419 , \1416 , \1414 );
nand \add_15_12_g7158/U$1 ( \1420 , \1418 , \1419 );
not \g4926/U$3 ( \1421 , \1420 );
not \g4926/U$4 ( \1422 , \1220 );
or \g4926/U$2 ( \1423 , \1421 , \1422 );
nor \add_14_12_g7224/U$1 ( \1424 , \1261 , \1253 );
not \add_14_12_g7158/U$3 ( \1425 , \1424 );
not \add_14_12_g7166/U$1 ( \1426 , \1252 );
not \add_14_12_g7158/U$4 ( \1427 , \1426 );
or \add_14_12_g7158/U$2 ( \1428 , \1425 , \1427 );
or \add_14_12_g7158/U$5 ( \1429 , \1426 , \1424 );
nand \add_14_12_g7158/U$1 ( \1430 , \1428 , \1429 );
and \g4950/U$2 ( \1431 , \1232 , \1430 );
not \g4977/U$3 ( \1432 , \d[4] );
not \g4977/U$4 ( \1433 , \1280 );
or \g4977/U$2 ( \1434 , \1432 , \1433 );
not \fopt35566/U$1 ( \1435 , \1323 );
and \g35871/U$2 ( \1436 , \1435 , \c[4] );
and \g35871/U$3 ( \1437 , \1293 , \b[4] );
nor \g35871/U$1 ( \1438 , \1436 , \1437 );
nand \g4977/U$1 ( \1439 , \1434 , \1438 );
nor \g4950/U$1 ( \1440 , \1431 , \1439 );
nand \g4926/U$1 ( \1441 , \1423 , \1440 );
nor \g4913/U$1 ( \1442 , \1413 , \1441 );
and \g4881/U$1 ( \1443 , \1407 , \1410 , \1442 );
nand \g4857/U$1 ( \1444 , \1405 , \1443 );
nor \g4844/U$1 ( \1445 , \1401 , \1444 );
nand \g4833/U$1 ( \1446 , \1399 , \1445 );
not \g5013/U$3 ( \1447 , \d[4] );
not \g5013/U$4 ( \1448 , \644 );
or \g5013/U$2 ( \1449 , \1447 , \1448 );
not \fopt35680/U$1 ( \1450 , \1341 );
nand \g5052/U$1 ( \1451 , \1450 , \a[4] );
nand \g5013/U$1 ( \1452 , \1449 , \1451 );
nor \g4811/U$1 ( \1453 , \1446 , \1452 );
not \g4810/U$1 ( \1454 , \1453 );
or \g5068/U$1 ( \1455 , \a[3] , \d[3] );
not \g4825/U$3 ( \1456 , \1455 );
not \fopt35681/U$1 ( \1457 , \1341 );
not \g4825/U$4 ( \1458 , \1457 );
or \g4825/U$2 ( \1459 , \1456 , \1458 );
and \g5047/U$1 ( \1460 , \b[3] , \c[3] );
and \g4845/U$2 ( \1461 , \1316 , \1460 );
not \g5080/U$2 ( \1462 , \a[3] );
not \g5157/U$1 ( \1463 , \b[3] );
nand \g5080/U$1 ( \1464 , \1462 , \1463 );
not \g4858/U$3 ( \1465 , \1464 );
not \g5116/U$1 ( \1466 , \1350 );
not \g4858/U$4 ( \1467 , \1466 );
or \g4858/U$2 ( \1468 , \1465 , \1467 );
not \g4882/U$3 ( \1469 , \917 );
nand \mul_17_13_g20232/U$1 ( \1470 , \868 , \842 );
xor \g35358/U$1 ( \1471 , \864 , \1470 );
not \g4882/U$4 ( \1472 , \1471 );
and \g4882/U$2 ( \1473 , \1469 , \1472 );
xor \g5033/U$1 ( \1474 , \c[3] , \d[3] );
not \g4892/U$3 ( \1475 , \1474 );
not \g4892/U$4 ( \1476 , \1320 );
or \g4892/U$2 ( \1477 , \1475 , \1476 );
not \fopt35535/U$1 ( \1478 , \1167 );
nand \mul_16_12_g20204/U$1 ( \1479 , \1071 , \1076 );
xnor \mul_16_12_g20701/U$1 ( \1480 , \1479 , \1050 );
and \g4915/U$2 ( \1481 , \1478 , \1480 );
not \add_15_12_g7235/U$1 ( \1482 , \1171 );
nand \add_15_12_g7225/U$1 ( \1483 , \1482 , \1184 );
not \add_15_12_g7162/U$3 ( \1484 , \1483 );
nand \add_15_12_g7183/U$1 ( \1485 , \1174 , \1180 );
not \add_15_12_g7240/U$1 ( \1486 , \1170 );
nand \add_15_12_g7181/U$1 ( \1487 , \1485 , \1177 , \1486 );
nand \add_15_12_g7170/U$1 ( \1488 , \1487 , \1186 );
not \add_15_12_g7162/U$4 ( \1489 , \1488 );
or \add_15_12_g7162/U$2 ( \1490 , \1484 , \1489 );
or \add_15_12_g7162/U$5 ( \1491 , \1488 , \1483 );
nand \add_15_12_g7162/U$1 ( \1492 , \1490 , \1491 );
not \g4927/U$3 ( \1493 , \1492 );
not \g4927/U$4 ( \1494 , \1220 );
or \g4927/U$2 ( \1495 , \1493 , \1494 );
not \add_14_12_g7235/U$1 ( \1496 , \1234 );
nand \add_14_12_g7225/U$1 ( \1497 , \1496 , \1247 );
not \add_14_12_g7162/U$3 ( \1498 , \1497 );
nand \add_14_12_g7183/U$1 ( \1499 , \1237 , \1243 );
not \add_14_12_g7240/U$1 ( \1500 , \1233 );
nand \add_14_12_g7181/U$1 ( \1501 , \1499 , \1240 , \1500 );
nand \add_14_12_g7170/U$1 ( \1502 , \1501 , \1249 );
not \add_14_12_g7162/U$4 ( \1503 , \1502 );
or \add_14_12_g7162/U$2 ( \1504 , \1498 , \1503 );
or \add_14_12_g7162/U$5 ( \1505 , \1502 , \1497 );
nand \add_14_12_g7162/U$1 ( \1506 , \1504 , \1505 );
and \g4953/U$2 ( \1507 , \1232 , \1506 );
not \g4980/U$3 ( \1508 , \d[3] );
not \g4980/U$4 ( \1509 , \1280 );
or \g4980/U$2 ( \1510 , \1508 , \1509 );
not \g5017/U$3 ( \1511 , \1324 );
not \g5017/U$4 ( \1512 , \1463 );
and \g5017/U$2 ( \1513 , \1511 , \1512 );
not \fopt35567/U$1 ( \1514 , \1323 );
and \g5017/U$5 ( \1515 , \1514 , \c[3] );
nor \g5017/U$1 ( \1516 , \1513 , \1515 );
nand \g4980/U$1 ( \1517 , \1510 , \1516 );
nor \g4953/U$1 ( \1518 , \1507 , \1517 );
nand \g4927/U$1 ( \1519 , \1495 , \1518 );
nor \g4915/U$1 ( \1520 , \1481 , \1519 );
nand \g4892/U$1 ( \1521 , \1477 , \1520 );
nor \g4882/U$1 ( \1522 , \1473 , \1521 );
nand \g4858/U$1 ( \1523 , \1468 , \1522 );
nor \g4845/U$1 ( \1524 , \1461 , \1523 );
nand \g4825/U$1 ( \1525 , \1459 , \1524 );
and \g4850/U$1 ( \1526 , \1338 , \a[3] );
nor \g4813/U$1 ( \1527 , \1525 , \1526 );
not \g4812/U$1 ( \1528 , \1527 );
buf \fopt35533/U$1 ( \1529 , \1478 );
not \g35631/U$3 ( \1530 , \1529 );
xor \mul_16_12_g20581/U$1 ( \1531 , \a[9] , \d[7] );
not \mul_16_12_g20338/U$3 ( \1532 , \1531 );
not \mul_16_12_g20338/U$4 ( \1533 , \958 );
or \mul_16_12_g20338/U$2 ( \1534 , \1532 , \1533 );
xor \mul_16_12_g20580/U$1 ( \1535 , \a[8] , \d[7] );
nand \mul_16_12_g20382/U$1 ( \1536 , \1128 , \1535 );
nand \mul_16_12_g20338/U$1 ( \1537 , \1534 , \1536 );
xor \mul_16_12_g20595/U$1 ( \1538 , \a[6] , \d[9] );
not \mul_16_12_g20325/U$3 ( \1539 , \1538 );
xnor \mul_16_12_g20685/U$1 ( \1540 , \d[9] , \d[8] );
xor \mul_16_12_g20669/U$1 ( \1541 , \d[8] , \d[7] );
nor \mul_16_12_g20671/U$1 ( \1542 , \1540 , \1541 );
not \mul_16_12_g20325/U$4 ( \1543 , \1542 );
or \mul_16_12_g20325/U$2 ( \1544 , \1539 , \1543 );
buf \mul_16_12_g20562/U$1 ( \1545 , \1541 );
xor \mul_16_12_g20596/U$1 ( \1546 , \a[7] , \d[9] );
nand \mul_16_12_g20457/U$1 ( \1547 , \1545 , \1546 );
nand \mul_16_12_g20325/U$1 ( \1548 , \1544 , \1547 );
xor \mul_16_12_g35502/U$1 ( \1549 , \1537 , \1548 );
xor \mul_16_12_g20635/U$1 ( \1550 , \a[2] , \d[13] );
not \mul_16_12_g20305/U$3 ( \1551 , \1550 );
xor \mul_16_12_g35704/U$1 ( \1552 , \d[12] , \d[11] );
xnor \mul_16_12_g20683/U$1 ( \1553 , \d[13] , \d[12] );
nor \mul_16_12_g20516/U$1 ( \1554 , \1552 , \1553 );
not \mul_16_12_g20305/U$4 ( \1555 , \1554 );
or \mul_16_12_g20305/U$2 ( \1556 , \1551 , \1555 );
xor \mul_16_12_g20634/U$1 ( \1557 , \a[3] , \d[13] );
nand \mul_16_12_g20442/U$1 ( \1558 , \1552 , \1557 );
nand \mul_16_12_g20305/U$1 ( \1559 , \1556 , \1558 );
xor \mul_16_12_g20608/U$1 ( \1560 , \d[15] , \d[14] );
xor \mul_16_12_g20564/U$1 ( \1561 , \a[0] , \d[15] );
nand \mul_16_12_g20478/U$1 ( \1562 , \1560 , \1561 );
xor \mul_16_12_g35960/U$1 ( \1563 , \d[14] , \d[13] );
or \mul_16_12_g20303/U$2 ( \1564 , \1562 , \1563 );
xor \mul_16_12_g20582/U$1 ( \1565 , \a[1] , \d[15] );
nand \mul_16_12_g20461/U$1 ( \1566 , \1563 , \1565 );
nand \mul_16_12_g20303/U$1 ( \1567 , \1564 , \1566 );
xor \mul_16_12_g20707/U$1 ( \1568 , \1559 , \1567 );
xor \mul_16_12_g35502/U$1_r1 ( \1569 , \1549 , \1568 );
not \mul_16_12_g20146/U$3 ( \1570 , \1569 );
and \mul_16_12_g20675/U$1 ( \1571 , \1563 , \a[0] );
xor \mul_16_12_g20543/U$1 ( \1572 , \a[13] , \d[1] );
not \mul_16_12_g20403/U$3 ( \1573 , \1572 );
not \mul_16_12_g20403/U$4 ( \1574 , \932 );
or \mul_16_12_g20403/U$2 ( \1575 , \1573 , \1574 );
xor \mul_16_12_g20545/U$1 ( \1576 , \a[14] , \d[1] );
nand \mul_16_12_g20483/U$1 ( \1577 , \1576 , \d[0] );
nand \mul_16_12_g20403/U$1 ( \1578 , \1575 , \1577 );
xor \mul_16_12_g20215/U$4 ( \1579 , \1571 , \1578 );
xor \mul_16_12_g20546/U$1 ( \1580 , \a[11] , \d[3] );
not \mul_16_12_g20381/U$3 ( \1581 , \1580 );
not \mul_16_12_g20381/U$4 ( \1582 , \973 );
or \mul_16_12_g20381/U$2 ( \1583 , \1581 , \1582 );
xor \mul_16_12_g20550/U$1 ( \1584 , \a[12] , \d[3] );
nand \mul_16_12_g20493/U$1 ( \1585 , \976 , \1584 );
nand \mul_16_12_g20381/U$1 ( \1586 , \1583 , \1585 );
and \mul_16_12_g20215/U$3 ( \1587 , \1579 , \1586 );
and \mul_16_12_g20215/U$5 ( \1588 , \1571 , \1578 );
or \mul_16_12_g20215/U$2 ( \1589 , \1587 , \1588 );
not \mul_16_12_g20174/U$3 ( \1590 , \1589 );
not \mul_16_12_g20380/U$3 ( \1591 , \1584 );
not \mul_16_12_g20380/U$4 ( \1592 , \973 );
or \mul_16_12_g20380/U$2 ( \1593 , \1591 , \1592 );
not \mul_16_12_g20645/U$2 ( \1594 , \d[3] );
nand \mul_16_12_g20645/U$1 ( \1595 , \1594 , \a[13] );
not \mul_16_12_g20494/U$3 ( \1596 , \1595 );
not \mul_16_12_g20639/U$2 ( \1597 , \a[13] );
nand \mul_16_12_g20639/U$1 ( \1598 , \1597 , \d[3] );
not \mul_16_12_g20494/U$4 ( \1599 , \1598 );
or \mul_16_12_g20494/U$2 ( \1600 , \1596 , \1599 );
nand \mul_16_12_g20494/U$1 ( \1601 , \1600 , \976 );
nand \mul_16_12_g20380/U$1 ( \1602 , \1593 , \1601 );
xor \mul_16_12_g20558/U$1 ( \1603 , \a[10] , \d[5] );
not \mul_16_12_g20365/U$3 ( \1604 , \1603 );
not \mul_16_12_g20365/U$4 ( \1605 , \1135 );
or \mul_16_12_g20365/U$2 ( \1606 , \1604 , \1605 );
not \mul_16_12_g20648/U$2 ( \1607 , \d[5] );
nand \mul_16_12_g20648/U$1 ( \1608 , \1607 , \a[11] );
not \mul_16_12_g20477/U$3 ( \1609 , \1608 );
not \mul_16_12_g20647/U$2 ( \1610 , \a[11] );
nand \mul_16_12_g20647/U$1 ( \1611 , \1610 , \d[5] );
not \mul_16_12_g20477/U$4 ( \1612 , \1611 );
or \mul_16_12_g20477/U$2 ( \1613 , \1609 , \1612 );
nand \mul_16_12_g20477/U$1 ( \1614 , \1613 , \951 );
nand \mul_16_12_g20365/U$1 ( \1615 , \1606 , \1614 );
not \mul_16_12_g35967/U$2 ( \1616 , \1615 );
xor \mul_16_12_g35967/U$1 ( \1617 , \1602 , \1616 );
not \mul_16_12_g20174/U$4 ( \1618 , \1617 );
and \mul_16_12_g20174/U$2 ( \1619 , \1590 , \1618 );
and \mul_16_12_g20174/U$5 ( \1620 , \1589 , \1617 );
nor \mul_16_12_g20174/U$1 ( \1621 , \1619 , \1620 );
not \mul_16_12_g20146/U$4 ( \1622 , \1621 );
or \mul_16_12_g20146/U$2 ( \1623 , \1570 , \1622 );
or \mul_16_12_g20146/U$5 ( \1624 , \1569 , \1621 );
nand \mul_16_12_g20146/U$1 ( \1625 , \1623 , \1624 );
not \mul_16_12_g20056/U$3 ( \1626 , \1625 );
xor \mul_16_12_g20630/U$1 ( \1627 , \a[1] , \d[13] );
not \mul_16_12_g20304/U$3 ( \1628 , \1627 );
not \mul_16_12_g20304/U$4 ( \1629 , \1554 );
or \mul_16_12_g20304/U$2 ( \1630 , \1628 , \1629 );
nand \mul_16_12_g20449/U$1 ( \1631 , \1552 , \1550 );
nand \mul_16_12_g20304/U$1 ( \1632 , \1630 , \1631 );
xor \mul_16_12_g20627/U$1 ( \1633 , \a[3] , \d[11] );
not \mul_16_12_g20312/U$3 ( \1634 , \1633 );
xor \mul_16_12_g35740/U$1 ( \1635 , \d[10] , \d[9] );
not \mul_16_12_g36020/U$2 ( \1636 , \d[10] );
xor \mul_16_12_g36020/U$1 ( \1637 , \d[11] , \1636 );
nor \mul_16_12_g20514/U$1 ( \1638 , \1635 , \1637 );
not \mul_16_12_g20312/U$4 ( \1639 , \1638 );
or \mul_16_12_g20312/U$2 ( \1640 , \1634 , \1639 );
xor \g35739/U$1 ( \1641 , \d[10] , \d[9] );
xor \mul_16_12_g20621/U$1 ( \1642 , \a[4] , \d[11] );
nand \mul_16_12_g20444/U$1 ( \1643 , \1641 , \1642 );
nand \mul_16_12_g20312/U$1 ( \1644 , \1640 , \1643 );
xor \mul_16_12_g20154/U$4 ( \1645 , \1632 , \1644 );
or \mul_16_12_g20519/U$2 ( \1646 , \a[0] , \d[12] );
nand \mul_16_12_g20519/U$1 ( \1647 , \1646 , \d[11] );
nand \mul_16_12_g20638/U$1 ( \1648 , \a[0] , \d[12] );
and \mul_16_12_g20680/U$1 ( \1649 , \1647 , \1648 , \d[13] );
xor \mul_16_12_g20540/U$1 ( \1650 , \a[12] , \d[1] );
not \mul_16_12_g20402/U$3 ( \1651 , \1650 );
not \mul_16_12_g20402/U$4 ( \1652 , \932 );
or \mul_16_12_g20402/U$2 ( \1653 , \1651 , \1652 );
nand \mul_16_12_g20482/U$1 ( \1654 , \1572 , \d[0] );
nand \mul_16_12_g20402/U$1 ( \1655 , \1653 , \1654 );
and \mul_16_12_g20275/U$2 ( \1656 , \1649 , \1655 );
and \mul_16_12_g20154/U$3 ( \1657 , \1645 , \1656 );
and \mul_16_12_g20154/U$5 ( \1658 , \1632 , \1644 );
or \mul_16_12_g20154/U$2 ( \1659 , \1657 , \1658 );
not \mul_16_12_g20404/U$3 ( \1660 , \1576 );
not \mul_16_12_g20404/U$4 ( \1661 , \932 );
or \mul_16_12_g20404/U$2 ( \1662 , \1660 , \1661 );
xor \mul_16_12_g20541/U$1 ( \1663 , \a[15] , \d[1] );
nand \mul_16_12_g20488/U$1 ( \1664 , \1663 , \d[0] );
nand \mul_16_12_g20404/U$1 ( \1665 , \1662 , \1664 );
or \mul_16_12_g20518/U$2 ( \1666 , \a[0] , \d[14] );
nand \mul_16_12_g20518/U$1 ( \1667 , \1666 , \d[13] );
nand \mul_16_12_g20644/U$1 ( \1668 , \a[0] , \d[14] );
nand \mul_16_12_g20512/U$1 ( \1669 , \1667 , \1668 , \d[15] );
xor \g36004/U$1 ( \1670 , \1665 , \1669 );
not \mul_16_12_g20315/U$3 ( \1671 , \1642 );
not \mul_16_12_g20315/U$4 ( \1672 , \1638 );
or \mul_16_12_g20315/U$2 ( \1673 , \1671 , \1672 );
xor \mul_16_12_g20620/U$1 ( \1674 , \a[5] , \d[11] );
nand \mul_16_12_g20447/U$1 ( \1675 , \1641 , \1674 );
nand \mul_16_12_g20315/U$1 ( \1676 , \1673 , \1675 );
xnor \g36004/U$1_r1 ( \1677 , \1670 , \1676 );
xor \mul_16_12_g20702/U$1 ( \1678 , \1659 , \1677 );
xor \mul_16_12_g20590/U$1 ( \1679 , \a[7] , \d[7] );
not \mul_16_12_g20330/U$3 ( \1680 , \1679 );
not \mul_16_12_g20330/U$4 ( \1681 , \1127 );
or \mul_16_12_g20330/U$2 ( \1682 , \1680 , \1681 );
nand \mul_16_12_g20453/U$1 ( \1683 , \958 , \1535 );
nand \mul_16_12_g20330/U$1 ( \1684 , \1682 , \1683 );
xor \mul_16_12_g20612/U$1 ( \1685 , \a[5] , \d[9] );
not \mul_16_12_g20319/U$3 ( \1686 , \1685 );
not \mul_16_12_g20319/U$4 ( \1687 , \1542 );
or \mul_16_12_g20319/U$2 ( \1688 , \1686 , \1687 );
nand \mul_16_12_g20455/U$1 ( \1689 , \1545 , \1538 );
nand \mul_16_12_g20319/U$1 ( \1690 , \1688 , \1689 );
xor \mul_16_12_g20217/U$4 ( \1691 , \1684 , \1690 );
xor \mul_16_12_g20578/U$1 ( \1692 , \a[9] , \d[5] );
not \mul_16_12_g20363/U$3 ( \1693 , \1692 );
not \mul_16_12_g20363/U$4 ( \1694 , \1135 );
or \mul_16_12_g20363/U$2 ( \1695 , \1693 , \1694 );
nand \mul_16_12_g20451/U$1 ( \1696 , \951 , \1603 );
nand \mul_16_12_g20363/U$1 ( \1697 , \1695 , \1696 );
and \mul_16_12_g20217/U$3 ( \1698 , \1691 , \1697 );
and \mul_16_12_g20217/U$5 ( \1699 , \1684 , \1690 );
or \mul_16_12_g20217/U$2 ( \1700 , \1698 , \1699 );
not \mul_16_12_g20216/U$1 ( \1701 , \1700 );
and \mul_16_12_g20082/U$2 ( \1702 , \1678 , \1701 );
not \mul_16_12_g20082/U$4 ( \1703 , \1678 );
and \mul_16_12_g20082/U$3 ( \1704 , \1703 , \1700 );
nor \mul_16_12_g20082/U$1 ( \1705 , \1702 , \1704 );
not \mul_16_12_g20056/U$4 ( \1706 , \1705 );
or \mul_16_12_g20056/U$2 ( \1707 , \1626 , \1706 );
or \mul_16_12_g20056/U$5 ( \1708 , \1705 , \1625 );
nand \mul_16_12_g20056/U$1 ( \1709 , \1707 , \1708 );
xor \mul_16_12_g20215/U$1 ( \1710 , \1571 , \1578 );
xor \mul_16_12_g20215/U$1_r1 ( \1711 , \1710 , \1586 );
xor \mul_16_12_g20599/U$1 ( \1712 , \a[0] , \d[13] );
not \mul_16_12_g20306/U$3 ( \1713 , \1712 );
nor \mul_16_12_g20515/U$1 ( \1714 , \1552 , \1553 );
not \mul_16_12_g20306/U$4 ( \1715 , \1714 );
or \mul_16_12_g20306/U$2 ( \1716 , \1713 , \1715 );
nand \mul_16_12_g20471/U$1 ( \1717 , \1552 , \1627 );
nand \mul_16_12_g20306/U$1 ( \1718 , \1716 , \1717 );
xor \mul_16_12_g20626/U$1 ( \1719 , \a[2] , \d[11] );
not \mul_16_12_g20316/U$3 ( \1720 , \1719 );
nor \mul_16_12_g20513/U$1 ( \1721 , \1637 , \1635 );
not \mul_16_12_g20316/U$4 ( \1722 , \1721 );
or \mul_16_12_g20316/U$2 ( \1723 , \1720 , \1722 );
nand \mul_16_12_g20475/U$1 ( \1724 , \1641 , \1633 );
nand \mul_16_12_g20316/U$1 ( \1725 , \1723 , \1724 );
xor \mul_16_12_g20225/U$4 ( \1726 , \1718 , \1725 );
xor \mul_16_12_g20577/U$1 ( \1727 , \a[8] , \d[5] );
not \mul_16_12_g20362/U$3 ( \1728 , \1727 );
not \mul_16_12_g20362/U$4 ( \1729 , \1135 );
or \mul_16_12_g20362/U$2 ( \1730 , \1728 , \1729 );
nand \mul_16_12_g20421/U$1 ( \1731 , \951 , \1692 );
nand \mul_16_12_g20362/U$1 ( \1732 , \1730 , \1731 );
and \mul_16_12_g20225/U$3 ( \1733 , \1726 , \1732 );
and \mul_16_12_g20225/U$5 ( \1734 , \1718 , \1725 );
or \mul_16_12_g20225/U$2 ( \1735 , \1733 , \1734 );
or \mul_16_12_g20143/U$2 ( \1736 , \1711 , \1735 );
xor \mul_16_12_g20611/U$1 ( \1737 , \a[4] , \d[9] );
not \mul_16_12_g20323/U$3 ( \1738 , \1737 );
not \mul_16_12_g20323/U$4 ( \1739 , \1542 );
or \mul_16_12_g20323/U$2 ( \1740 , \1738 , \1739 );
nand \mul_16_12_g20466/U$1 ( \1741 , \1545 , \1685 );
nand \mul_16_12_g20323/U$1 ( \1742 , \1740 , \1741 );
not \mul_16_12_g20208/U$3 ( \1743 , \1742 );
xor \mul_16_12_g20551/U$1 ( \1744 , \a[10] , \d[3] );
not \mul_16_12_g20377/U$3 ( \1745 , \1744 );
not \mul_16_12_g20377/U$4 ( \1746 , \1067 );
or \mul_16_12_g20377/U$2 ( \1747 , \1745 , \1746 );
nand \mul_16_12_g20473/U$1 ( \1748 , \976 , \1580 );
nand \mul_16_12_g20377/U$1 ( \1749 , \1747 , \1748 );
not \mul_16_12_g20208/U$4 ( \1750 , \1749 );
or \mul_16_12_g20208/U$2 ( \1751 , \1743 , \1750 );
or \mul_16_12_g20237/U$2 ( \1752 , \1749 , \1742 );
not \mul_16_12_g20333/U$3 ( \1753 , \1679 );
not \mul_16_12_g20333/U$4 ( \1754 , \958 );
or \mul_16_12_g20333/U$2 ( \1755 , \1753 , \1754 );
xor \mul_16_12_g20589/U$1 ( \1756 , \a[6] , \d[7] );
nand \mul_16_12_g20383/U$1 ( \1757 , \1127 , \1756 );
nand \mul_16_12_g20333/U$1 ( \1758 , \1755 , \1757 );
nand \mul_16_12_g20237/U$1 ( \1759 , \1752 , \1758 );
nand \mul_16_12_g20208/U$1 ( \1760 , \1751 , \1759 );
nand \mul_16_12_g20143/U$1 ( \1761 , \1736 , \1760 );
nand \mul_16_12_g20183/U$1 ( \1762 , \1711 , \1735 );
nand \mul_16_12_g20122/U$1 ( \1763 , \1761 , \1762 );
not \mul_16_12_g20107/U$1 ( \1764 , \1763 );
and \mul_16_12_g20040/U$2 ( \1765 , \1709 , \1764 );
not \mul_16_12_g20040/U$4 ( \1766 , \1709 );
and \mul_16_12_g20040/U$3 ( \1767 , \1766 , \1763 );
nor \mul_16_12_g20040/U$1 ( \1768 , \1765 , \1767 );
xor \mul_16_12_g20217/U$1 ( \1769 , \1684 , \1690 );
xor \mul_16_12_g20217/U$1_r1 ( \1770 , \1769 , \1697 );
xor \mul_16_12_g20154/U$1 ( \1771 , \1632 , \1644 );
xor \mul_16_12_g20154/U$1_r1 ( \1772 , \1771 , \1656 );
xor \mul_16_12_g20053/U$4 ( \1773 , \1770 , \1772 );
and \mul_16_12_g20480/U$1 ( \1774 , \1552 , \a[0] );
xor \g35457/U$1 ( \1775 , \d[7] , \a[5] );
not \mul_16_12_g20337/U$3 ( \1776 , \1775 );
not \mul_16_12_g20337/U$4 ( \1777 , \1127 );
or \mul_16_12_g20337/U$2 ( \1778 , \1776 , \1777 );
nand \mul_16_12_g20474/U$1 ( \1779 , \958 , \1756 );
nand \mul_16_12_g20337/U$1 ( \1780 , \1778 , \1779 );
xor \mul_16_12_g20193/U$4 ( \1781 , \1774 , \1780 );
xor \mul_16_12_g20575/U$1 ( \1782 , \a[9] , \d[3] );
not \mul_16_12_g20369/U$3 ( \1783 , \1782 );
not \mul_16_12_g20369/U$4 ( \1784 , \973 );
or \mul_16_12_g20369/U$2 ( \1785 , \1783 , \1784 );
nand \mul_16_12_g20454/U$1 ( \1786 , \976 , \1744 );
nand \mul_16_12_g20369/U$1 ( \1787 , \1785 , \1786 );
and \mul_16_12_g20193/U$3 ( \1788 , \1781 , \1787 );
and \mul_16_12_g20193/U$5 ( \1789 , \1774 , \1780 );
or \mul_16_12_g20193/U$2 ( \1790 , \1788 , \1789 );
xor \mul_16_12_g20275/U$1 ( \1791 , \1649 , \1655 );
or \mul_16_12_g20120/U$2 ( \1792 , \1790 , \1791 );
xor \mul_16_12_g35961/U$1 ( \1793 , \a[11] , \d[1] );
not \mul_16_12_g20405/U$3 ( \1794 , \1793 );
not \mul_16_12_g20405/U$4 ( \1795 , \932 );
or \mul_16_12_g20405/U$2 ( \1796 , \1794 , \1795 );
nand \mul_16_12_g20481/U$1 ( \1797 , \1650 , \d[0] );
nand \mul_16_12_g20405/U$1 ( \1798 , \1796 , \1797 );
xor \mul_16_12_g20622/U$1 ( \1799 , \a[3] , \d[9] );
not \mul_16_12_g20320/U$3 ( \1800 , \1799 );
not \mul_16_12_g20320/U$4 ( \1801 , \1542 );
or \mul_16_12_g20320/U$2 ( \1802 , \1800 , \1801 );
nand \mul_16_12_g20467/U$1 ( \1803 , \1545 , \1737 );
nand \mul_16_12_g20320/U$1 ( \1804 , \1802 , \1803 );
xor \mul_16_12_g20189/U$4 ( \1805 , \1798 , \1804 );
xor \mul_16_12_g20632/U$1 ( \1806 , \a[1] , \d[11] );
not \mul_16_12_g20313/U$3 ( \1807 , \1806 );
not \mul_16_12_g20313/U$4 ( \1808 , \1721 );
or \mul_16_12_g20313/U$2 ( \1809 , \1807 , \1808 );
nand \mul_16_12_g20470/U$1 ( \1810 , \1641 , \1719 );
nand \mul_16_12_g20313/U$1 ( \1811 , \1809 , \1810 );
and \mul_16_12_g20189/U$3 ( \1812 , \1805 , \1811 );
and \mul_16_12_g20189/U$5 ( \1813 , \1798 , \1804 );
or \mul_16_12_g20189/U$2 ( \1814 , \1812 , \1813 );
nand \mul_16_12_g20120/U$1 ( \1815 , \1792 , \1814 );
nand \mul_16_12_g20162/U$1 ( \1816 , \1790 , \1791 );
nand \mul_16_12_g20100/U$1 ( \1817 , \1815 , \1816 );
and \mul_16_12_g20053/U$3 ( \1818 , \1773 , \1817 );
and \mul_16_12_g20053/U$5 ( \1819 , \1770 , \1772 );
or \mul_16_12_g20053/U$2 ( \1820 , \1818 , \1819 );
not \mul_16_12_g20052/U$1 ( \1821 , \1820 );
and \mul_16_12_g20021/U$2 ( \1822 , \1768 , \1821 );
not \mul_16_12_g20021/U$4 ( \1823 , \1768 );
and \mul_16_12_g20021/U$3 ( \1824 , \1823 , \1820 );
nor \mul_16_12_g20021/U$1 ( \1825 , \1822 , \1824 );
xor \g35449/U$1 ( \1826 , \1735 , \1711 );
xnor \g35449/U$1_r1 ( \1827 , \1826 , \1760 );
not \mul_16_12_g35738/U$1 ( \1828 , \1827 );
not \mul_16_12_g19987/U$3 ( \1829 , \1828 );
xor \mul_16_12_g20053/U$1 ( \1830 , \1770 , \1772 );
xor \mul_16_12_g20053/U$1_r1 ( \1831 , \1830 , \1817 );
not \mul_16_12_g19987/U$4 ( \1832 , \1831 );
or \mul_16_12_g19987/U$2 ( \1833 , \1829 , \1832 );
or \mul_16_12_g20000/U$2 ( \1834 , \1831 , \1828 );
xor \mul_16_12_g20225/U$1 ( \1835 , \1718 , \1725 );
xor \mul_16_12_g20225/U$1_r1 ( \1836 , \1835 , \1732 );
not \mul_16_12_g20699/U$2 ( \1837 , \1836 );
xor \mul_16_12_g20710/U$1 ( \1838 , \1742 , \1758 );
xnor \mul_16_12_g20710/U$1_r1 ( \1839 , \1838 , \1749 );
nand \mul_16_12_g20699/U$1 ( \1840 , \1837 , \1839 );
not \mul_16_12_g20102/U$3 ( \1841 , \1840 );
xor \mul_16_12_g20588/U$1 ( \1842 , \a[7] , \d[5] );
not \mul_16_12_g20349/U$3 ( \1843 , \1842 );
not \mul_16_12_g20349/U$4 ( \1844 , \1135 );
or \mul_16_12_g20349/U$2 ( \1845 , \1843 , \1844 );
nand \mul_16_12_g20417/U$1 ( \1846 , \951 , \1727 );
nand \mul_16_12_g20349/U$1 ( \1847 , \1845 , \1846 );
not \mul_16_12_g20348/U$1 ( \1848 , \1847 );
not \mul_16_12_g20169/U$3 ( \1849 , \1848 );
xor \mul_16_12_g20576/U$1 ( \1850 , \a[8] , \d[3] );
not \mul_16_12_g20372/U$3 ( \1851 , \1850 );
not \mul_16_12_g20372/U$4 ( \1852 , \973 );
or \mul_16_12_g20372/U$2 ( \1853 , \1851 , \1852 );
nand \mul_16_12_g20437/U$1 ( \1854 , \976 , \1782 );
nand \mul_16_12_g20372/U$1 ( \1855 , \1853 , \1854 );
or \mul_16_12_g20520/U$2 ( \1856 , \a[0] , \d[10] );
nand \mul_16_12_g20520/U$1 ( \1857 , \1856 , \d[9] );
nand \mul_16_12_g20642/U$1 ( \1858 , \a[0] , \d[10] );
nand \mul_16_12_g20508/U$1 ( \1859 , \1857 , \1858 , \d[11] );
not \mul_16_12_g20507/U$1 ( \1860 , \1859 );
nand \mul_16_12_g20283/U$1 ( \1861 , \1855 , \1860 );
not \mul_16_12_g20169/U$4 ( \1862 , \1861 );
or \mul_16_12_g20169/U$2 ( \1863 , \1849 , \1862 );
xor \mul_16_12_g35962/U$1 ( \1864 , \a[10] , \d[1] );
not \mul_16_12_g20392/U$3 ( \1865 , \1864 );
not \mul_16_12_g20392/U$4 ( \1866 , \932 );
or \mul_16_12_g20392/U$2 ( \1867 , \1865 , \1866 );
nand \mul_16_12_g20445/U$1 ( \1868 , \1793 , \d[0] );
nand \mul_16_12_g20392/U$1 ( \1869 , \1867 , \1868 );
not \mul_16_12_g20252/U$3 ( \1870 , \1869 );
xor \g35459/U$1 ( \1871 , \d[9] , \a[2] );
not \mul_16_12_g20318/U$3 ( \1872 , \1871 );
not \mul_16_12_g20318/U$4 ( \1873 , \1542 );
or \mul_16_12_g20318/U$2 ( \1874 , \1872 , \1873 );
nand \mul_16_12_g20450/U$1 ( \1875 , \1545 , \1799 );
nand \mul_16_12_g20318/U$1 ( \1876 , \1874 , \1875 );
not \mul_16_12_g20252/U$4 ( \1877 , \1876 );
or \mul_16_12_g20252/U$2 ( \1878 , \1870 , \1877 );
or \mul_16_12_g20262/U$2 ( \1879 , \1876 , \1869 );
xor \g35458/U$1 ( \1880 , \d[7] , \a[4] );
not \mul_16_12_g20340/U$3 ( \1881 , \1880 );
xnor \g35768/U$1 ( \1882 , \d[7] , \d[6] );
nor \g35767/U$1 ( \1883 , \1882 , \957 );
not \mul_16_12_g20340/U$4 ( \1884 , \1883 );
or \mul_16_12_g20340/U$2 ( \1885 , \1881 , \1884 );
nand \mul_16_12_g20456/U$1 ( \1886 , \1775 , \957 );
nand \mul_16_12_g20340/U$1 ( \1887 , \1885 , \1886 );
nand \mul_16_12_g20262/U$1 ( \1888 , \1879 , \1887 );
nand \mul_16_12_g20252/U$1 ( \1889 , \1878 , \1888 );
nand \mul_16_12_g20169/U$1 ( \1890 , \1863 , \1889 );
not \mul_16_12_g20703/U$2 ( \1891 , \1861 );
nand \mul_16_12_g20703/U$1 ( \1892 , \1891 , \1847 );
nand \mul_16_12_g20149/U$1 ( \1893 , \1890 , \1892 );
not \mul_16_12_g20102/U$4 ( \1894 , \1893 );
or \mul_16_12_g20102/U$2 ( \1895 , \1841 , \1894 );
not \mul_16_12_g20697/U$2 ( \1896 , \1839 );
nand \mul_16_12_g20697/U$1 ( \1897 , \1896 , \1836 );
nand \mul_16_12_g20102/U$1 ( \1898 , \1895 , \1897 );
nand \mul_16_12_g20000/U$1 ( \1899 , \1834 , \1898 );
nand \mul_16_12_g19987/U$1 ( \1900 , \1833 , \1899 );
xnor \mul_16_12_g20686/U$1 ( \1901 , \1825 , \1900 );
not \mul_16_12_g19965/U$3 ( \1902 , \1901 );
xnor \g35737/U$1 ( \1903 , \1831 , \1827 );
not \fopt35586/U$1 ( \1904 , \1898 );
and \mul_16_12_g19990/U$2 ( \1905 , \1903 , \1904 );
not \mul_16_12_g19990/U$4 ( \1906 , \1903 );
and \mul_16_12_g19990/U$3 ( \1907 , \1906 , \1898 );
nor \mul_16_12_g19990/U$1 ( \1908 , \1905 , \1907 );
xor \mul_16_12_g20104/U$1 ( \1909 , \1791 , \1790 );
xnor \mul_16_12_g20104/U$1_r1 ( \1910 , \1909 , \1814 );
not \mul_16_12_g20088/U$1 ( \1911 , \1910 );
not \mul_16_12_g20063/U$2 ( \1912 , \1911 );
xor \g35904/U$1 ( \1913 , \1836 , \1839 );
xor \g35904/U$1_r1 ( \1914 , \1913 , \1893 );
nand \mul_16_12_g20063/U$1 ( \1915 , \1912 , \1914 );
xor \mul_16_12_g20193/U$1 ( \1916 , \1774 , \1780 );
xor \mul_16_12_g20193/U$1_r1 ( \1917 , \1916 , \1787 );
not \mul_16_12_g20696/U$2 ( \1918 , \1917 );
xor \mul_16_12_g20189/U$1 ( \1919 , \1798 , \1804 );
xor \mul_16_12_g20189/U$1_r1 ( \1920 , \1919 , \1811 );
not \mul_16_12_g20188/U$1 ( \1921 , \1920 );
nand \mul_16_12_g20696/U$1 ( \1922 , \1918 , \1921 );
not \g35733/U$3 ( \1923 , \1922 );
xor \mul_16_12_g20618/U$1 ( \1924 , \a[0] , \d[11] );
not \mul_16_12_g20311/U$3 ( \1925 , \1924 );
not \mul_16_12_g20311/U$4 ( \1926 , \1638 );
or \mul_16_12_g20311/U$2 ( \1927 , \1925 , \1926 );
nand \mul_16_12_g20414/U$1 ( \1928 , \1641 , \1806 );
nand \mul_16_12_g20311/U$1 ( \1929 , \1927 , \1928 );
not \mul_16_12_g20206/U$3 ( \1930 , \1929 );
xor \mul_16_12_g35963/U$1 ( \1931 , \a[6] , \d[5] );
not \mul_16_12_g20341/U$3 ( \1932 , \1931 );
not \mul_16_12_g20341/U$4 ( \1933 , \1135 );
or \mul_16_12_g20341/U$2 ( \1934 , \1932 , \1933 );
nand \mul_16_12_g20412/U$1 ( \1935 , \951 , \1842 );
nand \mul_16_12_g20341/U$1 ( \1936 , \1934 , \1935 );
not \mul_16_12_g20206/U$4 ( \1937 , \1936 );
or \mul_16_12_g20206/U$2 ( \1938 , \1930 , \1937 );
or \g35907/U$2 ( \1939 , \1936 , \1929 );
and \mul_16_12_g20715/U$2 ( \1940 , \1855 , \1860 );
not \mul_16_12_g20715/U$4 ( \1941 , \1855 );
and \mul_16_12_g20715/U$3 ( \1942 , \1941 , \1859 );
nor \mul_16_12_g20715/U$1 ( \1943 , \1940 , \1942 );
nand \g35907/U$1 ( \1944 , \1939 , \1943 );
nand \mul_16_12_g20206/U$1 ( \1945 , \1938 , \1944 );
not \g35733/U$4 ( \1946 , \1945 );
or \g35733/U$2 ( \1947 , \1923 , \1946 );
not \g35734/U$2 ( \1948 , \1921 );
nand \g35734/U$1 ( \1949 , \1948 , \1917 );
nand \g35733/U$1 ( \1950 , \1947 , \1949 );
and \mul_16_12_g20049/U$2 ( \1951 , \1915 , \1950 );
nor \mul_16_12_g20069/U$1 ( \1952 , \1914 , \1910 );
nor \mul_16_12_g20049/U$1 ( \1953 , \1951 , \1952 );
nand \mul_16_12_g19977/U$1 ( \1954 , \1908 , \1953 );
not \mul_16_12_g19971/U$2 ( \1955 , \1954 );
not \mul_16_12_g20060/U$3 ( \1956 , \1911 );
not \mul_16_12_g20091/U$1 ( \1957 , \1950 );
not \mul_16_12_g20060/U$4 ( \1958 , \1957 );
or \mul_16_12_g20060/U$2 ( \1959 , \1956 , \1958 );
nand \mul_16_12_g20068/U$1 ( \1960 , \1950 , \1910 );
nand \mul_16_12_g20060/U$1 ( \1961 , \1959 , \1960 );
xor \g35786/U$1 ( \1962 , \1914 , \1961 );
xor \mul_16_12_g20150/U$1 ( \1963 , \1848 , \1861 );
xnor \mul_16_12_g20150/U$1_r1 ( \1964 , \1963 , \1889 );
xor \mul_16_12_g20573/U$1 ( \1965 , \a[9] , \d[1] );
not \mul_16_12_g20394/U$3 ( \1966 , \1965 );
not \mul_16_12_g20394/U$4 ( \1967 , \932 );
or \mul_16_12_g20394/U$2 ( \1968 , \1966 , \1967 );
nand \mul_16_12_g20464/U$1 ( \1969 , \1864 , \d[0] );
nand \mul_16_12_g20394/U$1 ( \1970 , \1968 , \1969 );
xor \mul_16_12_g20629/U$1 ( \1971 , \a[1] , \d[9] );
not \mul_16_12_g20321/U$3 ( \1972 , \1971 );
not \mul_16_12_g20321/U$4 ( \1973 , \1542 );
or \mul_16_12_g20321/U$2 ( \1974 , \1972 , \1973 );
nand \mul_16_12_g20411/U$1 ( \1975 , \1541 , \1871 );
nand \mul_16_12_g20321/U$1 ( \1976 , \1974 , \1975 );
or \mul_16_12_g20238/U$2 ( \1977 , \1970 , \1976 );
xor \mul_16_12_g20598/U$1 ( \1978 , \a[5] , \d[5] );
not \mul_16_12_g20344/U$3 ( \1979 , \1978 );
not \mul_16_12_g20344/U$4 ( \1980 , \948 );
or \mul_16_12_g20344/U$2 ( \1981 , \1979 , \1980 );
nand \mul_16_12_g35964/U$1 ( \1982 , \951 , \1931 );
nand \mul_16_12_g20344/U$1 ( \1983 , \1981 , \1982 );
nand \mul_16_12_g20238/U$1 ( \1984 , \1977 , \1983 );
nand \mul_16_12_g20285/U$1 ( \1985 , \1976 , \1970 );
nand \mul_16_12_g20207/U$1 ( \1986 , \1984 , \1985 );
not \mul_16_12_g20200/U$1 ( \1987 , \1986 );
not \mul_16_12_g20121/U$3 ( \1988 , \1987 );
not \mul_16_12_g20266/U$3 ( \1989 , \1887 );
not \mul_16_12_g20391/U$1 ( \1990 , \1869 );
not \mul_16_12_g20266/U$4 ( \1991 , \1990 );
or \mul_16_12_g20266/U$2 ( \1992 , \1989 , \1991 );
not \mul_16_12_g20280/U$2 ( \1993 , \1887 );
nand \mul_16_12_g20280/U$1 ( \1994 , \1993 , \1869 );
nand \mul_16_12_g20266/U$1 ( \1995 , \1992 , \1994 );
not \mul_16_12_g20317/U$1 ( \1996 , \1876 );
and \mul_16_12_g20246/U$2 ( \1997 , \1995 , \1996 );
not \mul_16_12_g20246/U$4 ( \1998 , \1995 );
and \mul_16_12_g20246/U$3 ( \1999 , \1998 , \1876 );
nor \mul_16_12_g20246/U$1 ( \2000 , \1997 , \1999 );
not \mul_16_12_g20121/U$4 ( \2001 , \2000 );
or \mul_16_12_g20121/U$2 ( \2002 , \1988 , \2001 );
xor \g35456/U$1 ( \2003 , \d[3] , \a[7] );
not \mul_16_12_g20378/U$3 ( \2004 , \2003 );
not \mul_16_12_g20378/U$4 ( \2005 , \973 );
or \mul_16_12_g20378/U$2 ( \2006 , \2004 , \2005 );
nand \mul_16_12_g20472/U$1 ( \2007 , \976 , \1850 );
nand \mul_16_12_g20378/U$1 ( \2008 , \2006 , \2007 );
and \mul_16_12_g20677/U$1 ( \2009 , \1641 , \a[0] );
or \mul_16_12_g20718/U$1 ( \2010 , \2008 , \2009 );
xor \mul_16_12_g20617/U$1 ( \2011 , \a[3] , \d[7] );
not \mul_16_12_g20336/U$3 ( \2012 , \2011 );
not \mul_16_12_g20336/U$4 ( \2013 , \1127 );
or \mul_16_12_g20336/U$2 ( \2014 , \2012 , \2013 );
nand \mul_16_12_g20415/U$1 ( \2015 , \958 , \1880 );
nand \mul_16_12_g20336/U$1 ( \2016 , \2014 , \2015 );
and \mul_16_12_g20205/U$2 ( \2017 , \2010 , \2016 );
and \mul_16_12_g20674/U$1 ( \2018 , \2008 , \2009 );
nor \mul_16_12_g20205/U$1 ( \2019 , \2017 , \2018 );
not \mul_16_12_g20203/U$1 ( \2020 , \2019 );
nand \mul_16_12_g20121/U$1 ( \2021 , \2002 , \2020 );
not \mul_16_12_g20700/U$2 ( \2022 , \2000 );
nand \mul_16_12_g20700/U$1 ( \2023 , \2022 , \1986 );
and \mul_16_12_g2/U$1 ( \2024 , \2021 , \2023 );
xor \mul_16_12_g20031/U$4 ( \2025 , \1964 , \2024 );
xor \mul_16_12_g20114/U$1 ( \2026 , \1917 , \1920 );
xnor \mul_16_12_g20114/U$1_r1 ( \2027 , \2026 , \1945 );
and \mul_16_12_g20031/U$3 ( \2028 , \2025 , \2027 );
and \mul_16_12_g20031/U$5 ( \2029 , \1964 , \2024 );
or \mul_16_12_g20031/U$2 ( \2030 , \2028 , \2029 );
nand \mul_16_12_g20014/U$1 ( \2031 , \1962 , \2030 );
or \mul_16_12_g20521/U$2 ( \2032 , \a[0] , \d[8] );
nand \mul_16_12_g20521/U$1 ( \2033 , \2032 , \d[7] );
nand \mul_16_12_g20646/U$1 ( \2034 , \a[0] , \d[8] );
and \mul_16_12_g20679/U$1 ( \2035 , \2033 , \2034 , \d[9] );
xor \mul_16_12_g20586/U$1 ( \2036 , \a[6] , \d[3] );
not \mul_16_12_g20379/U$3 ( \2037 , \2036 );
not \mul_16_12_g20379/U$4 ( \2038 , \973 );
or \mul_16_12_g20379/U$2 ( \2039 , \2037 , \2038 );
nand \mul_16_12_g20435/U$1 ( \2040 , \976 , \2003 );
nand \mul_16_12_g20379/U$1 ( \2041 , \2039 , \2040 );
and \mul_16_12_g20260/U$2 ( \2042 , \2035 , \2041 );
xor \mul_16_12_g20574/U$1 ( \2043 , \a[8] , \d[1] );
not \mul_16_12_g20401/U$3 ( \2044 , \2043 );
not \mul_16_12_g20401/U$4 ( \2045 , \932 );
or \mul_16_12_g20401/U$2 ( \2046 , \2044 , \2045 );
nand \mul_16_12_g20479/U$1 ( \2047 , \1965 , \d[0] );
nand \mul_16_12_g20401/U$1 ( \2048 , \2046 , \2047 );
xor \mul_16_12_g20625/U$1 ( \2049 , \a[0] , \d[9] );
not \mul_16_12_g20324/U$3 ( \2050 , \2049 );
not \mul_16_12_g20324/U$4 ( \2051 , \1542 );
or \mul_16_12_g20324/U$2 ( \2052 , \2050 , \2051 );
nand \mul_16_12_g20419/U$1 ( \2053 , \1545 , \1971 );
nand \mul_16_12_g20324/U$1 ( \2054 , \2052 , \2053 );
or \mul_16_12_g20261/U$2 ( \2055 , \2048 , \2054 );
xor \mul_16_12_g20616/U$1 ( \2056 , \a[2] , \d[7] );
not \mul_16_12_g20328/U$3 ( \2057 , \2056 );
not \mul_16_12_g20328/U$4 ( \2058 , \1883 );
or \mul_16_12_g20328/U$2 ( \2059 , \2057 , \2058 );
nand \mul_16_12_g20420/U$1 ( \2060 , \958 , \2011 );
nand \mul_16_12_g20328/U$1 ( \2061 , \2059 , \2060 );
nand \mul_16_12_g20261/U$1 ( \2062 , \2055 , \2061 );
nand \mul_16_12_g20281/U$1 ( \2063 , \2048 , \2054 );
nand \mul_16_12_g20253/U$1 ( \2064 , \2062 , \2063 );
xor \mul_16_12_g20128/U$1 ( \2065 , \2042 , \2064 );
xor \mul_16_12_g35968/U$1 ( \2066 , \2009 , \2016 );
xor \mul_16_12_g35968/U$1_r1 ( \2067 , \2066 , \2008 );
xor \mul_16_12_g20128/U$1_r1 ( \2068 , \2065 , \2067 );
xor \mul_16_12_g20265/U$1 ( \2069 , \1976 , \1970 );
xor \mul_16_12_g20712/U$1 ( \2070 , \2069 , \1983 );
or \mul_16_12_g20692/U$2 ( \2071 , \2068 , \2070 );
xor \mul_16_12_g20597/U$1 ( \2072 , \a[4] , \d[5] );
not \mul_16_12_g20345/U$3 ( \2073 , \2072 );
not \mul_16_12_g20345/U$4 ( \2074 , \1135 );
or \mul_16_12_g20345/U$2 ( \2075 , \2073 , \2074 );
nand \mul_16_12_g20413/U$1 ( \2076 , \951 , \1978 );
nand \mul_16_12_g20345/U$1 ( \2077 , \2075 , \2076 );
and \mul_16_12_g20678/U$1 ( \2078 , \1541 , \a[0] );
not \mul_16_12_g20326/U$3 ( \2079 , \1131 );
not \mul_16_12_g20326/U$4 ( \2080 , \1127 );
or \mul_16_12_g20326/U$2 ( \2081 , \2079 , \2080 );
nand \mul_16_12_g20418/U$1 ( \2082 , \958 , \2056 );
nand \mul_16_12_g20326/U$1 ( \2083 , \2081 , \2082 );
xor \mul_16_12_g20211/U$4 ( \2084 , \2078 , \2083 );
not \mul_16_12_g20385/U$3 ( \2085 , \1106 );
not \mul_16_12_g20385/U$4 ( \2086 , \932 );
or \mul_16_12_g20385/U$2 ( \2087 , \2085 , \2086 );
nand \mul_16_12_g20416/U$1 ( \2088 , \2043 , \d[0] );
nand \mul_16_12_g20385/U$1 ( \2089 , \2087 , \2088 );
and \mul_16_12_g20211/U$3 ( \2090 , \2084 , \2089 );
and \mul_16_12_g20211/U$5 ( \2091 , \2078 , \2083 );
or \mul_16_12_g20211/U$2 ( \2092 , \2090 , \2091 );
xor \mul_16_12_g20130/U$4 ( \2093 , \2077 , \2092 );
xor \mul_16_12_g20260/U$1 ( \2094 , \2035 , \2041 );
and \mul_16_12_g20130/U$3 ( \2095 , \2093 , \2094 );
and \mul_16_12_g20130/U$5 ( \2096 , \2077 , \2092 );
or \mul_16_12_g20130/U$2 ( \2097 , \2095 , \2096 );
nand \mul_16_12_g20692/U$1 ( \2098 , \2071 , \2097 );
nand \mul_16_12_g20095/U$1 ( \2099 , \2068 , \2070 );
nand \mul_16_12_g20073/U$1 ( \2100 , \2098 , \2099 );
not \mul_16_12_g20005/U$2 ( \2101 , \2100 );
xor \g35976/U$1 ( \2102 , \1929 , \1936 );
xor \g35976/U$1_r1 ( \2103 , \2102 , \1943 );
xor \mul_16_12_g20112/U$1 ( \2104 , \1986 , \2000 );
xnor \mul_16_12_g20112/U$1_r1 ( \2105 , \2104 , \2019 );
xor \mul_16_12_g35758/U$1 ( \2106 , \2103 , \2105 );
xor \mul_16_12_g20128/U$4 ( \2107 , \2042 , \2064 );
and \mul_16_12_g20128/U$3 ( \2108 , \2107 , \2067 );
and \mul_16_12_g20128/U$5 ( \2109 , \2042 , \2064 );
or \mul_16_12_g20128/U$2 ( \2110 , \2108 , \2109 );
xor \mul_16_12_g35758/U$1_r1 ( \2111 , \2106 , \2110 );
nand \mul_16_12_g20005/U$1 ( \2112 , \2101 , \2111 );
nand \mul_16_12_g19996/U$1 ( \2113 , \2031 , \2112 );
nor \mul_16_12_g19971/U$1 ( \2114 , \1955 , \2113 );
not \mul_16_12_g19966/U$3 ( \2115 , \2114 );
or \mul_16_12_g20690/U$1 ( \2116 , \1149 , \1156 );
not \mul_16_12_g20673/U$3 ( \2117 , \2116 );
not \mul_16_12_g20673/U$4 ( \2118 , \1101 );
or \mul_16_12_g20673/U$2 ( \2119 , \2117 , \2118 );
nand \mul_16_12_g20673/U$1 ( \2120 , \2119 , \1158 );
not \g35901/U$3 ( \2121 , \2120 );
not \mul_16_12_g20352/U$3 ( \2122 , \1138 );
not \mul_16_12_g20352/U$4 ( \2123 , \948 );
or \mul_16_12_g20352/U$2 ( \2124 , \2122 , \2123 );
nand \mul_16_12_g20423/U$1 ( \2125 , \951 , \2072 );
nand \mul_16_12_g20352/U$1 ( \2126 , \2124 , \2125 );
not \mul_16_12_g20175/U$3 ( \2127 , \2126 );
nand \mul_16_12_g20297/U$1 ( \2128 , \1108 , \1113 );
not \mul_16_12_g20270/U$1 ( \2129 , \2128 );
not \mul_16_12_g20175/U$4 ( \2130 , \2129 );
or \mul_16_12_g20175/U$2 ( \2131 , \2127 , \2130 );
not \mul_16_12_g20351/U$1 ( \2132 , \2126 );
not \mul_16_12_g20185/U$3 ( \2133 , \2132 );
not \mul_16_12_g20185/U$4 ( \2134 , \2128 );
or \mul_16_12_g20185/U$2 ( \2135 , \2133 , \2134 );
not \mul_16_12_g20367/U$3 ( \2136 , \1145 );
not \mul_16_12_g20367/U$4 ( \2137 , \1067 );
or \mul_16_12_g20367/U$2 ( \2138 , \2136 , \2137 );
nand \mul_16_12_g20426/U$1 ( \2139 , \976 , \2036 );
nand \mul_16_12_g20367/U$1 ( \2140 , \2138 , \2139 );
nand \mul_16_12_g20185/U$1 ( \2141 , \2135 , \2140 );
nand \mul_16_12_g20175/U$1 ( \2142 , \2131 , \2141 );
not \mul_16_12_g20131/U$3 ( \2143 , \2142 );
xor \mul_16_12_g20717/U$1 ( \2144 , \2061 , \2048 );
xnor \mul_16_12_g20717/U$1_r1 ( \2145 , \2144 , \2054 );
not \mul_16_12_g20131/U$4 ( \2146 , \2145 );
or \mul_16_12_g20131/U$2 ( \2147 , \2143 , \2146 );
or \mul_16_12_g20131/U$5 ( \2148 , \2142 , \2145 );
nand \mul_16_12_g20131/U$1 ( \2149 , \2147 , \2148 );
xor \mul_16_12_g20130/U$1 ( \2150 , \2077 , \2092 );
xor \mul_16_12_g20130/U$1_r1 ( \2151 , \2150 , \2094 );
xor \mul_16_12_g20691/U$1 ( \2152 , \2149 , \2151 );
xor \mul_16_12_g20211/U$1 ( \2153 , \2078 , \2083 );
xor \mul_16_12_g20211/U$1_r1 ( \2154 , \2153 , \2089 );
xor \mul_16_12_g20202/U$4 ( \2155 , \1133 , \1140 );
and \mul_16_12_g20202/U$3 ( \2156 , \2155 , \1147 );
and \mul_16_12_g20202/U$5 ( \2157 , \1133 , \1140 );
or \mul_16_12_g20202/U$2 ( \2158 , \2156 , \2157 );
xor \mul_16_12_g20089/U$4 ( \2159 , \2154 , \2158 );
xor \mul_16_12_g20714/U$1 ( \2160 , \2126 , \2128 );
xnor \mul_16_12_g20714/U$1_r1 ( \2161 , \2160 , \2140 );
and \mul_16_12_g20089/U$3 ( \2162 , \2159 , \2161 );
and \mul_16_12_g20089/U$5 ( \2163 , \2154 , \2158 );
or \mul_16_12_g20089/U$2 ( \2164 , \2162 , \2163 );
nor \mul_16_12_g20043/U$1 ( \2165 , \2152 , \2164 );
xor \mul_16_12_g20109/U$4 ( \2166 , \1117 , \1121 );
and \mul_16_12_g20109/U$3 ( \2167 , \2166 , \1148 );
and \mul_16_12_g20109/U$5 ( \2168 , \1117 , \1121 );
or \mul_16_12_g20109/U$2 ( \2169 , \2167 , \2168 );
xor \mul_16_12_g20089/U$1 ( \2170 , \2154 , \2158 );
xor \mul_16_12_g20089/U$1_r1 ( \2171 , \2170 , \2161 );
nor \mul_16_12_g20065/U$1 ( \2172 , \2169 , \2171 );
nor \mul_16_12_g20036/U$1 ( \2173 , \2165 , \2172 );
not \g35901/U$4 ( \2174 , \2173 );
or \g35901/U$2 ( \2175 , \2121 , \2174 );
xor \mul_16_12_g20061/U$1 ( \2176 , \2070 , \2097 );
xnor \mul_16_12_g20061/U$1_r1 ( \2177 , \2176 , \2068 );
not \mul_16_12_g20132/U$2 ( \2178 , \2142 );
nand \mul_16_12_g20132/U$1 ( \2179 , \2178 , \2145 );
not \mul_16_12_g20072/U$3 ( \2180 , \2179 );
not \mul_16_12_g20072/U$4 ( \2181 , \2151 );
or \mul_16_12_g20072/U$2 ( \2182 , \2180 , \2181 );
not \mul_16_12_g20698/U$2 ( \2183 , \2145 );
nand \mul_16_12_g20698/U$1 ( \2184 , \2183 , \2142 );
nand \mul_16_12_g20072/U$1 ( \2185 , \2182 , \2184 );
not \mul_16_12_g20059/U$1 ( \2186 , \2185 );
nor \mul_16_12_g20039/U$1 ( \2187 , \2177 , \2186 );
nand \mul_16_12_g20067/U$1 ( \2188 , \2171 , \2169 );
or \mul_16_12_g20026/U$2 ( \2189 , \2165 , \2188 );
nand \mul_16_12_g20045/U$1 ( \2190 , \2152 , \2164 );
nand \mul_16_12_g20026/U$1 ( \2191 , \2189 , \2190 );
nor \mul_16_12_g20015/U$1 ( \2192 , \2187 , \2191 );
nand \g35901/U$1 ( \2193 , \2175 , \2192 );
not \mul_16_12_g19981/U$3 ( \2194 , \2193 );
xor \mul_16_12_g20031/U$1 ( \2195 , \1964 , \2024 );
xor \mul_16_12_g20031/U$1_r1 ( \2196 , \2195 , \2027 );
nand \mul_16_12_g20098/U$1 ( \2197 , \2110 , \2103 );
not \g36008/U$2 ( \2198 , \2197 );
not \g36009/U$3 ( \2199 , \2110 );
not \g36009/U$4 ( \2200 , \2103 );
and \g36009/U$2 ( \2201 , \2199 , \2200 );
buf \mul_16_12_g20092/U$1 ( \2202 , \2105 );
nor \g36009/U$1 ( \2203 , \2201 , \2202 );
nor \g36008/U$1 ( \2204 , \2198 , \2203 );
nand \mul_16_12_g20010/U$1 ( \2205 , \2196 , \2204 );
nand \mul_16_12_g20035/U$1 ( \2206 , \2177 , \2186 );
and \mul_16_12_g19998/U$1 ( \2207 , \2205 , \2206 );
not \mul_16_12_g19981/U$4 ( \2208 , \2207 );
or \mul_16_12_g19981/U$2 ( \2209 , \2194 , \2208 );
not \mul_16_12_g20007/U$2 ( \2210 , \2100 );
nor \mul_16_12_g20007/U$1 ( \2211 , \2210 , \2111 );
nand \mul_16_12_g19997/U$1 ( \2212 , \2205 , \2211 );
nand \mul_16_12_g19981/U$1 ( \2213 , \2209 , \2212 );
not \mul_16_12_g19966/U$4 ( \2214 , \2213 );
or \mul_16_12_g19966/U$2 ( \2215 , \2115 , \2214 );
not \mul_16_12_g20030/U$1 ( \2216 , \2030 );
not \mul_16_12_g19999/U$3 ( \2217 , \2216 );
not \fopt35505/U$1 ( \2218 , \1962 );
not \mul_16_12_g19999/U$4 ( \2219 , \2218 );
or \mul_16_12_g19999/U$2 ( \2220 , \2217 , \2219 );
nor \mul_16_12_g20017/U$1 ( \2221 , \2196 , \2204 );
not \fopt35672/U$1 ( \2222 , \2221 );
nand \mul_16_12_g19999/U$1 ( \2223 , \2220 , \2222 );
and \mul_16_12_g19968/U$2 ( \2224 , \1954 , \2223 , \2031 );
nor \mul_16_12_g19976/U$1 ( \2225 , \1908 , \1953 );
nor \mul_16_12_g19968/U$1 ( \2226 , \2224 , \2225 );
nand \mul_16_12_g19966/U$1 ( \2227 , \2215 , \2226 );
not \mul_16_12_g19965/U$4 ( \2228 , \2227 );
or \mul_16_12_g19965/U$2 ( \2229 , \1902 , \2228 );
or \mul_16_12_g19965/U$5 ( \2230 , \1901 , \2227 );
nand \mul_16_12_g19965/U$1 ( \2231 , \2229 , \2230 );
not \g35631/U$4 ( \2232 , \2231 );
or \g35631/U$2 ( \2233 , \1530 , \2232 );
xor \mul_17_13_g20655/U$1 ( \2234 , \b[2] , \c[11] );
not \mul_17_13_g20334/U$3 ( \2235 , \2234 );
xor \mul_17_13_g35711/U$1 ( \2236 , \c[10] , \c[9] );
xnor \g35473/U$1 ( \2237 , \c[11] , \c[10] );
nor \mul_17_13_g20540/U$1 ( \2238 , \2236 , \2237 );
not \mul_17_13_g20334/U$4 ( \2239 , \2238 );
or \mul_17_13_g20334/U$2 ( \2240 , \2235 , \2239 );
xor \g35479/U$1 ( \2241 , \c[11] , \b[3] );
nand \mul_17_13_g20493/U$1 ( \2242 , \2236 , \2241 );
nand \mul_17_13_g20334/U$1 ( \2243 , \2240 , \2242 );
xor \g35475/U$1 ( \2244 , \c[13] , \b[0] );
not \mul_17_13_g20323/U$3 ( \2245 , \2244 );
xor \mul_17_13_g20602/U$1 ( \2246 , \c[12] , \c[11] );
not \mul_17_13_g20554/U$3 ( \2247 , \c[12] );
not \mul_17_13_g20554/U$4 ( \2248 , \c[13] );
or \mul_17_13_g20554/U$2 ( \2249 , \2247 , \2248 );
or \mul_17_13_g20554/U$5 ( \2250 , \c[13] , \c[12] );
nand \mul_17_13_g20554/U$1 ( \2251 , \2249 , \2250 );
nor \mul_17_13_g20538/U$1 ( \2252 , \2246 , \2251 );
not \mul_17_13_g20323/U$4 ( \2253 , \2252 );
or \mul_17_13_g20323/U$2 ( \2254 , \2245 , \2253 );
xor \g35480/U$1 ( \2255 , \c[13] , \b[1] );
nand \mul_17_13_g20487/U$1 ( \2256 , \2246 , \2255 );
nand \mul_17_13_g20323/U$1 ( \2257 , \2254 , \2256 );
not \mul_17_13_g20322/U$1 ( \2258 , \2257 );
and \g36005/U$2 ( \2259 , \2243 , \2258 );
not \g36005/U$4 ( \2260 , \2243 );
and \g36005/U$3 ( \2261 , \2260 , \2257 );
or \g36005/U$1 ( \2262 , \2259 , \2261 );
xor \mul_17_13_g20607/U$1 ( \2263 , \b[8] , \c[5] );
not \mul_17_13_g20382/U$3 ( \2264 , \2263 );
buf \mul_17_13_g20447/U$1 ( \2265 , \736 );
not \mul_17_13_g20382/U$4 ( \2266 , \2265 );
or \mul_17_13_g20382/U$2 ( \2267 , \2264 , \2266 );
xor \mul_17_13_g20608/U$1 ( \2268 , \b[9] , \c[5] );
nand \mul_17_13_g20480/U$1 ( \2269 , \739 , \2268 );
nand \mul_17_13_g20382/U$1 ( \2270 , \2267 , \2269 );
not \mul_17_13_g20381/U$1 ( \2271 , \2270 );
and \mul_17_13_g20244/U$2 ( \2272 , \2262 , \2271 );
not \mul_17_13_g20244/U$4 ( \2273 , \2262 );
and \mul_17_13_g20244/U$3 ( \2274 , \2273 , \2270 );
nor \mul_17_13_g20244/U$1 ( \2275 , \2272 , \2274 );
not \mul_17_13_g20131/U$3 ( \2276 , \2275 );
xor \mul_17_13_g20642/U$1 ( \2277 , \b[4] , \c[9] );
not \mul_17_13_g20343/U$3 ( \2278 , \2277 );
xnor \mul_17_13_g20719/U$1 ( \2279 , \c[9] , \c[8] );
xor \mul_17_13_g35655/U$1 ( \2280 , \c[8] , \c[7] );
nor \mul_17_13_g20456/U$1 ( \2281 , \2279 , \2280 );
not \mul_17_13_g20343/U$4 ( \2282 , \2281 );
or \mul_17_13_g20343/U$2 ( \2283 , \2278 , \2282 );
buf \mul_17_13_g20591/U$1 ( \2284 , \2280 );
xor \mul_17_13_g20641/U$1 ( \2285 , \b[5] , \c[9] );
nand \mul_17_13_g20481/U$1 ( \2286 , \2284 , \2285 );
nand \mul_17_13_g20343/U$1 ( \2287 , \2283 , \2286 );
xor \mul_17_13_g20620/U$1 ( \2288 , \b[7] , \c[7] );
not \mul_17_13_g20351/U$3 ( \2289 , \2288 );
not \mul_17_13_g20351/U$4 ( \2290 , \714 );
or \mul_17_13_g20351/U$2 ( \2291 , \2289 , \2290 );
nor \mul_17_13_g20445/U$1 ( \2292 , \725 , \713 );
xor \mul_17_13_g20619/U$1 ( \2293 , \b[6] , \c[7] );
nand \mul_17_13_g20403/U$1 ( \2294 , \2292 , \2293 );
nand \mul_17_13_g20351/U$1 ( \2295 , \2291 , \2294 );
xor \mul_17_13_g20745/U$1 ( \2296 , \2287 , \2295 );
xor \mul_17_13_g20575/U$1 ( \2297 , \b[10] , \c[3] );
not \mul_17_13_g20398/U$3 ( \2298 , \2297 );
not \mul_17_13_g20398/U$4 ( \2299 , \746 );
or \mul_17_13_g20398/U$2 ( \2300 , \2298 , \2299 );
xor \mul_17_13_g20567/U$1 ( \2301 , \b[11] , \c[3] );
nand \mul_17_13_g20479/U$1 ( \2302 , \702 , \2301 );
nand \mul_17_13_g20398/U$1 ( \2303 , \2300 , \2302 );
xnor \mul_17_13_g20745/U$1_r1 ( \2304 , \2296 , \2303 );
not \mul_17_13_g20131/U$4 ( \2305 , \2304 );
or \mul_17_13_g20131/U$2 ( \2306 , \2276 , \2305 );
xor \mul_17_13_g20618/U$1 ( \2307 , \b[7] , \c[5] );
not \mul_17_13_g20364/U$3 ( \2308 , \2307 );
not \mul_17_13_g20364/U$4 ( \2309 , \2265 );
or \mul_17_13_g20364/U$2 ( \2310 , \2308 , \2309 );
nand \mul_17_13_g20441/U$1 ( \2311 , \739 , \2263 );
nand \mul_17_13_g20364/U$1 ( \2312 , \2310 , \2311 );
not \mul_17_13_g20165/U$3 ( \2313 , \2312 );
xor \mul_17_13_g20605/U$1 ( \2314 , \b[8] , \c[3] );
not \mul_17_13_g20390/U$3 ( \2315 , \2314 );
not \mul_17_13_g20390/U$4 ( \2316 , \746 );
or \mul_17_13_g20390/U$2 ( \2317 , \2315 , \2316 );
xor \mul_17_13_g20606/U$1 ( \2318 , \b[9] , \c[3] );
nand \mul_17_13_g20453/U$1 ( \2319 , \702 , \2318 );
nand \mul_17_13_g20390/U$1 ( \2320 , \2317 , \2319 );
or \mul_17_13_g20546/U$2 ( \2321 , \b[0] , \c[10] );
nand \mul_17_13_g20546/U$1 ( \2322 , \2321 , \c[9] );
nand \mul_17_13_g20672/U$1 ( \2323 , \b[0] , \c[10] );
nand \mul_17_13_g20532/U$1 ( \2324 , \2322 , \2323 , \c[11] );
not \mul_17_13_g20531/U$1 ( \2325 , \2324 );
and \mul_17_13_g20291/U$1 ( \2326 , \2320 , \2325 );
not \mul_17_13_g20165/U$4 ( \2327 , \2326 );
or \mul_17_13_g20165/U$2 ( \2328 , \2313 , \2327 );
or \g35841/U$2 ( \2329 , \2312 , \2326 );
xor \mul_17_13_g20556/U$1 ( \2330 , \b[10] , \c[1] );
not \mul_17_13_g20415/U$3 ( \2331 , \2330 );
not \mul_17_13_g20415/U$4 ( \2332 , \679 );
or \mul_17_13_g20415/U$2 ( \2333 , \2331 , \2332 );
xor \mul_17_13_g20557/U$1 ( \2334 , \b[11] , \c[1] );
nand \mul_17_13_g20443/U$1 ( \2335 , \2334 , \c[0] );
nand \mul_17_13_g20415/U$1 ( \2336 , \2333 , \2335 );
not \mul_17_13_g20254/U$3 ( \2337 , \2336 );
xor \mul_17_13_g20652/U$1 ( \2338 , \b[2] , \c[9] );
not \mul_17_13_g20336/U$3 ( \2339 , \2338 );
not \mul_17_13_g20336/U$4 ( \2340 , \2281 );
or \mul_17_13_g20336/U$2 ( \2341 , \2339 , \2340 );
xor \mul_17_13_g20651/U$1 ( \2342 , \b[3] , \c[9] );
nand \mul_17_13_g20488/U$1 ( \2343 , \2284 , \2342 );
nand \mul_17_13_g20336/U$1 ( \2344 , \2341 , \2343 );
not \mul_17_13_g20254/U$4 ( \2345 , \2344 );
or \mul_17_13_g20254/U$2 ( \2346 , \2337 , \2345 );
or \mul_17_13_g20264/U$2 ( \2347 , \2344 , \2336 );
xor \mul_17_13_g20632/U$1 ( \2348 , \b[4] , \c[7] );
not \mul_17_13_g20346/U$3 ( \2349 , \2348 );
not \mul_17_13_g20346/U$4 ( \2350 , \2292 );
or \mul_17_13_g20346/U$2 ( \2351 , \2349 , \2350 );
xor \mul_17_13_g20631/U$1 ( \2352 , \b[5] , \c[7] );
nand \mul_17_13_g20470/U$1 ( \2353 , \714 , \2352 );
nand \mul_17_13_g20346/U$1 ( \2354 , \2351 , \2353 );
nand \mul_17_13_g20264/U$1 ( \2355 , \2347 , \2354 );
nand \mul_17_13_g20254/U$1 ( \2356 , \2346 , \2355 );
nand \g35841/U$1 ( \2357 , \2329 , \2356 );
nand \mul_17_13_g20165/U$1 ( \2358 , \2328 , \2357 );
nand \mul_17_13_g20131/U$1 ( \2359 , \2306 , \2358 );
not \mul_17_13_g20736/U$2 ( \2360 , \2304 );
not \fopt35577/U$1 ( \2361 , \2275 );
nand \mul_17_13_g20736/U$1 ( \2362 , \2360 , \2361 );
nand \mul_17_13_g20117/U$1 ( \2363 , \2359 , \2362 );
xor \mul_17_13_g20609/U$1 ( \2364 , \c[14] , \c[13] );
and \mul_17_13_g20709/U$1 ( \2365 , \2364 , \b[0] );
xor \mul_17_13_g20565/U$1 ( \2366 , \b[13] , \c[1] );
not \mul_17_13_g20426/U$3 ( \2367 , \2366 );
not \mul_17_13_g20426/U$4 ( \2368 , \679 );
or \mul_17_13_g20426/U$2 ( \2369 , \2367 , \2368 );
xor \mul_17_13_g20566/U$1 ( \2370 , \b[14] , \c[1] );
nand \mul_17_13_g20503/U$1 ( \2371 , \2370 , \c[0] );
nand \mul_17_13_g20426/U$1 ( \2372 , \2369 , \2371 );
xor \mul_17_13_g20224/U$1 ( \2373 , \2365 , \2372 );
not \mul_17_13_g20402/U$3 ( \2374 , \2301 );
not \mul_17_13_g20402/U$4 ( \2375 , \746 );
or \mul_17_13_g20402/U$2 ( \2376 , \2374 , \2375 );
xor \mul_17_13_g20576/U$1 ( \2377 , \b[12] , \c[3] );
nand \mul_17_13_g20518/U$1 ( \2378 , \702 , \2377 );
nand \mul_17_13_g20402/U$1 ( \2379 , \2376 , \2378 );
xor \mul_17_13_g20224/U$1_r1 ( \2380 , \2373 , \2379 );
not \mul_17_13_g20216/U$3 ( \2381 , \2287 );
not \mul_17_13_g20216/U$4 ( \2382 , \2303 );
or \mul_17_13_g20216/U$2 ( \2383 , \2381 , \2382 );
or \mul_17_13_g20233/U$2 ( \2384 , \2303 , \2287 );
nand \mul_17_13_g20233/U$1 ( \2385 , \2384 , \2295 );
nand \mul_17_13_g20216/U$1 ( \2386 , \2383 , \2385 );
xor \mul_17_13_g20120/U$1 ( \2387 , \2380 , \2386 );
not \mul_17_13_g20263/U$3 ( \2388 , \2258 );
not \mul_17_13_g20263/U$4 ( \2389 , \2271 );
or \mul_17_13_g20263/U$2 ( \2390 , \2388 , \2389 );
nand \mul_17_13_g20263/U$1 ( \2391 , \2390 , \2243 );
nand \mul_17_13_g20287/U$1 ( \2392 , \2270 , \2257 );
nand \mul_17_13_g20257/U$1 ( \2393 , \2391 , \2392 );
xor \mul_17_13_g20120/U$1_r1 ( \2394 , \2387 , \2393 );
xor \mul_17_13_g20011/U$4 ( \2395 , \2363 , \2394 );
not \mul_17_13_g20348/U$3 ( \2396 , \2288 );
not \mul_17_13_g20348/U$4 ( \2397 , \2292 );
or \mul_17_13_g20348/U$2 ( \2398 , \2396 , \2397 );
xor \mul_17_13_g20610/U$1 ( \2399 , \b[8] , \c[7] );
nand \mul_17_13_g20466/U$1 ( \2400 , \714 , \2399 );
nand \mul_17_13_g20348/U$1 ( \2401 , \2398 , \2400 );
not \mul_17_13_g20337/U$3 ( \2402 , \2285 );
not \mul_17_13_g20337/U$4 ( \2403 , \2281 );
or \mul_17_13_g20337/U$2 ( \2404 , \2402 , \2403 );
xor \mul_17_13_g20626/U$1 ( \2405 , \b[6] , \c[9] );
nand \mul_17_13_g20467/U$1 ( \2406 , \2284 , \2405 );
nand \mul_17_13_g20337/U$1 ( \2407 , \2404 , \2406 );
xor \mul_17_13_g20226/U$1 ( \2408 , \2401 , \2407 );
not \mul_17_13_g20383/U$3 ( \2409 , \2268 );
not \mul_17_13_g20383/U$4 ( \2410 , \2265 );
or \mul_17_13_g20383/U$2 ( \2411 , \2409 , \2410 );
xor \mul_17_13_g20585/U$1 ( \2412 , \b[10] , \c[5] );
nand \mul_17_13_g20465/U$1 ( \2413 , \739 , \2412 );
nand \mul_17_13_g20383/U$1 ( \2414 , \2411 , \2413 );
xor \mul_17_13_g20226/U$1_r1 ( \2415 , \2408 , \2414 );
not \mul_17_13_g20318/U$3 ( \2416 , \2255 );
not \mul_17_13_g20318/U$4 ( \2417 , \2252 );
or \mul_17_13_g20318/U$2 ( \2418 , \2416 , \2417 );
xor \mul_17_13_g20663/U$1 ( \2419 , \b[2] , \c[13] );
nand \mul_17_13_g20463/U$1 ( \2420 , \2246 , \2419 );
nand \mul_17_13_g20318/U$1 ( \2421 , \2418 , \2420 );
not \mul_17_13_g20328/U$3 ( \2422 , \2241 );
not \mul_17_13_g20328/U$4 ( \2423 , \2238 );
or \mul_17_13_g20328/U$2 ( \2424 , \2422 , \2423 );
xor \mul_17_13_g20649/U$1 ( \2425 , \b[4] , \c[11] );
nand \mul_17_13_g20460/U$1 ( \2426 , \2236 , \2425 );
nand \mul_17_13_g20328/U$1 ( \2427 , \2424 , \2426 );
xor \mul_17_13_g20167/U$1 ( \2428 , \2421 , \2427 );
or \mul_17_13_g20545/U$2 ( \2429 , \b[0] , \c[12] );
nand \mul_17_13_g20545/U$1 ( \2430 , \2429 , \c[11] );
nand \mul_17_13_g20670/U$1 ( \2431 , \b[0] , \c[12] );
and \mul_17_13_g20715/U$1 ( \2432 , \2430 , \2431 , \c[13] );
xor \mul_17_13_g20555/U$1 ( \2433 , \b[12] , \c[1] );
not \mul_17_13_g20425/U$3 ( \2434 , \2433 );
not \mul_17_13_g20425/U$4 ( \2435 , \679 );
or \mul_17_13_g20425/U$2 ( \2436 , \2434 , \2435 );
nand \mul_17_13_g20502/U$1 ( \2437 , \2366 , \c[0] );
nand \mul_17_13_g20425/U$1 ( \2438 , \2436 , \2437 );
and \mul_17_13_g20278/U$2 ( \2439 , \2432 , \2438 );
xor \mul_17_13_g20167/U$1_r1 ( \2440 , \2428 , \2439 );
xor \mul_17_13_g20081/U$1 ( \2441 , \2415 , \2440 );
not \mul_17_13_g20428/U$3 ( \2442 , \2334 );
not \mul_17_13_g20428/U$4 ( \2443 , \679 );
or \mul_17_13_g20428/U$2 ( \2444 , \2442 , \2443 );
nand \mul_17_13_g20504/U$1 ( \2445 , \2433 , \c[0] );
nand \mul_17_13_g20428/U$1 ( \2446 , \2444 , \2445 );
not \mul_17_13_g20338/U$3 ( \2447 , \2342 );
nor \mul_17_13_g20457/U$1 ( \2448 , \2279 , \2280 );
not \mul_17_13_g20338/U$4 ( \2449 , \2448 );
or \mul_17_13_g20338/U$2 ( \2450 , \2447 , \2449 );
nand \mul_17_13_g20472/U$1 ( \2451 , \2284 , \2277 );
nand \mul_17_13_g20338/U$1 ( \2452 , \2450 , \2451 );
xor \mul_17_13_g20211/U$4 ( \2453 , \2446 , \2452 );
xor \mul_17_13_g20660/U$1 ( \2454 , \b[1] , \c[11] );
not \mul_17_13_g20329/U$3 ( \2455 , \2454 );
not \mul_17_13_g20329/U$4 ( \2456 , \2238 );
or \mul_17_13_g20329/U$2 ( \2457 , \2455 , \2456 );
nand \mul_17_13_g20473/U$1 ( \2458 , \2236 , \2234 );
nand \mul_17_13_g20329/U$1 ( \2459 , \2457 , \2458 );
and \mul_17_13_g20211/U$3 ( \2460 , \2453 , \2459 );
and \mul_17_13_g20211/U$5 ( \2461 , \2446 , \2452 );
or \mul_17_13_g20211/U$2 ( \2462 , \2460 , \2461 );
xor \mul_17_13_g20278/U$1 ( \2463 , \2432 , \2438 );
or \mul_17_13_g20163/U$2 ( \2464 , \2462 , \2463 );
and \mul_17_13_g20501/U$1 ( \2465 , \2246 , \b[0] );
not \mul_17_13_g20357/U$3 ( \2466 , \2352 );
not \mul_17_13_g20357/U$4 ( \2467 , \726 );
or \mul_17_13_g20357/U$2 ( \2468 , \2466 , \2467 );
nand \mul_17_13_g20492/U$1 ( \2469 , \714 , \2293 );
nand \mul_17_13_g20357/U$1 ( \2470 , \2468 , \2469 );
xor \mul_17_13_g20208/U$4 ( \2471 , \2465 , \2470 );
not \mul_17_13_g20393/U$3 ( \2472 , \2318 );
not \mul_17_13_g20393/U$4 ( \2473 , \699 );
or \mul_17_13_g20393/U$2 ( \2474 , \2472 , \2473 );
nand \mul_17_13_g20464/U$1 ( \2475 , \702 , \2297 );
nand \mul_17_13_g20393/U$1 ( \2476 , \2474 , \2475 );
and \mul_17_13_g20208/U$3 ( \2477 , \2471 , \2476 );
and \mul_17_13_g20208/U$5 ( \2478 , \2465 , \2470 );
or \mul_17_13_g20208/U$2 ( \2479 , \2477 , \2478 );
nand \mul_17_13_g20163/U$1 ( \2480 , \2464 , \2479 );
nand \mul_17_13_g20176/U$1 ( \2481 , \2462 , \2463 );
nand \mul_17_13_g20154/U$1 ( \2482 , \2480 , \2481 );
xor \mul_17_13_g20081/U$1_r1 ( \2483 , \2441 , \2482 );
and \mul_17_13_g20011/U$3 ( \2484 , \2395 , \2483 );
and \mul_17_13_g20011/U$5 ( \2485 , \2363 , \2394 );
or \mul_17_13_g20011/U$2 ( \2486 , \2484 , \2485 );
xor \mul_17_13_g20081/U$4 ( \2487 , \2415 , \2440 );
and \mul_17_13_g20081/U$3 ( \2488 , \2487 , \2482 );
and \mul_17_13_g20081/U$5 ( \2489 , \2415 , \2440 );
or \mul_17_13_g20081/U$2 ( \2490 , \2488 , \2489 );
not \mul_17_13_g20060/U$3 ( \2491 , \2490 );
xor \mul_17_13_g20120/U$4 ( \2492 , \2380 , \2386 );
and \mul_17_13_g20120/U$3 ( \2493 , \2492 , \2393 );
and \mul_17_13_g20120/U$5 ( \2494 , \2380 , \2386 );
or \mul_17_13_g20120/U$2 ( \2495 , \2493 , \2494 );
not \fopt35670/U$1 ( \2496 , \2495 );
not \mul_17_13_g20060/U$4 ( \2497 , \2496 );
and \mul_17_13_g20060/U$2 ( \2498 , \2491 , \2497 );
and \mul_17_13_g20060/U$5 ( \2499 , \2490 , \2496 );
nor \mul_17_13_g20060/U$1 ( \2500 , \2498 , \2499 );
not \mul_17_13_g20401/U$3 ( \2501 , \2377 );
not \mul_17_13_g20401/U$4 ( \2502 , \746 );
or \mul_17_13_g20401/U$2 ( \2503 , \2501 , \2502 );
xor \mul_17_13_g20569/U$1 ( \2504 , \b[13] , \c[3] );
nand \mul_17_13_g20517/U$1 ( \2505 , \702 , \2504 );
nand \mul_17_13_g20401/U$1 ( \2506 , \2503 , \2505 );
not \mul_17_13_g20385/U$3 ( \2507 , \2412 );
not \mul_17_13_g20385/U$4 ( \2508 , \2265 );
or \mul_17_13_g20385/U$2 ( \2509 , \2507 , \2508 );
xor \mul_17_13_g20584/U$1 ( \2510 , \b[11] , \c[5] );
nand \mul_17_13_g20497/U$1 ( \2511 , \739 , \2510 );
nand \mul_17_13_g20385/U$1 ( \2512 , \2509 , \2511 );
xor \g35463/U$1 ( \2513 , \2506 , \2512 );
xor \mul_17_13_g20224/U$4 ( \2514 , \2365 , \2372 );
and \mul_17_13_g20224/U$3 ( \2515 , \2514 , \2379 );
and \mul_17_13_g20224/U$5 ( \2516 , \2365 , \2372 );
or \mul_17_13_g20224/U$2 ( \2517 , \2515 , \2516 );
xor \g35463/U$1_r1 ( \2518 , \2513 , \2517 );
not \mul_17_13_g20358/U$3 ( \2519 , \2399 );
not \mul_17_13_g20358/U$4 ( \2520 , \2292 );
or \mul_17_13_g20358/U$2 ( \2521 , \2519 , \2520 );
not \mul_17_13_g20677/U$2 ( \2522 , \c[7] );
nand \mul_17_13_g20677/U$1 ( \2523 , \2522 , \b[9] );
not \mul_17_13_g20431/U$3 ( \2524 , \2523 );
not \mul_17_13_g20679/U$2 ( \2525 , \b[9] );
nand \mul_17_13_g20679/U$1 ( \2526 , \2525 , \c[7] );
not \mul_17_13_g20431/U$4 ( \2527 , \2526 );
or \mul_17_13_g20431/U$2 ( \2528 , \2524 , \2527 );
nand \mul_17_13_g20431/U$1 ( \2529 , \2528 , \714 );
nand \mul_17_13_g20358/U$1 ( \2530 , \2521 , \2529 );
not \mul_17_13_g20344/U$3 ( \2531 , \2405 );
not \mul_17_13_g20344/U$4 ( \2532 , \2281 );
or \mul_17_13_g20344/U$2 ( \2533 , \2531 , \2532 );
xor \mul_17_13_g20627/U$1 ( \2534 , \b[7] , \c[9] );
nand \mul_17_13_g20433/U$1 ( \2535 , \2284 , \2534 );
nand \mul_17_13_g20344/U$1 ( \2536 , \2533 , \2535 );
xor \mul_17_13_g20203/U$1 ( \2537 , \2530 , \2536 );
not \mul_17_13_g20319/U$3 ( \2538 , \2419 );
not \mul_17_13_g20319/U$4 ( \2539 , \2252 );
or \mul_17_13_g20319/U$2 ( \2540 , \2538 , \2539 );
xor \mul_17_13_g20662/U$1 ( \2541 , \b[3] , \c[13] );
nand \mul_17_13_g20500/U$1 ( \2542 , \2246 , \2541 );
nand \mul_17_13_g20319/U$1 ( \2543 , \2540 , \2542 );
not \mul_17_13_g20284/U$3 ( \2544 , \2543 );
xnor \mul_17_13_g20720/U$1 ( \2545 , \b[1] , \c[15] );
and \mul_17_13_g20708/U$2 ( \2546 , \2364 , \2545 );
not \mul_17_13_g20708/U$4 ( \2547 , \2364 );
xor \mul_17_13_g20638/U$1 ( \2548 , \c[15] , \c[14] );
xor \mul_17_13_g20593/U$1 ( \2549 , \b[0] , \c[15] );
nand \mul_17_13_g20498/U$1 ( \2550 , \2548 , \2549 );
and \mul_17_13_g20708/U$3 ( \2551 , \2547 , \2550 );
or \mul_17_13_g20708/U$1 ( \2552 , \2546 , \2551 );
not \mul_17_13_g20284/U$4 ( \2553 , \2552 );
and \mul_17_13_g20284/U$2 ( \2554 , \2544 , \2553 );
and \mul_17_13_g20284/U$5 ( \2555 , \2543 , \2552 );
nor \mul_17_13_g20284/U$1 ( \2556 , \2554 , \2555 );
xor \mul_17_13_g20203/U$1_r1 ( \2557 , \2537 , \2556 );
xnor \mul_17_13_g20735/U$1 ( \2558 , \2518 , \2557 );
not \mul_17_13_g20080/U$3 ( \2559 , \2558 );
xor \mul_17_13_g20167/U$4 ( \2560 , \2421 , \2427 );
and \mul_17_13_g20167/U$3 ( \2561 , \2560 , \2439 );
and \mul_17_13_g20167/U$5 ( \2562 , \2421 , \2427 );
or \mul_17_13_g20167/U$2 ( \2563 , \2561 , \2562 );
not \mul_17_13_g20134/U$3 ( \2564 , \2563 );
not \mul_17_13_g20427/U$3 ( \2565 , \2370 );
not \mul_17_13_g20427/U$4 ( \2566 , \679 );
or \mul_17_13_g20427/U$2 ( \2567 , \2565 , \2566 );
xor \mul_17_13_g20558/U$1 ( \2568 , \b[15] , \c[1] );
nand \mul_17_13_g20507/U$1 ( \2569 , \2568 , \c[0] );
nand \mul_17_13_g20427/U$1 ( \2570 , \2567 , \2569 );
or \mul_17_13_g20544/U$2 ( \2571 , \b[0] , \c[14] );
nand \mul_17_13_g20544/U$1 ( \2572 , \2571 , \c[13] );
nand \mul_17_13_g20675/U$1 ( \2573 , \b[0] , \c[14] );
nand \mul_17_13_g20536/U$1 ( \2574 , \2572 , \2573 , \c[15] );
xor \g35913/U$1 ( \2575 , \2570 , \2574 );
not \mul_17_13_g20331/U$3 ( \2576 , \2425 );
not \mul_17_13_g20331/U$4 ( \2577 , \2238 );
or \mul_17_13_g20331/U$2 ( \2578 , \2576 , \2577 );
xor \mul_17_13_g20650/U$1 ( \2579 , \b[5] , \c[11] );
nand \mul_17_13_g20458/U$1 ( \2580 , \2236 , \2579 );
nand \mul_17_13_g20331/U$1 ( \2581 , \2578 , \2580 );
xor \g35913/U$1_r1 ( \2582 , \2575 , \2581 );
not \mul_17_13_g20134/U$4 ( \2583 , \2582 );
and \mul_17_13_g20134/U$2 ( \2584 , \2564 , \2583 );
and \mul_17_13_g20134/U$5 ( \2585 , \2563 , \2582 );
nor \mul_17_13_g20134/U$1 ( \2586 , \2584 , \2585 );
xor \mul_17_13_g20226/U$4 ( \2587 , \2401 , \2407 );
and \mul_17_13_g20226/U$3 ( \2588 , \2587 , \2414 );
and \mul_17_13_g20226/U$5 ( \2589 , \2401 , \2407 );
or \mul_17_13_g20226/U$2 ( \2590 , \2588 , \2589 );
xor \mul_17_13_g20738/U$1 ( \2591 , \2586 , \2590 );
not \mul_17_13_g20080/U$4 ( \2592 , \2591 );
or \mul_17_13_g20080/U$2 ( \2593 , \2559 , \2592 );
or \mul_17_13_g20728/U$1 ( \2594 , \2591 , \2558 );
nand \mul_17_13_g20080/U$1 ( \2595 , \2593 , \2594 );
xor \mul_17_13_g20726/U$1 ( \2596 , \2500 , \2595 );
xor \mul_17_13_g20758/U$1 ( \2597 , \2486 , \2596 );
not \mul_17_13_g19986/U$3 ( \2598 , \2597 );
xor \mul_17_13_g20011/U$1 ( \2599 , \2363 , \2394 );
xor \mul_17_13_g20011/U$1_r1 ( \2600 , \2599 , \2483 );
not \g35908/U$3 ( \2601 , \2600 );
xor \mul_17_13_g20135/U$1 ( \2602 , \2463 , \2479 );
xnor \mul_17_13_g20135/U$1_r1 ( \2603 , \2602 , \2462 );
not \mul_17_13_g20121/U$1 ( \2604 , \2603 );
not \mul_17_13_g20068/U$3 ( \2605 , \2604 );
not \mul_17_13_g20175/U$3 ( \2606 , \2275 );
not \mul_17_13_g20209/U$1 ( \2607 , \2304 );
not \mul_17_13_g20175/U$4 ( \2608 , \2607 );
or \mul_17_13_g20175/U$2 ( \2609 , \2606 , \2608 );
nand \mul_17_13_g20177/U$1 ( \2610 , \2361 , \2304 );
nand \mul_17_13_g20175/U$1 ( \2611 , \2609 , \2610 );
and \mul_17_13_g20126/U$2 ( \2612 , \2611 , \2358 );
not \mul_17_13_g20126/U$4 ( \2613 , \2611 );
not \mul_17_13_g20162/U$1 ( \2614 , \2358 );
and \mul_17_13_g20126/U$3 ( \2615 , \2613 , \2614 );
nor \mul_17_13_g20126/U$1 ( \2616 , \2612 , \2615 );
not \mul_17_13_g20068/U$4 ( \2617 , \2616 );
or \mul_17_13_g20068/U$2 ( \2618 , \2605 , \2617 );
not \mul_17_13_g20073/U$3 ( \2619 , \2603 );
not \mul_17_13_g20104/U$1 ( \2620 , \2616 );
not \mul_17_13_g20073/U$4 ( \2621 , \2620 );
or \mul_17_13_g20073/U$2 ( \2622 , \2619 , \2621 );
xor \mul_17_13_g20208/U$1 ( \2623 , \2465 , \2470 );
xor \mul_17_13_g20208/U$1_r1 ( \2624 , \2623 , \2476 );
not \mul_17_13_g20116/U$3 ( \2625 , \2624 );
xor \mul_17_13_g20211/U$1 ( \2626 , \2446 , \2452 );
xor \mul_17_13_g20211/U$1_r1 ( \2627 , \2626 , \2459 );
not \mul_17_13_g20116/U$4 ( \2628 , \2627 );
or \mul_17_13_g20116/U$2 ( \2629 , \2625 , \2628 );
or \mul_17_13_g20130/U$2 ( \2630 , \2627 , \2624 );
xor \g35477/U$1 ( \2631 , \c[11] , \b[0] );
not \mul_17_13_g20327/U$3 ( \2632 , \2631 );
not \mul_17_13_g20327/U$4 ( \2633 , \2238 );
or \mul_17_13_g20327/U$2 ( \2634 , \2632 , \2633 );
nand \mul_17_13_g20437/U$1 ( \2635 , \2236 , \2454 );
nand \mul_17_13_g20327/U$1 ( \2636 , \2634 , \2635 );
not \g35851/U$2 ( \2637 , \2636 );
xor \mul_17_13_g20617/U$1 ( \2638 , \b[6] , \c[5] );
not \mul_17_13_g20360/U$3 ( \2639 , \2638 );
not \mul_17_13_g20360/U$4 ( \2640 , \2265 );
or \mul_17_13_g20360/U$2 ( \2641 , \2639 , \2640 );
nand \mul_17_13_g20435/U$1 ( \2642 , \739 , \2307 );
nand \mul_17_13_g20360/U$1 ( \2643 , \2641 , \2642 );
not \mul_17_13_g20359/U$1 ( \2644 , \2643 );
nand \g35851/U$1 ( \2645 , \2637 , \2644 );
not \mul_17_13_g20214/U$3 ( \2646 , \2645 );
and \mul_17_13_g20749/U$2 ( \2647 , \2320 , \2325 );
not \mul_17_13_g20749/U$4 ( \2648 , \2320 );
and \mul_17_13_g20749/U$3 ( \2649 , \2648 , \2324 );
nor \mul_17_13_g20749/U$1 ( \2650 , \2647 , \2649 );
not \mul_17_13_g20214/U$4 ( \2651 , \2650 );
or \mul_17_13_g20214/U$2 ( \2652 , \2646 , \2651 );
nand \mul_17_13_g20294/U$1 ( \2653 , \2643 , \2636 );
nand \mul_17_13_g20214/U$1 ( \2654 , \2652 , \2653 );
nand \mul_17_13_g20130/U$1 ( \2655 , \2630 , \2654 );
nand \mul_17_13_g20116/U$1 ( \2656 , \2629 , \2655 );
nand \mul_17_13_g20073/U$1 ( \2657 , \2622 , \2656 );
nand \mul_17_13_g20068/U$1 ( \2658 , \2618 , \2657 );
not \g35908/U$4 ( \2659 , \2658 );
and \g35908/U$2 ( \2660 , \2601 , \2659 );
not \mul_17_13_g20084/U$3 ( \2661 , \2603 );
not \mul_17_13_g20084/U$4 ( \2662 , \2656 );
or \mul_17_13_g20084/U$2 ( \2663 , \2661 , \2662 );
or \mul_17_13_g20084/U$5 ( \2664 , \2603 , \2656 );
nand \mul_17_13_g20084/U$1 ( \2665 , \2663 , \2664 );
and \mul_17_13_g20061/U$2 ( \2666 , \2665 , \2620 );
not \mul_17_13_g20061/U$4 ( \2667 , \2665 );
and \mul_17_13_g20061/U$3 ( \2668 , \2667 , \2616 );
nor \mul_17_13_g20061/U$1 ( \2669 , \2666 , \2668 );
xor \mul_17_13_g20166/U$1 ( \2670 , \2312 , \2326 );
xnor \mul_17_13_g20166/U$1_r1 ( \2671 , \2670 , \2356 );
not \mul_17_13_g20074/U$3 ( \2672 , \2671 );
xor \mul_17_13_g20127/U$1 ( \2673 , \2624 , \2627 );
xnor \mul_17_13_g20127/U$1_r1 ( \2674 , \2673 , \2654 );
not \mul_17_13_g20074/U$4 ( \2675 , \2674 );
or \mul_17_13_g20074/U$2 ( \2676 , \2672 , \2675 );
and \mul_17_13_g20711/U$1 ( \2677 , \2236 , \b[0] );
xor \mul_17_13_g20645/U$1 ( \2678 , \b[3] , \c[7] );
not \mul_17_13_g20352/U$3 ( \2679 , \2678 );
not \mul_17_13_g20352/U$4 ( \2680 , \726 );
or \mul_17_13_g20352/U$2 ( \2681 , \2679 , \2680 );
nand \mul_17_13_g20482/U$1 ( \2682 , \714 , \2348 );
nand \mul_17_13_g20352/U$1 ( \2683 , \2681 , \2682 );
xor \mul_17_13_g20212/U$4 ( \2684 , \2677 , \2683 );
xor \mul_17_13_g20616/U$1 ( \2685 , \b[7] , \c[3] );
not \mul_17_13_g20397/U$3 ( \2686 , \2685 );
not \mul_17_13_g20397/U$4 ( \2687 , \699 );
or \mul_17_13_g20397/U$2 ( \2688 , \2686 , \2687 );
nand \mul_17_13_g20439/U$1 ( \2689 , \702 , \2314 );
nand \mul_17_13_g20397/U$1 ( \2690 , \2688 , \2689 );
and \mul_17_13_g20212/U$3 ( \2691 , \2684 , \2690 );
and \mul_17_13_g20212/U$5 ( \2692 , \2677 , \2683 );
or \mul_17_13_g20212/U$2 ( \2693 , \2691 , \2692 );
xor \mul_17_13_g20657/U$1 ( \2694 , \b[1] , \c[9] );
not \mul_17_13_g20341/U$3 ( \2695 , \2694 );
not \mul_17_13_g20341/U$4 ( \2696 , \2448 );
or \mul_17_13_g20341/U$2 ( \2697 , \2695 , \2696 );
nand \mul_17_13_g20474/U$1 ( \2698 , \2280 , \2338 );
nand \mul_17_13_g20341/U$1 ( \2699 , \2697 , \2698 );
xor \mul_17_13_g20604/U$1 ( \2700 , \b[9] , \c[1] );
not \mul_17_13_g20419/U$3 ( \2701 , \2700 );
not \mul_17_13_g20419/U$4 ( \2702 , \679 );
or \mul_17_13_g20419/U$2 ( \2703 , \2701 , \2702 );
nand \mul_17_13_g20483/U$1 ( \2704 , \2330 , \c[0] );
nand \mul_17_13_g20419/U$1 ( \2705 , \2703 , \2704 );
or \mul_17_13_g20234/U$2 ( \2706 , \2699 , \2705 );
xor \mul_17_13_g20629/U$1 ( \2707 , \b[5] , \c[5] );
not \mul_17_13_g20378/U$3 ( \2708 , \2707 );
not \mul_17_13_g20378/U$4 ( \2709 , \736 );
or \mul_17_13_g20378/U$2 ( \2710 , \2708 , \2709 );
nand \mul_17_13_g20489/U$1 ( \2711 , \739 , \2638 );
nand \mul_17_13_g20378/U$1 ( \2712 , \2710 , \2711 );
nand \mul_17_13_g20234/U$1 ( \2713 , \2706 , \2712 );
nand \mul_17_13_g20293/U$1 ( \2714 , \2699 , \2705 );
nand \mul_17_13_g20215/U$1 ( \2715 , \2713 , \2714 );
nor \mul_17_13_g20180/U$1 ( \2716 , \2693 , \2715 );
xor \g35911/U$1 ( \2717 , \2354 , \2336 );
xnor \mul_17_13_g20744/U$1 ( \2718 , \2717 , \2344 );
or \mul_17_13_g20158/U$2 ( \2719 , \2716 , \2718 );
nand \mul_17_13_g20178/U$1 ( \2720 , \2693 , \2715 );
nand \mul_17_13_g20158/U$1 ( \2721 , \2719 , \2720 );
nand \mul_17_13_g20074/U$1 ( \2722 , \2676 , \2721 );
not \mul_17_13_g20733/U$2 ( \2723 , \2671 );
not \mul_17_13_g20107/U$1 ( \2724 , \2674 );
nand \mul_17_13_g20733/U$1 ( \2725 , \2723 , \2724 );
nand \mul_17_13_g20069/U$1 ( \2726 , \2722 , \2725 );
not \mul_17_13_g20059/U$1 ( \2727 , \2726 );
nand \mul_17_13_g20028/U$1 ( \2728 , \2669 , \2727 );
not \g35924/U$3 ( \2729 , \2644 );
not \g35924/U$4 ( \2730 , \2636 );
or \g35924/U$2 ( \2731 , \2729 , \2730 );
not \g35698/U$2 ( \2732 , \2636 );
nand \g35698/U$1 ( \2733 , \2732 , \2643 );
nand \g35924/U$1 ( \2734 , \2731 , \2733 );
xnor \mul_17_13_g20739/U$1 ( \2735 , \2734 , \2650 );
or \mul_17_13_g20547/U$2 ( \2736 , \b[0] , \c[8] );
nand \mul_17_13_g20547/U$1 ( \2737 , \2736 , \c[7] );
nand \mul_17_13_g20666/U$1 ( \2738 , \b[0] , \c[8] );
and \mul_17_13_g20714/U$1 ( \2739 , \2737 , \2738 , \c[9] );
xor \mul_17_13_g20615/U$1 ( \2740 , \b[6] , \c[3] );
not \mul_17_13_g20399/U$3 ( \2741 , \2740 );
not \mul_17_13_g20399/U$4 ( \2742 , \699 );
or \mul_17_13_g20399/U$2 ( \2743 , \2741 , \2742 );
nand \mul_17_13_g20494/U$1 ( \2744 , \702 , \2685 );
nand \mul_17_13_g20399/U$1 ( \2745 , \2743 , \2744 );
and \mul_17_13_g20258/U$2 ( \2746 , \2739 , \2745 );
xor \mul_17_13_g20212/U$1 ( \2747 , \2677 , \2683 );
xor \mul_17_13_g20212/U$1_r1 ( \2748 , \2747 , \2690 );
xor \mul_17_13_g20139/U$4 ( \2749 , \2746 , \2748 );
xor \g35478/U$1 ( \2750 , \c[9] , \b[0] );
not \mul_17_13_g20340/U$3 ( \2751 , \2750 );
not \mul_17_13_g20340/U$4 ( \2752 , \2281 );
or \mul_17_13_g20340/U$2 ( \2753 , \2751 , \2752 );
nand \mul_17_13_g20432/U$1 ( \2754 , \2284 , \2694 );
nand \mul_17_13_g20340/U$1 ( \2755 , \2753 , \2754 );
xor \g35474/U$1 ( \2756 , \c[1] , \b[8] );
not \mul_17_13_g20424/U$3 ( \2757 , \2756 );
not \mul_17_13_g20424/U$4 ( \2758 , \679 );
or \mul_17_13_g20424/U$2 ( \2759 , \2757 , \2758 );
nand \mul_17_13_g20499/U$1 ( \2760 , \2700 , \c[0] );
nand \mul_17_13_g20424/U$1 ( \2761 , \2759 , \2760 );
or \mul_17_13_g20262/U$2 ( \2762 , \2755 , \2761 );
xor \mul_17_13_g20646/U$1 ( \2763 , \b[2] , \c[7] );
not \mul_17_13_g20356/U$3 ( \2764 , \2763 );
not \mul_17_13_g20356/U$4 ( \2765 , \726 );
or \mul_17_13_g20356/U$2 ( \2766 , \2764 , \2765 );
nand \mul_17_13_g20430/U$1 ( \2767 , \714 , \2678 );
nand \mul_17_13_g20356/U$1 ( \2768 , \2766 , \2767 );
nand \mul_17_13_g20262/U$1 ( \2769 , \2762 , \2768 );
nand \mul_17_13_g20290/U$1 ( \2770 , \2755 , \2761 );
nand \mul_17_13_g20255/U$1 ( \2771 , \2769 , \2770 );
and \mul_17_13_g20139/U$3 ( \2772 , \2749 , \2771 );
and \mul_17_13_g20139/U$5 ( \2773 , \2746 , \2748 );
or \mul_17_13_g20139/U$2 ( \2774 , \2772 , \2773 );
not \mul_17_13_g20138/U$1 ( \2775 , \2774 );
xor \mul_17_13_g20058/U$1 ( \2776 , \2735 , \2775 );
xor \mul_17_13_g20144/U$1 ( \2777 , \2715 , \2693 );
xor \mul_17_13_g20144/U$1_r1 ( \2778 , \2777 , \2718 );
xor \mul_17_13_g20058/U$1_r1 ( \2779 , \2776 , \2778 );
xor \g35914/U$1 ( \2780 , \2705 , \2699 );
xor \g35914/U$1_r1 ( \2781 , \2780 , \2712 );
xor \mul_17_13_g20139/U$1 ( \2782 , \2746 , \2748 );
xor \mul_17_13_g20139/U$1_r1 ( \2783 , \2782 , \2771 );
or \g35945/U$2 ( \2784 , \2781 , \2783 );
xor \mul_17_13_g20628/U$1 ( \2785 , \b[4] , \c[5] );
not \mul_17_13_g20361/U$3 ( \2786 , \2785 );
not \mul_17_13_g20361/U$4 ( \2787 , \2265 );
or \mul_17_13_g20361/U$2 ( \2788 , \2786 , \2787 );
nand \mul_17_13_g20436/U$1 ( \2789 , \739 , \2707 );
nand \mul_17_13_g20361/U$1 ( \2790 , \2788 , \2789 );
xor \mul_17_13_g20258/U$1 ( \2791 , \2739 , \2745 );
xor \mul_17_13_g20141/U$4 ( \2792 , \2790 , \2791 );
not \mul_17_13_g20404/U$3 ( \2793 , \682 );
not \mul_17_13_g20404/U$4 ( \2794 , \679 );
or \mul_17_13_g20404/U$2 ( \2795 , \2793 , \2794 );
nand \mul_17_13_g20440/U$1 ( \2796 , \2756 , \c[0] );
nand \mul_17_13_g20404/U$1 ( \2797 , \2795 , \2796 );
and \mul_17_13_g20712/U$1 ( \2798 , \2280 , \b[0] );
or \mul_17_13_g20253/U$2 ( \2799 , \2797 , \2798 );
not \mul_17_13_g20345/U$3 ( \2800 , \729 );
not \mul_17_13_g20345/U$4 ( \2801 , \2292 );
or \mul_17_13_g20345/U$2 ( \2802 , \2800 , \2801 );
nand \mul_17_13_g20442/U$1 ( \2803 , \714 , \2763 );
nand \mul_17_13_g20345/U$1 ( \2804 , \2802 , \2803 );
nand \mul_17_13_g20253/U$1 ( \2805 , \2799 , \2804 );
nand \mul_17_13_g20304/U$1 ( \2806 , \2797 , \2798 );
nand \mul_17_13_g20236/U$1 ( \2807 , \2805 , \2806 );
and \mul_17_13_g20141/U$3 ( \2808 , \2792 , \2807 );
and \mul_17_13_g20141/U$5 ( \2809 , \2790 , \2791 );
or \mul_17_13_g20141/U$2 ( \2810 , \2808 , \2809 );
nand \g35945/U$1 ( \2811 , \2784 , \2810 );
nand \mul_17_13_g20110/U$1 ( \2812 , \2783 , \2781 );
and \g35944/U$1 ( \2813 , \2811 , \2812 );
nand \mul_17_13_g20037/U$1 ( \2814 , \2779 , \2813 );
nand \mul_17_13_g20017/U$1 ( \2815 , \2728 , \2814 );
nor \g35908/U$1 ( \2816 , \2660 , \2815 );
not \mul_17_13_g19988/U$3 ( \2817 , \2816 );
not \mul_17_13_g20096/U$3 ( \2818 , \2721 );
not \mul_17_13_g20096/U$4 ( \2819 , \2671 );
or \mul_17_13_g20096/U$2 ( \2820 , \2818 , \2819 );
or \mul_17_13_g20096/U$5 ( \2821 , \2671 , \2721 );
nand \mul_17_13_g20096/U$1 ( \2822 , \2820 , \2821 );
and \mul_17_13_g20071/U$2 ( \2823 , \2822 , \2674 );
not \mul_17_13_g20071/U$4 ( \2824 , \2822 );
and \mul_17_13_g20071/U$3 ( \2825 , \2824 , \2724 );
nor \mul_17_13_g20071/U$1 ( \2826 , \2823 , \2825 );
xor \mul_17_13_g20058/U$4 ( \2827 , \2735 , \2775 );
and \mul_17_13_g20058/U$3 ( \2828 , \2827 , \2778 );
and \mul_17_13_g20058/U$5 ( \2829 , \2735 , \2775 );
or \mul_17_13_g20058/U$2 ( \2830 , \2828 , \2829 );
nand \mul_17_13_g35647/U$1 ( \2831 , \2826 , \2830 );
xor \mul_17_13_g20085/U$1 ( \2832 , \2781 , \2810 );
xnor \mul_17_13_g20085/U$1_r1 ( \2833 , \2832 , \2783 );
not \mul_17_13_g20367/U$3 ( \2834 , \740 );
not \mul_17_13_g20367/U$4 ( \2835 , \736 );
or \mul_17_13_g20367/U$2 ( \2836 , \2834 , \2835 );
nand \mul_17_13_g20446/U$1 ( \2837 , \739 , \2785 );
nand \mul_17_13_g20367/U$1 ( \2838 , \2836 , \2837 );
not \mul_17_13_g20366/U$1 ( \2839 , \2838 );
not \mul_17_13_g20201/U$3 ( \2840 , \2839 );
not \mul_17_13_g20753/U$2 ( \2841 , \689 );
nand \mul_17_13_g20753/U$1 ( \2842 , \2841 , \684 );
not \mul_17_13_g20201/U$4 ( \2843 , \2842 );
or \mul_17_13_g20201/U$2 ( \2844 , \2840 , \2843 );
not \mul_17_13_g20386/U$3 ( \2845 , \749 );
not \mul_17_13_g20386/U$4 ( \2846 , \746 );
or \mul_17_13_g20386/U$2 ( \2847 , \2845 , \2846 );
nand \mul_17_13_g20429/U$1 ( \2848 , \702 , \2740 );
nand \mul_17_13_g20386/U$1 ( \2849 , \2847 , \2848 );
nand \mul_17_13_g20201/U$1 ( \2850 , \2844 , \2849 );
not \mul_17_13_g20245/U$2 ( \2851 , \2842 );
nand \mul_17_13_g20245/U$1 ( \2852 , \2851 , \2838 );
nand \mul_17_13_g20189/U$1 ( \2853 , \2850 , \2852 );
not \mul_17_13_g20170/U$1 ( \2854 , \2853 );
not \g35931/U$3 ( \2855 , \2854 );
xor \g35842/U$1 ( \2856 , \2761 , \2768 );
xnor \g35842/U$1_r1 ( \2857 , \2856 , \2755 );
not \g35931/U$4 ( \2858 , \2857 );
or \g35931/U$2 ( \2859 , \2855 , \2858 );
xor \mul_17_13_g20141/U$1 ( \2860 , \2790 , \2791 );
xor \mul_17_13_g20141/U$1_r1 ( \2861 , \2860 , \2807 );
nand \g35931/U$1 ( \2862 , \2859 , \2861 );
not \mul_17_13_g20221/U$1 ( \2863 , \2857 );
nand \mul_17_13_g20153/U$1 ( \2864 , \2863 , \2853 );
and \g35930/U$1 ( \2865 , \2862 , \2864 );
nand \mul_17_13_g20051/U$1 ( \2866 , \2833 , \2865 );
and \mul_17_13_g35646/U$1 ( \2867 , \2831 , \2866 );
not \g35909/U$3 ( \2868 , \2867 );
nand \mul_17_13_g20062/U$1 ( \2869 , \903 , \783 );
and \mul_17_13_g20143/U$2 ( \2870 , \2854 , \2863 );
not \mul_17_13_g20143/U$4 ( \2871 , \2854 );
and \mul_17_13_g20143/U$3 ( \2872 , \2871 , \2857 );
nor \mul_17_13_g20143/U$1 ( \2873 , \2870 , \2872 );
not \mul_17_13_g20097/U$3 ( \2874 , \2873 );
not \mul_17_13_g20097/U$4 ( \2875 , \2861 );
and \mul_17_13_g20097/U$2 ( \2876 , \2874 , \2875 );
and \mul_17_13_g20097/U$5 ( \2877 , \2861 , \2873 );
nor \mul_17_13_g20097/U$1 ( \2878 , \2876 , \2877 );
xor \mul_17_13_g20241/U$1 ( \2879 , \2798 , \2797 );
xnor \mul_17_13_g20241/U$1_r1 ( \2880 , \2879 , \2804 );
xor \mul_17_13_g20205/U$4 ( \2881 , \731 , \742 );
and \mul_17_13_g20205/U$3 ( \2882 , \2881 , \751 );
and \mul_17_13_g20205/U$5 ( \2883 , \731 , \742 );
or \mul_17_13_g20205/U$2 ( \2884 , \2882 , \2883 );
not \mul_17_13_g20204/U$1 ( \2885 , \2884 );
xor \mul_17_13_g20106/U$4 ( \2886 , \2880 , \2885 );
xor \mul_17_13_g35812/U$1 ( \2887 , \2838 , \2849 );
xor \mul_17_13_g35812/U$1_r1 ( \2888 , \2887 , \2842 );
and \mul_17_13_g20106/U$3 ( \2889 , \2886 , \2888 );
and \mul_17_13_g20106/U$5 ( \2890 , \2880 , \2885 );
or \mul_17_13_g20106/U$2 ( \2891 , \2889 , \2890 );
nand \mul_17_13_g20064/U$1 ( \2892 , \2878 , \2891 );
xor \mul_17_13_g20106/U$1 ( \2893 , \2880 , \2885 );
xor \mul_17_13_g20106/U$1_r1 ( \2894 , \2893 , \2888 );
not \mul_17_13_g20279/U$1 ( \2895 , \693 );
or \mul_17_13_g20164/U$2 ( \2896 , \752 , \2895 );
nand \mul_17_13_g20164/U$1 ( \2897 , \2896 , \721 );
nand \mul_17_13_g20179/U$1 ( \2898 , \752 , \2895 );
and \mul_17_13_g20155/U$1 ( \2899 , \2897 , \2898 );
nand \mul_17_13_g20089/U$1 ( \2900 , \2894 , \2899 );
nand \mul_17_13_g20032/U$1 ( \2901 , \2869 , \2892 , \2900 , \782 );
not \mul_17_13_g20046/U$3 ( \2902 , \2892 );
nor \mul_17_13_g20091/U$1 ( \2903 , \2894 , \2899 );
not \mul_17_13_g20046/U$4 ( \2904 , \2903 );
or \mul_17_13_g20046/U$2 ( \2905 , \2902 , \2904 );
or \mul_17_13_g20727/U$1 ( \2906 , \2878 , \2891 );
nand \mul_17_13_g20046/U$1 ( \2907 , \2905 , \2906 );
nor \mul_17_13_g20054/U$1 ( \2908 , \2833 , \2865 );
nor \mul_17_13_g20029/U$1 ( \2909 , \2907 , \2908 );
nand \mul_17_13_g20019/U$1 ( \2910 , \2901 , \2909 );
not \g35909/U$4 ( \2911 , \2910 );
or \g35909/U$2 ( \2912 , \2868 , \2911 );
buf \mul_17_13_g20041/U$1 ( \2913 , \2831 );
nor \mul_17_13_g20039/U$1 ( \2914 , \2779 , \2813 );
nand \mul_17_13_g20023/U$1 ( \2915 , \2913 , \2914 );
nand \g35909/U$1 ( \2916 , \2912 , \2915 );
not \mul_17_13_g19988/U$4 ( \2917 , \2916 );
or \mul_17_13_g19988/U$2 ( \2918 , \2817 , \2917 );
not \mul_17_13_g20010/U$1 ( \2919 , \2600 );
not \mul_17_13_g20048/U$1 ( \2920 , \2658 );
nand \mul_17_13_g20000/U$1 ( \2921 , \2919 , \2920 );
not \mul_17_13_g20018/U$3 ( \2922 , \2726 );
not \mul_17_13_g20047/U$1 ( \2923 , \2669 );
not \mul_17_13_g20018/U$4 ( \2924 , \2923 );
or \mul_17_13_g20018/U$2 ( \2925 , \2922 , \2924 );
or \mul_17_13_g20723/U$1 ( \2926 , \2826 , \2830 );
nand \mul_17_13_g20018/U$1 ( \2927 , \2925 , \2926 );
and \mul_17_13_g19991/U$2 ( \2928 , \2921 , \2927 , \2728 );
nor \mul_17_13_g19998/U$1 ( \2929 , \2920 , \2919 );
nor \mul_17_13_g19991/U$1 ( \2930 , \2928 , \2929 );
nand \mul_17_13_g19988/U$1 ( \2931 , \2918 , \2930 );
not \mul_17_13_g19986/U$4 ( \2932 , \2931 );
or \mul_17_13_g19986/U$2 ( \2933 , \2598 , \2932 );
or \mul_17_13_g19986/U$5 ( \2934 , \2931 , \2597 );
nand \mul_17_13_g19986/U$1 ( \2935 , \2933 , \2934 );
not \fopt5203/U$1 ( \2936 , \917 );
nand \g5082/U$1 ( \2937 , \2935 , \2936 );
nand \g35631/U$1 ( \2938 , \2233 , \2937 );
not \g4836/U$3 ( \2939 , \a[15] );
not \g4886/U$1 ( \2940 , \1331 );
not \g4852/U$3 ( \2941 , \2940 );
not \fopt35668/U$1 ( \2942 , \1316 );
not \g4852/U$4 ( \2943 , \2942 );
or \g4852/U$2 ( \2944 , \2941 , \2943 );
not \fopt35677/U$1 ( \2945 , \644 );
nand \g4852/U$1 ( \2946 , \2944 , \2945 );
not \g4836/U$4 ( \2947 , \2946 );
or \g4836/U$2 ( \2948 , \2939 , \2947 );
not \g4896/U$3 ( \2949 , \b[15] );
not \g35819/U$2 ( \2950 , \672 );
nand \g35819/U$1 ( \2951 , \2950 , \1324 );
not \g4896/U$4 ( \2952 , \2951 );
or \g4896/U$2 ( \2953 , \2949 , \2952 );
buf \g5115/U$1 ( \2954 , \1466 );
and \g4906/U$2 ( \2955 , \2954 , \a[15] );
xor \g5026/U$1 ( \2956 , \c[15] , \d[15] );
not \g4931/U$3 ( \2957 , \2956 );
not \g4931/U$4 ( \2958 , \925 );
or \g4931/U$2 ( \2959 , \2957 , \2958 );
not \fopt5215/U$1 ( \2960 , \1220 );
not \fopt5214/U$1 ( \2961 , \2960 );
and \add_15_12_g7226/U$2 ( \2962 , \b[15] , \d[15] );
nor \add_15_12_g7247/U$1 ( \2963 , \b[15] , \d[15] );
nor \add_15_12_g7226/U$1 ( \2964 , \2962 , \2963 );
not \add_15_12_g7137/U$3 ( \2965 , \2964 );
nand \g35881/U$1 ( \2966 , \1487 , \1186 , \1184 );
not \g36001/U$3 ( \2967 , \2966 );
nand \add_15_12_g7199/U$1 ( \2968 , \1209 , \1482 , \1202 );
nor \add_15_12_g7185/U$1 ( \2969 , \1193 , \2968 );
not \g36001/U$4 ( \2970 , \2969 );
or \g36001/U$2 ( \2971 , \2967 , \2970 );
and \add_15_12_g7198/U$1 ( \2972 , \1204 , \1210 , \1200 );
not \add_15_12_g7174/U$3 ( \2973 , \2972 );
not \add_15_12_g7174/U$4 ( \2974 , \1199 );
or \add_15_12_g7174/U$2 ( \2975 , \2973 , \2974 );
or \add_15_12_g7196/U$2 ( \2976 , \1208 , \1194 );
nand \add_15_12_g7196/U$1 ( \2977 , \2976 , \1210 );
nand \add_15_12_g7174/U$1 ( \2978 , \2975 , \2977 );
nand \g36001/U$1 ( \2979 , \2971 , \2978 );
nor \add_15_12_g7254/U$1 ( \2980 , \b[13] , \d[13] );
nor \add_15_12_g7270/U$1 ( \2981 , \b[12] , \d[12] );
nor \add_15_12_g7219/U$1 ( \2982 , \2980 , \2981 );
or \add_15_12_g7274/U$1 ( \2983 , \b[14] , \d[14] );
nand \add_15_12_g7191/U$1 ( \2984 , \2982 , \2983 );
not \add_15_12_g7190/U$1 ( \2985 , \2984 );
nor \add_15_12_g7250/U$1 ( \2986 , \b[11] , \d[11] );
nor \add_15_12_g7249/U$1 ( \2987 , \b[10] , \d[10] );
nor \add_15_12_g7222/U$1 ( \2988 , \2986 , \2987 );
nor \add_15_12_g7252/U$1 ( \2989 , \b[8] , \d[8] );
nor \add_15_12_g7271/U$1 ( \2990 , \b[9] , \d[9] );
nor \add_15_12_g7221/U$1 ( \2991 , \2989 , \2990 );
and \add_15_12_g7192/U$1 ( \2992 , \2988 , \2991 );
and \add_15_12_g7149/U$2 ( \2993 , \2979 , \2985 , \2992 );
nand \add_15_12_g7243/U$1 ( \2994 , \b[8] , \d[8] );
or \add_15_12_g7194/U$2 ( \2995 , \2990 , \2994 );
nand \add_15_12_g7255/U$1 ( \2996 , \b[9] , \d[9] );
nand \add_15_12_g7194/U$1 ( \2997 , \2995 , \2996 );
not \add_15_12_g7180/U$3 ( \2998 , \2997 );
not \add_15_12_g7180/U$4 ( \2999 , \2988 );
or \add_15_12_g7180/U$2 ( \3000 , \2998 , \2999 );
not \add_15_12_g7197/U$3 ( \3001 , \2986 );
nand \add_15_12_g7237/U$1 ( \3002 , \b[10] , \d[10] );
not \add_15_12_g7197/U$4 ( \3003 , \3002 );
and \add_15_12_g7197/U$2 ( \3004 , \3001 , \3003 );
and \add_15_12_g7264/U$1 ( \3005 , \b[11] , \d[11] );
nor \add_15_12_g7197/U$1 ( \3006 , \3004 , \3005 );
nand \add_15_12_g7180/U$1 ( \3007 , \3000 , \3006 );
not \add_15_12_g7179/U$1 ( \3008 , \3007 );
or \add_15_12_g7168/U$2 ( \3009 , \3008 , \2984 );
nand \add_15_12_g7253/U$1 ( \3010 , \b[12] , \d[12] );
or \add_15_12_g7193/U$2 ( \3011 , \2980 , \3010 );
nand \add_15_12_g7263/U$1 ( \3012 , \b[13] , \d[13] );
nand \add_15_12_g7193/U$1 ( \3013 , \3011 , \3012 );
and \add_15_12_g7178/U$2 ( \3014 , \3013 , \2983 );
and \add_15_12_g7246/U$1 ( \3015 , \b[14] , \d[14] );
nor \add_15_12_g7178/U$1 ( \3016 , \3014 , \3015 );
nand \add_15_12_g7168/U$1 ( \3017 , \3009 , \3016 );
nor \add_15_12_g7149/U$1 ( \3018 , \2993 , \3017 );
not \add_15_12_g7137/U$4 ( \3019 , \3018 );
or \add_15_12_g7137/U$2 ( \3020 , \2965 , \3019 );
or \add_15_12_g7137/U$5 ( \3021 , \3018 , \2964 );
nand \add_15_12_g7137/U$1 ( \3022 , \3020 , \3021 );
and \g4948/U$2 ( \3023 , \2961 , \3022 );
and \add_14_12_g7226/U$2 ( \3024 , \a[15] , \c[15] );
nor \add_14_12_g7247/U$1 ( \3025 , \a[15] , \c[15] );
nor \add_14_12_g7226/U$1 ( \3026 , \3024 , \3025 );
not \add_14_12_g7137/U$3 ( \3027 , \3026 );
nand \g35877/U$1 ( \3028 , \1501 , \1249 , \1247 );
not \g35876/U$3 ( \3029 , \3028 );
nand \add_14_12_g7199/U$1 ( \3030 , \1272 , \1496 , \1265 );
nor \add_14_12_g7185/U$1 ( \3031 , \1256 , \3030 );
not \g35876/U$4 ( \3032 , \3031 );
or \g35876/U$2 ( \3033 , \3029 , \3032 );
and \add_14_12_g7198/U$1 ( \3034 , \1267 , \1273 , \1263 );
not \add_14_12_g7174/U$3 ( \3035 , \3034 );
not \add_14_12_g7174/U$4 ( \3036 , \1262 );
or \add_14_12_g7174/U$2 ( \3037 , \3035 , \3036 );
or \add_14_12_g7196/U$2 ( \3038 , \1271 , \1257 );
nand \add_14_12_g7196/U$1 ( \3039 , \3038 , \1273 );
nand \add_14_12_g7174/U$1 ( \3040 , \3037 , \3039 );
nand \g35876/U$1 ( \3041 , \3033 , \3040 );
nor \add_14_12_g7254/U$1 ( \3042 , \a[13] , \c[13] );
nor \add_14_12_g7270/U$1 ( \3043 , \a[12] , \c[12] );
nor \add_14_12_g7219/U$1 ( \3044 , \3042 , \3043 );
or \add_14_12_g7274/U$1 ( \3045 , \a[14] , \c[14] );
nand \add_14_12_g7191/U$1 ( \3046 , \3044 , \3045 );
not \add_14_12_g7190/U$1 ( \3047 , \3046 );
nor \add_14_12_g7250/U$1 ( \3048 , \a[11] , \c[11] );
nor \add_14_12_g7249/U$1 ( \3049 , \a[10] , \c[10] );
nor \add_14_12_g7222/U$1 ( \3050 , \3048 , \3049 );
nor \add_14_12_g7252/U$1 ( \3051 , \a[8] , \c[8] );
nor \add_14_12_g7271/U$1 ( \3052 , \a[9] , \c[9] );
nor \add_14_12_g7221/U$1 ( \3053 , \3051 , \3052 );
and \add_14_12_g7192/U$1 ( \3054 , \3050 , \3053 );
and \add_14_12_g7149/U$2 ( \3055 , \3041 , \3047 , \3054 );
nand \add_14_12_g7243/U$1 ( \3056 , \a[8] , \c[8] );
or \add_14_12_g7194/U$2 ( \3057 , \3052 , \3056 );
nand \add_14_12_g7255/U$1 ( \3058 , \a[9] , \c[9] );
nand \add_14_12_g7194/U$1 ( \3059 , \3057 , \3058 );
not \add_14_12_g7180/U$3 ( \3060 , \3059 );
not \add_14_12_g7180/U$4 ( \3061 , \3050 );
or \add_14_12_g7180/U$2 ( \3062 , \3060 , \3061 );
not \add_14_12_g7197/U$3 ( \3063 , \3048 );
nand \add_14_12_g7237/U$1 ( \3064 , \a[10] , \c[10] );
not \add_14_12_g7197/U$4 ( \3065 , \3064 );
and \add_14_12_g7197/U$2 ( \3066 , \3063 , \3065 );
and \add_14_12_g7264/U$1 ( \3067 , \a[11] , \c[11] );
nor \add_14_12_g7197/U$1 ( \3068 , \3066 , \3067 );
nand \add_14_12_g7180/U$1 ( \3069 , \3062 , \3068 );
not \add_14_12_g7179/U$1 ( \3070 , \3069 );
or \add_14_12_g7168/U$2 ( \3071 , \3070 , \3046 );
nand \add_14_12_g7253/U$1 ( \3072 , \a[12] , \c[12] );
or \add_14_12_g7193/U$2 ( \3073 , \3042 , \3072 );
nand \add_14_12_g7263/U$1 ( \3074 , \a[13] , \c[13] );
nand \add_14_12_g7193/U$1 ( \3075 , \3073 , \3074 );
and \add_14_12_g7178/U$2 ( \3076 , \3075 , \3045 );
and \add_14_12_g7246/U$1 ( \3077 , \a[14] , \c[14] );
nor \add_14_12_g7178/U$1 ( \3078 , \3076 , \3077 );
nand \add_14_12_g7168/U$1 ( \3079 , \3071 , \3078 );
nor \add_14_12_g7149/U$1 ( \3080 , \3055 , \3079 );
not \add_14_12_g7137/U$4 ( \3081 , \3080 );
or \add_14_12_g7137/U$2 ( \3082 , \3027 , \3081 );
or \add_14_12_g7137/U$5 ( \3083 , \3080 , \3026 );
nand \add_14_12_g7137/U$1 ( \3084 , \3082 , \3083 );
not \g4975/U$3 ( \3085 , \3084 );
not \g5103/U$1 ( \3086 , \1232 );
not \g5100/U$1 ( \3087 , \3086 );
not \g4975/U$4 ( \3088 , \3087 );
or \g4975/U$2 ( \3089 , \3085 , \3088 );
and \g35870/U$2 ( \3090 , \1282 , \d[15] );
and \g35870/U$3 ( \3091 , \1435 , \c[15] );
nor \g35870/U$1 ( \3092 , \3090 , \3091 );
nand \g4975/U$1 ( \3093 , \3089 , \3092 );
nor \g4948/U$1 ( \3094 , \3023 , \3093 );
nand \g4931/U$1 ( \3095 , \2959 , \3094 );
nor \g4906/U$1 ( \3096 , \2955 , \3095 );
nand \g4896/U$1 ( \3097 , \2953 , \3096 );
not \g4979/U$3 ( \3098 , \d[15] );
not \g4979/U$4 ( \3099 , \1457 );
or \g4979/U$2 ( \3100 , \3098 , \3099 );
not \fopt35666/U$1 ( \3101 , \1316 );
not \fopt35665/U$1 ( \3102 , \3101 );
nand \g35860/U$1 ( \3103 , \3102 , \b[15] , \c[15] );
nand \g4979/U$1 ( \3104 , \3100 , \3103 );
nor \g4870/U$1 ( \3105 , \3097 , \3104 );
nand \g4836/U$1 ( \3106 , \2948 , \3105 );
nor \g4815/U$1 ( \3107 , \2938 , \3106 );
not \g4814/U$1 ( \3108 , \3107 );
not \g4837/U$3 ( \3109 , \a[11] );
not \g4851/U$3 ( \3110 , \2940 );
not \g4851/U$4 ( \3111 , \3101 );
or \g4851/U$2 ( \3112 , \3110 , \3111 );
not \fopt35673/U$1 ( \3113 , \644 );
nand \g4851/U$1 ( \3114 , \3112 , \3113 );
not \g4837/U$4 ( \3115 , \3114 );
or \g4837/U$2 ( \3116 , \3109 , \3115 );
not \g35934/U$3 ( \3117 , \d[11] );
not \g35934/U$4 ( \3118 , \1450 );
or \g35934/U$2 ( \3119 , \3117 , \3118 );
nand \g35935/U$1 ( \3120 , \1316 , \b[11] , \c[11] );
nand \g35934/U$1 ( \3121 , \3119 , \3120 );
not \g4897/U$3 ( \3122 , \b[11] );
not \g5252/U$2 ( \3123 , \671 );
nand \g5252/U$1 ( \3124 , \3123 , \1324 );
not \g4897/U$4 ( \3125 , \3124 );
or \g4897/U$2 ( \3126 , \3122 , \3125 );
not \g4910/U$3 ( \3127 , \a[11] );
not \g4910/U$4 ( \3128 , \672 );
or \g4910/U$2 ( \3129 , \3127 , \3128 );
xor \g5028/U$1 ( \3130 , \c[11] , \d[11] );
and \g4932/U$2 ( \3131 , \3130 , \925 );
nor \add_15_12_g7202/U$1 ( \3132 , \2986 , \3005 );
not \add_15_12_g7138/U$3 ( \3133 , \3132 );
not \add_15_12_g7248/U$1 ( \3134 , \2987 );
and \g35879/U$2 ( \3135 , \2979 , \2991 , \3134 );
not \add_15_12_g7177/U$3 ( \3136 , \3134 );
not \add_15_12_g7177/U$4 ( \3137 , \2997 );
or \add_15_12_g7177/U$2 ( \3138 , \3136 , \3137 );
nand \add_15_12_g7177/U$1 ( \3139 , \3138 , \3002 );
nor \g35879/U$1 ( \3140 , \3135 , \3139 );
not \add_15_12_g7138/U$4 ( \3141 , \3140 );
or \add_15_12_g7138/U$2 ( \3142 , \3133 , \3141 );
or \add_15_12_g7138/U$5 ( \3143 , \3140 , \3132 );
nand \add_15_12_g7138/U$1 ( \3144 , \3142 , \3143 );
not \g4947/U$3 ( \3145 , \3144 );
not \g4947/U$4 ( \3146 , \2961 );
or \g4947/U$2 ( \3147 , \3145 , \3146 );
nor \add_14_12_g7202/U$1 ( \3148 , \3048 , \3067 );
not \add_14_12_g7138/U$3 ( \3149 , \3148 );
not \add_14_12_g7248/U$1 ( \3150 , \3049 );
and \g35875/U$2 ( \3151 , \3041 , \3053 , \3150 );
not \add_14_12_g7177/U$3 ( \3152 , \3150 );
not \add_14_12_g7177/U$4 ( \3153 , \3059 );
or \add_14_12_g7177/U$2 ( \3154 , \3152 , \3153 );
nand \add_14_12_g7177/U$1 ( \3155 , \3154 , \3064 );
nor \g35875/U$1 ( \3156 , \3151 , \3155 );
not \add_14_12_g7138/U$4 ( \3157 , \3156 );
or \add_14_12_g7138/U$2 ( \3158 , \3149 , \3157 );
or \add_14_12_g7138/U$5 ( \3159 , \3156 , \3148 );
nand \add_14_12_g7138/U$1 ( \3160 , \3158 , \3159 );
and \g4973/U$2 ( \3161 , \3087 , \3160 );
not \g5009/U$3 ( \3162 , \d[11] );
not \g5009/U$4 ( \3163 , \1282 );
or \g5009/U$2 ( \3164 , \3162 , \3163 );
nand \g5077/U$1 ( \3165 , \1435 , \c[11] );
nand \g5009/U$1 ( \3166 , \3164 , \3165 );
nor \g4973/U$1 ( \3167 , \3161 , \3166 );
nand \g4947/U$1 ( \3168 , \3147 , \3167 );
nor \g4932/U$1 ( \3169 , \3131 , \3168 );
nand \g4910/U$1 ( \3170 , \3129 , \3169 );
not \g4909/U$1 ( \3171 , \3170 );
nand \g4897/U$1 ( \3172 , \3126 , \3171 );
nor \g4869/U$1 ( \3173 , \3121 , \3172 );
nand \g4837/U$1 ( \3174 , \3116 , \3173 );
not \g5004/U$3 ( \3175 , \1529 );
not \mul_16_12_g19994/U$2 ( \3176 , \2211 );
nand \mul_16_12_g19994/U$1 ( \3177 , \3176 , \2112 );
not \mul_16_12_g19979/U$3 ( \3178 , \3177 );
not \mul_16_12_g19985/U$3 ( \3179 , \2206 );
not \mul_16_12_g20002/U$3 ( \3180 , \2173 );
not \mul_16_12_g20002/U$4 ( \3181 , \2120 );
or \mul_16_12_g20002/U$2 ( \3182 , \3180 , \3181 );
not \mul_16_12_g20025/U$1 ( \3183 , \2191 );
nand \mul_16_12_g20002/U$1 ( \3184 , \3182 , \3183 );
not \mul_16_12_g19985/U$4 ( \3185 , \3184 );
or \mul_16_12_g19985/U$2 ( \3186 , \3179 , \3185 );
not \mul_16_12_g20038/U$1 ( \3187 , \2187 );
nand \mul_16_12_g19985/U$1 ( \3188 , \3186 , \3187 );
not \mul_16_12_g19979/U$4 ( \3189 , \3188 );
or \mul_16_12_g19979/U$2 ( \3190 , \3178 , \3189 );
or \mul_16_12_g19979/U$5 ( \3191 , \3188 , \3177 );
nand \mul_16_12_g19979/U$1 ( \3192 , \3190 , \3191 );
not \g5004/U$4 ( \3193 , \3192 );
or \g5004/U$2 ( \3194 , \3175 , \3193 );
not \g35623/U$2 ( \3195 , \2814 );
nor \g35623/U$1 ( \3196 , \3195 , \2914 );
not \mul_17_13_g20001/U$3 ( \3197 , \2866 );
not \g35648/U$2 ( \3198 , \2907 );
nand \g35648/U$1 ( \3199 , \3198 , \2901 );
not \mul_17_13_g20001/U$4 ( \3200 , \3199 );
or \mul_17_13_g20001/U$2 ( \3201 , \3197 , \3200 );
not \mul_17_13_g20052/U$1 ( \3202 , \2908 );
nand \mul_17_13_g20001/U$1 ( \3203 , \3201 , \3202 );
xor \g36024/U$1 ( \3204 , \3196 , \3203 );
nand \g5058/U$1 ( \3205 , \3204 , \2936 );
nand \g5004/U$1 ( \3206 , \3194 , \3205 );
nor \g4817/U$1 ( \3207 , \3174 , \3206 );
not \g4816/U$1 ( \3208 , \3207 );
not \g4818/U$3 ( \3209 , \a[6] );
not \g4818/U$4 ( \3210 , \3114 );
or \g4818/U$2 ( \3211 , \3209 , \3210 );
and \g36006/U$2 ( \3212 , \d[6] , \1342 );
nand \g35937/U$1 ( \3213 , \1316 , \b[6] , \c[6] );
or \g5067/U$1 ( \3214 , \a[6] , \b[6] );
nand \g4/U$1 ( \3215 , \3214 , \672 );
xor \g5027/U$1 ( \3216 , \c[6] , \d[6] );
not \g4890/U$3 ( \3217 , \3216 );
not \g4890/U$4 ( \3218 , \1320 );
or \g4890/U$2 ( \3219 , \3217 , \3218 );
not \mul_16_12_g20689/U$2 ( \3220 , \1090 );
nand \mul_16_12_g20689/U$1 ( \3221 , \3220 , \1095 );
not \mul_16_12_g20055/U$3 ( \3222 , \3221 );
nand \mul_16_12_g20694/U$1 ( \3223 , \1097 , \1008 );
not \mul_16_12_g20055/U$4 ( \3224 , \3223 );
or \mul_16_12_g20055/U$2 ( \3225 , \3222 , \3224 );
or \mul_16_12_g20055/U$5 ( \3226 , \3223 , \3221 );
nand \mul_16_12_g20055/U$1 ( \3227 , \3225 , \3226 );
and \g4908/U$2 ( \3228 , \3227 , \1353 );
not \add_15_12_g7205/U$1 ( \3229 , \1193 );
not \add_15_12_g7157/U$3 ( \3230 , \3229 );
not \add_15_12_g7157/U$4 ( \3231 , \1189 );
or \add_15_12_g7157/U$2 ( \3232 , \3230 , \3231 );
not \add_15_12_g7187/U$1 ( \3233 , \1201 );
nand \add_15_12_g7157/U$1 ( \3234 , \3232 , \3233 );
nand \add_15_12_g7214/U$1 ( \3235 , \1202 , \1204 );
xnor \add_15_12_g7146/U$1 ( \3236 , \3234 , \3235 );
not \g4924/U$3 ( \3237 , \3236 );
not \g4924/U$4 ( \3238 , \1220 );
or \g4924/U$2 ( \3239 , \3237 , \3238 );
not \add_14_12_g7205/U$1 ( \3240 , \1256 );
not \add_14_12_g7157/U$3 ( \3241 , \3240 );
not \add_14_12_g7157/U$4 ( \3242 , \1252 );
or \add_14_12_g7157/U$2 ( \3243 , \3241 , \3242 );
not \add_14_12_g7187/U$1 ( \3244 , \1264 );
nand \add_14_12_g7157/U$1 ( \3245 , \3243 , \3244 );
nand \add_14_12_g7214/U$1 ( \3246 , \1265 , \1267 );
xnor \add_14_12_g7146/U$1 ( \3247 , \3245 , \3246 );
not \g4946/U$3 ( \3248 , \3247 );
not \g4946/U$4 ( \3249 , \1232 );
or \g4946/U$2 ( \3250 , \3248 , \3249 );
and \g4972/U$2 ( \3251 , \1280 , \d[6] );
not \g5007/U$3 ( \3252 , \c[6] );
not \g5007/U$4 ( \3253 , \1287 );
or \g5007/U$2 ( \3254 , \3252 , \3253 );
nand \g5034/U$1 ( \3255 , \1293 , \b[6] );
nand \g5007/U$1 ( \3256 , \3254 , \3255 );
nor \g4972/U$1 ( \3257 , \3251 , \3256 );
nand \g4946/U$1 ( \3258 , \3250 , \3257 );
not \g4945/U$1 ( \3259 , \3258 );
nand \g4924/U$1 ( \3260 , \3239 , \3259 );
nor \g4908/U$1 ( \3261 , \3228 , \3260 );
nand \g4890/U$1 ( \3262 , \3219 , \3261 );
not \g35354/U$2 ( \3263 , \916 );
not \mul_17_13_g20128/U$2 ( \3264 , \895 );
nand \mul_17_13_g20128/U$1 ( \3265 , \3264 , \901 );
nand \mul_17_13_g20086/U$1 ( \3266 , \880 , \899 );
xor \g35355/U$1 ( \3267 , \3265 , \3266 );
nor \g35354/U$1 ( \3268 , \3263 , \3267 );
nor \g4879/U$1 ( \3269 , \3262 , \3268 );
nand \g36007/U$1 ( \3270 , \3213 , \3215 , \3269 );
nor \g36006/U$1 ( \3271 , \3212 , \3270 );
nand \g4818/U$1 ( \3272 , \3211 , \3271 );
not \mul_17_13_g19994/U$2 ( \3273 , \2929 );
nand \mul_17_13_g19994/U$1 ( \3274 , \3273 , \2921 );
not \mul_17_13_g19987/U$3 ( \3275 , \3274 );
not \mul_17_13_g20016/U$1 ( \3276 , \2815 );
not \mul_17_13_g19990/U$3 ( \3277 , \3276 );
not \mul_17_13_g19990/U$4 ( \3278 , \2916 );
or \mul_17_13_g19990/U$2 ( \3279 , \3277 , \3278 );
buf \fopt35596/U$1 ( \3280 , \2728 );
nand \mul_17_13_g20007/U$1 ( \3281 , \2927 , \3280 );
nand \mul_17_13_g19990/U$1 ( \3282 , \3279 , \3281 );
not \mul_17_13_g19987/U$4 ( \3283 , \3282 );
or \mul_17_13_g19987/U$2 ( \3284 , \3275 , \3283 );
or \mul_17_13_g19987/U$5 ( \3285 , \3282 , \3274 );
nand \mul_17_13_g19987/U$1 ( \3286 , \3284 , \3285 );
nand \g5036/U$1 ( \3287 , \3286 , \2936 );
nand \g4848/U$1 ( \3288 , \a[14] , \1338 );
or \g5061/U$1 ( \3289 , \a[14] , \d[14] );
not \g4959/U$3 ( \3290 , \3289 );
not \g4959/U$4 ( \3291 , \1457 );
or \g4959/U$2 ( \3292 , \3290 , \3291 );
nand \g35861/U$1 ( \3293 , \3102 , \b[14] , \c[14] );
nand \g4959/U$1 ( \3294 , \3292 , \3293 );
not \g4895/U$3 ( \3295 , \b[14] );
not \g4895/U$4 ( \3296 , \2951 );
or \g4895/U$2 ( \3297 , \3295 , \3296 );
and \g4905/U$2 ( \3298 , \a[14] , \1351 );
and \g5023/U$2 ( \3299 , \d[14] , \c[14] );
not \g5023/U$4 ( \3300 , \d[14] );
not \g5158/U$1 ( \3301 , \c[14] );
and \g5023/U$3 ( \3302 , \3300 , \3301 );
nor \g5023/U$1 ( \3303 , \3299 , \3302 );
not \g4930/U$3 ( \3304 , \3303 );
buf \fopt5182/U$1 ( \3305 , \1320 );
not \g4930/U$4 ( \3306 , \3305 );
or \g4930/U$2 ( \3307 , \3304 , \3306 );
not \add_15_12_g7281/U$2 ( \3308 , \2983 );
nor \add_15_12_g7281/U$1 ( \3309 , \3308 , \3015 );
not \add_15_12_g7141/U$3 ( \3310 , \3309 );
and \add_15_12_g7153/U$2 ( \3311 , \2979 , \2992 , \2982 );
not \add_15_12_g7164/U$2 ( \3312 , \3013 );
nand \add_15_12_g7171/U$1 ( \3313 , \3007 , \2982 );
nand \add_15_12_g7164/U$1 ( \3314 , \3312 , \3313 );
nor \add_15_12_g7153/U$1 ( \3315 , \3311 , \3314 );
not \add_15_12_g7141/U$4 ( \3316 , \3315 );
or \add_15_12_g7141/U$2 ( \3317 , \3310 , \3316 );
or \add_15_12_g7141/U$5 ( \3318 , \3315 , \3309 );
nand \add_15_12_g7141/U$1 ( \3319 , \3317 , \3318 );
and \g4944/U$2 ( \3320 , \2961 , \3319 );
not \add_14_12_g7281/U$2 ( \3321 , \3045 );
nor \add_14_12_g7281/U$1 ( \3322 , \3321 , \3077 );
not \add_14_12_g7141/U$3 ( \3323 , \3322 );
and \add_14_12_g7153/U$2 ( \3324 , \3041 , \3054 , \3044 );
not \add_14_12_g7164/U$2 ( \3325 , \3075 );
nand \add_14_12_g7171/U$1 ( \3326 , \3069 , \3044 );
nand \add_14_12_g7164/U$1 ( \3327 , \3325 , \3326 );
nor \add_14_12_g7153/U$1 ( \3328 , \3324 , \3327 );
not \add_14_12_g7141/U$4 ( \3329 , \3328 );
or \add_14_12_g7141/U$2 ( \3330 , \3323 , \3329 );
or \add_14_12_g7141/U$5 ( \3331 , \3328 , \3322 );
nand \add_14_12_g7141/U$1 ( \3332 , \3330 , \3331 );
not \g4970/U$3 ( \3333 , \3332 );
not \g4970/U$4 ( \3334 , \3087 );
or \g4970/U$2 ( \3335 , \3333 , \3334 );
not \g5006/U$3 ( \3336 , \1323 );
not \g5006/U$4 ( \3337 , \3301 );
and \g5006/U$2 ( \3338 , \3336 , \3337 );
and \g5006/U$5 ( \3339 , \1282 , \d[14] );
nor \g5006/U$1 ( \3340 , \3338 , \3339 );
nand \g4970/U$1 ( \3341 , \3335 , \3340 );
nor \g4944/U$1 ( \3342 , \3320 , \3341 );
nand \g4930/U$1 ( \3343 , \3307 , \3342 );
nor \g4905/U$1 ( \3344 , \3298 , \3343 );
nand \g4895/U$1 ( \3345 , \3297 , \3344 );
nor \g4872/U$1 ( \3346 , \3294 , \3345 );
not \mul_16_12_g20028/U$1 ( \3347 , \1953 );
not \mul_16_12_g19972/U$3 ( \3348 , \3347 );
not \mul_16_12_g19983/U$1 ( \3349 , \1908 );
not \mul_16_12_g19972/U$4 ( \3350 , \3349 );
or \mul_16_12_g19972/U$2 ( \3351 , \3348 , \3350 );
or \mul_16_12_g19972/U$5 ( \3352 , \3349 , \3347 );
nand \mul_16_12_g19972/U$1 ( \3353 , \3351 , \3352 );
not \mul_16_12_g19967/U$3 ( \3354 , \3353 );
not \mul_16_12_g19995/U$1 ( \3355 , \2113 );
not \mul_16_12_g19973/U$3 ( \3356 , \3355 );
not \mul_16_12_g19973/U$4 ( \3357 , \2213 );
or \mul_16_12_g19973/U$2 ( \3358 , \3356 , \3357 );
nand \mul_16_12_g19986/U$1 ( \3359 , \2223 , \2031 );
nand \mul_16_12_g19973/U$1 ( \3360 , \3358 , \3359 );
not \mul_16_12_g19967/U$4 ( \3361 , \3360 );
or \mul_16_12_g19967/U$2 ( \3362 , \3354 , \3361 );
or \mul_16_12_g19967/U$5 ( \3363 , \3353 , \3360 );
nand \mul_16_12_g19967/U$1 ( \3364 , \3362 , \3363 );
nand \g5065/U$1 ( \3365 , \3364 , \1529 );
nand \g4819/U$1 ( \3366 , \3287 , \3288 , \3346 , \3365 );
not \g4820/U$3 ( \3367 , \a[2] );
not \g4820/U$4 ( \3368 , \3114 );
or \g4820/U$2 ( \3369 , \3367 , \3368 );
not \g5234/U$3 ( \3370 , \d[2] );
not \g5234/U$4 ( \3371 , \1457 );
or \g5234/U$2 ( \3372 , \3370 , \3371 );
not \fopt35667/U$1 ( \3373 , \2942 );
and \g5059/U$1 ( \3374 , \b[2] , \c[2] );
and \g5235/U$2 ( \3375 , \3373 , \3374 );
or \g5055/U$1 ( \3376 , \a[2] , \b[2] );
not \g4859/U$3 ( \3377 , \3376 );
not \g4859/U$4 ( \3378 , \1351 );
or \g4859/U$2 ( \3379 , \3377 , \3378 );
xor \g5019/U$1 ( \3380 , \c[2] , \d[2] );
not \g4893/U$3 ( \3381 , \3380 );
not \g4893/U$4 ( \3382 , \1383 );
or \g4893/U$2 ( \3383 , \3381 , \3382 );
not \mul_16_12_g20243/U$3 ( \3384 , \1046 );
not \mul_16_12_g20284/U$2 ( \3385 , \1049 );
nor \mul_16_12_g20284/U$1 ( \3386 , \3385 , \1037 );
not \mul_16_12_g20243/U$4 ( \3387 , \3386 );
or \mul_16_12_g20243/U$2 ( \3388 , \3384 , \3387 );
or \mul_16_12_g20243/U$5 ( \3389 , \3386 , \1046 );
nand \mul_16_12_g20243/U$1 ( \3390 , \3388 , \3389 );
and \g4900/U$2 ( \3391 , \1478 , \3390 );
nand \add_15_12_g7209/U$1 ( \3392 , \1486 , \1186 );
not \add_15_12_g7169/U$3 ( \3393 , \3392 );
not \add_15_12_g7169/U$4 ( \3394 , \1181 );
or \add_15_12_g7169/U$2 ( \3395 , \3393 , \3394 );
or \add_15_12_g7169/U$5 ( \3396 , \1181 , \3392 );
nand \add_15_12_g7169/U$1 ( \3397 , \3395 , \3396 );
not \g4918/U$3 ( \3398 , \3397 );
not \g4918/U$4 ( \3399 , \1220 );
or \g4918/U$2 ( \3400 , \3398 , \3399 );
nand \add_14_12_g7209/U$1 ( \3401 , \1500 , \1249 );
not \add_14_12_g7169/U$3 ( \3402 , \3401 );
not \add_14_12_g7169/U$4 ( \3403 , \1244 );
or \add_14_12_g7169/U$2 ( \3404 , \3402 , \3403 );
or \add_14_12_g7169/U$5 ( \3405 , \1244 , \3401 );
nand \add_14_12_g7169/U$1 ( \3406 , \3404 , \3405 );
not \g4937/U$3 ( \3407 , \3406 );
not \g4937/U$4 ( \3408 , \1232 );
or \g4937/U$2 ( \3409 , \3407 , \3408 );
and \g4960/U$2 ( \3410 , \1282 , \d[2] );
not \g4996/U$3 ( \3411 , \c[2] );
not \g4996/U$4 ( \3412 , \1287 );
or \g4996/U$2 ( \3413 , \3411 , \3412 );
nand \g5038/U$1 ( \3414 , \1293 , \b[2] );
nand \g4996/U$1 ( \3415 , \3413 , \3414 );
nor \g4960/U$1 ( \3416 , \3410 , \3415 );
nand \g4937/U$1 ( \3417 , \3409 , \3416 );
not \g4936/U$1 ( \3418 , \3417 );
nand \g4918/U$1 ( \3419 , \3400 , \3418 );
nor \g4900/U$1 ( \3420 , \3391 , \3419 );
nand \g4893/U$1 ( \3421 , \3383 , \3420 );
not \g35352/U$2 ( \3422 , \916 );
not \mul_17_13_g20292/U$2 ( \3423 , \863 );
nor \mul_17_13_g20292/U$1 ( \3424 , \3423 , \851 );
xor \g35353/U$1 ( \3425 , \861 , \3424 );
nor \g35352/U$1 ( \3426 , \3422 , \3425 );
nor \g4883/U$1 ( \3427 , \3421 , \3426 );
nand \g4859/U$1 ( \3428 , \3379 , \3427 );
nor \g5235/U$1 ( \3429 , \3375 , \3428 );
nand \g5234/U$1 ( \3430 , \3372 , \3429 );
not \g10/U$1 ( \3431 , \3430 );
nand \g4820/U$1 ( \3432 , \3369 , \3431 );
not \g4821/U$3 ( \3433 , \a[10] );
not \g4821/U$4 ( \3434 , \2946 );
or \g4821/U$2 ( \3435 , \3433 , \3434 );
not \g4912/U$3 ( \3436 , \a[10] );
not \g4912/U$4 ( \3437 , \1466 );
or \g4912/U$2 ( \3438 , \3436 , \3437 );
xor \g5031/U$1 ( \3439 , \c[10] , \d[10] );
and \g4933/U$2 ( \3440 , \3305 , \3439 );
and \add_15_12_g7204/U$1 ( \3441 , \3134 , \3002 );
not \add_15_12_g7139/U$3 ( \3442 , \3441 );
and \add_15_12_g7147/U$2 ( \3443 , \2979 , \2991 );
nor \add_15_12_g7147/U$1 ( \3444 , \3443 , \2997 );
not \add_15_12_g7139/U$4 ( \3445 , \3444 );
or \add_15_12_g7139/U$2 ( \3446 , \3442 , \3445 );
or \add_15_12_g7139/U$5 ( \3447 , \3444 , \3441 );
nand \add_15_12_g7139/U$1 ( \3448 , \3446 , \3447 );
not \g4951/U$3 ( \3449 , \3448 );
not \g4951/U$4 ( \3450 , \2961 );
or \g4951/U$2 ( \3451 , \3449 , \3450 );
and \add_14_12_g7204/U$1 ( \3452 , \3150 , \3064 );
not \add_14_12_g7139/U$3 ( \3453 , \3452 );
and \add_14_12_g7147/U$2 ( \3454 , \3041 , \3053 );
nor \add_14_12_g7147/U$1 ( \3455 , \3454 , \3059 );
not \add_14_12_g7139/U$4 ( \3456 , \3455 );
or \add_14_12_g7139/U$2 ( \3457 , \3453 , \3456 );
or \add_14_12_g7139/U$5 ( \3458 , \3455 , \3452 );
nand \add_14_12_g7139/U$1 ( \3459 , \3457 , \3458 );
and \g4978/U$2 ( \3460 , \3087 , \3459 );
not \g5015/U$3 ( \3461 , \d[10] );
not \g5015/U$4 ( \3462 , \1282 );
or \g5015/U$2 ( \3463 , \3461 , \3462 );
nand \g5090/U$1 ( \3464 , \1435 , \c[10] );
nand \g5015/U$1 ( \3465 , \3463 , \3464 );
nor \g4978/U$1 ( \3466 , \3460 , \3465 );
nand \g4951/U$1 ( \3467 , \3451 , \3466 );
nor \g4933/U$1 ( \3468 , \3440 , \3467 );
nand \g4912/U$1 ( \3469 , \3438 , \3468 );
not \g4873/U$2 ( \3470 , \3469 );
not \mul_17_13_g20035/U$2 ( \3471 , \2908 );
nand \mul_17_13_g20035/U$1 ( \3472 , \3471 , \2866 );
xnor \g35460/U$1 ( \3473 , \3472 , \3199 );
and \g5012/U$2 ( \3474 , \3473 , \2936 );
nand \mul_16_12_g20023/U$1 ( \3475 , \3187 , \2206 );
xnor \mul_16_12_g20687/U$1 ( \3476 , \3184 , \3475 );
and \g5012/U$3 ( \3477 , \3476 , \1529 );
nor \g5012/U$1 ( \3478 , \3474 , \3477 );
nand \g35866/U$1 ( \3479 , \3102 , \b[10] , \c[10] );
nand \g4873/U$1 ( \3480 , \3470 , \3478 , \3479 );
not \g4982/U$3 ( \3481 , \d[10] );
not \g4982/U$4 ( \3482 , \1342 );
or \g4982/U$2 ( \3483 , \3481 , \3482 );
nand \g4983/U$1 ( \3484 , \2951 , \b[10] );
nand \g4982/U$1 ( \3485 , \3483 , \3484 );
nor \g4863/U$1 ( \3486 , \3480 , \3485 );
nand \g4821/U$1 ( \3487 , \3435 , \3486 );
nor \mul_16_12_g20003/U$1 ( \3488 , \2030 , \1962 );
not \mul_16_12_g19991/U$2 ( \3489 , \3488 );
nand \mul_16_12_g19991/U$1 ( \3490 , \3489 , \2031 );
not \mul_16_12_g19969/U$3 ( \3491 , \3490 );
not \mul_16_12_g19978/U$3 ( \3492 , \2193 );
and \mul_16_12_g19984/U$1 ( \3493 , \2205 , \2112 , \2206 );
not \mul_16_12_g19978/U$4 ( \3494 , \3493 );
or \mul_16_12_g19978/U$2 ( \3495 , \3492 , \3494 );
and \g35442/U$2 ( \3496 , \2205 , \2211 );
nor \g35442/U$1 ( \3497 , \3496 , \2221 );
nand \mul_16_12_g19978/U$1 ( \3498 , \3495 , \3497 );
not \mul_16_12_g19969/U$4 ( \3499 , \3498 );
or \mul_16_12_g19969/U$2 ( \3500 , \3491 , \3499 );
or \mul_16_12_g19969/U$5 ( \3501 , \3490 , \3498 );
nand \mul_16_12_g19969/U$1 ( \3502 , \3500 , \3501 );
nand \g5076/U$1 ( \3503 , \3502 , \1529 );
nor \mul_17_13_g20022/U$1 ( \3504 , \2669 , \2727 );
not \mul_17_13_g20013/U$2 ( \3505 , \3504 );
nand \mul_17_13_g20013/U$1 ( \3506 , \3505 , \3280 );
not \mul_17_13_g19992/U$3 ( \3507 , \3506 );
nand \g35461/U$1 ( \3508 , \2913 , \2914 );
not \g35645/U$3 ( \3509 , \2826 );
not \g35645/U$4 ( \3510 , \2830 );
or \g35645/U$2 ( \3511 , \3509 , \3510 );
nand \g35645/U$1 ( \3512 , \3511 , \2866 );
not \g35644/U$2 ( \3513 , \3512 );
nand \g35644/U$1 ( \3514 , \3513 , \2910 , \2814 );
nand \mul_17_13_g20003/U$1 ( \3515 , \3508 , \3514 , \2926 );
not \mul_17_13_g19992/U$4 ( \3516 , \3515 );
or \mul_17_13_g19992/U$2 ( \3517 , \3507 , \3516 );
or \mul_17_13_g19992/U$5 ( \3518 , \3515 , \3506 );
nand \mul_17_13_g19992/U$1 ( \3519 , \3517 , \3518 );
nand \g5083/U$1 ( \3520 , \3519 , \2936 );
nand \g5008/U$1 ( \3521 , \3503 , \3520 );
not \g4899/U$3 ( \3522 , \b[13] );
not \g4899/U$4 ( \3523 , \3124 );
or \g4899/U$2 ( \3524 , \3522 , \3523 );
and \g4914/U$2 ( \3525 , \a[13] , \1466 );
xor \g5032/U$1 ( \3526 , \c[13] , \d[13] );
not \g4934/U$3 ( \3527 , \3526 );
not \g4934/U$4 ( \3528 , \1383 );
or \g4934/U$2 ( \3529 , \3527 , \3528 );
not \add_15_12_g7223/U$2 ( \3530 , \3012 );
nor \add_15_12_g7223/U$1 ( \3531 , \3530 , \2980 );
not \add_15_12_g7142/U$3 ( \3532 , \3531 );
not \add_15_12_g7269/U$1 ( \3533 , \2981 );
and \g35878/U$2 ( \3534 , \2979 , \2992 , \3533 );
nand \add_15_12_g7172/U$1 ( \3535 , \3007 , \3533 );
nand \add_15_12_g7165/U$1 ( \3536 , \3535 , \3010 );
nor \g35878/U$1 ( \3537 , \3534 , \3536 );
not \add_15_12_g7142/U$4 ( \3538 , \3537 );
or \add_15_12_g7142/U$2 ( \3539 , \3532 , \3538 );
or \add_15_12_g7142/U$5 ( \3540 , \3537 , \3531 );
nand \add_15_12_g7142/U$1 ( \3541 , \3539 , \3540 );
and \g4952/U$2 ( \3542 , \2961 , \3541 );
not \add_14_12_g7223/U$2 ( \3543 , \3074 );
nor \add_14_12_g7223/U$1 ( \3544 , \3543 , \3042 );
not \add_14_12_g7142/U$3 ( \3545 , \3544 );
not \add_14_12_g7269/U$1 ( \3546 , \3043 );
and \g35874/U$2 ( \3547 , \3041 , \3054 , \3546 );
nand \add_14_12_g7172/U$1 ( \3548 , \3069 , \3546 );
nand \add_14_12_g7165/U$1 ( \3549 , \3548 , \3072 );
nor \g35874/U$1 ( \3550 , \3547 , \3549 );
not \add_14_12_g7142/U$4 ( \3551 , \3550 );
or \add_14_12_g7142/U$2 ( \3552 , \3545 , \3551 );
or \add_14_12_g7142/U$5 ( \3553 , \3550 , \3544 );
nand \add_14_12_g7142/U$1 ( \3554 , \3552 , \3553 );
not \g4981/U$3 ( \3555 , \3554 );
not \g4981/U$4 ( \3556 , \3087 );
or \g4981/U$2 ( \3557 , \3555 , \3556 );
and \g35868/U$2 ( \3558 , \1282 , \d[13] );
and \g35868/U$3 ( \3559 , \1514 , \c[13] );
nor \g35868/U$1 ( \3560 , \3558 , \3559 );
nand \g4981/U$1 ( \3561 , \3557 , \3560 );
nor \g4952/U$1 ( \3562 , \3542 , \3561 );
nand \g4934/U$1 ( \3563 , \3529 , \3562 );
nor \g4914/U$1 ( \3564 , \3525 , \3563 );
nand \g4899/U$1 ( \3565 , \3524 , \3564 );
not \g35818/U$2 ( \3566 , \3565 );
nand \g4849/U$1 ( \3567 , \1338 , \a[13] );
not \g4958/U$3 ( \3568 , \3101 );
nand \g5086/U$1 ( \3569 , \b[13] , \c[13] );
not \g4958/U$4 ( \3570 , \3569 );
and \g4958/U$2 ( \3571 , \3568 , \3570 );
or \g5073/U$1 ( \3572 , \a[13] , \d[13] );
and \g4958/U$5 ( \3573 , \1457 , \3572 );
nor \g4958/U$1 ( \3574 , \3571 , \3573 );
nand \g35818/U$1 ( \3575 , \3566 , \3567 , \3574 );
nor \g4823/U$1 ( \3576 , \3521 , \3575 );
not \g4822/U$1 ( \3577 , \3576 );
not \g4826/U$3 ( \3578 , \a[0] );
not \g4826/U$4 ( \3579 , \2946 );
or \g4826/U$2 ( \3580 , \3578 , \3579 );
not \g4877/U$3 ( \3581 , \d[0] );
not \g4877/U$4 ( \3582 , \1457 );
or \g4877/U$2 ( \3583 , \3581 , \3582 );
xor \g5025/U$1 ( \3584 , \c[0] , \d[0] );
and \g4888/U$2 ( \3585 , \3305 , \3584 );
not \mul_16_12_g20651/U$1 ( \3586 , \1044 );
not \g4903/U$3 ( \3587 , \3586 );
not \g4903/U$4 ( \3588 , \1529 );
or \g4903/U$2 ( \3589 , \3587 , \3588 );
xor \add_15_12_g7227/U$1 ( \3590 , \b[0] , \d[0] );
and \g4922/U$2 ( \3591 , \2961 , \3590 );
xor \add_14_12_g7227/U$1 ( \3592 , \a[0] , \c[0] );
not \g4940/U$3 ( \3593 , \3592 );
not \g4940/U$4 ( \3594 , \3087 );
or \g4940/U$2 ( \3595 , \3593 , \3594 );
nand \g5062/U$1 ( \3596 , \1282 , \d[0] );
and \g5000/U$2 ( \3597 , \1293 , \b[0] );
and \g5000/U$3 ( \3598 , \1435 , \c[0] );
nor \g5000/U$1 ( \3599 , \3597 , \3598 );
and \g4965/U$1 ( \3600 , \3596 , \3599 );
nand \g4940/U$1 ( \3601 , \3595 , \3600 );
nor \g4922/U$1 ( \3602 , \3591 , \3601 );
nand \g4903/U$1 ( \3603 , \3589 , \3602 );
nor \g4888/U$1 ( \3604 , \3585 , \3603 );
nand \g4877/U$1 ( \3605 , \3583 , \3604 );
and \g5037/U$1 ( \3606 , \b[0] , \c[0] );
not \g4955/U$3 ( \3607 , \3606 );
not \g4955/U$4 ( \3608 , \3102 );
or \g4955/U$2 ( \3609 , \3607 , \3608 );
or \g5044/U$1 ( \3610 , \a[0] , \b[0] );
and \g4964/U$2 ( \3611 , \2954 , \3610 );
not \mul_17_13_g20680/U$1 ( \3612 , \852 );
and \g5072/U$1 ( \3613 , \2936 , \3612 );
nor \g4964/U$1 ( \3614 , \3611 , \3613 );
nand \g4955/U$1 ( \3615 , \3609 , \3614 );
nor \g4861/U$1 ( \3616 , \3605 , \3615 );
nand \g4826/U$1 ( \3617 , \3580 , \3616 );
not \g4827/U$3 ( \3618 , \a[8] );
not \g4827/U$4 ( \3619 , \2946 );
or \g4827/U$2 ( \3620 , \3618 , \3619 );
not \fopt35674/U$1 ( \3621 , \645 );
and \g4840/U$2 ( \3622 , \3621 , \d[8] );
not \mul_17_13_g20055/U$3 ( \3623 , \782 );
not \mul_17_13_g20055/U$4 ( \3624 , \904 );
or \mul_17_13_g20055/U$2 ( \3625 , \3623 , \3624 );
nand \mul_17_13_g20055/U$1 ( \3626 , \3625 , \783 );
not \mul_17_13_g20072/U$2 ( \3627 , \2903 );
nand \mul_17_13_g20072/U$1 ( \3628 , \3627 , \2900 );
xnor \g35462/U$1 ( \3629 , \3626 , \3628 );
not \g4999/U$3 ( \3630 , \3629 );
not \g4999/U$4 ( \3631 , \916 );
or \g4999/U$2 ( \3632 , \3630 , \3631 );
not \mul_16_12_g20054/U$2 ( \3633 , \2172 );
nand \mul_16_12_g20054/U$1 ( \3634 , \3633 , \2188 );
not \mul_16_12_g20019/U$3 ( \3635 , \3634 );
not \mul_16_12_g20019/U$4 ( \3636 , \2120 );
or \mul_16_12_g20019/U$2 ( \3637 , \3635 , \3636 );
or \mul_16_12_g20019/U$5 ( \3638 , \2120 , \3634 );
nand \mul_16_12_g20019/U$1 ( \3639 , \3637 , \3638 );
nand \g5046/U$1 ( \3640 , \3639 , \1478 );
nand \g4999/U$1 ( \3641 , \3632 , \3640 );
xor \g5021/U$1 ( \3642 , \c[8] , \d[8] );
not \g4916/U$3 ( \3643 , \3642 );
not \g4916/U$4 ( \3644 , \1320 );
or \g4916/U$2 ( \3645 , \3643 , \3644 );
not \add_15_12_g7251/U$1 ( \3646 , \2989 );
nand \add_15_12_g7217/U$1 ( \3647 , \3646 , \2994 );
not \add_15_12_g7154/U$3 ( \3648 , \3647 );
not \add_15_12_g7154/U$4 ( \3649 , \2979 );
or \add_15_12_g7154/U$2 ( \3650 , \3648 , \3649 );
or \add_15_12_g7154/U$5 ( \3651 , \2979 , \3647 );
nand \add_15_12_g7154/U$1 ( \3652 , \3650 , \3651 );
and \g4921/U$2 ( \3653 , \2961 , \3652 );
not \add_14_12_g7251/U$1 ( \3654 , \3051 );
nand \add_14_12_g7217/U$1 ( \3655 , \3654 , \3056 );
not \add_14_12_g7154/U$3 ( \3656 , \3655 );
not \add_14_12_g7154/U$4 ( \3657 , \3041 );
or \add_14_12_g7154/U$2 ( \3658 , \3656 , \3657 );
or \add_14_12_g7154/U$5 ( \3659 , \3041 , \3655 );
nand \add_14_12_g7154/U$1 ( \3660 , \3658 , \3659 );
not \g4941/U$3 ( \3661 , \3660 );
not \g4941/U$4 ( \3662 , \3087 );
or \g4941/U$2 ( \3663 , \3661 , \3662 );
and \g35857/U$2 ( \3664 , \1282 , \d[8] );
and \g35857/U$3 ( \3665 , \c[8] , \1514 );
and \g35857/U$4 ( \3666 , \1293 , \b[8] );
nor \g35857/U$1 ( \3667 , \3664 , \3665 , \3666 );
nand \g4941/U$1 ( \3668 , \3663 , \3667 );
nor \g4921/U$1 ( \3669 , \3653 , \3668 );
nand \g4916/U$1 ( \3670 , \3645 , \3669 );
nor \g4885/U$1 ( \3671 , \3641 , \3670 );
or \g35736/U$2 ( \3672 , \a[8] , \b[8] );
nand \g35736/U$1 ( \3673 , \3672 , \1351 );
and \g5056/U$1 ( \3674 , \b[8] , \c[8] );
nand \g4986/U$1 ( \3675 , \1316 , \3674 );
nand \g35735/U$1 ( \3676 , \3671 , \3673 , \3675 );
nor \g4840/U$1 ( \3677 , \3622 , \3676 );
nand \g4827/U$1 ( \3678 , \3620 , \3677 );
not \g4828/U$3 ( \3679 , \a[9] );
not \g4828/U$4 ( \3680 , \3114 );
or \g4828/U$2 ( \3681 , \3679 , \3680 );
and \g5253/U$1 ( \3682 , \644 , \d[9] );
nand \mul_17_13_g20724/U$1 ( \3683 , \2906 , \2892 );
not \mul_17_13_g20009/U$3 ( \3684 , \3683 );
not \mul_17_13_g20030/U$3 ( \3685 , \2900 );
not \mul_17_13_g20030/U$4 ( \3686 , \3626 );
or \mul_17_13_g20030/U$2 ( \3687 , \3685 , \3686 );
not \mul_17_13_g20090/U$1 ( \3688 , \2903 );
nand \mul_17_13_g20030/U$1 ( \3689 , \3687 , \3688 );
not \mul_17_13_g20009/U$4 ( \3690 , \3689 );
or \mul_17_13_g20009/U$2 ( \3691 , \3684 , \3690 );
or \mul_17_13_g20009/U$5 ( \3692 , \3689 , \3683 );
nand \mul_17_13_g20009/U$1 ( \3693 , \3691 , \3692 );
and \g5016/U$2 ( \3694 , \3693 , \2936 );
not \mul_16_12_g20033/U$2 ( \3695 , \2165 );
nand \mul_16_12_g20033/U$1 ( \3696 , \3695 , \2190 );
not \mul_16_12_g19989/U$3 ( \3697 , \3696 );
not \mul_16_12_g20064/U$1 ( \3698 , \2172 );
not \mul_16_12_g20018/U$3 ( \3699 , \3698 );
not \mul_16_12_g20018/U$4 ( \3700 , \2120 );
or \mul_16_12_g20018/U$2 ( \3701 , \3699 , \3700 );
nand \mul_16_12_g20018/U$1 ( \3702 , \3701 , \2188 );
not \mul_16_12_g19989/U$4 ( \3703 , \3702 );
or \mul_16_12_g19989/U$2 ( \3704 , \3697 , \3703 );
or \mul_16_12_g19989/U$5 ( \3705 , \3702 , \3696 );
nand \mul_16_12_g19989/U$1 ( \3706 , \3704 , \3705 );
and \g5016/U$3 ( \3707 , \3706 , \1478 );
nor \g5016/U$1 ( \3708 , \3694 , \3707 );
and \g5092/U$1 ( \3709 , \b[9] , \c[9] );
nand \g4992/U$1 ( \3710 , \1316 , \3709 );
or \g5057/U$1 ( \3711 , \a[9] , \b[9] );
and \g4884/U$2 ( \3712 , \672 , \3711 );
xor \g5018/U$1 ( \3713 , \c[9] , \d[9] );
not \g4917/U$3 ( \3714 , \3713 );
not \g4917/U$4 ( \3715 , \925 );
or \g4917/U$2 ( \3716 , \3714 , \3715 );
not \add_15_12_g7150/U$3 ( \3717 , \3646 );
not \add_15_12_g7150/U$4 ( \3718 , \2979 );
or \add_15_12_g7150/U$2 ( \3719 , \3717 , \3718 );
nand \add_15_12_g7150/U$1 ( \3720 , \3719 , \2994 );
not \add_15_12_g7208/U$2 ( \3721 , \2990 );
nand \add_15_12_g7208/U$1 ( \3722 , \3721 , \2996 );
xnor \add_15_12_g7277/U$1 ( \3723 , \3720 , \3722 );
and \g4919/U$2 ( \3724 , \2961 , \3723 );
not \add_14_12_g7150/U$3 ( \3725 , \3654 );
not \add_14_12_g7150/U$4 ( \3726 , \3041 );
or \add_14_12_g7150/U$2 ( \3727 , \3725 , \3726 );
nand \add_14_12_g7150/U$1 ( \3728 , \3727 , \3056 );
not \add_14_12_g7208/U$2 ( \3729 , \3052 );
nand \add_14_12_g7208/U$1 ( \3730 , \3729 , \3058 );
xnor \add_14_12_g7277/U$1 ( \3731 , \3728 , \3730 );
not \g4938/U$3 ( \3732 , \3731 );
not \g4938/U$4 ( \3733 , \3087 );
or \g4938/U$2 ( \3734 , \3732 , \3733 );
and \g35855/U$2 ( \3735 , \1282 , \d[9] );
and \g35855/U$3 ( \3736 , \c[9] , \1435 );
and \g35855/U$4 ( \3737 , \1293 , \b[9] );
nor \g35855/U$1 ( \3738 , \3735 , \3736 , \3737 );
nand \g4938/U$1 ( \3739 , \3734 , \3738 );
nor \g4919/U$1 ( \3740 , \3724 , \3739 );
nand \g4917/U$1 ( \3741 , \3716 , \3740 );
nor \g4884/U$1 ( \3742 , \3712 , \3741 );
nand \g4864/U$1 ( \3743 , \3708 , \3710 , \3742 );
nor \g4839/U$1 ( \3744 , \3682 , \3743 );
nand \g4828/U$1 ( \3745 , \3681 , \3744 );
not \mul_17_13_g20004/U$3 ( \3746 , \2866 );
not \mul_17_13_g20004/U$4 ( \3747 , \2910 );
or \mul_17_13_g20004/U$2 ( \3748 , \3746 , \3747 );
not \mul_17_13_g20038/U$1 ( \3749 , \2914 );
nand \mul_17_13_g20004/U$1 ( \3750 , \3748 , \3749 );
nand \mul_17_13_g19996/U$1 ( \3751 , \3750 , \2814 );
nand \mul_17_13_g20722/U$1 ( \3752 , \2926 , \2913 );
xor \mul_17_13_g19989/U$1 ( \3753 , \3751 , \3752 );
and \g4995/U$2 ( \3754 , \3753 , \2936 );
not \mul_16_12_g19980/U$3 ( \3755 , \2206 );
not \mul_16_12_g19980/U$4 ( \3756 , \2193 );
or \mul_16_12_g19980/U$2 ( \3757 , \3755 , \3756 );
not \mul_16_12_g20006/U$1 ( \3758 , \2211 );
nand \mul_16_12_g19980/U$1 ( \3759 , \3757 , \3758 );
nand \mul_16_12_g19975/U$1 ( \3760 , \3759 , \2112 );
not \mul_16_12_g19993/U$2 ( \3761 , \2221 );
nand \mul_16_12_g19993/U$1 ( \3762 , \3761 , \2205 );
and \mul_16_12_g19970/U$2 ( \3763 , \3760 , \3762 );
not \mul_16_12_g19970/U$4 ( \3764 , \3760 );
not \mul_16_12_g19992/U$1 ( \3765 , \3762 );
and \mul_16_12_g19970/U$3 ( \3766 , \3764 , \3765 );
nor \mul_16_12_g19970/U$1 ( \3767 , \3763 , \3766 );
and \g4995/U$3 ( \3768 , \3767 , \1529 );
nor \g4995/U$1 ( \3769 , \3754 , \3768 );
nand \g4838/U$1 ( \3770 , \2946 , \a[12] );
not \g4963/U$3 ( \3771 , \d[12] );
not \g4963/U$4 ( \3772 , \1457 );
or \g4963/U$2 ( \3773 , \3771 , \3772 );
and \g5049/U$1 ( \3774 , \b[12] , \c[12] );
nand \g4987/U$1 ( \3775 , \1316 , \3774 );
nand \g4963/U$1 ( \3776 , \3773 , \3775 );
not \g4894/U$3 ( \3777 , \b[12] );
not \g4894/U$4 ( \3778 , \3124 );
or \g4894/U$2 ( \3779 , \3777 , \3778 );
and \g4904/U$2 ( \3780 , \1351 , \a[12] );
xor \g5022/U$1 ( \3781 , \c[12] , \d[12] );
not \g4928/U$3 ( \3782 , \3781 );
not \g4928/U$4 ( \3783 , \3305 );
or \g4928/U$2 ( \3784 , \3782 , \3783 );
nand \add_15_12_g7213/U$1 ( \3785 , \3533 , \3010 );
not \add_15_12_g7143/U$3 ( \3786 , \3785 );
not \add_15_12_g7151/U$3 ( \3787 , \2992 );
not \add_15_12_g7151/U$4 ( \3788 , \2979 );
or \add_15_12_g7151/U$2 ( \3789 , \3787 , \3788 );
nand \add_15_12_g7151/U$1 ( \3790 , \3789 , \3008 );
not \add_15_12_g7143/U$4 ( \3791 , \3790 );
or \add_15_12_g7143/U$2 ( \3792 , \3786 , \3791 );
or \add_15_12_g7143/U$5 ( \3793 , \3790 , \3785 );
nand \add_15_12_g7143/U$1 ( \3794 , \3792 , \3793 );
and \g4942/U$2 ( \3795 , \3794 , \2961 );
nand \add_14_12_g7213/U$1 ( \3796 , \3546 , \3072 );
not \add_14_12_g7143/U$3 ( \3797 , \3796 );
not \add_14_12_g7151/U$3 ( \3798 , \3054 );
not \add_14_12_g7151/U$4 ( \3799 , \3041 );
or \add_14_12_g7151/U$2 ( \3800 , \3798 , \3799 );
nand \add_14_12_g7151/U$1 ( \3801 , \3800 , \3070 );
not \add_14_12_g7143/U$4 ( \3802 , \3801 );
or \add_14_12_g7143/U$2 ( \3803 , \3797 , \3802 );
or \add_14_12_g7143/U$5 ( \3804 , \3801 , \3796 );
nand \add_14_12_g7143/U$1 ( \3805 , \3803 , \3804 );
not \g4967/U$3 ( \3806 , \3805 );
not \g4967/U$4 ( \3807 , \3087 );
or \g4967/U$2 ( \3808 , \3806 , \3807 );
and \g35869/U$2 ( \3809 , \1282 , \d[12] );
and \g35869/U$3 ( \3810 , \1435 , \c[12] );
nor \g35869/U$1 ( \3811 , \3809 , \3810 );
nand \g4967/U$1 ( \3812 , \3808 , \3811 );
nor \g4942/U$1 ( \3813 , \3795 , \3812 );
nand \g4928/U$1 ( \3814 , \3784 , \3813 );
nor \g4904/U$1 ( \3815 , \3780 , \3814 );
nand \g4894/U$1 ( \3816 , \3779 , \3815 );
nor \g4868/U$1 ( \3817 , \3776 , \3816 );
nand \g4829/U$1 ( \3818 , \3769 , \3770 , \3817 );
not \g4841/U$3 ( \3819 , \a[5] );
not \g4841/U$4 ( \3820 , \1338 );
or \g4841/U$2 ( \3821 , \3819 , \3820 );
or \g5081/U$1 ( \3822 , \a[5] , \d[5] );
not \g4954/U$3 ( \3823 , \3822 );
not \g4954/U$4 ( \3824 , \644 );
or \g4954/U$2 ( \3825 , \3823 , \3824 );
not \g4974/U$3 ( \3826 , \917 );
nand \mul_17_13_g20129/U$1 ( \3827 , \899 , \819 );
xor \g35814/U$1 ( \3828 , \3827 , \879 );
not \g4974/U$4 ( \3829 , \3828 );
and \g4974/U$2 ( \3830 , \3826 , \3829 );
or \g5078/U$1 ( \3831 , \a[5] , \b[5] );
and \g4974/U$5 ( \3832 , \672 , \3831 );
nor \g4974/U$1 ( \3833 , \3830 , \3832 );
nand \g4954/U$1 ( \3834 , \3825 , \3833 );
and \g5093/U$1 ( \3835 , \b[5] , \c[5] );
not \g4880/U$3 ( \3836 , \3835 );
not \g4880/U$4 ( \3837 , \1316 );
or \g4880/U$2 ( \3838 , \3836 , \3837 );
xor \g5029/U$1 ( \3839 , \c[5] , \d[5] );
and \g4891/U$2 ( \3840 , \3305 , \3839 );
not \mul_16_12_g20081/U$3 ( \3841 , \1089 );
nand \mul_16_12_g20115/U$1 ( \3842 , \1095 , \1027 );
not \mul_16_12_g20081/U$4 ( \3843 , \3842 );
or \mul_16_12_g20081/U$2 ( \3844 , \3841 , \3843 );
or \mul_16_12_g20081/U$5 ( \3845 , \3842 , \1089 );
nand \mul_16_12_g20081/U$1 ( \3846 , \3844 , \3845 );
not \g4911/U$3 ( \3847 , \3846 );
not \g4911/U$4 ( \3848 , \1478 );
or \g4911/U$2 ( \3849 , \3847 , \3848 );
nand \add_15_12_g7215/U$1 ( \3850 , \1192 , \1200 );
not \add_15_12_g7145/U$3 ( \3851 , \3850 );
or \add_15_12_g7155/U$2 ( \3852 , \1416 , \1190 );
nand \add_15_12_g7155/U$1 ( \3853 , \3852 , \1197 );
not \add_15_12_g7145/U$4 ( \3854 , \3853 );
or \add_15_12_g7145/U$2 ( \3855 , \3851 , \3854 );
or \add_15_12_g7145/U$5 ( \3856 , \3853 , \3850 );
nand \add_15_12_g7145/U$1 ( \3857 , \3855 , \3856 );
and \g4925/U$2 ( \3858 , \2961 , \3857 );
nand \add_14_12_g7215/U$1 ( \3859 , \1255 , \1263 );
not \add_14_12_g7145/U$3 ( \3860 , \3859 );
or \add_14_12_g7155/U$2 ( \3861 , \1426 , \1253 );
nand \add_14_12_g7155/U$1 ( \3862 , \3861 , \1260 );
not \add_14_12_g7145/U$4 ( \3863 , \3862 );
or \add_14_12_g7145/U$2 ( \3864 , \3860 , \3863 );
or \add_14_12_g7145/U$5 ( \3865 , \3862 , \3859 );
nand \add_14_12_g7145/U$1 ( \3866 , \3864 , \3865 );
not \g4949/U$3 ( \3867 , \3866 );
not \g4949/U$4 ( \3868 , \3087 );
or \g4949/U$2 ( \3869 , \3867 , \3868 );
and \g35859/U$2 ( \3870 , \1282 , \d[5] );
and \g35859/U$3 ( \3871 , \c[5] , \1514 );
and \g35859/U$4 ( \3872 , \1293 , \b[5] );
nor \g35859/U$1 ( \3873 , \3870 , \3871 , \3872 );
nand \g4949/U$1 ( \3874 , \3869 , \3873 );
nor \g4925/U$1 ( \3875 , \3858 , \3874 );
nand \g4911/U$1 ( \3876 , \3849 , \3875 );
nor \g4891/U$1 ( \3877 , \3840 , \3876 );
nand \g4880/U$1 ( \3878 , \3838 , \3877 );
nor \g4862/U$1 ( \3879 , \3834 , \3878 );
nand \g4841/U$1 ( \3880 , \3821 , \3879 );
nor \add_7_12_g9771/U$1 ( \3881 , \c[14] , \d[14] );
not \add_7_12_g9733/U$2 ( \3882 , \3881 );
nand \add_7_12_g9768/U$1 ( \3883 , \c[14] , \d[14] );
nand \add_7_12_g9733/U$1 ( \3884 , \3882 , \3883 );
nand \add_7_12_g9743/U$1 ( \3885 , \c[1] , \d[1] );
nand \add_7_12_g9772/U$1 ( \3886 , \c[0] , \d[0] );
and \add_7_12_g9698/U$2 ( \3887 , \3885 , \3886 );
nor \add_7_12_g9750/U$1 ( \3888 , \c[1] , \d[1] );
nor \add_7_12_g9753/U$1 ( \3889 , \c[2] , \d[2] );
nor \add_7_12_g9698/U$1 ( \3890 , \3887 , \3888 , \3889 );
not \add_7_12_g9780/U$2 ( \3891 , \3890 );
nand \add_7_12_g9747/U$1 ( \3892 , \c[3] , \d[3] );
nand \add_7_12_g9738/U$1 ( \3893 , \c[2] , \d[2] );
nand \add_7_12_g9780/U$1 ( \3894 , \3891 , \3892 , \3893 );
nor \add_7_12_g9748/U$1 ( \3895 , \c[5] , \d[5] );
nor \add_7_12_g9757/U$1 ( \3896 , \c[4] , \d[4] );
nor \add_7_12_g9730/U$1 ( \3897 , \3895 , \3896 );
nor \add_7_12_g9741/U$1 ( \3898 , \c[7] , \d[7] );
nor \add_7_12_g9739/U$1 ( \3899 , \c[6] , \d[6] );
nor \add_7_12_g9735/U$1 ( \3900 , \3898 , \3899 );
nor \add_7_12_g9756/U$1 ( \3901 , \c[3] , \d[3] );
not \add_7_12_g9755/U$1 ( \3902 , \3901 );
nand \add_7_12_g9683/U$1 ( \3903 , \3894 , \3897 , \3900 , \3902 );
nand \add_7_12_g9759/U$1 ( \3904 , \c[4] , \d[4] );
nor \add_7_12_g9713/U$1 ( \3905 , \3895 , \3904 );
nand \add_7_12_g9749/U$1 ( \3906 , \c[6] , \d[6] );
nand \add_7_12_g9752/U$1 ( \3907 , \c[7] , \d[7] );
nand \add_7_12_g9765/U$1 ( \3908 , \c[5] , \d[5] );
nand \add_7_12_g9712/U$1 ( \3909 , \3906 , \3907 , \3908 );
or \add_7_12_g9694/U$2 ( \3910 , \3905 , \3909 );
not \add_7_12_g9751/U$1 ( \3911 , \3907 );
or \add_7_12_g9694/U$3 ( \3912 , \3900 , \3911 );
nand \add_7_12_g9694/U$1 ( \3913 , \3910 , \3912 );
nand \add_7_12_g9677/U$1 ( \3914 , \3903 , \3913 );
nor \add_7_12_g9742/U$1 ( \3915 , \c[11] , \d[11] );
nor \add_7_12_g9762/U$1 ( \3916 , \c[10] , \d[10] );
nor \add_7_12_g9724/U$1 ( \3917 , \3915 , \3916 );
nor \add_7_12_g9745/U$1 ( \3918 , \c[9] , \d[9] );
nor \add_7_12_g9769/U$1 ( \3919 , \c[8] , \d[8] );
nor \add_7_12_g9728/U$1 ( \3920 , \3918 , \3919 );
and \add_7_12_g9705/U$1 ( \3921 , \3917 , \3920 );
nor \add_7_12_g9770/U$1 ( \3922 , \c[13] , \d[13] );
nor \add_7_12_g9767/U$1 ( \3923 , \c[12] , \d[12] );
nor \add_7_12_g9729/U$1 ( \3924 , \3922 , \3923 );
and \add_7_12_g9660/U$2 ( \3925 , \3914 , \3921 , \3924 );
nand \add_7_12_g9744/U$1 ( \3926 , \c[12] , \d[12] );
or \add_7_12_g9708/U$2 ( \3927 , \3922 , \3926 );
nand \add_7_12_g9746/U$1 ( \3928 , \c[13] , \d[13] );
nand \add_7_12_g9708/U$1 ( \3929 , \3927 , \3928 );
not \add_7_12_g9679/U$2 ( \3930 , \3929 );
nand \add_7_12_g9764/U$1 ( \3931 , \c[10] , \d[10] );
or \add_7_12_g9696/U$2 ( \3932 , \3915 , \3931 );
nand \add_7_12_g9740/U$1 ( \3933 , \c[8] , \d[8] );
or \add_7_12_g9711/U$2 ( \3934 , \3918 , \3933 );
nand \add_7_12_g9760/U$1 ( \3935 , \c[9] , \d[9] );
nand \add_7_12_g9711/U$1 ( \3936 , \3934 , \3935 );
nand \add_7_12_g9700/U$1 ( \3937 , \3917 , \3936 );
nand \add_7_12_g9758/U$1 ( \3938 , \c[11] , \d[11] );
nand \add_7_12_g9696/U$1 ( \3939 , \3932 , \3937 , \3938 );
nand \add_7_12_g9689/U$1 ( \3940 , \3939 , \3924 );
nand \add_7_12_g9679/U$1 ( \3941 , \3930 , \3940 );
nor \add_7_12_g9660/U$1 ( \3942 , \3925 , \3941 );
xor \add_7_12_g9651/U$1 ( \3943 , \3884 , \3942 );
not \add_7_12_g9723/U$2 ( \3944 , \3899 );
nand \add_7_12_g9723/U$1 ( \3945 , \3944 , \3906 );
or \add_7_12_g9692/U$2 ( \3946 , \3888 , \3886 );
nand \add_7_12_g9692/U$1 ( \3947 , \3946 , \3885 );
nor \add_7_12_g9719/U$1 ( \3948 , \3901 , \3889 );
and \add_7_12_g9682/U$2 ( \3949 , \3947 , \3948 );
or \add_7_12_g9709/U$2 ( \3950 , \3901 , \3893 );
nand \add_7_12_g9709/U$1 ( \3951 , \3950 , \3892 );
nor \add_7_12_g9682/U$1 ( \3952 , \3949 , \3951 );
not \add_7_12_g9779/U$2 ( \3953 , \3952 );
nand \add_7_12_g9779/U$1 ( \3954 , \3953 , \3897 );
not \add_7_12_g9702/U$2 ( \3955 , \3908 );
nor \add_7_12_g9702/U$1 ( \3956 , \3955 , \3905 );
and \add_7_12_g9673/U$1 ( \3957 , \3954 , \3956 );
xor \add_7_12_g9654/U$1 ( \3958 , \3945 , \3957 );
not \add_7_12_g9716/U$2 ( \3959 , \3908 );
nor \add_7_12_g9716/U$1 ( \3960 , \3959 , \3895 );
or \add_7_12_g9670/U$2 ( \3961 , \3952 , \3896 );
nand \add_7_12_g9670/U$1 ( \3962 , \3961 , \3904 );
xor \add_7_12_g9655/U$1 ( \3963 , \3960 , \3962 );
and \add_7_12_g9657/U$2 ( \3964 , \3914 , \3920 );
nor \add_7_12_g9657/U$1 ( \3965 , \3964 , \3936 );
not \add_7_12_g9766/U$1 ( \3966 , \3923 );
and \add_7_12_g9659/U$2 ( \3967 , \3914 , \3921 , \3966 );
not \add_7_12_g9695/U$1 ( \3968 , \3939 );
or \add_7_12_g9680/U$2 ( \3969 , \3968 , \3923 );
nand \add_7_12_g9680/U$1 ( \3970 , \3969 , \3926 );
nor \add_7_12_g9659/U$1 ( \3971 , \3967 , \3970 );
not \add_7_12_g9676/U$1 ( \3972 , \3914 );
or \add_7_12_g9662/U$2 ( \3973 , \3972 , \3919 );
nand \add_7_12_g9662/U$1 ( \3974 , \3973 , \3933 );
not \add_7_12_g9706/U$2 ( \3975 , \3924 );
nor \add_7_12_g9706/U$1 ( \3976 , \3975 , \3881 );
and \add_7_12_g9664/U$2 ( \3977 , \3914 , \3921 , \3976 );
nand \add_7_12_g9690/U$1 ( \3978 , \3939 , \3976 );
not \add_7_12_g9701/U$2 ( \3979 , \3881 );
nand \add_7_12_g9701/U$1 ( \3980 , \3979 , \3929 );
nand \add_7_12_g9686/U$1 ( \3981 , \3978 , \3980 , \3883 );
nor \add_7_12_g9664/U$1 ( \3982 , \3977 , \3981 );
not \add_7_12_g9704/U$1 ( \3983 , \3921 );
nor \add_7_12_g9763/U$1 ( \3984 , \c[15] , \d[15] );
nor \add_7_12_g9731/U$1 ( \3985 , \3881 , \3984 );
nand \add_7_12_g9707/U$1 ( \3986 , \3985 , \3924 );
or \add_7_12_g9665/U$2 ( \3987 , \3972 , \3983 , \3986 );
and \add_7_12_g9684/U$2 ( \3988 , \3929 , \3985 );
nor \add_7_12_g9688/U$1 ( \3989 , \3968 , \3986 );
or \add_7_12_g9710/U$2 ( \3990 , \3984 , \3883 );
nand \add_7_12_g9754/U$1 ( \3991 , \c[15] , \d[15] );
nand \add_7_12_g9710/U$1 ( \3992 , \3990 , \3991 );
nor \add_7_12_g9684/U$1 ( \3993 , \3988 , \3989 , \3992 );
nand \add_7_12_g9665/U$1 ( \3994 , \3987 , \3993 );
not \add_7_12_g9761/U$1 ( \3995 , \3916 );
and \add_7_12_g9667/U$2 ( \3996 , \3914 , \3920 , \3995 );
not \add_7_12_g9693/U$3 ( \3997 , \3995 );
not \add_7_12_g9693/U$4 ( \3998 , \3936 );
or \add_7_12_g9693/U$2 ( \3999 , \3997 , \3998 );
nand \add_7_12_g9693/U$1 ( \4000 , \3999 , \3931 );
nor \add_7_12_g9667/U$1 ( \4001 , \3996 , \4000 );
not \add_7_12_g9668/U$3 ( \4002 , \3921 );
not \add_7_12_g9668/U$4 ( \4003 , \3914 );
or \add_7_12_g9668/U$2 ( \4004 , \4002 , \4003 );
nand \add_7_12_g9668/U$1 ( \4005 , \4004 , \3968 );
not \add_7_12_g9721/U$2 ( \4006 , \3919 );
nand \add_7_12_g9721/U$1 ( \4007 , \4006 , \3933 );
and \add_7_12_g9669/U$2 ( \4008 , \4007 , \3914 );
not \add_7_12_g9669/U$4 ( \4009 , \4007 );
and \add_7_12_g9669/U$3 ( \4010 , \4009 , \3972 );
or \add_7_12_g9669/U$1 ( \4011 , \4008 , \4010 );
not \add_7_12_g9703/U$2 ( \4012 , \3899 );
nand \add_7_12_g9703/U$1 ( \4013 , \4012 , \3897 );
or \add_7_12_g9672/U$2 ( \4014 , \3952 , \4013 );
or \add_7_12_g9672/U$3 ( \4015 , \3899 , \3956 );
nand \add_7_12_g9672/U$1 ( \4016 , \4014 , \4015 , \3906 );
not \add_7_12_g9725/U$2 ( \4017 , \3896 );
nand \add_7_12_g9725/U$1 ( \4018 , \4017 , \3904 );
xor \add_7_12_g9674/U$1 ( \4019 , \4018 , \3952 );
and \add_7_12_g9734/U$1 ( \4020 , \3902 , \3892 );
not \add_7_12_g9687/U$2 ( \4021 , \3890 );
nand \add_7_12_g9687/U$1 ( \4022 , \4021 , \3893 );
xor \add_7_12_g9678/U$1 ( \4023 , \4020 , \4022 );
not \add_7_12_g9726/U$2 ( \4024 , \3893 );
nor \add_7_12_g9726/U$1 ( \4025 , \4024 , \3889 );
xor \add_7_12_g9685/U$1 ( \4026 , \4025 , \3947 );
not \add_7_12_g9732/U$2 ( \4027 , \3888 );
nand \add_7_12_g9732/U$1 ( \4028 , \4027 , \3885 );
xor \add_7_12_g9699/U$1 ( \4029 , \3886 , \4028 );
nand \add_7_12_g9715/U$1 ( \4030 , \3966 , \3926 );
not \add_7_12_g9717/U$2 ( \4031 , \3915 );
nand \add_7_12_g9717/U$1 ( \4032 , \4031 , \3938 );
and \add_7_12_g9718/U$1 ( \4033 , \3995 , \3931 );
not \add_7_12_g9720/U$2 ( \4034 , \3935 );
nor \add_7_12_g9720/U$1 ( \4035 , \4034 , \3918 );
or \add_7_12_g9722/U$1 ( \4036 , \3911 , \3898 );
not \add_7_12_g9727/U$2 ( \4037 , \3991 );
nor \add_7_12_g9727/U$1 ( \4038 , \4037 , \3984 );
not \add_7_12_g9736/U$2 ( \4039 , \3922 );
nand \add_7_12_g9736/U$1 ( \4040 , \4039 , \3928 );
xnor \add_7_12_g2/U$1 ( \4041 , \4033 , \3965 );
xor \add_7_12_g9774/U$1 ( \4042 , \4040 , \3971 );
xor \add_7_12_g9775/U$1 ( \4043 , \4035 , \3974 );
xnor \add_7_12_g9776/U$1 ( \4044 , \4038 , \3982 );
xor \add_7_12_g9777/U$1 ( \4045 , \4032 , \4001 );
xnor \add_7_12_g9778/U$1 ( \4046 , \4036 , \4016 );
xnor \add_7_12_g9781/U$1 ( \4047 , \4005 , \4030 );
xor \add_7_12_g9782/U$1 ( \4048 , \d[0] , \c[0] );
not \mul_7_15_g35030/U$1 ( \4049 , \1454 );
and \mul_7_15_g34585/U$2 ( \4050 , \1528 , \4049 );
not \mul_7_15_g34585/U$4 ( \4051 , \1528 );
and \mul_7_15_g34585/U$3 ( \4052 , \4051 , \1454 );
nor \mul_7_15_g34585/U$1 ( \4053 , \4050 , \4052 );
not \mul_7_15_g34579/U$1 ( \4054 , \4053 );
buf \mul_7_15_g34578/U$1 ( \4055 , \4054 );
not \mul_7_15_g34581/U$1 ( \4056 , \4055 );
not \mul_7_15_g34133/U$3 ( \4057 , \4056 );
not \mul_7_15_g34574/U$3 ( \4058 , \4049 );
not \mul_7_15_g34574/U$4 ( \4059 , \3880 );
or \mul_7_15_g34574/U$2 ( \4060 , \4058 , \4059 );
not \mul_7_15_fopt35204/U$1 ( \4061 , \3880 );
nand \mul_7_15_g34822/U$1 ( \4062 , \4061 , \1454 );
nand \mul_7_15_g34574/U$1 ( \4063 , \4060 , \4062 );
nand \mul_7_15_g34479/U$1 ( \4064 , \4053 , \4063 );
not \fopt35526/U$1 ( \4065 , \4064 );
not \fopt35525/U$1 ( \4066 , \4065 );
not \mul_7_15_g34133/U$4 ( \4067 , \4066 );
or \mul_7_15_g34133/U$2 ( \4068 , \4057 , \4067 );
buf \mul_7_15_fopt35193/U$1 ( \4069 , \4061 );
not \mul_7_15_fopt35187/U$1 ( \4070 , \4069 );
nand \mul_7_15_g34133/U$1 ( \4071 , \4068 , \4070 );
not \mul_7_15_g34132/U$1 ( \4072 , \4071 );
not \mul_7_15_g34023/U$3 ( \4073 , \4072 );
and \mul_7_15_g34621/U$2 ( \4074 , \4061 , \3272 );
not \mul_7_15_g34621/U$4 ( \4075 , \4061 );
not \mul_7_15_g35060/U$1 ( \4076 , \3272 );
and \mul_7_15_g34621/U$3 ( \4077 , \4075 , \4076 );
nor \mul_7_15_g34621/U$1 ( \4078 , \4074 , \4077 );
not \mul_7_15_g34623/U$3 ( \4079 , \1336 );
not \mul_7_15_g34623/U$4 ( \4080 , \4076 );
or \mul_7_15_g34623/U$2 ( \4081 , \4079 , \4080 );
not \mul_7_15_g35337/U$2 ( \4082 , \1336 );
nand \mul_7_15_g35337/U$1 ( \4083 , \4082 , \3272 );
nand \mul_7_15_g34623/U$1 ( \4084 , \4081 , \4083 );
and \mul_7_15_g34467/U$1 ( \4085 , \4078 , \4084 );
buf \mul_7_15_g34464/U$1 ( \4086 , \4085 );
not \mul_7_15_g34710/U$3 ( \4087 , \4044 );
buf \mul_7_15_g35024/U$1 ( \4088 , \1336 );
not \mul_7_15_g35011/U$1 ( \4089 , \4088 );
not \mul_7_15_g34710/U$4 ( \4090 , \4089 );
or \mul_7_15_g34710/U$2 ( \4091 , \4087 , \4090 );
not \mul_7_15_g35006/U$1 ( \4092 , \4044 );
nand \mul_7_15_g34912/U$1 ( \4093 , \4088 , \4092 );
nand \mul_7_15_g34710/U$1 ( \4094 , \4091 , \4093 );
and \mul_7_15_g35323/U$2 ( \4095 , \4086 , \4094 );
not \mul_7_15_g34673/U$3 ( \4096 , \3994 );
not \mul_7_15_g34673/U$4 ( \4097 , \4089 );
or \mul_7_15_g34673/U$2 ( \4098 , \4096 , \4097 );
not \mul_7_15_g35059/U$1 ( \4099 , \3994 );
nand \mul_7_15_g34837/U$1 ( \4100 , \4088 , \4099 );
nand \mul_7_15_g34673/U$1 ( \4101 , \4098 , \4100 );
not \mul_7_15_g35333/U$2 ( \4102 , \4101 );
buf \fopt35519/U$1 ( \4103 , \4078 );
nor \mul_7_15_g35333/U$1 ( \4104 , \4102 , \4103 );
nor \mul_7_15_g35323/U$1 ( \4105 , \4095 , \4104 );
not \mul_7_15_g34023/U$4 ( \4106 , \4105 );
or \mul_7_15_g34023/U$2 ( \4107 , \4073 , \4106 );
not \mul_7_15_g34693/U$3 ( \4108 , \4042 );
buf \fopt35556/U$1 ( \4109 , \3745 );
not \fopt35555/U$1 ( \4110 , \4109 );
not \mul_7_15_g34693/U$4 ( \4111 , \4110 );
or \mul_7_15_g34693/U$2 ( \4112 , \4108 , \4111 );
buf \fopt35563/U$1 ( \4113 , \3745 );
not \fopt35543/U$1 ( \4114 , \4113 );
not \fopt35542/U$1 ( \4115 , \4114 );
not \mul_7_15_g35176/U$1 ( \4116 , \4042 );
nand \mul_7_15_g34930/U$1 ( \4117 , \4115 , \4116 );
nand \mul_7_15_g34693/U$1 ( \4118 , \4112 , \4117 );
not \mul_7_15_g34251/U$3 ( \4119 , \4118 );
not \mul_7_15_g34607/U$3 ( \4120 , \1336 );
not \mul_7_15_g35169/U$1 ( \4121 , \3678 );
not \mul_7_15_g34607/U$4 ( \4122 , \4121 );
or \mul_7_15_g34607/U$2 ( \4123 , \4120 , \4122 );
not \mul_7_15_g35026/U$1 ( \4124 , \1336 );
nand \mul_7_15_g34821/U$1 ( \4125 , \4124 , \3678 );
nand \mul_7_15_g34607/U$1 ( \4126 , \4123 , \4125 );
not \mul_7_15_g34596/U$1 ( \4127 , \4126 );
not \mul_7_15_g35168/U$1 ( \4128 , \3678 );
not \mul_7_15_g34646/U$3 ( \4129 , \4128 );
not \mul_7_15_g34646/U$4 ( \4130 , \3745 );
or \mul_7_15_g34646/U$2 ( \4131 , \4129 , \4130 );
not \fopt35557/U$1 ( \4132 , \3745 );
nand \mul_7_15_g34818/U$1 ( \4133 , \4132 , \3678 );
nand \mul_7_15_g34646/U$1 ( \4134 , \4131 , \4133 );
nand \mul_7_15_g34455/U$1 ( \4135 , \4127 , \4134 );
not \mul_7_15_g34453/U$1 ( \4136 , \4135 );
not \mul_7_15_g34251/U$4 ( \4137 , \4136 );
or \mul_7_15_g34251/U$2 ( \4138 , \4119 , \4137 );
buf \mul_7_15_g34606/U$1 ( \4139 , \4126 );
buf \mul_7_15_g34602/U$1 ( \4140 , \4139 );
not \mul_7_15_g34705/U$3 ( \4141 , \3943 );
not \fopt35560/U$1 ( \4142 , \4113 );
not \mul_7_15_g34705/U$4 ( \4143 , \4142 );
or \mul_7_15_g34705/U$2 ( \4144 , \4141 , \4143 );
not \fopt35545/U$1 ( \4145 , \4113 );
not \fopt35544/U$1 ( \4146 , \4145 );
not \mul_7_15_g35107/U$1 ( \4147 , \3943 );
nand \mul_7_15_g34845/U$1 ( \4148 , \4146 , \4147 );
nand \mul_7_15_g34705/U$1 ( \4149 , \4144 , \4148 );
nand \mul_7_15_g34461/U$1 ( \4150 , \4140 , \4149 );
nand \mul_7_15_g34251/U$1 ( \4151 , \4138 , \4150 );
nand \mul_7_15_g34023/U$1 ( \4152 , \4107 , \4151 );
not \mul_7_15_g34136/U$1 ( \4153 , \4105 );
nand \mul_7_15_g34067/U$1 ( \4154 , \4153 , \4071 );
nand \mul_7_15_g33995/U$1 ( \4155 , \4152 , \4154 );
buf \mul_7_15_g35098/U$1 ( \4156 , \3108 );
nand \mul_7_15_g34832/U$1 ( \4157 , \4156 , \4046 );
not \mul_7_15_g34263/U$3 ( \4158 , \4136 );
not \mul_7_15_g34263/U$4 ( \4159 , \4149 );
or \mul_7_15_g34263/U$2 ( \4160 , \4158 , \4159 );
not \mul_7_15_g34727/U$3 ( \4161 , \4044 );
not \mul_7_15_g34727/U$4 ( \4162 , \4110 );
or \mul_7_15_g34727/U$2 ( \4163 , \4161 , \4162 );
nand \mul_7_15_g34853/U$1 ( \4164 , \4109 , \4092 );
nand \mul_7_15_g34727/U$1 ( \4165 , \4163 , \4164 );
nand \mul_7_15_g34391/U$1 ( \4166 , \4140 , \4165 );
nand \mul_7_15_g34263/U$1 ( \4167 , \4160 , \4166 );
not \mul_7_15_g34259/U$1 ( \4168 , \4167 );
xor \mul_7_15_g33978/U$1 ( \4169 , \4157 , \4168 );
not \mul_7_15_g34785/U$3 ( \4170 , \4047 );
buf \mul_7_15_g35140/U$1 ( \4171 , \3208 );
buf \mul_7_15_g35132/U$1 ( \4172 , \4171 );
not \mul_7_15_g35127/U$1 ( \4173 , \4172 );
not \mul_7_15_g34785/U$4 ( \4174 , \4173 );
or \mul_7_15_g34785/U$2 ( \4175 , \4170 , \4174 );
not \mul_7_15_g35116/U$1 ( \4176 , \4171 );
not \mul_7_15_g35115/U$1 ( \4177 , \4176 );
not \mul_7_15_g35057/U$1 ( \4178 , \4047 );
nand \mul_7_15_g34863/U$1 ( \4179 , \4177 , \4178 );
nand \mul_7_15_g34785/U$1 ( \4180 , \4175 , \4179 );
not \mul_7_15_g34121/U$3 ( \4181 , \4180 );
and \mul_7_15_g34569/U$2 ( \4182 , \3487 , \4171 );
not \mul_7_15_g34569/U$4 ( \4183 , \3487 );
not \mul_7_15_g35139/U$1 ( \4184 , \4171 );
and \mul_7_15_g34569/U$3 ( \4185 , \4183 , \4184 );
nor \mul_7_15_g34569/U$1 ( \4186 , \4182 , \4185 );
not \fopt35547/U$1 ( \4187 , \3745 );
and \mul_7_15_g34634/U$2 ( \4188 , \4187 , \3487 );
not \mul_7_15_g34634/U$4 ( \4189 , \4187 );
not \fopt35574/U$1 ( \4190 , \3487 );
and \mul_7_15_g34634/U$3 ( \4191 , \4189 , \4190 );
nor \mul_7_15_g34634/U$1 ( \4192 , \4188 , \4191 );
nand \mul_7_15_g34509/U$1 ( \4193 , \4186 , \4192 );
not \mul_7_15_g34508/U$1 ( \4194 , \4193 );
buf \mul_7_15_g34506/U$1 ( \4195 , \4194 );
not \mul_7_15_g34121/U$4 ( \4196 , \4195 );
or \mul_7_15_g34121/U$2 ( \4197 , \4181 , \4196 );
and \mul_7_15_g34734/U$2 ( \4198 , \4116 , \4172 );
not \mul_7_15_g34734/U$4 ( \4199 , \4116 );
and \mul_7_15_g34734/U$3 ( \4200 , \4199 , \4173 );
nor \mul_7_15_g34734/U$1 ( \4201 , \4198 , \4200 );
not \mul_7_15_g35335/U$2 ( \4202 , \4201 );
buf \mul_7_15_g34632/U$1 ( \4203 , \4192 );
not \mul_7_15_g34629/U$1 ( \4204 , \4203 );
buf \mul_7_15_g34628/U$1 ( \4205 , \4204 );
nand \mul_7_15_g35335/U$1 ( \4206 , \4202 , \4205 );
nand \mul_7_15_g34121/U$1 ( \4207 , \4197 , \4206 );
xnor \mul_7_15_g33978/U$1_r1 ( \4208 , \4169 , \4207 );
xor \mul_7_15_g33719/U$4 ( \4209 , \4155 , \4208 );
not \mul_7_15_g34783/U$3 ( \4210 , \4043 );
not \mul_7_15_g35075/U$1 ( \4211 , \3577 );
buf \mul_7_15_g35074/U$1 ( \4212 , \4211 );
buf \mul_7_15_g35069/U$1 ( \4213 , \4212 );
not \mul_7_15_g34783/U$4 ( \4214 , \4213 );
or \mul_7_15_g34783/U$2 ( \4215 , \4210 , \4214 );
not \mul_7_15_g35071/U$1 ( \4216 , \4212 );
not \mul_7_15_g35058/U$1 ( \4217 , \4043 );
nand \mul_7_15_g34913/U$1 ( \4218 , \4216 , \4217 );
nand \mul_7_15_g34783/U$1 ( \4219 , \4215 , \4218 );
not \mul_7_15_g34219/U$3 ( \4220 , \4219 );
xor \g35897/U$1 ( \4221 , \3208 , \3818 );
not \mul_7_15_g34409/U$2 ( \4222 , \4221 );
not \mul_7_15_g34635/U$3 ( \4223 , \3577 );
not \mul_7_15_g35034/U$1 ( \4224 , \3818 );
not \mul_7_15_g34635/U$4 ( \4225 , \4224 );
or \mul_7_15_g34635/U$2 ( \4226 , \4223 , \4225 );
not \mul_7_15_g35339/U$2 ( \4227 , \3577 );
nand \mul_7_15_g35339/U$1 ( \4228 , \4227 , \3818 );
nand \mul_7_15_g34635/U$1 ( \4229 , \4226 , \4228 );
nand \mul_7_15_g34409/U$1 ( \4230 , \4222 , \4229 );
not \mul_7_15_g34408/U$1 ( \4231 , \4230 );
not \mul_7_15_g34219/U$4 ( \4232 , \4231 );
or \mul_7_15_g34219/U$2 ( \4233 , \4220 , \4232 );
buf \mul_7_15_g34591/U$1 ( \4234 , \4221 );
not \mul_7_15_g34701/U$3 ( \4235 , \4041 );
not \mul_7_15_g34701/U$4 ( \4236 , \4213 );
or \mul_7_15_g34701/U$2 ( \4237 , \4235 , \4236 );
not \mul_7_15_g35007/U$1 ( \4238 , \4041 );
nand \mul_7_15_g34923/U$1 ( \4239 , \4216 , \4238 );
nand \mul_7_15_g34701/U$1 ( \4240 , \4237 , \4239 );
nand \mul_7_15_g34491/U$1 ( \4241 , \4234 , \4240 );
nand \mul_7_15_g34219/U$1 ( \4242 , \4233 , \4241 );
not \mul_7_15_g34007/U$3 ( \4243 , \4242 );
not \mul_7_15_g34954/U$1 ( \4244 , \3366 );
not \mul_7_15_g34953/U$1 ( \4245 , \4244 );
not \mul_7_15_g34570/U$3 ( \4246 , \4245 );
not \mul_7_15_g35082/U$1 ( \4247 , \3108 );
not \mul_7_15_g34570/U$4 ( \4248 , \4247 );
or \mul_7_15_g34570/U$2 ( \4249 , \4246 , \4248 );
nand \mul_7_15_g34820/U$1 ( \4250 , \3108 , \4244 );
nand \mul_7_15_g34570/U$1 ( \4251 , \4249 , \4250 );
xnor \g35430/U$1 ( \4252 , \3577 , \3366 );
and \mul_7_15_g34419/U$1 ( \4253 , \4251 , \4252 );
not \mul_7_15_g34418/U$1 ( \4254 , \4253 );
not \mul_7_15_g34165/U$3 ( \4255 , \4254 );
not \mul_7_15_g34947/U$1 ( \4256 , \4046 );
not \mul_7_15_g34663/U$3 ( \4257 , \4256 );
not \mul_7_15_g34663/U$4 ( \4258 , \4156 );
or \mul_7_15_g34663/U$2 ( \4259 , \4257 , \4258 );
not \mul_7_15_g35103/U$1 ( \4260 , \3108 );
nand \mul_7_15_g34865/U$1 ( \4261 , \4260 , \4046 );
nand \mul_7_15_g34663/U$1 ( \4262 , \4259 , \4261 );
not \mul_7_15_g34552/U$1 ( \4263 , \4262 );
not \mul_7_15_g34165/U$4 ( \4264 , \4263 );
and \mul_7_15_g34165/U$2 ( \4265 , \4255 , \4264 );
not \mul_7_15_g34667/U$3 ( \4266 , \4011 );
not \mul_7_15_g35084/U$1 ( \4267 , \4156 );
not \mul_7_15_g34667/U$4 ( \4268 , \4267 );
or \mul_7_15_g34667/U$2 ( \4269 , \4266 , \4268 );
not \mul_7_15_g34948/U$1 ( \4270 , \4011 );
nand \mul_7_15_g34852/U$1 ( \4271 , \4156 , \4270 );
nand \mul_7_15_g34667/U$1 ( \4272 , \4269 , \4271 );
not \mul_7_15_g34644/U$1 ( \4273 , \4252 );
buf \mul_7_15_g34643/U$1 ( \4274 , \4273 );
and \mul_7_15_g35329/U$1 ( \4275 , \4272 , \4274 );
nor \mul_7_15_g34165/U$1 ( \4276 , \4265 , \4275 );
not \mul_7_15_g34164/U$1 ( \4277 , \4276 );
not \mul_7_15_g34007/U$4 ( \4278 , \4277 );
or \mul_7_15_g34007/U$2 ( \4279 , \4243 , \4278 );
or \mul_7_15_g34016/U$2 ( \4280 , \4277 , \4242 );
not \mul_7_15_g34781/U$3 ( \4281 , \4045 );
not \mul_7_15_g34781/U$4 ( \4282 , \4176 );
or \mul_7_15_g34781/U$2 ( \4283 , \4281 , \4282 );
not \mul_7_15_g35135/U$1 ( \4284 , \4171 );
not \mul_7_15_g35133/U$1 ( \4285 , \4284 );
not \mul_7_15_g35029/U$1 ( \4286 , \4045 );
nand \mul_7_15_g34932/U$1 ( \4287 , \4285 , \4286 );
nand \mul_7_15_g34781/U$1 ( \4288 , \4283 , \4287 );
not \mul_7_15_g34117/U$3 ( \4289 , \4288 );
not \mul_7_15_g34117/U$4 ( \4290 , \4195 );
or \mul_7_15_g34117/U$2 ( \4291 , \4289 , \4290 );
nand \mul_7_15_g34494/U$1 ( \4292 , \4205 , \4180 );
nand \mul_7_15_g34117/U$1 ( \4293 , \4291 , \4292 );
nand \mul_7_15_g34016/U$1 ( \4294 , \4280 , \4293 );
nand \mul_7_15_g34007/U$1 ( \4295 , \4279 , \4294 );
and \mul_7_15_g33719/U$3 ( \4296 , \4209 , \4295 );
and \mul_7_15_g33719/U$5 ( \4297 , \4155 , \4208 );
or \mul_7_15_g33719/U$2 ( \4298 , \4296 , \4297 );
not \mul_7_15_g34028/U$3 ( \4299 , \4157 );
not \mul_7_15_g34028/U$4 ( \4300 , \4167 );
or \mul_7_15_g34028/U$2 ( \4301 , \4299 , \4300 );
nand \mul_7_15_g34028/U$1 ( \4302 , \4301 , \4207 );
not \mul_7_15_g35330/U$2 ( \4303 , \4157 );
nand \mul_7_15_g35330/U$1 ( \4304 , \4303 , \4168 );
nand \mul_7_15_g34010/U$1 ( \4305 , \4302 , \4304 );
not \mul_7_15_g34009/U$1 ( \4306 , \4305 );
and \mul_7_15_g34831/U$1 ( \4307 , \4156 , \4011 );
not \mul_7_15_g35102/U$1 ( \4308 , \4260 );
xor \mul_7_15_g34546/U$1 ( \4309 , \4043 , \4308 );
not \mul_7_15_g34186/U$3 ( \4310 , \4309 );
not \mul_7_15_g34186/U$4 ( \4311 , \4253 );
or \mul_7_15_g34186/U$2 ( \4312 , \4310 , \4311 );
xor \mul_7_15_g34549/U$1 ( \4313 , \4041 , \4156 );
nand \mul_7_15_g34298/U$1 ( \4314 , \4313 , \4274 );
nand \mul_7_15_g34186/U$1 ( \4315 , \4312 , \4314 );
xor \mul_7_15_g33917/U$1 ( \4316 , \4307 , \4315 );
not \mul_7_15_g34503/U$1 ( \4317 , \4195 );
or \mul_7_15_g34114/U$2 ( \4318 , \4317 , \4201 );
not \mul_7_15_g34626/U$1 ( \4319 , \4205 );
and \mul_7_15_g34708/U$2 ( \4320 , \4147 , \4172 );
not \mul_7_15_g34708/U$4 ( \4321 , \4147 );
and \mul_7_15_g34708/U$3 ( \4322 , \4321 , \4173 );
nor \mul_7_15_g34708/U$1 ( \4323 , \4320 , \4322 );
or \mul_7_15_g34114/U$3 ( \4324 , \4319 , \4323 );
nand \mul_7_15_g34114/U$1 ( \4325 , \4318 , \4324 );
xor \mul_7_15_g33917/U$1_r1 ( \4326 , \4316 , \4325 );
xor \g35380/U$1 ( \4327 , \4306 , \4326 );
not \mul_7_15_g34292/U$3 ( \4328 , \4101 );
not \mul_7_15_g34292/U$4 ( \4329 , \4086 );
or \mul_7_15_g34292/U$2 ( \4330 , \4328 , \4329 );
not \fopt35516/U$1 ( \4331 , \4103 );
nand \mul_7_15_g34528/U$1 ( \4332 , \4331 , \4088 );
nand \mul_7_15_g34292/U$1 ( \4333 , \4330 , \4332 );
not \mul_7_15_g33997/U$3 ( \4334 , \4333 );
not \mul_7_15_g34191/U$3 ( \4335 , \4240 );
not \mul_7_15_g34191/U$4 ( \4336 , \4231 );
or \mul_7_15_g34191/U$2 ( \4337 , \4335 , \4336 );
not \mul_7_15_g34744/U$3 ( \4338 , \4045 );
not \mul_7_15_g34744/U$4 ( \4339 , \4212 );
or \mul_7_15_g34744/U$2 ( \4340 , \4338 , \4339 );
nand \mul_7_15_g34893/U$1 ( \4341 , \4216 , \4286 );
nand \mul_7_15_g34744/U$1 ( \4342 , \4340 , \4341 );
nand \mul_7_15_g34460/U$1 ( \4343 , \4234 , \4342 );
nand \mul_7_15_g34191/U$1 ( \4344 , \4337 , \4343 );
not \mul_7_15_g33997/U$4 ( \4345 , \4344 );
or \mul_7_15_g33997/U$2 ( \4346 , \4334 , \4345 );
or \mul_7_15_g34025/U$2 ( \4347 , \4344 , \4333 );
not \mul_7_15_g34195/U$3 ( \4348 , \4272 );
not \mul_7_15_g34195/U$4 ( \4349 , \4253 );
or \mul_7_15_g34195/U$2 ( \4350 , \4348 , \4349 );
nand \mul_7_15_g34306/U$1 ( \4351 , \4274 , \4309 );
nand \mul_7_15_g34195/U$1 ( \4352 , \4350 , \4351 );
nand \mul_7_15_g34025/U$1 ( \4353 , \4347 , \4352 );
nand \mul_7_15_g33997/U$1 ( \4354 , \4346 , \4353 );
xor \mul_7_15_g33781/U$1 ( \4355 , \4168 , \4354 );
not \mul_7_15_g34622/U$1 ( \4356 , \4084 );
not \mul_7_15_g34310/U$3 ( \4357 , \4356 );
not \mul_7_15_g34310/U$4 ( \4358 , \4103 );
or \mul_7_15_g34310/U$2 ( \4359 , \4357 , \4358 );
nand \mul_7_15_g34310/U$1 ( \4360 , \4359 , \4088 );
not \mul_7_15_g34309/U$1 ( \4361 , \4360 );
not \mul_7_15_g34255/U$3 ( \4362 , \4165 );
not \mul_7_15_g34255/U$4 ( \4363 , \4136 );
or \mul_7_15_g34255/U$2 ( \4364 , \4362 , \4363 );
not \mul_7_15_g34671/U$3 ( \4365 , \3994 );
not \mul_7_15_g34671/U$4 ( \4366 , \4142 );
or \mul_7_15_g34671/U$2 ( \4367 , \4365 , \4366 );
not \fopt35558/U$1 ( \4368 , \4142 );
nand \mul_7_15_g34841/U$1 ( \4369 , \4368 , \4099 );
nand \mul_7_15_g34671/U$1 ( \4370 , \4367 , \4369 );
nand \mul_7_15_g34376/U$1 ( \4371 , \4140 , \4370 );
nand \mul_7_15_g34255/U$1 ( \4372 , \4364 , \4371 );
xor \mul_7_15_g33905/U$1 ( \4373 , \4361 , \4372 );
not \mul_7_15_g34178/U$3 ( \4374 , \4342 );
not \mul_7_15_g34178/U$4 ( \4375 , \4231 );
or \mul_7_15_g34178/U$2 ( \4376 , \4374 , \4375 );
buf \mul_7_15_g34589/U$1 ( \4377 , \4234 );
not \mul_7_15_g34756/U$3 ( \4378 , \4047 );
not \mul_7_15_g34756/U$4 ( \4379 , \4212 );
or \mul_7_15_g34756/U$2 ( \4380 , \4378 , \4379 );
nand \mul_7_15_g34849/U$1 ( \4381 , \4216 , \4178 );
nand \mul_7_15_g34756/U$1 ( \4382 , \4380 , \4381 );
nand \mul_7_15_g34459/U$1 ( \4383 , \4377 , \4382 );
nand \mul_7_15_g34178/U$1 ( \4384 , \4376 , \4383 );
xnor \mul_7_15_g33905/U$1_r1 ( \4385 , \4373 , \4384 );
xnor \mul_7_15_g33781/U$1_r1 ( \4386 , \4355 , \4385 );
xnor \g35380/U$1_r1 ( \4387 , \4327 , \4386 );
xor \mul_7_15_g33493/U$1 ( \4388 , \4298 , \4387 );
and \mul_7_15_g34031/U$2 ( \4389 , \4352 , \4333 );
not \mul_7_15_g34031/U$4 ( \4390 , \4352 );
not \mul_7_15_g34291/U$1 ( \4391 , \4333 );
and \mul_7_15_g34031/U$3 ( \4392 , \4390 , \4391 );
nor \mul_7_15_g34031/U$1 ( \4393 , \4389 , \4392 );
buf \mul_7_15_g34190/U$1 ( \4394 , \4344 );
xnor \g35835/U$1 ( \4395 , \4393 , \4394 );
not \mul_7_15_g33950/U$1 ( \4396 , \4395 );
not \mul_7_15_g33614/U$3 ( \4397 , \4396 );
not \g35942/U$3 ( \4398 , \4056 );
not \mul_7_15_fopt35186/U$1 ( \4399 , \4070 );
not \g35942/U$4 ( \4400 , \4399 );
and \g35942/U$2 ( \4401 , \4398 , \4400 );
not \mul_7_15_g34675/U$3 ( \4402 , \3994 );
buf \mul_7_15_fopt35181/U$1 ( \4403 , \3880 );
not \mul_7_15_fopt35179/U$1 ( \4404 , \4403 );
not \mul_7_15_g34675/U$4 ( \4405 , \4404 );
or \mul_7_15_g34675/U$2 ( \4406 , \4402 , \4405 );
not \mul_7_15_fopt35183/U$1 ( \4407 , \4069 );
nand \mul_7_15_g35971/U$1 ( \4408 , \4407 , \4099 );
nand \mul_7_15_g34675/U$1 ( \4409 , \4406 , \4408 );
not \g35943/U$2 ( \4410 , \4409 );
not \fopt35522/U$1 ( \4411 , \4065 );
nor \g35943/U$1 ( \4412 , \4410 , \4411 );
nor \g35942/U$1 ( \4413 , \4401 , \4412 );
not \mul_7_15_g34287/U$1 ( \4414 , \4413 );
not \g35616/U$2 ( \4415 , \4414 );
nand \mul_7_15_g34830/U$1 ( \4416 , \4156 , \3958 );
nand \g35616/U$1 ( \4417 , \4415 , \4416 );
not \g35615/U$3 ( \4418 , \4417 );
not \mul_7_15_g34694/U$3 ( \4419 , \4047 );
not \mul_7_15_g34694/U$4 ( \4420 , \4110 );
or \mul_7_15_g34694/U$2 ( \4421 , \4419 , \4420 );
nand \mul_7_15_g34919/U$1 ( \4422 , \4109 , \4178 );
nand \mul_7_15_g34694/U$1 ( \4423 , \4421 , \4422 );
not \mul_7_15_g34249/U$3 ( \4424 , \4423 );
not \mul_7_15_g34447/U$1 ( \4425 , \4135 );
not \mul_7_15_g34249/U$4 ( \4426 , \4425 );
or \mul_7_15_g34249/U$2 ( \4427 , \4424 , \4426 );
not \mul_7_15_g34599/U$1 ( \4428 , \4139 );
not \mul_7_15_g34597/U$1 ( \4429 , \4428 );
nand \mul_7_15_g34382/U$1 ( \4430 , \4118 , \4429 );
nand \mul_7_15_g34249/U$1 ( \4431 , \4427 , \4430 );
and \mul_7_15_g34711/U$2 ( \4432 , \3943 , \4088 );
not \mul_7_15_g34711/U$4 ( \4433 , \3943 );
and \mul_7_15_g34711/U$3 ( \4434 , \4433 , \4089 );
nor \mul_7_15_g34711/U$1 ( \4435 , \4432 , \4434 );
not \mul_7_15_g34139/U$3 ( \4436 , \4435 );
buf \mul_7_15_g34466/U$1 ( \4437 , \4085 );
not \mul_7_15_g34139/U$4 ( \4438 , \4437 );
or \mul_7_15_g34139/U$2 ( \4439 , \4436 , \4438 );
nand \mul_7_15_g34355/U$1 ( \4440 , \4331 , \4094 );
nand \mul_7_15_g34139/U$1 ( \4441 , \4439 , \4440 );
xor \mul_7_15_g33893/U$4 ( \4442 , \4431 , \4441 );
and \mul_7_15_g34700/U$2 ( \4443 , \4041 , \4285 );
not \mul_7_15_g34700/U$4 ( \4444 , \4041 );
and \mul_7_15_g34700/U$3 ( \4445 , \4444 , \4176 );
nor \mul_7_15_g34700/U$1 ( \4446 , \4443 , \4445 );
not \mul_7_15_g34113/U$3 ( \4447 , \4446 );
not \mul_7_15_g34113/U$4 ( \4448 , \4195 );
or \mul_7_15_g34113/U$2 ( \4449 , \4447 , \4448 );
nand \mul_7_15_g34410/U$1 ( \4450 , \4205 , \4288 );
nand \mul_7_15_g34113/U$1 ( \4451 , \4449 , \4450 );
and \mul_7_15_g33893/U$3 ( \4452 , \4442 , \4451 );
and \mul_7_15_g33893/U$5 ( \4453 , \4431 , \4441 );
or \mul_7_15_g33893/U$2 ( \4454 , \4452 , \4453 );
not \g35615/U$4 ( \4455 , \4454 );
or \g35615/U$2 ( \4456 , \4418 , \4455 );
not \mul_7_15_g34076/U$2 ( \4457 , \4416 );
nand \mul_7_15_g34076/U$1 ( \4458 , \4457 , \4414 );
nand \g35615/U$1 ( \4459 , \4456 , \4458 );
not \mul_7_15_g33614/U$4 ( \4460 , \4459 );
or \mul_7_15_g33614/U$2 ( \4461 , \4397 , \4460 );
not \mul_7_15_g34218/U$1 ( \4462 , \4242 );
xor \g35709/U$1 ( \4463 , \4293 , \4462 );
xor \g35709/U$1_r1 ( \4464 , \4463 , \4276 );
and \g35397/U$2 ( \4465 , \4151 , \4072 );
not \g35397/U$4 ( \4466 , \4151 );
and \g35397/U$3 ( \4467 , \4466 , \4071 );
or \g35397/U$1 ( \4468 , \4465 , \4467 );
and \g35396/U$2 ( \4469 , \4468 , \4105 );
not \g35396/U$4 ( \4470 , \4468 );
and \g35396/U$3 ( \4471 , \4470 , \4153 );
nor \g35396/U$1 ( \4472 , \4469 , \4471 );
not \mul_7_15_g35174/U$1 ( \4473 , \3958 );
not \mul_7_15_g34665/U$3 ( \4474 , \4473 );
not \mul_7_15_g34665/U$4 ( \4475 , \4156 );
or \mul_7_15_g34665/U$2 ( \4476 , \4474 , \4475 );
nand \mul_7_15_g34937/U$1 ( \4477 , \4267 , \3958 );
nand \mul_7_15_g34665/U$1 ( \4478 , \4476 , \4477 );
not \mul_7_15_g34174/U$3 ( \4479 , \4478 );
and \mul_7_15_g34420/U$1 ( \4480 , \4251 , \4252 );
not \mul_7_15_g34174/U$4 ( \4481 , \4480 );
or \mul_7_15_g34174/U$2 ( \4482 , \4479 , \4481 );
nand \mul_7_15_g34297/U$1 ( \4483 , \4262 , \4273 );
nand \mul_7_15_g34174/U$1 ( \4484 , \4482 , \4483 );
not \mul_7_15_g34834/U$2 ( \4485 , \4156 );
not \mul_7_15_g35028/U$1 ( \4486 , \3963 );
nor \mul_7_15_g34834/U$1 ( \4487 , \4485 , \4486 );
nor \mul_7_15_g34056/U$1 ( \4488 , \4484 , \4487 );
not \mul_7_15_g34714/U$3 ( \4489 , \4011 );
not \mul_7_15_g34714/U$4 ( \4490 , \4212 );
or \mul_7_15_g34714/U$2 ( \4491 , \4489 , \4490 );
buf \mul_7_15_g35080/U$1 ( \4492 , \3577 );
nand \mul_7_15_g34844/U$1 ( \4493 , \4492 , \4270 );
nand \mul_7_15_g34714/U$1 ( \4494 , \4491 , \4493 );
not \mul_7_15_g34183/U$3 ( \4495 , \4494 );
buf \mul_7_15_g34404/U$1 ( \4496 , \4231 );
not \mul_7_15_g34183/U$4 ( \4497 , \4496 );
or \mul_7_15_g34183/U$2 ( \4498 , \4495 , \4497 );
nand \mul_7_15_g34458/U$1 ( \4499 , \4377 , \4219 );
nand \mul_7_15_g34183/U$1 ( \4500 , \4498 , \4499 );
not \mul_7_15_g34182/U$1 ( \4501 , \4500 );
or \mul_7_15_g33998/U$2 ( \4502 , \4488 , \4501 );
nand \mul_7_15_g34054/U$1 ( \4503 , \4484 , \4487 );
nand \mul_7_15_g33998/U$1 ( \4504 , \4502 , \4503 );
not \mul_7_15_g33948/U$1 ( \4505 , \4504 );
nand \mul_7_15_g33867/U$1 ( \4506 , \4472 , \4505 );
and \mul_7_15_g33741/U$2 ( \4507 , \4464 , \4506 );
nor \mul_7_15_g33875/U$1 ( \4508 , \4472 , \4505 );
nor \mul_7_15_g33741/U$1 ( \4509 , \4507 , \4508 );
not \fopt35576/U$1 ( \4510 , \4509 );
not \mul_7_15_g33733/U$2 ( \4511 , \4459 );
nand \mul_7_15_g33733/U$1 ( \4512 , \4511 , \4395 );
nand \mul_7_15_g33641/U$1 ( \4513 , \4510 , \4512 );
nand \mul_7_15_g33614/U$1 ( \4514 , \4461 , \4513 );
xor \mul_7_15_g33493/U$1_r1 ( \4515 , \4388 , \4514 );
not \mul_7_15_g33491/U$1 ( \4516 , \4515 );
xor \mul_7_15_g33719/U$1 ( \4517 , \4155 , \4208 );
xor \mul_7_15_g33719/U$1_r1 ( \4518 , \4517 , \4295 );
not \mul_7_15_g33471/U$3 ( \4519 , \4518 );
not \mul_7_15_g35813/U$3 ( \4520 , \4510 );
not \mul_7_15_g33726/U$3 ( \4521 , \4395 );
not \mul_7_15_g33726/U$4 ( \4522 , \4459 );
or \mul_7_15_g33726/U$2 ( \4523 , \4521 , \4522 );
or \mul_7_15_g33726/U$5 ( \4524 , \4459 , \4395 );
nand \mul_7_15_g33726/U$1 ( \4525 , \4523 , \4524 );
not \mul_7_15_g33673/U$1 ( \4526 , \4525 );
not \mul_7_15_g35813/U$4 ( \4527 , \4526 );
or \mul_7_15_g35813/U$2 ( \4528 , \4520 , \4527 );
nand \mul_7_15_g33634/U$1 ( \4529 , \4525 , \4509 );
nand \mul_7_15_g35813/U$1 ( \4530 , \4528 , \4529 );
not \mul_7_15_g33471/U$4 ( \4531 , \4530 );
or \mul_7_15_g33471/U$2 ( \4532 , \4519 , \4531 );
or \mul_7_15_g33485/U$2 ( \4533 , \4530 , \4518 );
not \mul_7_15_g34573/U$3 ( \4534 , \1528 );
not \mul_7_15_g35172/U$1 ( \4535 , \3432 );
not \mul_7_15_g34573/U$4 ( \4536 , \4535 );
or \mul_7_15_g34573/U$2 ( \4537 , \4534 , \4536 );
not \mul_7_15_g35345/U$2 ( \4538 , \1528 );
nand \mul_7_15_g35345/U$1 ( \4539 , \4538 , \3432 );
nand \mul_7_15_g34573/U$1 ( \4540 , \4537 , \4539 );
buf \mul_7_15_g34572/U$1 ( \4541 , \4540 );
not \mul_7_15_g34571/U$1 ( \4542 , \4541 );
not \mul_7_15_g34312/U$3 ( \4543 , \4542 );
xnor \g35837/U$1 ( \4544 , \1395 , \3432 );
buf \mul_7_15_g34656/U$1 ( \4545 , \4544 );
not \mul_7_15_g34312/U$4 ( \4546 , \4545 );
or \mul_7_15_g34312/U$2 ( \4547 , \4543 , \4546 );
buf \mul_7_15_g35165/U$1 ( \4548 , \1528 );
nand \mul_7_15_g34312/U$1 ( \4549 , \4547 , \4548 );
buf \mul_7_15_g34311/U$1 ( \4550 , \4549 );
not \mul_7_15_g33904/U$3 ( \4551 , \4550 );
not \mul_7_15_g34768/U$3 ( \4552 , \4044 );
not \mul_7_15_g34768/U$4 ( \4553 , \4069 );
or \mul_7_15_g34768/U$2 ( \4554 , \4552 , \4553 );
nand \mul_7_15_g34906/U$1 ( \4555 , \4407 , \4092 );
nand \mul_7_15_g34768/U$1 ( \4556 , \4554 , \4555 );
not \mul_7_15_g34176/U$3 ( \4557 , \4556 );
and \mul_7_15_g35266/U$1 ( \4558 , \4063 , \4053 );
not \mul_7_15_g34176/U$4 ( \4559 , \4558 );
or \mul_7_15_g34176/U$2 ( \4560 , \4557 , \4559 );
buf \mul_7_15_g34577/U$1 ( \4561 , \4053 );
not \mul_7_15_g34576/U$1 ( \4562 , \4561 );
nand \mul_7_15_g34371/U$1 ( \4563 , \4562 , \4409 );
nand \mul_7_15_g34176/U$1 ( \4564 , \4560 , \4563 );
not \mul_7_15_g33904/U$4 ( \4565 , \4564 );
or \mul_7_15_g33904/U$2 ( \4566 , \4551 , \4565 );
or \mul_7_15_g33960/U$2 ( \4567 , \4550 , \4564 );
not \mul_7_15_g34763/U$3 ( \4568 , \4045 );
not \fopt35552/U$1 ( \4569 , \4109 );
not \mul_7_15_g34763/U$4 ( \4570 , \4569 );
or \mul_7_15_g34763/U$2 ( \4571 , \4568 , \4570 );
nand \mul_7_15_g34851/U$1 ( \4572 , \4109 , \4286 );
nand \mul_7_15_g34763/U$1 ( \4573 , \4571 , \4572 );
not \g35925/U$3 ( \4574 , \4573 );
not \g35925/U$4 ( \4575 , \4136 );
or \g35925/U$2 ( \4576 , \4574 , \4575 );
nand \mul_7_15_g34486/U$1 ( \4577 , \4429 , \4423 );
nand \g35925/U$1 ( \4578 , \4576 , \4577 );
nand \mul_7_15_g33960/U$1 ( \4579 , \4567 , \4578 );
nand \mul_7_15_g33904/U$1 ( \4580 , \4566 , \4579 );
not \g36017/U$2 ( \4581 , \4580 );
nand \g36017/U$1 ( \4582 , \4581 , \4414 );
not \g36016/U$3 ( \4583 , \4582 );
not \mul_7_15_g34829/U$2 ( \4584 , \4156 );
not \mul_7_15_g35175/U$1 ( \4585 , \4019 );
nor \mul_7_15_g34829/U$1 ( \4586 , \4584 , \4585 );
not \mul_7_15_g33899/U$3 ( \4587 , \4586 );
not \g35923/U$3 ( \4588 , \4042 );
not \g35923/U$4 ( \4589 , \4089 );
or \g35923/U$2 ( \4590 , \4588 , \4589 );
nand \mul_7_15_g34890/U$1 ( \4591 , \4088 , \4116 );
nand \g35923/U$1 ( \4592 , \4590 , \4591 );
not \mul_7_15_g34143/U$3 ( \4593 , \4592 );
not \mul_7_15_g34143/U$4 ( \4594 , \4437 );
or \mul_7_15_g34143/U$2 ( \4595 , \4593 , \4594 );
not \fopt35510/U$1 ( \4596 , \4103 );
nand \mul_7_15_g34374/U$1 ( \4597 , \4596 , \4435 );
nand \mul_7_15_g34143/U$1 ( \4598 , \4595 , \4597 );
not \mul_7_15_g33899/U$4 ( \4599 , \4598 );
or \mul_7_15_g33899/U$2 ( \4600 , \4587 , \4599 );
or \g35921/U$2 ( \4601 , \4598 , \4586 );
and \mul_7_15_g34771/U$2 ( \4602 , \4043 , \4172 );
not \mul_7_15_g34771/U$4 ( \4603 , \4043 );
and \mul_7_15_g34771/U$3 ( \4604 , \4603 , \4173 );
nor \mul_7_15_g34771/U$1 ( \4605 , \4602 , \4604 );
not \mul_7_15_g34116/U$3 ( \4606 , \4605 );
not \mul_7_15_g34116/U$4 ( \4607 , \4195 );
or \mul_7_15_g34116/U$2 ( \4608 , \4606 , \4607 );
nand \mul_7_15_g34363/U$1 ( \4609 , \4205 , \4446 );
nand \mul_7_15_g34116/U$1 ( \4610 , \4608 , \4609 );
nand \g35921/U$1 ( \4611 , \4601 , \4610 );
nand \mul_7_15_g33899/U$1 ( \4612 , \4600 , \4611 );
not \g36016/U$4 ( \4613 , \4612 );
or \g36016/U$2 ( \4614 , \4583 , \4613 );
not \g35848/U$2 ( \4615 , \4414 );
nand \g35848/U$1 ( \4616 , \4615 , \4580 );
nand \g36016/U$1 ( \4617 , \4614 , \4616 );
not \mul_7_15_g33635/U$2 ( \4618 , \4617 );
not \mul_7_15_g33803/U$3 ( \4619 , \4454 );
and \mul_7_15_g35319/U$2 ( \4620 , \4416 , \4414 );
not \mul_7_15_g35319/U$4 ( \4621 , \4416 );
and \mul_7_15_g35319/U$3 ( \4622 , \4621 , \4413 );
nor \mul_7_15_g35319/U$1 ( \4623 , \4620 , \4622 );
not \mul_7_15_g33803/U$4 ( \4624 , \4623 );
and \mul_7_15_g33803/U$2 ( \4625 , \4619 , \4624 );
and \mul_7_15_g33803/U$5 ( \4626 , \4454 , \4623 );
nor \mul_7_15_g33803/U$1 ( \4627 , \4625 , \4626 );
nand \mul_7_15_g33635/U$1 ( \4628 , \4618 , \4627 );
not \mul_7_15_g33538/U$3 ( \4629 , \4628 );
xor \mul_7_15_g33893/U$1 ( \4630 , \4431 , \4441 );
xor \mul_7_15_g33893/U$1_r1 ( \4631 , \4630 , \4451 );
not \g35606/U$2 ( \4632 , \4631 );
not \mul_7_15_g34014/U$2 ( \4633 , \4488 );
nand \mul_7_15_g34014/U$1 ( \4634 , \4633 , \4503 );
and \mul_7_15_g33967/U$2 ( \4635 , \4634 , \4500 );
not \mul_7_15_g33967/U$4 ( \4636 , \4634 );
and \mul_7_15_g33967/U$3 ( \4637 , \4636 , \4501 );
nor \mul_7_15_g33967/U$1 ( \4638 , \4635 , \4637 );
nand \g35606/U$1 ( \4639 , \4632 , \4638 );
not \mul_7_15_g34664/U$3 ( \4640 , \3963 );
not \mul_7_15_g34664/U$4 ( \4641 , \4260 );
or \mul_7_15_g34664/U$2 ( \4642 , \4640 , \4641 );
nand \mul_7_15_g34915/U$1 ( \4643 , \4156 , \4486 );
nand \mul_7_15_g34664/U$1 ( \4644 , \4642 , \4643 );
not \mul_7_15_g34181/U$3 ( \4645 , \4644 );
not \mul_7_15_g34181/U$4 ( \4646 , \4253 );
or \mul_7_15_g34181/U$2 ( \4647 , \4645 , \4646 );
nand \mul_7_15_g34301/U$1 ( \4648 , \4273 , \4478 );
nand \mul_7_15_g34181/U$1 ( \4649 , \4647 , \4648 );
not \mul_7_15_g34695/U$3 ( \4650 , \4046 );
not \mul_7_15_g34695/U$4 ( \4651 , \4212 );
or \mul_7_15_g34695/U$2 ( \4652 , \4650 , \4651 );
nand \mul_7_15_g34899/U$1 ( \4653 , \4492 , \4256 );
nand \mul_7_15_g34695/U$1 ( \4654 , \4652 , \4653 );
not \mul_7_15_g34185/U$3 ( \4655 , \4654 );
not \mul_7_15_g34185/U$4 ( \4656 , \4231 );
or \mul_7_15_g34185/U$2 ( \4657 , \4655 , \4656 );
nand \mul_7_15_g34352/U$1 ( \4658 , \4234 , \4494 );
nand \mul_7_15_g34185/U$1 ( \4659 , \4657 , \4658 );
or \mul_7_15_g34029/U$2 ( \4660 , \4649 , \4659 );
and \mul_7_15_g34400/U$1 ( \4661 , \4540 , \4544 );
buf \mul_7_15_g34399/U$1 ( \4662 , \4661 );
not \mul_7_15_g34398/U$1 ( \4663 , \4662 );
not \mul_7_15_g34282/U$3 ( \4664 , \4663 );
buf \mul_7_15_g35152/U$1 ( \4665 , \1528 );
not \mul_7_15_g35146/U$1 ( \4666 , \4665 );
and \mul_7_15_g34677/U$2 ( \4667 , \4666 , \3994 );
and \mul_7_15_g34677/U$3 ( \4668 , \4548 , \4099 );
nor \mul_7_15_g34677/U$1 ( \4669 , \4667 , \4668 );
not \mul_7_15_g34282/U$4 ( \4670 , \4669 );
and \mul_7_15_g34282/U$2 ( \4671 , \4664 , \4670 );
not \mul_7_15_g34654/U$1 ( \4672 , \4545 );
not \mul_7_15_g35332/U$2 ( \4673 , \4672 );
nor \mul_7_15_g35332/U$1 ( \4674 , \4673 , \4666 );
nor \mul_7_15_g34282/U$1 ( \4675 , \4671 , \4674 );
not \mul_7_15_g34281/U$1 ( \4676 , \4675 );
nand \mul_7_15_g34029/U$1 ( \4677 , \4660 , \4676 );
nand \mul_7_15_g34059/U$1 ( \4678 , \4659 , \4649 );
and \mul_7_15_g33994/U$1 ( \4679 , \4677 , \4678 );
not \mul_7_15_g33946/U$1 ( \4680 , \4679 );
and \mul_7_15_g33780/U$2 ( \4681 , \4639 , \4680 );
not \mul_7_15_g35607/U$1 ( \4682 , \4631 );
nor \mul_7_15_g33825/U$1 ( \4683 , \4638 , \4682 );
nor \mul_7_15_g33780/U$1 ( \4684 , \4681 , \4683 );
not \fopt35541/U$1 ( \4685 , \4684 );
not \mul_7_15_g33538/U$4 ( \4686 , \4685 );
or \mul_7_15_g33538/U$2 ( \4687 , \4629 , \4686 );
not \mul_7_15_g35293/U$2 ( \4688 , \4627 );
nand \mul_7_15_g35293/U$1 ( \4689 , \4688 , \4617 );
nand \mul_7_15_g33538/U$1 ( \4690 , \4687 , \4689 );
nand \mul_7_15_g33485/U$1 ( \4691 , \4533 , \4690 );
nand \mul_7_15_g33471/U$1 ( \4692 , \4532 , \4691 );
not \mul_7_15_g33457/U$1 ( \4693 , \4692 );
nand \mul_7_15_g33413/U$1 ( \4694 , \4516 , \4693 );
xor \mul_7_15_g33493/U$4 ( \4695 , \4298 , \4387 );
and \mul_7_15_g33493/U$3 ( \4696 , \4695 , \4514 );
and \mul_7_15_g33493/U$5 ( \4697 , \4298 , \4387 );
or \mul_7_15_g33493/U$2 ( \4698 , \4696 , \4697 );
not \mul_7_15_g33492/U$1 ( \4699 , \4698 );
not \mul_7_15_g34202/U$3 ( \4700 , \4382 );
not \mul_7_15_g34202/U$4 ( \4701 , \4496 );
or \mul_7_15_g34202/U$2 ( \4702 , \4700 , \4701 );
not \mul_7_15_g34720/U$3 ( \4703 , \4042 );
not \mul_7_15_g34720/U$4 ( \4704 , \4212 );
or \mul_7_15_g34720/U$2 ( \4705 , \4703 , \4704 );
nand \mul_7_15_g34850/U$1 ( \4706 , \4216 , \4116 );
nand \mul_7_15_g34720/U$1 ( \4707 , \4705 , \4706 );
nand \mul_7_15_g34345/U$1 ( \4708 , \4377 , \4707 );
nand \mul_7_15_g34202/U$1 ( \4709 , \4702 , \4708 );
not \mul_7_15_g34280/U$3 ( \4710 , \4370 );
not \mul_7_15_g34280/U$4 ( \4711 , \4136 );
or \mul_7_15_g34280/U$2 ( \4712 , \4710 , \4711 );
not \g35847/U$2 ( \4713 , \4110 );
nand \g35847/U$1 ( \4714 , \4713 , \4140 );
nand \mul_7_15_g34280/U$1 ( \4715 , \4712 , \4714 );
not \mul_7_15_g34279/U$1 ( \4716 , \4715 );
xor \mul_7_15_g33817/U$1 ( \4717 , \4709 , \4716 );
xor \mul_7_15_g33917/U$4 ( \4718 , \4307 , \4315 );
and \mul_7_15_g33917/U$3 ( \4719 , \4718 , \4325 );
and \mul_7_15_g33917/U$5 ( \4720 , \4307 , \4315 );
or \mul_7_15_g33917/U$2 ( \4721 , \4719 , \4720 );
xor \mul_7_15_g33817/U$1_r1 ( \4722 , \4717 , \4721 );
not \mul_7_15_g33664/U$3 ( \4723 , \4386 );
not \mul_7_15_g35349/U$2 ( \4724 , \4326 );
nand \mul_7_15_g35349/U$1 ( \4725 , \4724 , \4306 );
not \mul_7_15_g33664/U$4 ( \4726 , \4725 );
or \mul_7_15_g33664/U$2 ( \4727 , \4723 , \4726 );
nand \mul_7_15_g33873/U$1 ( \4728 , \4326 , \4305 );
nand \mul_7_15_g33664/U$1 ( \4729 , \4727 , \4728 );
xor \mul_7_15_g33490/U$1 ( \4730 , \4722 , \4729 );
not \mul_7_15_g34072/U$2 ( \4731 , \4372 );
nand \mul_7_15_g34072/U$1 ( \4732 , \4731 , \4361 );
nand \mul_7_15_g33961/U$1 ( \4733 , \4732 , \4384 );
not \mul_7_15_g34071/U$2 ( \4734 , \4361 );
nand \mul_7_15_g34071/U$1 ( \4735 , \4734 , \4372 );
and \mul_7_15_g33903/U$1 ( \4736 , \4733 , \4735 );
and \mul_7_15_g34546/U$2 ( \4737 , \4043 , \4308 );
not \mul_7_15_g34167/U$3 ( \4738 , \4313 );
not \mul_7_15_g34167/U$4 ( \4739 , \4253 );
or \mul_7_15_g34167/U$2 ( \4740 , \4738 , \4739 );
xor \mul_7_15_g34550/U$1 ( \4741 , \4045 , \4156 );
buf \mul_7_15_g34641/U$1 ( \4742 , \4273 );
nand \mul_7_15_g34294/U$1 ( \4743 , \4741 , \4742 );
nand \mul_7_15_g34167/U$1 ( \4744 , \4740 , \4743 );
xor \mul_7_15_g33920/U$1 ( \4745 , \4737 , \4744 );
not \mul_7_15_g34707/U$1 ( \4746 , \4323 );
not \mul_7_15_g34111/U$3 ( \4747 , \4746 );
not \mul_7_15_g34111/U$4 ( \4748 , \4195 );
or \mul_7_15_g34111/U$2 ( \4749 , \4747 , \4748 );
not \mul_7_15_g34719/U$3 ( \4750 , \4044 );
not \mul_7_15_g34719/U$4 ( \4751 , \4173 );
or \mul_7_15_g34719/U$2 ( \4752 , \4750 , \4751 );
nand \mul_7_15_g34858/U$1 ( \4753 , \4172 , \4092 );
nand \mul_7_15_g34719/U$1 ( \4754 , \4752 , \4753 );
nand \mul_7_15_g34344/U$1 ( \4755 , \4205 , \4754 );
nand \mul_7_15_g34111/U$1 ( \4756 , \4749 , \4755 );
xor \mul_7_15_g33920/U$1_r1 ( \4757 , \4745 , \4756 );
xor \g35887/U$1 ( \4758 , \4736 , \4757 );
or \mul_7_15_g33799/U$2 ( \4759 , \4385 , \4167 );
nand \mul_7_15_g33799/U$1 ( \4760 , \4759 , \4354 );
nand \mul_7_15_g33828/U$1 ( \4761 , \4385 , \4167 );
nand \mul_7_15_g33779/U$1 ( \4762 , \4760 , \4761 );
xnor \g35887/U$1_r1 ( \4763 , \4758 , \4762 );
xor \mul_7_15_g33490/U$1_r1 ( \4764 , \4730 , \4763 );
not \mul_7_15_g33488/U$1 ( \4765 , \4764 );
nand \mul_7_15_g33466/U$1 ( \4766 , \4699 , \4765 );
nand \mul_7_15_g33402/U$1 ( \4767 , \4694 , \4766 );
xor \mul_7_15_g33490/U$4 ( \4768 , \4722 , \4729 );
and \mul_7_15_g33490/U$3 ( \4769 , \4768 , \4763 );
and \mul_7_15_g33490/U$5 ( \4770 , \4722 , \4729 );
or \mul_7_15_g33490/U$2 ( \4771 , \4769 , \4770 );
not \mul_7_15_g33489/U$1 ( \4772 , \4771 );
xor \mul_7_15_g33817/U$4 ( \4773 , \4709 , \4716 );
and \mul_7_15_g33817/U$3 ( \4774 , \4773 , \4721 );
and \mul_7_15_g33817/U$5 ( \4775 , \4709 , \4716 );
or \mul_7_15_g33817/U$2 ( \4776 , \4774 , \4775 );
and \mul_7_15_g34549/U$2 ( \4777 , \4041 , \4156 );
xor \mul_7_15_g33931/U$1 ( \4778 , \4777 , \4715 );
not \mul_7_15_g34199/U$3 ( \4779 , \4707 );
not \mul_7_15_g34199/U$4 ( \4780 , \4496 );
or \mul_7_15_g34199/U$2 ( \4781 , \4779 , \4780 );
not \mul_7_15_g34703/U$3 ( \4782 , \3943 );
not \mul_7_15_g34703/U$4 ( \4783 , \4212 );
or \mul_7_15_g34703/U$2 ( \4784 , \4782 , \4783 );
nand \mul_7_15_g34914/U$1 ( \4785 , \4216 , \4147 );
nand \mul_7_15_g34703/U$1 ( \4786 , \4784 , \4785 );
nand \mul_7_15_g34386/U$1 ( \4787 , \4377 , \4786 );
nand \mul_7_15_g34199/U$1 ( \4788 , \4781 , \4787 );
xor \mul_7_15_g33931/U$1_r1 ( \4789 , \4778 , \4788 );
xor \mul_7_15_g33920/U$4 ( \4790 , \4737 , \4744 );
and \mul_7_15_g33920/U$3 ( \4791 , \4790 , \4756 );
and \mul_7_15_g33920/U$5 ( \4792 , \4737 , \4744 );
or \mul_7_15_g33920/U$2 ( \4793 , \4791 , \4792 );
xor \mul_7_15_g33759/U$1 ( \4794 , \4789 , \4793 );
not \mul_7_15_g34120/U$3 ( \4795 , \4754 );
not \mul_7_15_g34120/U$4 ( \4796 , \4195 );
or \mul_7_15_g34120/U$2 ( \4797 , \4795 , \4796 );
not \mul_7_15_g34669/U$3 ( \4798 , \3994 );
not \mul_7_15_g34669/U$4 ( \4799 , \4173 );
or \mul_7_15_g34669/U$2 ( \4800 , \4798 , \4799 );
nand \mul_7_15_g34838/U$1 ( \4801 , \4172 , \4099 );
nand \mul_7_15_g34669/U$1 ( \4802 , \4800 , \4801 );
nand \mul_7_15_g34443/U$1 ( \4803 , \4802 , \4205 );
nand \mul_7_15_g34120/U$1 ( \4804 , \4797 , \4803 );
not \mul_7_15_g35322/U$3 ( \4805 , \4136 );
not \mul_7_15_g35322/U$4 ( \4806 , \4140 );
and \mul_7_15_g35322/U$2 ( \4807 , \4805 , \4806 );
nor \mul_7_15_g35322/U$1 ( \4808 , \4807 , \4110 );
not \mul_7_15_g34127/U$1 ( \4809 , \4808 );
and \mul_7_15_g34036/U$2 ( \4810 , \4804 , \4809 );
not \mul_7_15_g34036/U$4 ( \4811 , \4804 );
and \mul_7_15_g34036/U$3 ( \4812 , \4811 , \4808 );
nor \mul_7_15_g34036/U$1 ( \4813 , \4810 , \4812 );
not \mul_7_15_g34204/U$3 ( \4814 , \4741 );
not \mul_7_15_g34417/U$1 ( \4815 , \4254 );
not \mul_7_15_g34204/U$4 ( \4816 , \4815 );
or \mul_7_15_g34204/U$2 ( \4817 , \4814 , \4816 );
xor \mul_7_15_g34545/U$1 ( \4818 , \4047 , \4156 );
nand \mul_7_15_g34303/U$1 ( \4819 , \4818 , \4742 );
nand \mul_7_15_g34204/U$1 ( \4820 , \4817 , \4819 );
xor \mul_7_15_g35314/U$1 ( \4821 , \4813 , \4820 );
xor \mul_7_15_g33759/U$1_r1 ( \4822 , \4794 , \4821 );
xor \mul_7_15_g33574/U$1 ( \4823 , \4776 , \4822 );
not \mul_7_15_g35305/U$2 ( \4824 , \4757 );
nand \mul_7_15_g35305/U$1 ( \4825 , \4824 , \4736 );
not \mul_7_15_g33665/U$3 ( \4826 , \4825 );
not \mul_7_15_g33665/U$4 ( \4827 , \4762 );
or \mul_7_15_g33665/U$2 ( \4828 , \4826 , \4827 );
not \mul_7_15_g35299/U$2 ( \4829 , \4736 );
nand \mul_7_15_g35299/U$1 ( \4830 , \4829 , \4757 );
nand \mul_7_15_g33665/U$1 ( \4831 , \4828 , \4830 );
xor \mul_7_15_g33574/U$1_r1 ( \4832 , \4823 , \4831 );
not \mul_7_15_g33572/U$1 ( \4833 , \4832 );
nand \mul_7_15_g33465/U$1 ( \4834 , \4772 , \4833 );
not \mul_7_15_g33464/U$1 ( \4835 , \4834 );
nor \mul_7_15_g33385/U$1 ( \4836 , \4767 , \4835 );
xor \mul_7_15_g33574/U$4 ( \4837 , \4776 , \4822 );
and \mul_7_15_g33574/U$3 ( \4838 , \4837 , \4831 );
and \mul_7_15_g33574/U$5 ( \4839 , \4776 , \4822 );
or \mul_7_15_g33574/U$2 ( \4840 , \4838 , \4839 );
not \mul_7_15_g33573/U$1 ( \4841 , \4840 );
and \mul_7_15_g34550/U$2 ( \4842 , \4045 , \4156 );
not \mul_7_15_g34213/U$3 ( \4843 , \4786 );
not \mul_7_15_g34213/U$4 ( \4844 , \4496 );
or \mul_7_15_g34213/U$2 ( \4845 , \4843 , \4844 );
not \mul_7_15_g34755/U$3 ( \4846 , \4044 );
not \mul_7_15_g34755/U$4 ( \4847 , \4213 );
or \mul_7_15_g34755/U$2 ( \4848 , \4846 , \4847 );
not \mul_7_15_g35067/U$1 ( \4849 , \4213 );
nand \mul_7_15_g34924/U$1 ( \4850 , \4849 , \4092 );
nand \mul_7_15_g34755/U$1 ( \4851 , \4848 , \4850 );
nand \mul_7_15_g34488/U$1 ( \4852 , \4377 , \4851 );
nand \mul_7_15_g34213/U$1 ( \4853 , \4845 , \4852 );
xor \mul_7_15_g33884/U$1 ( \4854 , \4842 , \4853 );
not \mul_7_15_g34221/U$3 ( \4855 , \4818 );
not \mul_7_15_g34221/U$4 ( \4856 , \4815 );
or \mul_7_15_g34221/U$2 ( \4857 , \4855 , \4856 );
xor \mul_7_15_g34559/U$1 ( \4858 , \4042 , \4156 );
buf \mul_7_15_g34640/U$1 ( \4859 , \4742 );
nand \mul_7_15_g34299/U$1 ( \4860 , \4858 , \4859 );
nand \mul_7_15_g34221/U$1 ( \4861 , \4857 , \4860 );
xor \mul_7_15_g33884/U$1_r1 ( \4862 , \4854 , \4861 );
and \mul_7_15_g34278/U$2 ( \4863 , \4195 , \4802 );
and \mul_7_15_g34278/U$3 ( \4864 , \4205 , \4172 );
nor \mul_7_15_g34278/U$1 ( \4865 , \4863 , \4864 );
xor \mul_7_15_g33931/U$4 ( \4866 , \4777 , \4715 );
and \mul_7_15_g33931/U$3 ( \4867 , \4866 , \4788 );
and \mul_7_15_g33931/U$5 ( \4868 , \4777 , \4715 );
or \mul_7_15_g33931/U$2 ( \4869 , \4867 , \4868 );
xor \mul_7_15_g33754/U$1 ( \4870 , \4865 , \4869 );
not \mul_7_15_g33996/U$3 ( \4871 , \4809 );
not \mul_7_15_g33996/U$4 ( \4872 , \4820 );
or \mul_7_15_g33996/U$2 ( \4873 , \4871 , \4872 );
or \mul_7_15_g34015/U$2 ( \4874 , \4820 , \4809 );
nand \mul_7_15_g34015/U$1 ( \4875 , \4874 , \4804 );
nand \mul_7_15_g33996/U$1 ( \4876 , \4873 , \4875 );
xor \mul_7_15_g33754/U$1_r1 ( \4877 , \4870 , \4876 );
xor \mul_7_15_g33602/U$1 ( \4878 , \4862 , \4877 );
xor \mul_7_15_g33759/U$4 ( \4879 , \4789 , \4793 );
and \mul_7_15_g33759/U$3 ( \4880 , \4879 , \4821 );
and \mul_7_15_g33759/U$5 ( \4881 , \4789 , \4793 );
or \mul_7_15_g33759/U$2 ( \4882 , \4880 , \4881 );
xor \mul_7_15_g33602/U$1_r1 ( \4883 , \4878 , \4882 );
not \mul_7_15_g33570/U$1 ( \4884 , \4883 );
nand \mul_7_15_g33518/U$1 ( \4885 , \4841 , \4884 );
and \mul_7_15_g34545/U$2 ( \4886 , \4047 , \4156 );
not \mul_7_15_g34168/U$3 ( \4887 , \4851 );
not \mul_7_15_g34168/U$4 ( \4888 , \4496 );
or \mul_7_15_g34168/U$2 ( \4889 , \4887 , \4888 );
and \mul_7_15_g34670/U$2 ( \4890 , \4213 , \3994 );
and \mul_7_15_g34670/U$3 ( \4891 , \4849 , \4099 );
nor \mul_7_15_g34670/U$1 ( \4892 , \4890 , \4891 );
not \mul_7_15_g34384/U$2 ( \4893 , \4892 );
nand \mul_7_15_g34384/U$1 ( \4894 , \4893 , \4377 );
nand \mul_7_15_g34168/U$1 ( \4895 , \4889 , \4894 );
xor \mul_7_15_g33940/U$1 ( \4896 , \4886 , \4895 );
not \mul_7_15_g34109/U$3 ( \4897 , \4319 );
not \mul_7_15_g34109/U$4 ( \4898 , \4317 );
or \mul_7_15_g34109/U$2 ( \4899 , \4897 , \4898 );
nand \mul_7_15_g34109/U$1 ( \4900 , \4899 , \4172 );
xor \mul_7_15_g33940/U$1_r1 ( \4901 , \4896 , \4900 );
not \mul_7_15_g34277/U$1 ( \4902 , \4865 );
not \mul_7_15_g34208/U$3 ( \4903 , \4858 );
not \mul_7_15_g34208/U$4 ( \4904 , \4815 );
or \mul_7_15_g34208/U$2 ( \4905 , \4903 , \4904 );
xor \mul_7_15_g34555/U$1 ( \4906 , \3943 , \4156 );
nand \mul_7_15_g34304/U$1 ( \4907 , \4906 , \4859 );
nand \mul_7_15_g34208/U$1 ( \4908 , \4905 , \4907 );
xor \mul_7_15_g33783/U$1 ( \4909 , \4902 , \4908 );
xor \mul_7_15_g33884/U$4 ( \4910 , \4842 , \4853 );
and \mul_7_15_g33884/U$3 ( \4911 , \4910 , \4861 );
and \mul_7_15_g33884/U$5 ( \4912 , \4842 , \4853 );
or \mul_7_15_g33884/U$2 ( \4913 , \4911 , \4912 );
xor \mul_7_15_g33783/U$1_r1 ( \4914 , \4909 , \4913 );
xor \mul_7_15_g33617/U$1 ( \4915 , \4901 , \4914 );
xor \mul_7_15_g33754/U$4 ( \4916 , \4865 , \4869 );
and \mul_7_15_g33754/U$3 ( \4917 , \4916 , \4876 );
and \mul_7_15_g33754/U$5 ( \4918 , \4865 , \4869 );
or \mul_7_15_g33754/U$2 ( \4919 , \4917 , \4918 );
xnor \mul_7_15_g33617/U$1_r1 ( \4920 , \4915 , \4919 );
not \mul_7_15_g33753/U$1 ( \4921 , \4877 );
not \mul_7_15_g33883/U$1 ( \4922 , \4862 );
nand \mul_7_15_g33688/U$1 ( \4923 , \4921 , \4922 );
and \mul_7_15_g33594/U$2 ( \4924 , \4923 , \4882 );
nor \mul_7_15_g33691/U$1 ( \4925 , \4921 , \4922 );
nor \mul_7_15_g33594/U$1 ( \4926 , \4924 , \4925 );
nand \mul_7_15_g33532/U$1 ( \4927 , \4920 , \4926 );
nand \g35618/U$1 ( \4928 , \4836 , \4885 , \4927 );
or \mul_7_15_g35292/U$2 ( \4929 , \4901 , \4914 );
nand \mul_7_15_g35292/U$1 ( \4930 , \4929 , \4919 );
nand \mul_7_15_g33735/U$1 ( \4931 , \4914 , \4901 );
nand \mul_7_15_g33613/U$1 ( \4932 , \4930 , \4931 );
xor \mul_7_15_g33940/U$4 ( \4933 , \4886 , \4895 );
and \mul_7_15_g33940/U$3 ( \4934 , \4933 , \4900 );
and \mul_7_15_g33940/U$5 ( \4935 , \4886 , \4895 );
or \mul_7_15_g33940/U$2 ( \4936 , \4934 , \4935 );
and \mul_7_15_g34559/U$2 ( \4937 , \4042 , \4156 );
not \mul_7_15_g34290/U$3 ( \4938 , \4892 );
not \mul_7_15_g34401/U$1 ( \4939 , \4496 );
not \mul_7_15_g34290/U$4 ( \4940 , \4939 );
and \mul_7_15_g34290/U$2 ( \4941 , \4938 , \4940 );
and \mul_7_15_g34290/U$5 ( \4942 , \4377 , \4849 );
nor \mul_7_15_g34290/U$1 ( \4943 , \4941 , \4942 );
xor \mul_7_15_g33918/U$1 ( \4944 , \4937 , \4943 );
not \mul_7_15_g34554/U$1 ( \4945 , \4906 );
or \mul_7_15_g34179/U$2 ( \4946 , \4254 , \4945 );
and \mul_7_15_g34666/U$2 ( \4947 , \4267 , \4044 );
and \mul_7_15_g34666/U$3 ( \4948 , \4156 , \4092 );
nor \mul_7_15_g34666/U$1 ( \4949 , \4947 , \4948 );
not \mul_7_15_g34638/U$1 ( \4950 , \4859 );
or \mul_7_15_g34179/U$3 ( \4951 , \4949 , \4950 );
nand \mul_7_15_g34179/U$1 ( \4952 , \4946 , \4951 );
xor \mul_7_15_g33918/U$1_r1 ( \4953 , \4944 , \4952 );
xor \mul_7_15_g33674/U$1 ( \4954 , \4936 , \4953 );
xor \mul_7_15_g33783/U$4 ( \4955 , \4902 , \4908 );
and \mul_7_15_g33783/U$3 ( \4956 , \4955 , \4913 );
and \mul_7_15_g33783/U$5 ( \4957 , \4902 , \4908 );
or \mul_7_15_g33783/U$2 ( \4958 , \4956 , \4957 );
xor \mul_7_15_g33674/U$1_r1 ( \4959 , \4954 , \4958 );
nor \mul_7_15_g33562/U$1 ( \4960 , \4932 , \4959 );
xor \mul_7_15_g33674/U$4 ( \4961 , \4936 , \4953 );
and \mul_7_15_g33674/U$3 ( \4962 , \4961 , \4958 );
and \mul_7_15_g33674/U$5 ( \4963 , \4936 , \4953 );
or \mul_7_15_g33674/U$2 ( \4964 , \4962 , \4963 );
xor \mul_7_15_g33918/U$4 ( \4965 , \4937 , \4943 );
and \mul_7_15_g33918/U$3 ( \4966 , \4965 , \4952 );
and \mul_7_15_g33918/U$5 ( \4967 , \4937 , \4943 );
or \mul_7_15_g33918/U$2 ( \4968 , \4966 , \4967 );
not \mul_7_15_g34289/U$1 ( \4969 , \4943 );
xor \mul_7_15_g33743/U$1 ( \4970 , \4968 , \4969 );
or \mul_7_15_g34129/U$2 ( \4971 , \4496 , \4377 );
nand \mul_7_15_g34129/U$1 ( \4972 , \4971 , \4849 );
and \mul_7_15_g34555/U$2 ( \4973 , \3943 , \4156 );
xor \mul_7_15_g33941/U$1 ( \4974 , \4972 , \4973 );
or \mul_7_15_g34161/U$2 ( \4975 , \4254 , \4949 );
and \mul_7_15_g34659/U$2 ( \4976 , \4267 , \3994 );
and \mul_7_15_g34659/U$3 ( \4977 , \4156 , \4099 );
nor \mul_7_15_g34659/U$1 ( \4978 , \4976 , \4977 );
or \mul_7_15_g34161/U$3 ( \4979 , \4978 , \4950 );
nand \mul_7_15_g34161/U$1 ( \4980 , \4975 , \4979 );
xor \mul_7_15_g33941/U$1_r1 ( \4981 , \4974 , \4980 );
xor \mul_7_15_g33743/U$1_r1 ( \4982 , \4970 , \4981 );
nor \mul_7_15_g33637/U$1 ( \4983 , \4964 , \4982 );
nor \mul_7_15_g33318/U$1 ( \4984 , \4928 , \4960 , \4983 );
not \mul_7_15_g33290/U$3 ( \4985 , \4984 );
xor \mul_7_15_g33901/U$1 ( \4986 , \4586 , \4598 );
xnor \mul_7_15_g33901/U$1_r1 ( \4987 , \4986 , \4610 );
not \mul_7_15_g34032/U$3 ( \4988 , \4676 );
not \mul_7_15_g34184/U$1 ( \4989 , \4659 );
not \mul_7_15_g34032/U$4 ( \4990 , \4989 );
or \mul_7_15_g34032/U$2 ( \4991 , \4988 , \4990 );
nand \mul_7_15_g34052/U$1 ( \4992 , \4675 , \4659 );
nand \mul_7_15_g34032/U$1 ( \4993 , \4991 , \4992 );
not \mul_7_15_g33968/U$3 ( \4994 , \4993 );
not \mul_7_15_g34180/U$1 ( \4995 , \4649 );
not \mul_7_15_g33968/U$4 ( \4996 , \4995 );
and \mul_7_15_g33968/U$2 ( \4997 , \4994 , \4996 );
and \mul_7_15_g33968/U$5 ( \4998 , \4993 , \4995 );
nor \mul_7_15_g33968/U$1 ( \4999 , \4997 , \4998 );
xor \mul_7_15_g33724/U$4 ( \5000 , \4987 , \4999 );
not \mul_7_15_g34685/U$3 ( \5001 , \4045 );
not \mul_7_15_g34685/U$4 ( \5002 , \4089 );
or \mul_7_15_g34685/U$2 ( \5003 , \5001 , \5002 );
nand \mul_7_15_g34921/U$1 ( \5004 , \4088 , \4286 );
nand \mul_7_15_g34685/U$1 ( \5005 , \5003 , \5004 );
not \mul_7_15_g34148/U$3 ( \5006 , \5005 );
not \mul_7_15_g34148/U$4 ( \5007 , \4437 );
or \mul_7_15_g34148/U$2 ( \5008 , \5006 , \5007 );
not \mul_7_15_g34702/U$3 ( \5009 , \4047 );
not \mul_7_15_g34702/U$4 ( \5010 , \4089 );
or \mul_7_15_g34702/U$2 ( \5011 , \5009 , \5010 );
nand \mul_7_15_g34928/U$1 ( \5012 , \4088 , \4178 );
nand \mul_7_15_g34702/U$1 ( \5013 , \5011 , \5012 );
nand \mul_7_15_g34423/U$1 ( \5014 , \4596 , \5013 );
nand \mul_7_15_g34148/U$1 ( \5015 , \5008 , \5014 );
buf \mul_7_15_g35045/U$1 ( \5016 , \1395 );
not \mul_7_15_g35037/U$1 ( \5017 , \5016 );
nor \mul_7_15_g34941/U$1 ( \5018 , \5017 , \3617 );
buf \mul_7_15_g34940/U$1 ( \5019 , \5018 );
buf \mul_7_15_g34939/U$1 ( \5020 , \5019 );
buf \mul_7_15_g34981/U$1 ( \5021 , \3617 );
or \mul_7_15_g34542/U$2 ( \5022 , \5020 , \5021 );
not \mul_7_15_g35042/U$1 ( \5023 , \5016 );
not \mul_7_15_g35041/U$1 ( \5024 , \5023 );
nand \mul_7_15_g34542/U$1 ( \5025 , \5022 , \5024 );
nor \mul_7_15_g34062/U$1 ( \5026 , \5015 , \5025 );
not \mul_7_15_g34661/U$3 ( \5027 , \4019 );
not \mul_7_15_g34661/U$4 ( \5028 , \4267 );
or \mul_7_15_g34661/U$2 ( \5029 , \5027 , \5028 );
nand \mul_7_15_g34909/U$1 ( \5030 , \4308 , \4585 );
nand \mul_7_15_g34661/U$1 ( \5031 , \5029 , \5030 );
not \mul_7_15_g34171/U$3 ( \5032 , \5031 );
not \mul_7_15_g34171/U$4 ( \5033 , \4253 );
or \mul_7_15_g34171/U$2 ( \5034 , \5032 , \5033 );
nand \mul_7_15_g34302/U$1 ( \5035 , \4644 , \4742 );
nand \mul_7_15_g34171/U$1 ( \5036 , \5034 , \5035 );
not \mul_7_15_g34170/U$1 ( \5037 , \5036 );
xor \mul_7_15_g33894/U$4 ( \5038 , \5026 , \5037 );
and \mul_7_15_g33894/U$3 ( \5039 , \5038 , \4676 );
and \mul_7_15_g33894/U$5 ( \5040 , \5026 , \5037 );
or \mul_7_15_g33894/U$2 ( \5041 , \5039 , \5040 );
and \mul_7_15_g33724/U$3 ( \5042 , \5000 , \5041 );
and \mul_7_15_g33724/U$5 ( \5043 , \4987 , \4999 );
or \mul_7_15_g33724/U$2 ( \5044 , \5042 , \5043 );
xor \mul_7_15_g33698/U$1 ( \5045 , \4413 , \4580 );
xnor \mul_7_15_g33698/U$1_r1 ( \5046 , \5045 , \4612 );
xor \mul_7_15_g33906/U$1 ( \5047 , \4549 , \4564 );
xnor \mul_7_15_g33906/U$1_r1 ( \5048 , \5047 , \4578 );
not \mul_7_15_g33880/U$1 ( \5049 , \5048 );
not \mul_7_15_g33694/U$3 ( \5050 , \5049 );
not \mul_7_15_g34155/U$3 ( \5051 , \5013 );
not \mul_7_15_g34155/U$4 ( \5052 , \4437 );
or \mul_7_15_g34155/U$2 ( \5053 , \5051 , \5052 );
nand \mul_7_15_g34359/U$1 ( \5054 , \4331 , \4592 );
nand \mul_7_15_g34155/U$1 ( \5055 , \5053 , \5054 );
not \mul_7_15_g34002/U$3 ( \5056 , \5055 );
not \mul_7_15_g34780/U$3 ( \5057 , \3943 );
not \mul_7_15_g34780/U$4 ( \5058 , \4069 );
or \mul_7_15_g34780/U$2 ( \5059 , \5057 , \5058 );
not \mul_7_15_fopt35199/U$1 ( \5060 , \4069 );
nand \mul_7_15_g34886/U$1 ( \5061 , \5060 , \4147 );
nand \mul_7_15_g34780/U$1 ( \5062 , \5059 , \5061 );
not \mul_7_15_g34214/U$3 ( \5063 , \5062 );
not \mul_7_15_g34214/U$4 ( \5064 , \4065 );
or \mul_7_15_g34214/U$2 ( \5065 , \5063 , \5064 );
nand \mul_7_15_g34366/U$1 ( \5066 , \4055 , \4556 );
nand \mul_7_15_g34214/U$1 ( \5067 , \5065 , \5066 );
not \mul_7_15_g34002/U$4 ( \5068 , \5067 );
or \mul_7_15_g34002/U$2 ( \5069 , \5056 , \5068 );
or \mul_7_15_g34021/U$2 ( \5070 , \5067 , \5055 );
not \mul_7_15_g34767/U$3 ( \5071 , \4041 );
not \mul_7_15_g34767/U$4 ( \5072 , \4142 );
or \mul_7_15_g34767/U$2 ( \5073 , \5071 , \5072 );
nand \mul_7_15_g34895/U$1 ( \5074 , \4109 , \4238 );
nand \mul_7_15_g34767/U$1 ( \5075 , \5073 , \5074 );
not \mul_7_15_g34276/U$3 ( \5076 , \5075 );
not \mul_7_15_g34276/U$4 ( \5077 , \4136 );
or \mul_7_15_g34276/U$2 ( \5078 , \5076 , \5077 );
nand \mul_7_15_g34489/U$1 ( \5079 , \4140 , \4573 );
nand \mul_7_15_g34276/U$1 ( \5080 , \5078 , \5079 );
nand \mul_7_15_g34021/U$1 ( \5081 , \5070 , \5080 );
nand \mul_7_15_g34002/U$1 ( \5082 , \5069 , \5081 );
not \mul_7_15_g33694/U$4 ( \5083 , \5082 );
or \mul_7_15_g33694/U$2 ( \5084 , \5050 , \5083 );
not \mul_7_15_g33922/U$1 ( \5085 , \5082 );
not \mul_7_15_g33736/U$3 ( \5086 , \5085 );
not \mul_7_15_g33736/U$4 ( \5087 , \5048 );
or \mul_7_15_g33736/U$2 ( \5088 , \5086 , \5087 );
and \mul_7_15_g34827/U$1 ( \5089 , \4156 , \4023 );
not \mul_7_15_g33999/U$3 ( \5090 , \5089 );
and \mul_7_15_g34757/U$2 ( \5091 , \3958 , \4216 );
not \mul_7_15_g34757/U$4 ( \5092 , \3958 );
and \mul_7_15_g34757/U$3 ( \5093 , \5092 , \4213 );
nor \mul_7_15_g34757/U$1 ( \5094 , \5091 , \5093 );
not \mul_7_15_g34201/U$3 ( \5095 , \5094 );
not \mul_7_15_g34201/U$4 ( \5096 , \4231 );
or \mul_7_15_g34201/U$2 ( \5097 , \5095 , \5096 );
nand \mul_7_15_g34437/U$1 ( \5098 , \4234 , \4654 );
nand \mul_7_15_g34201/U$1 ( \5099 , \5097 , \5098 );
not \mul_7_15_g33999/U$4 ( \5100 , \5099 );
or \mul_7_15_g33999/U$2 ( \5101 , \5090 , \5100 );
or \mul_7_15_g34026/U$2 ( \5102 , \5099 , \5089 );
not \mul_7_15_g34772/U$3 ( \5103 , \4011 );
not \mul_7_15_g34772/U$4 ( \5104 , \4176 );
or \mul_7_15_g34772/U$2 ( \5105 , \5103 , \5104 );
nand \mul_7_15_g34891/U$1 ( \5106 , \4172 , \4270 );
nand \mul_7_15_g34772/U$1 ( \5107 , \5105 , \5106 );
not \mul_7_15_g34110/U$3 ( \5108 , \5107 );
not \mul_7_15_g34110/U$4 ( \5109 , \4194 );
or \mul_7_15_g34110/U$2 ( \5110 , \5108 , \5109 );
not \mul_7_15_g34631/U$1 ( \5111 , \4203 );
nand \mul_7_15_g34433/U$1 ( \5112 , \4605 , \5111 );
nand \mul_7_15_g34110/U$1 ( \5113 , \5110 , \5112 );
nand \mul_7_15_g34026/U$1 ( \5114 , \5102 , \5113 );
nand \mul_7_15_g33999/U$1 ( \5115 , \5101 , \5114 );
nand \mul_7_15_g33736/U$1 ( \5116 , \5088 , \5115 );
nand \mul_7_15_g33694/U$1 ( \5117 , \5084 , \5116 );
xor \g35369/U$1 ( \5118 , \5046 , \5117 );
xor \g35659/U$1 ( \5119 , \4679 , \4631 );
not \mul_7_15_g33947/U$1 ( \5120 , \4638 );
and \g35620/U$2 ( \5121 , \5119 , \5120 );
not \g35620/U$4 ( \5122 , \5119 );
and \g35620/U$3 ( \5123 , \5122 , \4638 );
nor \g35620/U$1 ( \5124 , \5121 , \5123 );
xnor \g35369/U$1_r1 ( \5125 , \5118 , \5124 );
xor \mul_7_15_g33409/U$1 ( \5126 , \5044 , \5125 );
not \mul_7_15_g34209/U$3 ( \5127 , \4480 );
not \mul_7_15_g34668/U$3 ( \5128 , \4023 );
not \mul_7_15_g34668/U$4 ( \5129 , \4267 );
or \mul_7_15_g34668/U$2 ( \5130 , \5128 , \5129 );
not \mul_7_15_g35081/U$1 ( \5131 , \4023 );
nand \mul_7_15_g34922/U$1 ( \5132 , \4156 , \5131 );
nand \mul_7_15_g34668/U$1 ( \5133 , \5130 , \5132 );
not \mul_7_15_g34209/U$4 ( \5134 , \5133 );
or \mul_7_15_g34209/U$2 ( \5135 , \5127 , \5134 );
nand \mul_7_15_g34296/U$1 ( \5136 , \5031 , \4273 );
nand \mul_7_15_g34209/U$1 ( \5137 , \5135 , \5136 );
and \mul_7_15_g35267/U$1 ( \5138 , \4156 , \4026 );
or \mul_7_15_g33959/U$2 ( \5139 , \5137 , \5138 );
not \mul_7_15_g34746/U$3 ( \5140 , \4046 );
not \mul_7_15_g34746/U$4 ( \5141 , \4284 );
or \mul_7_15_g34746/U$2 ( \5142 , \5140 , \5141 );
nand \mul_7_15_g34900/U$1 ( \5143 , \4177 , \4256 );
nand \mul_7_15_g34746/U$1 ( \5144 , \5142 , \5143 );
not \mul_7_15_g34124/U$3 ( \5145 , \5144 );
not \mul_7_15_g34124/U$4 ( \5146 , \4194 );
or \mul_7_15_g34124/U$2 ( \5147 , \5145 , \5146 );
nand \mul_7_15_g34368/U$1 ( \5148 , \5107 , \4204 );
nand \mul_7_15_g34124/U$1 ( \5149 , \5147 , \5148 );
nand \mul_7_15_g33959/U$1 ( \5150 , \5139 , \5149 );
nand \mul_7_15_g34069/U$1 ( \5151 , \5137 , \5138 );
nand \mul_7_15_g33900/U$1 ( \5152 , \5150 , \5151 );
not \mul_7_15_g34689/U$3 ( \5153 , \4042 );
not \mul_7_15_g34689/U$4 ( \5154 , \4069 );
or \mul_7_15_g34689/U$2 ( \5155 , \5153 , \5154 );
nand \mul_7_15_g34878/U$1 ( \5156 , \5060 , \4116 );
nand \mul_7_15_g34689/U$1 ( \5157 , \5155 , \5156 );
not \mul_7_15_g34215/U$3 ( \5158 , \5157 );
not \mul_7_15_g34215/U$4 ( \5159 , \4558 );
or \mul_7_15_g34215/U$2 ( \5160 , \5158 , \5159 );
nand \mul_7_15_g34347/U$1 ( \5161 , \4054 , \5062 );
nand \mul_7_15_g34215/U$1 ( \5162 , \5160 , \5161 );
not \mul_7_15_g34006/U$3 ( \5163 , \5162 );
not \g35940/U$3 ( \5164 , \4140 );
not \g35940/U$4 ( \5165 , \5075 );
or \g35940/U$2 ( \5166 , \5164 , \5165 );
and \mul_7_15_g34681/U$2 ( \5167 , \4217 , \4109 );
not \mul_7_15_g34681/U$4 ( \5168 , \4217 );
and \mul_7_15_g34681/U$3 ( \5169 , \5168 , \4569 );
nor \mul_7_15_g34681/U$1 ( \5170 , \5167 , \5169 );
not \g35941/U$2 ( \5171 , \5170 );
nand \g35941/U$1 ( \5172 , \5171 , \4136 );
nand \g35940/U$1 ( \5173 , \5166 , \5172 );
not \mul_7_15_g34006/U$4 ( \5174 , \5173 );
or \mul_7_15_g34006/U$2 ( \5175 , \5163 , \5174 );
or \mul_7_15_g34020/U$2 ( \5176 , \5173 , \5162 );
not \mul_7_15_g34739/U$3 ( \5177 , \4044 );
not \mul_7_15_g35161/U$1 ( \5178 , \4548 );
not \mul_7_15_g34739/U$4 ( \5179 , \5178 );
or \mul_7_15_g34739/U$2 ( \5180 , \5177 , \5179 );
nand \mul_7_15_g34933/U$1 ( \5181 , \4548 , \4092 );
nand \mul_7_15_g34739/U$1 ( \5182 , \5180 , \5181 );
not \mul_7_15_g34246/U$3 ( \5183 , \5182 );
not \mul_7_15_g34246/U$4 ( \5184 , \4661 );
or \mul_7_15_g34246/U$2 ( \5185 , \5183 , \5184 );
not \mul_7_15_g34385/U$2 ( \5186 , \4669 );
not \mul_7_15_g34650/U$1 ( \5187 , \4545 );
nand \mul_7_15_g34385/U$1 ( \5188 , \5186 , \5187 );
nand \mul_7_15_g34246/U$1 ( \5189 , \5185 , \5188 );
nand \mul_7_15_g34020/U$1 ( \5190 , \5176 , \5189 );
nand \mul_7_15_g34006/U$1 ( \5191 , \5175 , \5190 );
or \mul_7_15_g35300/U$1 ( \5192 , \5152 , \5191 );
xor \g35399/U$1 ( \5193 , \5067 , \5080 );
xor \g35399/U$1_r1 ( \5194 , \5193 , \5055 );
and \mul_7_15_g33693/U$2 ( \5195 , \5192 , \5194 );
and \mul_7_15_g33784/U$2 ( \5196 , \5152 , \5191 );
nor \mul_7_15_g33693/U$1 ( \5197 , \5195 , \5196 );
xor \g35392/U$1 ( \5198 , \5082 , \5048 );
xor \g35392/U$1_r1 ( \5199 , \5198 , \5115 );
xor \mul_7_15_g33549/U$4 ( \5200 , \5197 , \5199 );
xor \mul_7_15_g33724/U$1 ( \5201 , \4987 , \4999 );
xor \mul_7_15_g33724/U$1_r1 ( \5202 , \5201 , \5041 );
and \mul_7_15_g33549/U$3 ( \5203 , \5200 , \5202 );
and \mul_7_15_g33549/U$5 ( \5204 , \5197 , \5199 );
or \mul_7_15_g33549/U$2 ( \5205 , \5203 , \5204 );
xor \mul_7_15_g33409/U$1_r1 ( \5206 , \5126 , \5205 );
xor \mul_7_15_g33974/U$1 ( \5207 , \5089 , \5113 );
xnor \mul_7_15_g33974/U$1_r1 ( \5208 , \5207 , \5099 );
nand \mul_7_15_g34454/U$1 ( \5209 , \4127 , \4134 );
not \mul_7_15_g34254/U$3 ( \5210 , \5209 );
not \mul_7_15_g34748/U$3 ( \5211 , \4011 );
not \mul_7_15_g34748/U$4 ( \5212 , \4145 );
or \mul_7_15_g34748/U$2 ( \5213 , \5211 , \5212 );
nand \mul_7_15_g34905/U$1 ( \5214 , \4109 , \4270 );
nand \mul_7_15_g34748/U$1 ( \5215 , \5213 , \5214 );
not \mul_7_15_g34747/U$1 ( \5216 , \5215 );
not \mul_7_15_g34254/U$4 ( \5217 , \5216 );
and \mul_7_15_g34254/U$2 ( \5218 , \5210 , \5217 );
nor \mul_7_15_g34434/U$1 ( \5219 , \5170 , \4428 );
nor \mul_7_15_g34254/U$1 ( \5220 , \5218 , \5219 );
not \mul_7_15_g34758/U$3 ( \5221 , \3943 );
not \mul_7_15_g34758/U$4 ( \5222 , \5178 );
or \mul_7_15_g34758/U$2 ( \5223 , \5221 , \5222 );
nand \mul_7_15_g34907/U$1 ( \5224 , \4665 , \4147 );
nand \mul_7_15_g34758/U$1 ( \5225 , \5223 , \5224 );
not \mul_7_15_g34241/U$3 ( \5226 , \5225 );
not \mul_7_15_g34241/U$4 ( \5227 , \4662 );
or \mul_7_15_g34241/U$2 ( \5228 , \5226 , \5227 );
nand \mul_7_15_g34436/U$1 ( \5229 , \4672 , \5182 );
nand \mul_7_15_g34241/U$1 ( \5230 , \5228 , \5229 );
not \mul_7_15_g34240/U$1 ( \5231 , \5230 );
xor \mul_7_15_g33925/U$4 ( \5232 , \5220 , \5231 );
not \mul_7_15_g34750/U$3 ( \5233 , \4041 );
not \mul_7_15_g35020/U$1 ( \5234 , \4088 );
not \mul_7_15_g34750/U$4 ( \5235 , \5234 );
or \mul_7_15_g34750/U$2 ( \5236 , \5233 , \5235 );
nand \mul_7_15_g34842/U$1 ( \5237 , \4088 , \4238 );
nand \mul_7_15_g34750/U$1 ( \5238 , \5236 , \5237 );
and \mul_7_15_g35324/U$2 ( \5239 , \4437 , \5238 );
not \mul_7_15_g35334/U$2 ( \5240 , \5005 );
buf \fopt35518/U$1 ( \5241 , \4103 );
nor \mul_7_15_g35334/U$1 ( \5242 , \5240 , \5241 );
nor \mul_7_15_g35324/U$1 ( \5243 , \5239 , \5242 );
and \mul_7_15_g33925/U$3 ( \5244 , \5232 , \5243 );
and \mul_7_15_g33925/U$5 ( \5245 , \5220 , \5231 );
or \mul_7_15_g33925/U$2 ( \5246 , \5244 , \5245 );
not \mul_7_15_g35306/U$2 ( \5247 , \5246 );
not \mul_7_15_g34765/U$3 ( \5248 , \3963 );
not \mul_7_15_g34765/U$4 ( \5249 , \4212 );
or \mul_7_15_g34765/U$2 ( \5250 , \5248 , \5249 );
nand \mul_7_15_g34856/U$1 ( \5251 , \4492 , \4486 );
nand \mul_7_15_g34765/U$1 ( \5252 , \5250 , \5251 );
not \mul_7_15_g34198/U$3 ( \5253 , \5252 );
not \mul_7_15_g34198/U$4 ( \5254 , \4496 );
or \mul_7_15_g34198/U$2 ( \5255 , \5253 , \5254 );
nand \mul_7_15_g34348/U$1 ( \5256 , \4377 , \5094 );
nand \mul_7_15_g34198/U$1 ( \5257 , \5255 , \5256 );
nand \mul_7_15_g35306/U$1 ( \5258 , \5247 , \5257 );
xor \mul_7_15_g33652/U$4 ( \5259 , \5208 , \5258 );
xor \mul_7_15_g33894/U$1 ( \5260 , \5026 , \5037 );
xor \mul_7_15_g33894/U$1_r1 ( \5261 , \5260 , \4676 );
and \mul_7_15_g33652/U$3 ( \5262 , \5259 , \5261 );
and \mul_7_15_g33652/U$5 ( \5263 , \5208 , \5258 );
or \mul_7_15_g33652/U$2 ( \5264 , \5262 , \5263 );
not \mul_7_15_g34980/U$1 ( \5265 , \5021 );
not \mul_7_15_g34339/U$3 ( \5266 , \5265 );
not \mul_7_15_g34339/U$4 ( \5267 , \5023 );
and \mul_7_15_g34339/U$2 ( \5268 , \5266 , \5267 );
not \mul_7_15_g34678/U$3 ( \5269 , \3994 );
not \mul_7_15_g35036/U$1 ( \5270 , \1395 );
not \mul_7_15_g34678/U$4 ( \5271 , \5270 );
or \mul_7_15_g34678/U$2 ( \5272 , \5269 , \5271 );
buf \mul_7_15_g35056/U$1 ( \5273 , \1395 );
nand \mul_7_15_g34839/U$1 ( \5274 , \5273 , \4099 );
nand \mul_7_15_g34678/U$1 ( \5275 , \5272 , \5274 );
and \mul_7_15_g34339/U$5 ( \5276 , \5019 , \5275 );
nor \mul_7_15_g34339/U$1 ( \5277 , \5268 , \5276 );
not \mul_7_15_g34027/U$3 ( \5278 , \5277 );
not \mul_7_15_g34778/U$3 ( \5279 , \4019 );
not \mul_7_15_g34778/U$4 ( \5280 , \4211 );
or \mul_7_15_g34778/U$2 ( \5281 , \5279 , \5280 );
nand \mul_7_15_g34848/U$1 ( \5282 , \4585 , \3577 );
nand \mul_7_15_g34778/U$1 ( \5283 , \5281 , \5282 );
not \mul_7_15_g34207/U$3 ( \5284 , \5283 );
not \mul_7_15_g34207/U$4 ( \5285 , \4231 );
or \mul_7_15_g34207/U$2 ( \5286 , \5284 , \5285 );
nand \mul_7_15_g34440/U$1 ( \5287 , \4234 , \5252 );
nand \mul_7_15_g34207/U$1 ( \5288 , \5286 , \5287 );
not \mul_7_15_g34206/U$1 ( \5289 , \5288 );
not \mul_7_15_g34027/U$4 ( \5290 , \5289 );
or \mul_7_15_g34027/U$2 ( \5291 , \5278 , \5290 );
not \mul_7_15_g34713/U$3 ( \5292 , \3958 );
not \mul_7_15_g34713/U$4 ( \5293 , \4176 );
or \mul_7_15_g34713/U$2 ( \5294 , \5292 , \5293 );
nand \mul_7_15_g34911/U$1 ( \5295 , \4172 , \4473 );
nand \mul_7_15_g34713/U$1 ( \5296 , \5294 , \5295 );
not \mul_7_15_g34123/U$3 ( \5297 , \5296 );
not \mul_7_15_g34123/U$4 ( \5298 , \4194 );
or \mul_7_15_g34123/U$2 ( \5299 , \5297 , \5298 );
nand \mul_7_15_g34442/U$1 ( \5300 , \5144 , \4204 );
nand \mul_7_15_g34123/U$1 ( \5301 , \5299 , \5300 );
nand \mul_7_15_g34027/U$1 ( \5302 , \5291 , \5301 );
not \mul_7_15_g34068/U$2 ( \5303 , \5277 );
nand \mul_7_15_g34068/U$1 ( \5304 , \5303 , \5288 );
nand \mul_7_15_g34000/U$1 ( \5305 , \5302 , \5304 );
not \mul_7_15_g33930/U$1 ( \5306 , \5305 );
xor \mul_7_15_g33902/U$1 ( \5307 , \5138 , \5149 );
xnor \mul_7_15_g33902/U$1_r1 ( \5308 , \5307 , \5137 );
nand \mul_7_15_g35762/U$1 ( \5309 , \5306 , \5308 );
not \mul_7_15_g33858/U$3 ( \5310 , \5257 );
not \mul_7_15_g33858/U$4 ( \5311 , \5246 );
or \mul_7_15_g33858/U$2 ( \5312 , \5310 , \5311 );
or \mul_7_15_g33858/U$5 ( \5313 , \5246 , \5257 );
nand \mul_7_15_g33858/U$1 ( \5314 , \5312 , \5313 );
and \mul_7_15_g33695/U$2 ( \5315 , \5309 , \5314 );
nor \mul_7_15_g33837/U$1 ( \5316 , \5306 , \5308 );
nor \mul_7_15_g33695/U$1 ( \5317 , \5315 , \5316 );
not \mul_7_15_g33612/U$3 ( \5318 , \5317 );
xor \mul_7_15_g33784/U$1 ( \5319 , \5152 , \5191 );
and \mul_7_15_g33730/U$2 ( \5320 , \5319 , \5194 );
not \mul_7_15_g33730/U$4 ( \5321 , \5319 );
not \mul_7_15_g33921/U$1 ( \5322 , \5194 );
and \mul_7_15_g33730/U$3 ( \5323 , \5321 , \5322 );
nor \mul_7_15_g33730/U$1 ( \5324 , \5320 , \5323 );
not \mul_7_15_g33681/U$1 ( \5325 , \5324 );
not \mul_7_15_g33612/U$4 ( \5326 , \5325 );
or \mul_7_15_g33612/U$2 ( \5327 , \5318 , \5326 );
not \mul_7_15_g34017/U$2 ( \5328 , \5026 );
nand \mul_7_15_g34066/U$1 ( \5329 , \5015 , \5025 );
nand \mul_7_15_g34017/U$1 ( \5330 , \5328 , \5329 );
not \mul_7_15_g33871/U$2 ( \5331 , \5330 );
xor \g35402/U$1 ( \5332 , \5162 , \5189 );
not \mul_7_15_g34271/U$1 ( \5333 , \5173 );
and \mul_7_15_g33983/U$2 ( \5334 , \5332 , \5333 );
not \mul_7_15_g33983/U$4 ( \5335 , \5332 );
and \mul_7_15_g33983/U$3 ( \5336 , \5335 , \5173 );
nor \mul_7_15_g33983/U$1 ( \5337 , \5334 , \5336 );
nand \mul_7_15_g33871/U$1 ( \5338 , \5331 , \5337 );
not \mul_7_15_g34949/U$1 ( \5339 , \4029 );
nor \mul_7_15_g34828/U$1 ( \5340 , \4267 , \5339 );
and \mul_7_15_g34662/U$2 ( \5341 , \4260 , \4026 );
not \mul_7_15_g35106/U$1 ( \5342 , \3108 );
not \mul_7_15_g35105/U$1 ( \5343 , \5342 );
not \mul_7_15_g35027/U$1 ( \5344 , \4026 );
and \mul_7_15_g34662/U$3 ( \5345 , \5343 , \5344 );
nor \mul_7_15_g34662/U$1 ( \5346 , \5341 , \5345 );
not \mul_7_15_g34556/U$1 ( \5347 , \5346 );
not \mul_7_15_g34175/U$3 ( \5348 , \5347 );
not \mul_7_15_g34175/U$4 ( \5349 , \4480 );
or \mul_7_15_g34175/U$2 ( \5350 , \5348 , \5349 );
nand \mul_7_15_g34300/U$1 ( \5351 , \5133 , \4273 );
nand \mul_7_15_g34175/U$1 ( \5352 , \5350 , \5351 );
xor \mul_7_15_g33928/U$4 ( \5353 , \5340 , \5352 );
not \mul_7_15_g34774/U$3 ( \5354 , \4047 );
not \mul_7_15_g34774/U$4 ( \5355 , \4404 );
or \mul_7_15_g34774/U$2 ( \5356 , \5354 , \5355 );
not \mul_7_15_fopt35203/U$1 ( \5357 , \4061 );
nand \mul_7_15_g34854/U$1 ( \5358 , \5357 , \4178 );
nand \mul_7_15_g34774/U$1 ( \5359 , \5356 , \5358 );
not \mul_7_15_g34210/U$3 ( \5360 , \5359 );
not \fopt35523/U$1 ( \5361 , \4066 );
not \mul_7_15_g34210/U$4 ( \5362 , \5361 );
or \mul_7_15_g34210/U$2 ( \5363 , \5360 , \5362 );
nand \mul_7_15_g34429/U$1 ( \5364 , \4562 , \5157 );
nand \mul_7_15_g34210/U$1 ( \5365 , \5363 , \5364 );
and \mul_7_15_g33928/U$3 ( \5366 , \5353 , \5365 );
and \mul_7_15_g33928/U$5 ( \5367 , \5340 , \5352 );
or \mul_7_15_g33928/U$2 ( \5368 , \5366 , \5367 );
and \mul_7_15_g33767/U$2 ( \5369 , \5338 , \5368 );
not \g35834/U$2 ( \5370 , \5330 );
nor \g35834/U$1 ( \5371 , \5370 , \5337 );
nor \mul_7_15_g33767/U$1 ( \5372 , \5369 , \5371 );
not \mul_7_15_g33704/U$1 ( \5373 , \5372 );
nand \mul_7_15_g33612/U$1 ( \5374 , \5327 , \5373 );
or \mul_7_15_g35284/U$1 ( \5375 , \5325 , \5317 );
and \mul_7_15_g35263/U$1 ( \5376 , \5374 , \5375 );
xor \mul_7_15_g33434/U$4 ( \5377 , \5264 , \5376 );
xor \mul_7_15_g33549/U$1 ( \5378 , \5197 , \5199 );
xor \mul_7_15_g33549/U$1_r1 ( \5379 , \5378 , \5202 );
and \mul_7_15_g33434/U$3 ( \5380 , \5377 , \5379 );
and \mul_7_15_g33434/U$5 ( \5381 , \5264 , \5376 );
or \mul_7_15_g33434/U$2 ( \5382 , \5380 , \5381 );
nand \mul_7_15_g33372/U$1 ( \5383 , \5206 , \5382 );
xor \mul_7_15_g33434/U$1 ( \5384 , \5264 , \5376 );
xor \mul_7_15_g33434/U$1_r1 ( \5385 , \5384 , \5379 );
xor \mul_7_15_g33652/U$1 ( \5386 , \5208 , \5258 );
xor \mul_7_15_g33652/U$1_r1 ( \5387 , \5386 , \5261 );
not \mul_7_15_g35061/U$1 ( \5388 , \4048 );
nor \mul_7_15_g34943/U$1 ( \5389 , \5342 , \5388 );
nor \mul_7_15_g34942/U$1 ( \5390 , \3617 , \5270 );
not \mul_7_15_g34335/U$3 ( \5391 , \5390 );
not \mul_7_15_g34789/U$3 ( \5392 , \4044 );
not \mul_7_15_g34789/U$4 ( \5393 , \5270 );
or \mul_7_15_g34789/U$2 ( \5394 , \5392 , \5393 );
nand \mul_7_15_g34908/U$1 ( \5395 , \5273 , \4092 );
nand \mul_7_15_g34789/U$1 ( \5396 , \5394 , \5395 );
not \mul_7_15_g34335/U$4 ( \5397 , \5396 );
or \mul_7_15_g34335/U$2 ( \5398 , \5391 , \5397 );
nand \mul_7_15_g34482/U$1 ( \5399 , \5275 , \5021 );
nand \mul_7_15_g34335/U$1 ( \5400 , \5398 , \5399 );
xor \mul_7_15_g33934/U$4 ( \5401 , \5389 , \5400 );
not \mul_7_15_g34692/U$3 ( \5402 , \4042 );
not \mul_7_15_g34692/U$4 ( \5403 , \5178 );
or \mul_7_15_g34692/U$2 ( \5404 , \5402 , \5403 );
nand \mul_7_15_g34855/U$1 ( \5405 , \4665 , \4116 );
nand \mul_7_15_g34692/U$1 ( \5406 , \5404 , \5405 );
not \mul_7_15_g34248/U$3 ( \5407 , \5406 );
not \mul_7_15_g34248/U$4 ( \5408 , \4661 );
or \mul_7_15_g34248/U$2 ( \5409 , \5407 , \5408 );
nand \mul_7_15_g34354/U$1 ( \5410 , \5225 , \5187 );
nand \mul_7_15_g34248/U$1 ( \5411 , \5409 , \5410 );
and \mul_7_15_g33934/U$3 ( \5412 , \5401 , \5411 );
and \mul_7_15_g33934/U$5 ( \5413 , \5389 , \5400 );
or \mul_7_15_g33934/U$2 ( \5414 , \5412 , \5413 );
not \mul_7_15_g34107/U$3 ( \5415 , \4054 );
not \mul_7_15_g34107/U$4 ( \5416 , \5359 );
or \mul_7_15_g34107/U$2 ( \5417 , \5415 , \5416 );
and \mul_7_15_g34752/U$2 ( \5418 , \4045 , \4403 );
not \mul_7_15_g34752/U$4 ( \5419 , \4045 );
not \mul_7_15_fopt35202/U$1 ( \5420 , \5357 );
and \mul_7_15_g34752/U$3 ( \5421 , \5419 , \5420 );
nor \mul_7_15_g34752/U$1 ( \5422 , \5418 , \5421 );
nand \mul_7_15_g34313/U$1 ( \5423 , \4063 , \4053 , \5422 );
nand \mul_7_15_g34107/U$1 ( \5424 , \5417 , \5423 );
not \mul_7_15_g34704/U$3 ( \5425 , \4046 );
not \mul_7_15_g34704/U$4 ( \5426 , \4145 );
or \mul_7_15_g34704/U$2 ( \5427 , \5425 , \5426 );
nand \mul_7_15_g35974/U$1 ( \5428 , \4109 , \4256 );
nand \mul_7_15_g34704/U$1 ( \5429 , \5427 , \5428 );
not \mul_7_15_g34269/U$3 ( \5430 , \5429 );
not \fopt35686/U$1 ( \5431 , \5209 );
not \mul_7_15_g34269/U$4 ( \5432 , \5431 );
or \mul_7_15_g34269/U$2 ( \5433 , \5430 , \5432 );
nand \mul_7_15_g34495/U$1 ( \5434 , \4139 , \5215 );
nand \mul_7_15_g34269/U$1 ( \5435 , \5433 , \5434 );
xor \mul_7_15_g33952/U$4 ( \5436 , \5424 , \5435 );
not \mul_7_15_g34784/U$3 ( \5437 , \4043 );
not \mul_7_15_g34784/U$4 ( \5438 , \4089 );
or \mul_7_15_g34784/U$2 ( \5439 , \5437 , \5438 );
nand \mul_7_15_g34904/U$1 ( \5440 , \4088 , \4217 );
nand \mul_7_15_g34784/U$1 ( \5441 , \5439 , \5440 );
not \mul_7_15_g34156/U$3 ( \5442 , \5441 );
not \mul_7_15_g34156/U$4 ( \5443 , \4085 );
or \mul_7_15_g34156/U$2 ( \5444 , \5442 , \5443 );
nand \mul_7_15_g34372/U$1 ( \5445 , \4331 , \5238 );
nand \mul_7_15_g34156/U$1 ( \5446 , \5444 , \5445 );
and \mul_7_15_g33952/U$3 ( \5447 , \5436 , \5446 );
and \mul_7_15_g33952/U$5 ( \5448 , \5424 , \5435 );
or \mul_7_15_g33952/U$2 ( \5449 , \5447 , \5448 );
xor \mul_7_15_g33708/U$4 ( \5450 , \5414 , \5449 );
xor \g35437/U$1 ( \5451 , \4023 , \3577 );
nand \mul_7_15_g34499/U$1 ( \5452 , \4229 , \5451 );
or \mul_7_15_g34108/U$2 ( \5453 , \5452 , \4221 );
nand \mul_7_15_g34411/U$1 ( \5454 , \4221 , \5283 );
nand \mul_7_15_g34108/U$1 ( \5455 , \5453 , \5454 );
or \mul_7_15_g34079/U$2 ( \5456 , \5346 , \4252 );
and \g35436/U$2 ( \5457 , \3108 , \5339 );
not \g35436/U$4 ( \5458 , \3108 );
and \g35436/U$3 ( \5459 , \5458 , \4029 );
or \g35436/U$1 ( \5460 , \5457 , \5459 );
nand \mul_7_15_g34103/U$1 ( \5461 , \5460 , \4252 , \4251 );
nand \mul_7_15_g34079/U$1 ( \5462 , \5456 , \5461 );
xor \mul_7_15_g33926/U$4 ( \5463 , \5455 , \5462 );
not \mul_7_15_g34764/U$3 ( \5464 , \3963 );
not \mul_7_15_g34764/U$4 ( \5465 , \4176 );
or \mul_7_15_g34764/U$2 ( \5466 , \5464 , \5465 );
nand \mul_7_15_g34868/U$1 ( \5467 , \4171 , \4486 );
nand \mul_7_15_g34764/U$1 ( \5468 , \5466 , \5467 );
not \mul_7_15_g34112/U$3 ( \5469 , \5468 );
not \mul_7_15_g34112/U$4 ( \5470 , \4194 );
or \mul_7_15_g34112/U$2 ( \5471 , \5469 , \5470 );
nand \mul_7_15_g34481/U$1 ( \5472 , \4204 , \5296 );
nand \mul_7_15_g34112/U$1 ( \5473 , \5471 , \5472 );
and \mul_7_15_g33926/U$3 ( \5474 , \5463 , \5473 );
and \mul_7_15_g33926/U$5 ( \5475 , \5455 , \5462 );
or \mul_7_15_g33926/U$2 ( \5476 , \5474 , \5475 );
and \mul_7_15_g33708/U$3 ( \5477 , \5450 , \5476 );
and \mul_7_15_g33708/U$5 ( \5478 , \5414 , \5449 );
or \mul_7_15_g33708/U$2 ( \5479 , \5477 , \5478 );
not \mul_7_15_g33706/U$1 ( \5480 , \5479 );
not \mul_7_15_g33591/U$3 ( \5481 , \5480 );
xor \mul_7_15_g33977/U$1 ( \5482 , \5277 , \5301 );
xnor \mul_7_15_g33977/U$1_r1 ( \5483 , \5482 , \5288 );
not \mul_7_15_g33804/U$3 ( \5484 , \5483 );
xor \mul_7_15_g33925/U$1 ( \5485 , \5220 , \5231 );
xor \mul_7_15_g33925/U$1_r1 ( \5486 , \5485 , \5243 );
not \mul_7_15_g33923/U$1 ( \5487 , \5486 );
not \mul_7_15_g33804/U$4 ( \5488 , \5487 );
or \mul_7_15_g33804/U$2 ( \5489 , \5484 , \5488 );
or \mul_7_15_g33835/U$2 ( \5490 , \5487 , \5483 );
xor \mul_7_15_g33928/U$1 ( \5491 , \5340 , \5352 );
xor \mul_7_15_g33928/U$1_r1 ( \5492 , \5491 , \5365 );
nand \mul_7_15_g33835/U$1 ( \5493 , \5490 , \5492 );
nand \mul_7_15_g33804/U$1 ( \5494 , \5489 , \5493 );
not \mul_7_15_g33762/U$1 ( \5495 , \5494 );
not \mul_7_15_g33591/U$4 ( \5496 , \5495 );
or \mul_7_15_g33591/U$2 ( \5497 , \5481 , \5496 );
xor \g35833/U$1 ( \5498 , \5330 , \5337 );
xnor \g35833/U$1_r1 ( \5499 , \5498 , \5368 );
nand \mul_7_15_g33591/U$1 ( \5500 , \5497 , \5499 );
not \mul_7_15_g35291/U$2 ( \5501 , \5495 );
nand \mul_7_15_g35291/U$1 ( \5502 , \5501 , \5479 );
and \g35817/U$1 ( \5503 , \5500 , \5502 );
xor \mul_7_15_g33429/U$4 ( \5504 , \5387 , \5503 );
xor \mul_7_15_g33568/U$1 ( \5505 , \5372 , \5324 );
xnor \mul_7_15_g33568/U$1_r1 ( \5506 , \5505 , \5317 );
and \mul_7_15_g33429/U$3 ( \5507 , \5504 , \5506 );
and \mul_7_15_g33429/U$5 ( \5508 , \5387 , \5503 );
or \mul_7_15_g33429/U$2 ( \5509 , \5507 , \5508 );
nand \mul_7_15_g33400/U$1 ( \5510 , \5385 , \5509 );
and \mul_7_15_g33361/U$1 ( \5511 , \5383 , \5510 );
and \g35891/U$2 ( \5512 , \4472 , \4504 );
not \g35891/U$4 ( \5513 , \4472 );
and \g35891/U$3 ( \5514 , \5513 , \4505 );
or \g35891/U$1 ( \5515 , \5512 , \5514 );
and \mul_7_15_g33770/U$2 ( \5516 , \5515 , \4464 );
not \mul_7_15_g33770/U$4 ( \5517 , \5515 );
not \mul_7_15_g33938/U$1 ( \5518 , \4464 );
and \mul_7_15_g33770/U$3 ( \5519 , \5517 , \5518 );
nor \mul_7_15_g33770/U$1 ( \5520 , \5516 , \5519 );
not \mul_7_15_g33623/U$3 ( \5521 , \4617 );
not \mul_7_15_g33623/U$4 ( \5522 , \4627 );
or \mul_7_15_g33623/U$2 ( \5523 , \5521 , \5522 );
or \mul_7_15_g33623/U$5 ( \5524 , \4617 , \4627 );
nand \mul_7_15_g33623/U$1 ( \5525 , \5523 , \5524 );
and \mul_7_15_g33550/U$2 ( \5526 , \4684 , \5525 );
not \mul_7_15_g33550/U$4 ( \5527 , \4684 );
not \mul_7_15_g33598/U$1 ( \5528 , \5525 );
and \mul_7_15_g33550/U$3 ( \5529 , \5527 , \5528 );
nor \mul_7_15_g33550/U$1 ( \5530 , \5526 , \5529 );
xor \g35504/U$1 ( \5531 , \5520 , \5530 );
not \mul_7_15_g33611/U$3 ( \5532 , \5124 );
not \mul_7_15_g33611/U$4 ( \5533 , \5046 );
or \mul_7_15_g33611/U$2 ( \5534 , \5532 , \5533 );
nand \mul_7_15_g33611/U$1 ( \5535 , \5534 , \5117 );
or \mul_7_15_g35283/U$1 ( \5536 , \5124 , \5046 );
nand \mul_7_15_g33597/U$1 ( \5537 , \5535 , \5536 );
xor \g35504/U$1_r1 ( \5538 , \5531 , \5537 );
xor \mul_7_15_g33409/U$4 ( \5539 , \5044 , \5125 );
and \mul_7_15_g33409/U$3 ( \5540 , \5539 , \5205 );
and \mul_7_15_g33409/U$5 ( \5541 , \5044 , \5125 );
or \mul_7_15_g33409/U$2 ( \5542 , \5540 , \5541 );
nand \mul_7_15_g33358/U$1 ( \5543 , \5538 , \5542 );
not \mul_7_15_g33406/U$3 ( \5544 , \5520 );
not \mul_7_15_g33516/U$1 ( \5545 , \5530 );
not \mul_7_15_g33406/U$4 ( \5546 , \5545 );
or \mul_7_15_g33406/U$2 ( \5547 , \5544 , \5546 );
not \mul_7_15_g33722/U$1 ( \5548 , \5520 );
not \mul_7_15_g33423/U$3 ( \5549 , \5548 );
not \mul_7_15_g33423/U$4 ( \5550 , \5530 );
or \mul_7_15_g33423/U$2 ( \5551 , \5549 , \5550 );
nand \mul_7_15_g33423/U$1 ( \5552 , \5551 , \5537 );
nand \mul_7_15_g33406/U$1 ( \5553 , \5547 , \5552 );
not \mul_7_15_g33356/U$2 ( \5554 , \5553 );
xor \mul_7_15_g33480/U$1 ( \5555 , \4518 , \4530 );
xnor \mul_7_15_g33480/U$1_r1 ( \5556 , \5555 , \4690 );
nand \mul_7_15_g33356/U$1 ( \5557 , \5554 , \5556 );
nand \mul_7_15_g33332/U$1 ( \5558 , \5543 , \5557 );
not \mul_7_15_g33331/U$1 ( \5559 , \5558 );
and \mul_7_15_g33321/U$1 ( \5560 , \5511 , \5559 );
not \mul_7_15_g33302/U$3 ( \5561 , \5560 );
xor \mul_7_15_g33429/U$1 ( \5562 , \5387 , \5503 );
xor \mul_7_15_g33429/U$1_r1 ( \5563 , \5562 , \5506 );
and \g35890/U$2 ( \5564 , \5308 , \5305 );
not \g35890/U$4 ( \5565 , \5308 );
and \g35890/U$3 ( \5566 , \5565 , \5306 );
or \g35890/U$1 ( \5567 , \5564 , \5566 );
xnor \mul_7_15_g35296/U$1 ( \5568 , \5567 , \5314 );
not \mul_7_15_g34563/U$3 ( \5569 , \5388 );
not \mul_7_15_g34563/U$4 ( \5570 , \4244 );
or \mul_7_15_g34563/U$2 ( \5571 , \5569 , \5570 );
nand \mul_7_15_g34563/U$1 ( \5572 , \5571 , \4492 );
nand \mul_7_15_g34816/U$1 ( \5573 , \4245 , \4048 );
and \mul_7_15_g34530/U$1 ( \5574 , \5572 , \4156 , \5573 );
not \mul_7_15_g34797/U$3 ( \5575 , \3943 );
not \mul_7_15_g35044/U$1 ( \5576 , \5016 );
not \mul_7_15_g34797/U$4 ( \5577 , \5576 );
or \mul_7_15_g34797/U$2 ( \5578 , \5575 , \5577 );
nand \mul_7_15_g34936/U$1 ( \5579 , \5016 , \4147 );
nand \mul_7_15_g34797/U$1 ( \5580 , \5578 , \5579 );
not \mul_7_15_g34321/U$3 ( \5581 , \5580 );
not \mul_7_15_g34321/U$4 ( \5582 , \5019 );
or \mul_7_15_g34321/U$2 ( \5583 , \5581 , \5582 );
nand \mul_7_15_g34370/U$1 ( \5584 , \5396 , \5021 );
nand \mul_7_15_g34321/U$1 ( \5585 , \5583 , \5584 );
and \mul_7_15_g35265/U$1 ( \5586 , \5574 , \5585 );
xor \mul_7_15_g33934/U$1 ( \5587 , \5389 , \5400 );
xor \mul_7_15_g33934/U$1_r1 ( \5588 , \5587 , \5411 );
xor \mul_7_15_g33744/U$4 ( \5589 , \5586 , \5588 );
not \mul_7_15_g34723/U$3 ( \5590 , \4011 );
not \mul_7_15_g34723/U$4 ( \5591 , \5234 );
or \mul_7_15_g34723/U$2 ( \5592 , \5590 , \5591 );
nand \mul_7_15_g34877/U$1 ( \5593 , \4088 , \4270 );
nand \mul_7_15_g34723/U$1 ( \5594 , \5592 , \5593 );
not \mul_7_15_g34142/U$3 ( \5595 , \5594 );
not \mul_7_15_g34142/U$4 ( \5596 , \4437 );
or \mul_7_15_g34142/U$2 ( \5597 , \5595 , \5596 );
nand \mul_7_15_g34373/U$1 ( \5598 , \4596 , \5441 );
nand \mul_7_15_g34142/U$1 ( \5599 , \5597 , \5598 );
not \mul_7_15_g34712/U$3 ( \5600 , \3958 );
not \mul_7_15_g34712/U$4 ( \5601 , \4142 );
or \mul_7_15_g34712/U$2 ( \5602 , \5600 , \5601 );
nand \mul_7_15_g34910/U$1 ( \5603 , \4109 , \4473 );
nand \mul_7_15_g34712/U$1 ( \5604 , \5602 , \5603 );
not \mul_7_15_g34253/U$3 ( \5605 , \5604 );
not \mul_7_15_g34253/U$4 ( \5606 , \4425 );
or \mul_7_15_g34253/U$2 ( \5607 , \5605 , \5606 );
nand \mul_7_15_g34387/U$1 ( \5608 , \4139 , \5429 );
nand \mul_7_15_g34253/U$1 ( \5609 , \5607 , \5608 );
nor \mul_7_15_g34058/U$1 ( \5610 , \5599 , \5609 );
not \mul_7_15_g34736/U$3 ( \5611 , \4047 );
not \mul_7_15_g34736/U$4 ( \5612 , \4666 );
or \mul_7_15_g34736/U$2 ( \5613 , \5611 , \5612 );
nand \mul_7_15_g34869/U$1 ( \5614 , \4548 , \4178 );
nand \mul_7_15_g34736/U$1 ( \5615 , \5613 , \5614 );
not \mul_7_15_g34232/U$3 ( \5616 , \5615 );
not \mul_7_15_g34232/U$4 ( \5617 , \4661 );
or \mul_7_15_g34232/U$2 ( \5618 , \5616 , \5617 );
nand \mul_7_15_g34393/U$1 ( \5619 , \4672 , \5406 );
nand \mul_7_15_g34232/U$1 ( \5620 , \5618 , \5619 );
not \fopt35793/U$1 ( \5621 , \5620 );
or \mul_7_15_g34001/U$2 ( \5622 , \5610 , \5621 );
nand \mul_7_15_g34057/U$1 ( \5623 , \5599 , \5609 );
nand \mul_7_15_g34001/U$1 ( \5624 , \5622 , \5623 );
and \mul_7_15_g33744/U$3 ( \5625 , \5589 , \5624 );
and \mul_7_15_g33744/U$5 ( \5626 , \5586 , \5588 );
or \mul_7_15_g33744/U$2 ( \5627 , \5625 , \5626 );
xor \mul_7_15_g33708/U$1 ( \5628 , \5414 , \5449 );
xor \mul_7_15_g33708/U$1_r1 ( \5629 , \5628 , \5476 );
xor \mul_7_15_g33543/U$4 ( \5630 , \5627 , \5629 );
xor \mul_7_15_g33952/U$1 ( \5631 , \5424 , \5435 );
xor \mul_7_15_g33952/U$1_r1 ( \5632 , \5631 , \5446 );
xor \mul_7_15_g33926/U$1 ( \5633 , \5455 , \5462 );
xor \mul_7_15_g33926/U$1_r1 ( \5634 , \5633 , \5473 );
xor \mul_7_15_g33672/U$4 ( \5635 , \5632 , \5634 );
not \mul_7_15_g34766/U$3 ( \5636 , \4041 );
not \mul_7_15_g34766/U$4 ( \5637 , \4069 );
or \mul_7_15_g34766/U$2 ( \5638 , \5636 , \5637 );
nand \mul_7_15_g34882/U$1 ( \5639 , \5060 , \4238 );
nand \mul_7_15_g34766/U$1 ( \5640 , \5638 , \5639 );
not \mul_7_15_g34169/U$3 ( \5641 , \5640 );
not \mul_7_15_g34169/U$4 ( \5642 , \4065 );
or \mul_7_15_g34169/U$2 ( \5643 , \5641 , \5642 );
nand \mul_7_15_g34361/U$1 ( \5644 , \5422 , \4055 );
nand \mul_7_15_g34169/U$1 ( \5645 , \5643 , \5644 );
not \mul_7_15_g34679/U$3 ( \5646 , \4585 );
not \mul_7_15_g34679/U$4 ( \5647 , \4171 );
or \mul_7_15_g34679/U$2 ( \5648 , \5646 , \5647 );
nand \mul_7_15_g34847/U$1 ( \5649 , \4284 , \4019 );
nand \mul_7_15_g34679/U$1 ( \5650 , \5648 , \5649 );
not \mul_7_15_g34115/U$3 ( \5651 , \5650 );
not \mul_7_15_g34115/U$4 ( \5652 , \4194 );
or \mul_7_15_g34115/U$2 ( \5653 , \5651 , \5652 );
nand \mul_7_15_g35969/U$1 ( \5654 , \5111 , \5468 );
nand \mul_7_15_g34115/U$1 ( \5655 , \5653 , \5654 );
xor \mul_7_15_g33882/U$4 ( \5656 , \5645 , \5655 );
and \mul_7_15_g34803/U$2 ( \5657 , \5388 , \4267 );
not \mul_7_15_g34803/U$4 ( \5658 , \5388 );
and \mul_7_15_g34803/U$3 ( \5659 , \5658 , \4156 );
nor \mul_7_15_g34803/U$1 ( \5660 , \5657 , \5659 );
not \mul_7_15_g34166/U$3 ( \5661 , \5660 );
not \mul_7_15_g34166/U$4 ( \5662 , \4253 );
or \mul_7_15_g34166/U$2 ( \5663 , \5661 , \5662 );
nand \mul_7_15_g34305/U$1 ( \5664 , \4273 , \5460 );
nand \mul_7_15_g34166/U$1 ( \5665 , \5663 , \5664 );
and \mul_7_15_g33882/U$3 ( \5666 , \5656 , \5665 );
and \mul_7_15_g33882/U$5 ( \5667 , \5645 , \5655 );
or \mul_7_15_g33882/U$2 ( \5668 , \5666 , \5667 );
and \mul_7_15_g33672/U$3 ( \5669 , \5635 , \5668 );
and \mul_7_15_g33672/U$5 ( \5670 , \5632 , \5634 );
or \mul_7_15_g33672/U$2 ( \5671 , \5669 , \5670 );
and \mul_7_15_g33543/U$3 ( \5672 , \5630 , \5671 );
and \mul_7_15_g33543/U$5 ( \5673 , \5627 , \5629 );
or \mul_7_15_g33543/U$2 ( \5674 , \5672 , \5673 );
not \mul_7_15_g33542/U$1 ( \5675 , \5674 );
xor \mul_7_15_g33431/U$4 ( \5676 , \5568 , \5675 );
xor \mul_7_15_g33582/U$1 ( \5677 , \5479 , \5494 );
xnor \mul_7_15_g33582/U$1_r1 ( \5678 , \5677 , \5499 );
and \mul_7_15_g33431/U$3 ( \5679 , \5676 , \5678 );
and \mul_7_15_g33431/U$5 ( \5680 , \5568 , \5675 );
or \mul_7_15_g33431/U$2 ( \5681 , \5679 , \5680 );
nand \mul_7_15_g33397/U$1 ( \5682 , \5563 , \5681 );
xor \mul_7_15_g33431/U$1 ( \5683 , \5568 , \5675 );
xor \mul_7_15_g33431/U$1_r1 ( \5684 , \5683 , \5678 );
xor \mul_7_15_g33543/U$1 ( \5685 , \5627 , \5629 );
xor \mul_7_15_g33543/U$1_r1 ( \5686 , \5685 , \5671 );
buf \mul_7_15_fopt35209/U$1 ( \5687 , \5686 );
not \mul_7_15_fopt35207/U$1 ( \5688 , \5687 );
xor \g35501/U$1 ( \5689 , \5486 , \5492 );
xor \g35501/U$1_r1 ( \5690 , \5689 , \5483 );
buf \mul_7_15_g33760/U$1 ( \5691 , \5690 );
nand \mul_7_15_g33507/U$1 ( \5692 , \5688 , \5691 );
xor \mul_7_15_g35340/U$1 ( \5693 , \5344 , \4492 );
not \mul_7_15_g34759/U$1 ( \5694 , \5693 );
not \mul_7_15_g34177/U$3 ( \5695 , \5694 );
not \mul_7_15_g34177/U$4 ( \5696 , \4231 );
or \mul_7_15_g34177/U$2 ( \5697 , \5695 , \5696 );
nand \mul_7_15_g34375/U$1 ( \5698 , \4234 , \5451 );
nand \mul_7_15_g34177/U$1 ( \5699 , \5697 , \5698 );
xor \g35424/U$1 ( \5700 , \5574 , \5585 );
xor \mul_7_15_g33812/U$4 ( \5701 , \5699 , \5700 );
not \mul_7_15_g34788/U$3 ( \5702 , \4042 );
not \mul_7_15_g34788/U$4 ( \5703 , \5270 );
or \mul_7_15_g34788/U$2 ( \5704 , \5702 , \5703 );
nand \mul_7_15_g34864/U$1 ( \5705 , \5273 , \4116 );
nand \mul_7_15_g34788/U$1 ( \5706 , \5704 , \5705 );
and \mul_7_15_g34323/U$2 ( \5707 , \5019 , \5706 );
and \mul_7_15_g34323/U$3 ( \5708 , \5580 , \5021 );
nor \mul_7_15_g34323/U$1 ( \5709 , \5707 , \5708 );
not \mul_7_15_g34322/U$1 ( \5710 , \5709 );
not \mul_7_15_g33963/U$3 ( \5711 , \5710 );
not \mul_7_15_g34517/U$2 ( \5712 , \4252 );
nand \mul_7_15_g34517/U$1 ( \5713 , \5712 , \4048 );
not \mul_7_15_g34515/U$1 ( \5714 , \5713 );
not \mul_7_15_g33963/U$4 ( \5715 , \5714 );
or \mul_7_15_g33963/U$2 ( \5716 , \5711 , \5715 );
not \mul_7_15_g34728/U$3 ( \5717 , \4045 );
not \mul_7_15_g34728/U$4 ( \5718 , \5178 );
or \mul_7_15_g34728/U$2 ( \5719 , \5717 , \5718 );
nand \mul_7_15_g34862/U$1 ( \5720 , \4665 , \4286 );
nand \mul_7_15_g34728/U$1 ( \5721 , \5719 , \5720 );
not \mul_7_15_g34234/U$3 ( \5722 , \5721 );
not \mul_7_15_g34234/U$4 ( \5723 , \4662 );
or \mul_7_15_g34234/U$2 ( \5724 , \5722 , \5723 );
nand \mul_7_15_g34377/U$1 ( \5725 , \4672 , \5615 );
nand \mul_7_15_g34234/U$1 ( \5726 , \5724 , \5725 );
nand \mul_7_15_g34095/U$1 ( \5727 , \5713 , \5709 );
nand \mul_7_15_g33992/U$1 ( \5728 , \5726 , \5727 );
nand \mul_7_15_g33963/U$1 ( \5729 , \5716 , \5728 );
and \mul_7_15_g33812/U$3 ( \5730 , \5701 , \5729 );
and \mul_7_15_g33812/U$5 ( \5731 , \5699 , \5700 );
or \mul_7_15_g33812/U$2 ( \5732 , \5730 , \5731 );
xor \mul_7_15_g33744/U$1 ( \5733 , \5586 , \5588 );
xor \mul_7_15_g33744/U$1_r1 ( \5734 , \5733 , \5624 );
xor \mul_7_15_g33569/U$4 ( \5735 , \5732 , \5734 );
xor \mul_7_15_g33672/U$1 ( \5736 , \5632 , \5634 );
xor \mul_7_15_g33672/U$1_r1 ( \5737 , \5736 , \5668 );
and \mul_7_15_g33569/U$3 ( \5738 , \5735 , \5737 );
and \mul_7_15_g33569/U$5 ( \5739 , \5732 , \5734 );
or \mul_7_15_g33569/U$2 ( \5740 , \5738 , \5739 );
and \mul_7_15_g33426/U$2 ( \5741 , \5692 , \5740 );
nor \mul_7_15_g33512/U$1 ( \5742 , \5688 , \5691 );
nor \mul_7_15_g33426/U$1 ( \5743 , \5741 , \5742 );
nand \mul_7_15_g33383/U$1 ( \5744 , \5684 , \5743 );
and \mul_7_15_g33359/U$1 ( \5745 , \5682 , \5744 );
not \mul_7_15_g34687/U$3 ( \5746 , \4011 );
not \mul_7_15_g34687/U$4 ( \5747 , \4404 );
or \mul_7_15_g34687/U$2 ( \5748 , \5746 , \5747 );
not \mul_7_15_fopt35191/U$1 ( \5749 , \4069 );
nand \mul_7_15_g34898/U$1 ( \5750 , \5749 , \4270 );
nand \mul_7_15_g34687/U$1 ( \5751 , \5748 , \5750 );
not \mul_7_15_g34197/U$3 ( \5752 , \5751 );
not \mul_7_15_g34197/U$4 ( \5753 , \4558 );
or \mul_7_15_g34197/U$2 ( \5754 , \5752 , \5753 );
not \mul_7_15_g34738/U$3 ( \5755 , \4043 );
not \mul_7_15_g34738/U$4 ( \5756 , \4069 );
or \mul_7_15_g34738/U$2 ( \5757 , \5755 , \5756 );
nand \mul_7_15_g34917/U$1 ( \5758 , \5749 , \4217 );
nand \mul_7_15_g34738/U$1 ( \5759 , \5757 , \5758 );
nand \mul_7_15_g34431/U$1 ( \5760 , \4562 , \5759 );
nand \mul_7_15_g34197/U$1 ( \5761 , \5754 , \5760 );
not \mul_7_15_g34809/U$3 ( \5762 , \4048 );
not \mul_7_15_g34809/U$4 ( \5763 , \4212 );
or \mul_7_15_g34809/U$2 ( \5764 , \5762 , \5763 );
nand \mul_7_15_g34945/U$1 ( \5765 , \4492 , \5388 );
nand \mul_7_15_g34809/U$1 ( \5766 , \5764 , \5765 );
not \mul_7_15_g34196/U$3 ( \5767 , \5766 );
not \mul_7_15_g34196/U$4 ( \5768 , \4231 );
or \mul_7_15_g34196/U$2 ( \5769 , \5767 , \5768 );
not \mul_7_15_g34697/U$3 ( \5770 , \4029 );
not \mul_7_15_g34697/U$4 ( \5771 , \4212 );
or \mul_7_15_g34697/U$2 ( \5772 , \5770 , \5771 );
nand \mul_7_15_g34925/U$1 ( \5773 , \4492 , \5339 );
nand \mul_7_15_g34697/U$1 ( \5774 , \5772 , \5773 );
nand \mul_7_15_g34425/U$1 ( \5775 , \4234 , \5774 );
nand \mul_7_15_g34196/U$1 ( \5776 , \5769 , \5775 );
xor \mul_7_15_g33914/U$4 ( \5777 , \5761 , \5776 );
not \mul_7_15_g34745/U$3 ( \5778 , \4026 );
not \mul_7_15_g34745/U$4 ( \5779 , \4173 );
or \mul_7_15_g34745/U$2 ( \5780 , \5778 , \5779 );
nand \mul_7_15_g34867/U$1 ( \5781 , \4177 , \5344 );
nand \mul_7_15_g34745/U$1 ( \5782 , \5780 , \5781 );
not \mul_7_15_g34118/U$3 ( \5783 , \5782 );
not \mul_7_15_g34118/U$4 ( \5784 , \4194 );
or \mul_7_15_g34118/U$2 ( \5785 , \5783 , \5784 );
not \mul_7_15_g34779/U$3 ( \5786 , \4023 );
not \mul_7_15_g34779/U$4 ( \5787 , \4184 );
or \mul_7_15_g34779/U$2 ( \5788 , \5786 , \5787 );
nand \mul_7_15_g34903/U$1 ( \5789 , \4171 , \5131 );
nand \mul_7_15_g34779/U$1 ( \5790 , \5788 , \5789 );
nand \mul_7_15_g34490/U$1 ( \5791 , \5111 , \5790 );
nand \mul_7_15_g34118/U$1 ( \5792 , \5785 , \5791 );
and \mul_7_15_g33914/U$3 ( \5793 , \5777 , \5792 );
and \mul_7_15_g33914/U$5 ( \5794 , \5761 , \5776 );
or \mul_7_15_g33914/U$2 ( \5795 , \5793 , \5794 );
not \mul_7_15_g33913/U$1 ( \5796 , \5795 );
nand \mul_7_15_g34817/U$1 ( \5797 , \4224 , \5388 );
and \mul_7_15_g34535/U$2 ( \5798 , \5797 , \4172 );
not \mul_7_15_g34566/U$3 ( \5799 , \4048 );
not \mul_7_15_g35033/U$1 ( \5800 , \4224 );
not \mul_7_15_g34566/U$4 ( \5801 , \5800 );
or \mul_7_15_g34566/U$2 ( \5802 , \5799 , \5801 );
nand \mul_7_15_g34566/U$1 ( \5803 , \5802 , \4492 );
nor \mul_7_15_g34535/U$1 ( \5804 , \5798 , \5803 );
not \mul_7_15_g34791/U$3 ( \5805 , \4047 );
not \mul_7_15_g34791/U$4 ( \5806 , \5270 );
or \mul_7_15_g34791/U$2 ( \5807 , \5805 , \5806 );
nand \mul_7_15_g34896/U$1 ( \5808 , \5016 , \4178 );
nand \mul_7_15_g34791/U$1 ( \5809 , \5807 , \5808 );
not \mul_7_15_g34326/U$3 ( \5810 , \5809 );
not \mul_7_15_g34326/U$4 ( \5811 , \5390 );
or \mul_7_15_g34326/U$2 ( \5812 , \5810 , \5811 );
nand \mul_7_15_g34422/U$1 ( \5813 , \5706 , \5021 );
nand \mul_7_15_g34326/U$1 ( \5814 , \5812 , \5813 );
nand \mul_7_15_g34100/U$1 ( \5815 , \5804 , \5814 );
not \mul_7_15_g34633/U$1 ( \5816 , \4192 );
and \g36018/U$2 ( \5817 , \5816 , \5650 );
not \g36018/U$4 ( \5818 , \5816 );
and \g36019/U$1 ( \5819 , \5790 , \4186 );
and \g36018/U$3 ( \5820 , \5818 , \5819 );
nor \g36018/U$1 ( \5821 , \5817 , \5820 );
xor \mul_7_15_g33852/U$1 ( \5822 , \5815 , \5821 );
not \mul_7_15_g34192/U$3 ( \5823 , \4230 );
not \mul_7_15_g34696/U$1 ( \5824 , \5774 );
not \mul_7_15_g34192/U$4 ( \5825 , \5824 );
and \mul_7_15_g34192/U$2 ( \5826 , \5823 , \5825 );
not \g35836/U$2 ( \5827 , \4234 );
nor \g35836/U$1 ( \5828 , \5827 , \5693 );
nor \mul_7_15_g34192/U$1 ( \5829 , \5826 , \5828 );
xor \mul_7_15_g33852/U$1_r1 ( \5830 , \5822 , \5829 );
nand \mul_7_15_g33798/U$1 ( \5831 , \5796 , \5830 );
not \mul_7_15_g33648/U$3 ( \5832 , \5831 );
xor \g35425/U$1 ( \5833 , \5804 , \5814 );
and \g35743/U$1 ( \5834 , \4234 , \4048 );
not \mul_7_15_g34762/U$3 ( \5835 , \3963 );
not \mul_7_15_g34762/U$4 ( \5836 , \5234 );
or \mul_7_15_g34762/U$2 ( \5837 , \5835 , \5836 );
nand \mul_7_15_g34927/U$1 ( \5838 , \4088 , \4486 );
nand \mul_7_15_g34762/U$1 ( \5839 , \5837 , \5838 );
not \mul_7_15_g34149/U$3 ( \5840 , \5839 );
not \mul_7_15_g34149/U$4 ( \5841 , \4085 );
or \mul_7_15_g34149/U$2 ( \5842 , \5840 , \5841 );
not \mul_7_15_g34721/U$3 ( \5843 , \3958 );
not \mul_7_15_g34721/U$4 ( \5844 , \5234 );
or \mul_7_15_g34721/U$2 ( \5845 , \5843 , \5844 );
nand \mul_7_15_g34884/U$1 ( \5846 , \4088 , \4473 );
nand \mul_7_15_g34721/U$1 ( \5847 , \5845 , \5846 );
nand \mul_7_15_g34432/U$1 ( \5848 , \4596 , \5847 );
nand \mul_7_15_g34149/U$1 ( \5849 , \5842 , \5848 );
or \g35742/U$2 ( \5850 , \5834 , \5849 );
not \mul_7_15_g34717/U$3 ( \5851 , \4043 );
not \mul_7_15_g34717/U$4 ( \5852 , \5178 );
or \mul_7_15_g34717/U$2 ( \5853 , \5851 , \5852 );
nand \mul_7_15_g34873/U$1 ( \5854 , \4548 , \4217 );
nand \mul_7_15_g34717/U$1 ( \5855 , \5853 , \5854 );
not \mul_7_15_g34239/U$3 ( \5856 , \5855 );
not \mul_7_15_g34239/U$4 ( \5857 , \4662 );
or \mul_7_15_g34239/U$2 ( \5858 , \5856 , \5857 );
not \mul_7_15_g34730/U$3 ( \5859 , \4041 );
not \mul_7_15_g34730/U$4 ( \5860 , \4666 );
or \mul_7_15_g34730/U$2 ( \5861 , \5859 , \5860 );
nand \mul_7_15_g34860/U$1 ( \5862 , \4665 , \4238 );
nand \mul_7_15_g34730/U$1 ( \5863 , \5861 , \5862 );
nand \mul_7_15_g34496/U$1 ( \5864 , \4672 , \5863 );
nand \mul_7_15_g34239/U$1 ( \5865 , \5858 , \5864 );
nand \g35742/U$1 ( \5866 , \5850 , \5865 );
nand \mul_7_15_g35745/U$1 ( \5867 , \4234 , \4048 );
not \g35852/U$2 ( \5868 , \5867 );
nand \g35852/U$1 ( \5869 , \5868 , \5849 );
nand \mul_7_15_g33993/U$1 ( \5870 , \5866 , \5869 );
xor \mul_7_15_g33703/U$4 ( \5871 , \5833 , \5870 );
not \mul_7_15_g34800/U$3 ( \5872 , \4045 );
buf \mul_7_15_g35054/U$1 ( \5873 , \1395 );
not \mul_7_15_g35053/U$1 ( \5874 , \5873 );
not \mul_7_15_g34800/U$4 ( \5875 , \5874 );
or \mul_7_15_g34800/U$2 ( \5876 , \5872 , \5875 );
nand \mul_7_15_g34901/U$1 ( \5877 , \5273 , \4286 );
nand \mul_7_15_g34800/U$1 ( \5878 , \5876 , \5877 );
not \mul_7_15_g34328/U$3 ( \5879 , \5878 );
not \mul_7_15_g34328/U$4 ( \5880 , \5019 );
or \mul_7_15_g34328/U$2 ( \5881 , \5879 , \5880 );
nand \mul_7_15_g34483/U$1 ( \5882 , \5809 , \5021 );
nand \mul_7_15_g34328/U$1 ( \5883 , \5881 , \5882 );
not \mul_7_15_g33896/U$3 ( \5884 , \5883 );
not \mul_7_15_g34742/U$3 ( \5885 , \4023 );
not \mul_7_15_g34742/U$4 ( \5886 , \4110 );
or \mul_7_15_g34742/U$2 ( \5887 , \5885 , \5886 );
nand \mul_7_15_g34875/U$1 ( \5888 , \4109 , \5131 );
nand \mul_7_15_g34742/U$1 ( \5889 , \5887 , \5888 );
not \mul_7_15_g34268/U$3 ( \5890 , \5889 );
not \mul_7_15_g34268/U$4 ( \5891 , \5431 );
or \mul_7_15_g34268/U$2 ( \5892 , \5890 , \5891 );
not \mul_7_15_g34737/U$3 ( \5893 , \4019 );
not \mul_7_15_g34737/U$4 ( \5894 , \4142 );
or \mul_7_15_g34737/U$2 ( \5895 , \5893 , \5894 );
nand \mul_7_15_g34885/U$1 ( \5896 , \4109 , \4585 );
nand \mul_7_15_g34737/U$1 ( \5897 , \5895 , \5896 );
nand \mul_7_15_g34435/U$1 ( \5898 , \5897 , \4139 );
nand \mul_7_15_g34268/U$1 ( \5899 , \5892 , \5898 );
not \mul_7_15_g33896/U$4 ( \5900 , \5899 );
or \mul_7_15_g33896/U$2 ( \5901 , \5884 , \5900 );
or \mul_7_15_g33956/U$2 ( \5902 , \5899 , \5883 );
not \mul_7_15_g34686/U$3 ( \5903 , \4046 );
buf \mul_7_15_fopt35196/U$1 ( \5904 , \4069 );
not \mul_7_15_g34686/U$4 ( \5905 , \5904 );
or \mul_7_15_g34686/U$2 ( \5906 , \5903 , \5905 );
nand \mul_7_15_g34887/U$1 ( \5907 , \5060 , \4256 );
nand \mul_7_15_g34686/U$1 ( \5908 , \5906 , \5907 );
not \mul_7_15_g34200/U$3 ( \5909 , \5908 );
not \mul_7_15_g34200/U$4 ( \5910 , \5361 );
or \mul_7_15_g34200/U$2 ( \5911 , \5909 , \5910 );
nand \mul_7_15_g34439/U$1 ( \5912 , \4055 , \5751 );
nand \mul_7_15_g34200/U$1 ( \5913 , \5911 , \5912 );
nand \mul_7_15_g33956/U$1 ( \5914 , \5902 , \5913 );
nand \mul_7_15_g33896/U$1 ( \5915 , \5901 , \5914 );
and \mul_7_15_g33703/U$3 ( \5916 , \5871 , \5915 );
and \mul_7_15_g33703/U$5 ( \5917 , \5833 , \5870 );
or \mul_7_15_g33703/U$2 ( \5918 , \5916 , \5917 );
not \mul_7_15_g33648/U$4 ( \5919 , \5918 );
or \mul_7_15_g33648/U$2 ( \5920 , \5832 , \5919 );
or \g35999/U$1 ( \5921 , \5830 , \5796 );
nand \mul_7_15_g33648/U$1 ( \5922 , \5920 , \5921 );
not \mul_7_15_g33579/U$3 ( \5923 , \5922 );
not \mul_7_15_g34188/U$3 ( \5924 , \5759 );
not \mul_7_15_g34188/U$4 ( \5925 , \4558 );
or \mul_7_15_g34188/U$2 ( \5926 , \5924 , \5925 );
nand \mul_7_15_g34364/U$1 ( \5927 , \4055 , \5640 );
nand \mul_7_15_g34188/U$1 ( \5928 , \5926 , \5927 );
not \mul_7_15_g34003/U$3 ( \5929 , \5928 );
not \mul_7_15_g34718/U$3 ( \5930 , \4046 );
not \mul_7_15_g34718/U$4 ( \5931 , \4089 );
or \mul_7_15_g34718/U$2 ( \5932 , \5930 , \5931 );
nand \mul_7_15_g34861/U$1 ( \5933 , \4088 , \4256 );
nand \mul_7_15_g34718/U$1 ( \5934 , \5932 , \5933 );
not \mul_7_15_g34145/U$3 ( \5935 , \5934 );
not \mul_7_15_g34145/U$4 ( \5936 , \4086 );
or \mul_7_15_g34145/U$2 ( \5937 , \5935 , \5936 );
nand \mul_7_15_g34392/U$1 ( \5938 , \4596 , \5594 );
nand \mul_7_15_g34145/U$1 ( \5939 , \5937 , \5938 );
not \mul_7_15_g34003/U$4 ( \5940 , \5939 );
or \mul_7_15_g34003/U$2 ( \5941 , \5929 , \5940 );
or \mul_7_15_g34022/U$2 ( \5942 , \5939 , \5928 );
not \mul_7_15_g34735/U$3 ( \5943 , \3963 );
not \mul_7_15_g34735/U$4 ( \5944 , \4110 );
or \mul_7_15_g34735/U$2 ( \5945 , \5943 , \5944 );
nand \mul_7_15_g34871/U$1 ( \5946 , \4115 , \4486 );
nand \mul_7_15_g34735/U$1 ( \5947 , \5945 , \5946 );
not \mul_7_15_g34265/U$3 ( \5948 , \5947 );
not \mul_7_15_g34265/U$4 ( \5949 , \4425 );
or \mul_7_15_g34265/U$2 ( \5950 , \5948 , \5949 );
nand \mul_7_15_g34383/U$1 ( \5951 , \4429 , \5604 );
nand \mul_7_15_g34265/U$1 ( \5952 , \5950 , \5951 );
nand \mul_7_15_g34022/U$1 ( \5953 , \5942 , \5952 );
nand \mul_7_15_g34003/U$1 ( \5954 , \5941 , \5953 );
xor \g35398/U$1 ( \5955 , \5609 , \5621 );
xnor \g35398/U$1_r1 ( \5956 , \5955 , \5599 );
xor \mul_7_15_g2/U$1 ( \5957 , \5954 , \5956 );
xor \mul_7_15_g33882/U$1 ( \5958 , \5645 , \5655 );
xor \mul_7_15_g33882/U$1_r1 ( \5959 , \5958 , \5665 );
xnor \mul_7_15_g2/U$1_r1 ( \5960 , \5957 , \5959 );
not \mul_7_15_g33579/U$4 ( \5961 , \5960 );
or \mul_7_15_g33579/U$2 ( \5962 , \5923 , \5961 );
not \g35828/U$2 ( \5963 , \5922 );
xor \mul_7_15_g35206/U$1 ( \5964 , \5954 , \5956 );
xor \mul_7_15_g35206/U$1_r1 ( \5965 , \5964 , \5959 );
nand \g35828/U$1 ( \5966 , \5963 , \5965 );
nand \mul_7_15_g33579/U$1 ( \5967 , \5962 , \5966 );
xor \g35894/U$1 ( \5968 , \5928 , \5952 );
not \mul_7_15_g34144/U$1 ( \5969 , \5939 );
and \mul_7_15_g33980/U$2 ( \5970 , \5968 , \5969 );
not \mul_7_15_g33980/U$4 ( \5971 , \5968 );
and \mul_7_15_g33980/U$3 ( \5972 , \5971 , \5939 );
nor \mul_7_15_g33980/U$1 ( \5973 , \5970 , \5972 );
xor \g35893/U$1 ( \5974 , \5709 , \5714 );
xor \g35893/U$1_r1 ( \5975 , \5974 , \5726 );
nand \mul_7_15_g33866/U$1 ( \5976 , \5973 , \5975 );
not \mul_7_15_g34147/U$3 ( \5977 , \5847 );
not \mul_7_15_g34147/U$4 ( \5978 , \4086 );
or \mul_7_15_g34147/U$2 ( \5979 , \5977 , \5978 );
nand \mul_7_15_g34341/U$1 ( \5980 , \4596 , \5934 );
nand \mul_7_15_g34147/U$1 ( \5981 , \5979 , \5980 );
not \mul_7_15_g34004/U$3 ( \5982 , \5981 );
not \mul_7_15_g34267/U$3 ( \5983 , \4425 );
not \mul_7_15_g34267/U$4 ( \5984 , \5897 );
or \mul_7_15_g34267/U$2 ( \5985 , \5983 , \5984 );
nand \mul_7_15_g34497/U$1 ( \5986 , \4140 , \5947 );
nand \mul_7_15_g34267/U$1 ( \5987 , \5985 , \5986 );
not \mul_7_15_g34004/U$4 ( \5988 , \5987 );
or \mul_7_15_g34004/U$2 ( \5989 , \5982 , \5988 );
or \mul_7_15_g34019/U$2 ( \5990 , \5981 , \5987 );
not \mul_7_15_g34238/U$3 ( \5991 , \5863 );
not \mul_7_15_g34238/U$4 ( \5992 , \4662 );
or \mul_7_15_g34238/U$2 ( \5993 , \5991 , \5992 );
nand \mul_7_15_g34412/U$1 ( \5994 , \4672 , \5721 );
nand \mul_7_15_g34238/U$1 ( \5995 , \5993 , \5994 );
nand \mul_7_15_g34019/U$1 ( \5996 , \5990 , \5995 );
nand \mul_7_15_g34004/U$1 ( \5997 , \5989 , \5996 );
and \mul_7_15_g33805/U$2 ( \5998 , \5976 , \5997 );
nor \mul_7_15_g33864/U$1 ( \5999 , \5973 , \5975 );
nor \mul_7_15_g33805/U$1 ( \6000 , \5998 , \5999 );
not \mul_7_15_g33752/U$1 ( \6001 , \6000 );
not \mul_7_15_g33654/U$3 ( \6002 , \6001 );
xor \mul_7_15_g33852/U$4 ( \6003 , \5815 , \5821 );
and \mul_7_15_g33852/U$3 ( \6004 , \6003 , \5829 );
and \mul_7_15_g33852/U$5 ( \6005 , \5815 , \5821 );
or \mul_7_15_g33852/U$2 ( \6006 , \6004 , \6005 );
not \mul_7_15_g33764/U$3 ( \6007 , \6006 );
xor \mul_7_15_g33812/U$1 ( \6008 , \5699 , \5700 );
xor \mul_7_15_g33812/U$1_r1 ( \6009 , \6008 , \5729 );
not \mul_7_15_g33764/U$4 ( \6010 , \6009 );
or \mul_7_15_g33764/U$2 ( \6011 , \6007 , \6010 );
or \mul_7_15_g33764/U$5 ( \6012 , \6009 , \6006 );
nand \mul_7_15_g33764/U$1 ( \6013 , \6011 , \6012 );
not \mul_7_15_g33705/U$1 ( \6014 , \6013 );
not \mul_7_15_g33654/U$4 ( \6015 , \6014 );
or \mul_7_15_g33654/U$2 ( \6016 , \6002 , \6015 );
nand \mul_7_15_g33656/U$1 ( \6017 , \6013 , \6000 );
nand \mul_7_15_g33654/U$1 ( \6018 , \6016 , \6017 );
not \mul_7_15_g33621/U$1 ( \6019 , \6018 );
and \mul_7_15_g33517/U$2 ( \6020 , \5967 , \6019 );
not \mul_7_15_g33517/U$4 ( \6021 , \5967 );
and \mul_7_15_g33517/U$3 ( \6022 , \6021 , \6018 );
nor \mul_7_15_g33517/U$1 ( \6023 , \6020 , \6022 );
not \mul_7_15_g33790/U$3 ( \6024 , \5795 );
not \mul_7_15_g33790/U$4 ( \6025 , \5830 );
or \mul_7_15_g33790/U$2 ( \6026 , \6024 , \6025 );
or \mul_7_15_g33790/U$5 ( \6027 , \5795 , \5830 );
nand \mul_7_15_g33790/U$1 ( \6028 , \6026 , \6027 );
xor \g35886/U$1 ( \6029 , \6028 , \5918 );
not \mul_7_15_g33856/U$3 ( \6030 , \5975 );
not \mul_7_15_g33856/U$4 ( \6031 , \5997 );
or \mul_7_15_g33856/U$2 ( \6032 , \6030 , \6031 );
or \mul_7_15_g33856/U$5 ( \6033 , \5997 , \5975 );
nand \mul_7_15_g33856/U$1 ( \6034 , \6032 , \6033 );
not \mul_7_15_g33915/U$1 ( \6035 , \5973 );
and \mul_7_15_g33792/U$2 ( \6036 , \6034 , \6035 );
not \mul_7_15_g33792/U$4 ( \6037 , \6034 );
and \mul_7_15_g33792/U$3 ( \6038 , \6037 , \5973 );
nor \mul_7_15_g33792/U$1 ( \6039 , \6036 , \6038 );
or \mul_7_15_g35280/U$1 ( \6040 , \6029 , \6039 );
xor \mul_7_15_g33914/U$1 ( \6041 , \5761 , \5776 );
xor \mul_7_15_g33914/U$1_r1 ( \6042 , \6041 , \5792 );
not \mul_7_15_g35304/U$2 ( \6043 , \6042 );
and \mul_7_15_g34040/U$2 ( \6044 , \5995 , \5987 );
not \mul_7_15_g34040/U$4 ( \6045 , \5995 );
not \mul_7_15_g34266/U$1 ( \6046 , \5987 );
and \mul_7_15_g34040/U$3 ( \6047 , \6045 , \6046 );
nor \mul_7_15_g34040/U$1 ( \6048 , \6044 , \6047 );
not \mul_7_15_g34146/U$1 ( \6049 , \5981 );
and \mul_7_15_g33981/U$2 ( \6050 , \6048 , \6049 );
not \mul_7_15_g33981/U$4 ( \6051 , \6048 );
and \mul_7_15_g33981/U$3 ( \6052 , \6051 , \5981 );
nor \mul_7_15_g33981/U$1 ( \6053 , \6050 , \6052 );
buf \mul_7_15_g33909/U$1 ( \6054 , \6053 );
nand \mul_7_15_g35304/U$1 ( \6055 , \6043 , \6054 );
not \mul_7_15_g33666/U$3 ( \6056 , \6055 );
and \mul_7_15_g34706/U$2 ( \6057 , \4029 , \4177 );
not \mul_7_15_g34706/U$4 ( \6058 , \4029 );
and \mul_7_15_g34706/U$3 ( \6059 , \6058 , \4176 );
nor \mul_7_15_g34706/U$1 ( \6060 , \6057 , \6059 );
not \mul_7_15_g34119/U$3 ( \6061 , \6060 );
not \mul_7_15_g34119/U$4 ( \6062 , \4195 );
or \mul_7_15_g34119/U$2 ( \6063 , \6061 , \6062 );
nand \mul_7_15_g34369/U$1 ( \6064 , \5111 , \5782 );
nand \mul_7_15_g34119/U$1 ( \6065 , \6063 , \6064 );
not \mul_7_15_g34564/U$3 ( \6066 , \5388 );
not \mul_7_15_g34564/U$4 ( \6067 , \4190 );
or \mul_7_15_g34564/U$2 ( \6068 , \6066 , \6067 );
nand \mul_7_15_g34564/U$1 ( \6069 , \6068 , \4368 );
nand \mul_7_15_g34811/U$1 ( \6070 , \3487 , \4048 );
and \mul_7_15_g34538/U$1 ( \6071 , \6069 , \4172 , \6070 );
not \mul_7_15_g34715/U$3 ( \6072 , \4011 );
not \mul_7_15_g34715/U$4 ( \6073 , \5178 );
or \mul_7_15_g34715/U$2 ( \6074 , \6072 , \6073 );
nand \mul_7_15_g34918/U$1 ( \6075 , \4665 , \4270 );
nand \mul_7_15_g34715/U$1 ( \6076 , \6074 , \6075 );
not \mul_7_15_g34242/U$3 ( \6077 , \6076 );
not \mul_7_15_g34242/U$4 ( \6078 , \4662 );
or \mul_7_15_g34242/U$2 ( \6079 , \6077 , \6078 );
nand \mul_7_15_g34380/U$1 ( \6080 , \4672 , \5855 );
nand \mul_7_15_g34242/U$1 ( \6081 , \6079 , \6080 );
and \mul_7_15_g34011/U$2 ( \6082 , \6071 , \6081 );
xor \mul_7_15_g33757/U$4 ( \6083 , \6065 , \6082 );
and \mul_7_15_g34799/U$2 ( \6084 , \4238 , \5873 );
not \mul_7_15_g34799/U$4 ( \6085 , \4238 );
and \mul_7_15_g34799/U$3 ( \6086 , \6085 , \5874 );
nor \mul_7_15_g34799/U$1 ( \6087 , \6084 , \6086 );
not \mul_7_15_g34798/U$1 ( \6088 , \6087 );
not \mul_7_15_g34329/U$3 ( \6089 , \6088 );
not \mul_7_15_g34329/U$4 ( \6090 , \5019 );
or \mul_7_15_g34329/U$2 ( \6091 , \6089 , \6090 );
nand \mul_7_15_g34441/U$1 ( \6092 , \5878 , \5021 );
nand \mul_7_15_g34329/U$1 ( \6093 , \6091 , \6092 );
and \mul_7_15_g34775/U$2 ( \6094 , \5344 , \4142 );
not \mul_7_15_g34775/U$4 ( \6095 , \5344 );
and \mul_7_15_g34775/U$3 ( \6096 , \6095 , \4109 );
nor \mul_7_15_g34775/U$1 ( \6097 , \6094 , \6096 );
not \mul_7_15_g34270/U$3 ( \6098 , \6097 );
not \mul_7_15_g34270/U$4 ( \6099 , \4425 );
or \mul_7_15_g34270/U$2 ( \6100 , \6098 , \6099 );
nand \mul_7_15_g34457/U$1 ( \6101 , \4429 , \5889 );
nand \mul_7_15_g34270/U$1 ( \6102 , \6100 , \6101 );
xor \mul_7_15_g33895/U$4 ( \6103 , \6093 , \6102 );
and \mul_7_15_g34722/U$2 ( \6104 , \4019 , \4088 );
not \mul_7_15_g34722/U$4 ( \6105 , \4019 );
and \mul_7_15_g34722/U$3 ( \6106 , \6105 , \5234 );
nor \mul_7_15_g34722/U$1 ( \6107 , \6104 , \6106 );
not \mul_7_15_g34151/U$3 ( \6108 , \6107 );
not \mul_7_15_g34151/U$4 ( \6109 , \4437 );
or \mul_7_15_g34151/U$2 ( \6110 , \6108 , \6109 );
nand \mul_7_15_g34357/U$1 ( \6111 , \4331 , \5839 );
nand \mul_7_15_g34151/U$1 ( \6112 , \6110 , \6111 );
and \mul_7_15_g33895/U$3 ( \6113 , \6103 , \6112 );
and \mul_7_15_g33895/U$5 ( \6114 , \6093 , \6102 );
or \mul_7_15_g33895/U$2 ( \6115 , \6113 , \6114 );
and \mul_7_15_g33757/U$3 ( \6116 , \6083 , \6115 );
and \mul_7_15_g33757/U$5 ( \6117 , \6065 , \6082 );
or \mul_7_15_g33757/U$2 ( \6118 , \6116 , \6117 );
not \mul_7_15_g33666/U$4 ( \6119 , \6118 );
or \mul_7_15_g33666/U$2 ( \6120 , \6056 , \6119 );
not \mul_7_15_g35303/U$2 ( \6121 , \6054 );
nand \mul_7_15_g35303/U$1 ( \6122 , \6121 , \6042 );
nand \mul_7_15_g33666/U$1 ( \6123 , \6120 , \6122 );
and \mul_7_15_g33487/U$2 ( \6124 , \6040 , \6123 );
and \mul_7_15_g33544/U$2 ( \6125 , \6039 , \6029 );
nor \mul_7_15_g33487/U$1 ( \6126 , \6124 , \6125 );
nand \mul_7_15_g33451/U$1 ( \6127 , \6023 , \6126 );
xor \mul_7_15_g33544/U$1 ( \6128 , \6039 , \6029 );
not \mul_7_15_g33651/U$1 ( \6129 , \6123 );
and \mul_7_15_g33497/U$2 ( \6130 , \6128 , \6129 );
not \mul_7_15_g33497/U$4 ( \6131 , \6128 );
and \mul_7_15_g33497/U$3 ( \6132 , \6131 , \6123 );
nor \mul_7_15_g33497/U$1 ( \6133 , \6130 , \6132 );
xor \mul_7_15_g33703/U$1 ( \6134 , \5833 , \5870 );
xor \mul_7_15_g33703/U$1_r1 ( \6135 , \6134 , \5915 );
not \mul_7_15_g33610/U$2 ( \6136 , \6135 );
not \mul_7_15_g33857/U$3 ( \6137 , \6042 );
not \mul_7_15_g33857/U$4 ( \6138 , \6053 );
or \mul_7_15_g33857/U$2 ( \6139 , \6137 , \6138 );
or \mul_7_15_g33857/U$5 ( \6140 , \6053 , \6042 );
nand \mul_7_15_g33857/U$1 ( \6141 , \6139 , \6140 );
not \mul_7_15_g33756/U$1 ( \6142 , \6118 );
and \mul_7_15_g33687/U$2 ( \6143 , \6141 , \6142 );
not \mul_7_15_g33687/U$4 ( \6144 , \6141 );
and \mul_7_15_g33687/U$3 ( \6145 , \6144 , \6118 );
nor \mul_7_15_g33687/U$1 ( \6146 , \6143 , \6145 );
nand \mul_7_15_g33610/U$1 ( \6147 , \6136 , \6146 );
xor \mul_7_15_g33970/U$1 ( \6148 , \5867 , \5849 );
xor \mul_7_15_g33970/U$1_r1 ( \6149 , \6148 , \5865 );
not \mul_7_15_g33738/U$3 ( \6150 , \6149 );
xor \mul_7_15_g33954/U$1 ( \6151 , \5883 , \5899 );
xnor \mul_7_15_g33954/U$1_r1 ( \6152 , \6151 , \5913 );
not \mul_7_15_g33738/U$4 ( \6153 , \6152 );
or \mul_7_15_g33738/U$2 ( \6154 , \6150 , \6153 );
not \mul_7_15_g34773/U$3 ( \6155 , \3958 );
not \mul_7_15_g34773/U$4 ( \6156 , \4069 );
or \mul_7_15_g34773/U$2 ( \6157 , \6155 , \6156 );
not \mul_7_15_g35347/U$2 ( \6158 , \5904 );
nand \mul_7_15_g35347/U$1 ( \6159 , \6158 , \4473 );
nand \mul_7_15_g34773/U$1 ( \6160 , \6157 , \6159 );
not \mul_7_15_g34194/U$3 ( \6161 , \6160 );
not \fopt35521/U$1 ( \6162 , \4411 );
not \mul_7_15_g34194/U$4 ( \6163 , \6162 );
or \mul_7_15_g34194/U$2 ( \6164 , \6161 , \6163 );
nand \mul_7_15_g34379/U$1 ( \6165 , \4562 , \5908 );
nand \mul_7_15_g34194/U$1 ( \6166 , \6164 , \6165 );
not \mul_7_15_g34064/U$2 ( \6167 , \6166 );
and \mul_7_15_g34806/U$2 ( \6168 , \4048 , \4177 );
not \mul_7_15_g34806/U$4 ( \6169 , \4048 );
and \mul_7_15_g34806/U$3 ( \6170 , \6169 , \4284 );
nor \mul_7_15_g34806/U$1 ( \6171 , \6168 , \6170 );
not \mul_7_15_g34126/U$3 ( \6172 , \6171 );
not \mul_7_15_g34126/U$4 ( \6173 , \4194 );
or \mul_7_15_g34126/U$2 ( \6174 , \6172 , \6173 );
nand \mul_7_15_g34390/U$1 ( \6175 , \6060 , \5111 );
nand \mul_7_15_g34126/U$1 ( \6176 , \6174 , \6175 );
not \mul_7_15_g34125/U$1 ( \6177 , \6176 );
nand \mul_7_15_g34064/U$1 ( \6178 , \6167 , \6177 );
not \mul_7_15_g33898/U$3 ( \6179 , \6178 );
xor \mul_7_15_g34011/U$1 ( \6180 , \6071 , \6081 );
not \mul_7_15_g33898/U$4 ( \6181 , \6180 );
or \mul_7_15_g33898/U$2 ( \6182 , \6179 , \6181 );
nand \mul_7_15_g34065/U$1 ( \6183 , \6166 , \6176 );
nand \mul_7_15_g33898/U$1 ( \6184 , \6182 , \6183 );
nand \mul_7_15_g33738/U$1 ( \6185 , \6154 , \6184 );
not \mul_7_15_g33885/U$1 ( \6186 , \6152 );
not \mul_7_15_g33927/U$1 ( \6187 , \6149 );
nand \mul_7_15_g33838/U$1 ( \6188 , \6186 , \6187 );
nand \mul_7_15_g33696/U$1 ( \6189 , \6185 , \6188 );
not \mul_7_15_g33678/U$1 ( \6190 , \6189 );
not \mul_7_15_g33677/U$1 ( \6191 , \6190 );
and \mul_7_15_g33567/U$2 ( \6192 , \6147 , \6191 );
not \mul_7_15_g35287/U$2 ( \6193 , \6135 );
nor \mul_7_15_g35287/U$1 ( \6194 , \6193 , \6146 );
nor \mul_7_15_g33567/U$1 ( \6195 , \6192 , \6194 );
nand \mul_7_15_g33449/U$1 ( \6196 , \6133 , \6195 );
nand \mul_7_15_g33422/U$1 ( \6197 , \6127 , \6196 );
not \mul_7_15_g35272/U$2 ( \6198 , \6197 );
xor \mul_7_15_g35350/U$1 ( \6199 , \6166 , \6176 );
xor \mul_7_15_g35350/U$1_r1 ( \6200 , \6199 , \6180 );
not \mul_7_15_g35167/U$1 ( \6201 , \4128 );
nor \mul_7_15_g34814/U$1 ( \6202 , \6201 , \4048 );
not \mul_7_15_g34541/U$3 ( \6203 , \6202 );
not \mul_7_15_g34541/U$4 ( \6204 , \4089 );
and \mul_7_15_g34541/U$2 ( \6205 , \6203 , \6204 );
not \mul_7_15_g34567/U$3 ( \6206 , \4048 );
not \mul_7_15_g34567/U$4 ( \6207 , \6201 );
or \mul_7_15_g34567/U$2 ( \6208 , \6206 , \6207 );
nand \mul_7_15_g34567/U$1 ( \6209 , \6208 , \4109 );
nor \mul_7_15_g34541/U$1 ( \6210 , \6205 , \6209 );
and \mul_7_15_g34741/U$2 ( \6211 , \4473 , \5178 );
not \mul_7_15_g34741/U$4 ( \6212 , \4473 );
and \mul_7_15_g34741/U$3 ( \6213 , \6212 , \4665 );
nor \mul_7_15_g34741/U$1 ( \6214 , \6211 , \6213 );
nand \mul_7_15_g34353/U$1 ( \6215 , \4541 , \6214 );
or \mul_7_15_g34105/U$2 ( \6216 , \6215 , \5187 );
not \mul_7_15_g34753/U$3 ( \6217 , \4046 );
not \mul_7_15_g34753/U$4 ( \6218 , \5178 );
or \mul_7_15_g34753/U$2 ( \6219 , \6217 , \6218 );
nand \mul_7_15_g35809/U$1 ( \6220 , \4665 , \4256 );
nand \mul_7_15_g34753/U$1 ( \6221 , \6219 , \6220 );
nand \mul_7_15_g34367/U$1 ( \6222 , \5187 , \6221 );
nand \mul_7_15_g34105/U$1 ( \6223 , \6216 , \6222 );
and \mul_7_15_g34013/U$2 ( \6224 , \6210 , \6223 );
not \mul_7_15_g34334/U$3 ( \6225 , \5390 );
not \mul_7_15_g34792/U$3 ( \6226 , \4011 );
not \mul_7_15_g35055/U$1 ( \6227 , \5273 );
not \mul_7_15_g34792/U$4 ( \6228 , \6227 );
or \mul_7_15_g34792/U$2 ( \6229 , \6226 , \6228 );
nand \mul_7_15_g34881/U$1 ( \6230 , \5873 , \4270 );
nand \mul_7_15_g34792/U$1 ( \6231 , \6229 , \6230 );
not \mul_7_15_g34334/U$4 ( \6232 , \6231 );
or \mul_7_15_g34334/U$2 ( \6233 , \6225 , \6232 );
not \mul_7_15_g34795/U$3 ( \6234 , \4043 );
not \mul_7_15_g34795/U$4 ( \6235 , \5576 );
or \mul_7_15_g34795/U$2 ( \6236 , \6234 , \6235 );
nand \mul_7_15_g34859/U$1 ( \6237 , \4217 , \5873 );
nand \mul_7_15_g34795/U$1 ( \6238 , \6236 , \6237 );
nand \mul_7_15_g34381/U$1 ( \6239 , \6238 , \5021 );
nand \mul_7_15_g34334/U$1 ( \6240 , \6233 , \6239 );
and \mul_7_15_g34682/U$2 ( \6241 , \4114 , \4029 );
and \mul_7_15_g34682/U$3 ( \6242 , \4109 , \5339 );
nor \mul_7_15_g34682/U$1 ( \6243 , \6241 , \6242 );
not \mul_7_15_g34605/U$1 ( \6244 , \4139 );
or \mul_7_15_g34106/U$2 ( \6245 , \6243 , \6244 );
not \mul_7_15_g34603/U$1 ( \6246 , \4139 );
and \mul_7_15_g34805/U$2 ( \6247 , \4048 , \4146 );
not \mul_7_15_g34805/U$4 ( \6248 , \4048 );
and \mul_7_15_g34805/U$3 ( \6249 , \6248 , \4145 );
nor \mul_7_15_g34805/U$1 ( \6250 , \6247 , \6249 );
nand \mul_7_15_g34307/U$1 ( \6251 , \6246 , \6250 , \4134 );
nand \mul_7_15_g34106/U$1 ( \6252 , \6245 , \6251 );
xor \mul_7_15_g33891/U$4 ( \6253 , \6240 , \6252 );
not \mul_7_15_g34690/U$3 ( \6254 , \4026 );
not \mul_7_15_g34690/U$4 ( \6255 , \4089 );
or \mul_7_15_g34690/U$2 ( \6256 , \6254 , \6255 );
nand \mul_7_15_g34888/U$1 ( \6257 , \4088 , \5344 );
nand \mul_7_15_g34690/U$1 ( \6258 , \6256 , \6257 );
not \mul_7_15_g34153/U$3 ( \6259 , \6258 );
not \mul_7_15_g34153/U$4 ( \6260 , \4437 );
or \mul_7_15_g34153/U$2 ( \6261 , \6259 , \6260 );
not \mul_7_15_g34724/U$3 ( \6262 , \4023 );
not \mul_7_15_g34724/U$4 ( \6263 , \5234 );
or \mul_7_15_g34724/U$2 ( \6264 , \6262 , \6263 );
nand \mul_7_15_g34892/U$1 ( \6265 , \4088 , \5131 );
nand \mul_7_15_g34724/U$1 ( \6266 , \6264 , \6265 );
nand \mul_7_15_g34349/U$1 ( \6267 , \4331 , \6266 );
nand \mul_7_15_g34153/U$1 ( \6268 , \6261 , \6267 );
and \mul_7_15_g33891/U$3 ( \6269 , \6253 , \6268 );
and \mul_7_15_g33891/U$5 ( \6270 , \6240 , \6252 );
or \mul_7_15_g33891/U$2 ( \6271 , \6269 , \6270 );
xor \mul_7_15_g33715/U$4 ( \6272 , \6224 , \6271 );
and \mul_7_15_g34521/U$1 ( \6273 , \5816 , \4048 );
not \mul_7_15_g34152/U$3 ( \6274 , \6266 );
not \mul_7_15_g34152/U$4 ( \6275 , \4437 );
or \mul_7_15_g34152/U$2 ( \6276 , \6274 , \6275 );
nand \mul_7_15_g34500/U$1 ( \6277 , \4331 , \6107 );
nand \mul_7_15_g34152/U$1 ( \6278 , \6276 , \6277 );
xor \mul_7_15_g33936/U$1 ( \6279 , \6273 , \6278 );
not \mul_7_15_g34235/U$3 ( \6280 , \6221 );
not \mul_7_15_g34235/U$4 ( \6281 , \4662 );
or \mul_7_15_g34235/U$2 ( \6282 , \6280 , \6281 );
nand \mul_7_15_g34356/U$1 ( \6283 , \4672 , \6076 );
nand \mul_7_15_g34235/U$1 ( \6284 , \6282 , \6283 );
xor \mul_7_15_g33936/U$1_r1 ( \6285 , \6279 , \6284 );
and \mul_7_15_g33715/U$3 ( \6286 , \6272 , \6285 );
and \mul_7_15_g33715/U$5 ( \6287 , \6224 , \6271 );
or \mul_7_15_g33715/U$2 ( \6288 , \6286 , \6287 );
xor \mul_7_15_g33601/U$1 ( \6289 , \6200 , \6288 );
not \mul_7_15_g34333/U$3 ( \6290 , \6087 );
not \mul_7_15_g34333/U$4 ( \6291 , \5265 );
and \mul_7_15_g34333/U$2 ( \6292 , \6290 , \6291 );
and \mul_7_15_g34333/U$5 ( \6293 , \5019 , \6238 );
nor \mul_7_15_g34333/U$1 ( \6294 , \6292 , \6293 );
not \mul_7_15_g34332/U$1 ( \6295 , \6294 );
not \mul_7_15_g33897/U$3 ( \6296 , \6295 );
not \mul_7_15_g34104/U$3 ( \6297 , \6244 );
not \mul_7_15_g34462/U$2 ( \6298 , \4134 );
nor \mul_7_15_g34462/U$1 ( \6299 , \6298 , \6243 );
not \mul_7_15_g34104/U$4 ( \6300 , \6299 );
or \mul_7_15_g34104/U$2 ( \6301 , \6297 , \6300 );
nand \mul_7_15_g34351/U$1 ( \6302 , \4139 , \6097 );
nand \mul_7_15_g34104/U$1 ( \6303 , \6301 , \6302 );
not \mul_7_15_g33897/U$4 ( \6304 , \6303 );
or \mul_7_15_g33897/U$2 ( \6305 , \6296 , \6304 );
or \mul_7_15_g33957/U$2 ( \6306 , \6303 , \6295 );
not \mul_7_15_g34726/U$3 ( \6307 , \3963 );
not \mul_7_15_g34726/U$4 ( \6308 , \5904 );
or \mul_7_15_g34726/U$2 ( \6309 , \6307 , \6308 );
nand \mul_7_15_g34916/U$1 ( \6310 , \4403 , \4486 );
nand \mul_7_15_g34726/U$1 ( \6311 , \6309 , \6310 );
not \mul_7_15_g34212/U$3 ( \6312 , \6311 );
not \mul_7_15_g34212/U$4 ( \6313 , \6162 );
or \mul_7_15_g34212/U$2 ( \6314 , \6312 , \6313 );
nand \mul_7_15_g34484/U$1 ( \6315 , \4055 , \6160 );
nand \mul_7_15_g34212/U$1 ( \6316 , \6314 , \6315 );
nand \mul_7_15_g33957/U$1 ( \6317 , \6306 , \6316 );
nand \mul_7_15_g33897/U$1 ( \6318 , \6305 , \6317 );
xor \mul_7_15_g33936/U$4 ( \6319 , \6273 , \6278 );
and \mul_7_15_g33936/U$3 ( \6320 , \6319 , \6284 );
and \mul_7_15_g33936/U$5 ( \6321 , \6273 , \6278 );
or \mul_7_15_g33936/U$2 ( \6322 , \6320 , \6321 );
xor \mul_7_15_g33711/U$1 ( \6323 , \6318 , \6322 );
xor \mul_7_15_g33895/U$1 ( \6324 , \6093 , \6102 );
xor \mul_7_15_g33895/U$1_r1 ( \6325 , \6324 , \6112 );
xor \mul_7_15_g33711/U$1_r1 ( \6326 , \6323 , \6325 );
xnor \mul_7_15_g33601/U$1_r1 ( \6327 , \6289 , \6326 );
xor \mul_7_15_g33715/U$1 ( \6328 , \6224 , \6271 );
xor \mul_7_15_g33715/U$1_r1 ( \6329 , \6328 , \6285 );
not \mul_7_15_g33712/U$1 ( \6330 , \6329 );
not \mul_7_15_g33615/U$3 ( \6331 , \6330 );
not \mul_7_15_g34729/U$3 ( \6332 , \4019 );
not \mul_7_15_g34729/U$4 ( \6333 , \4069 );
or \mul_7_15_g34729/U$2 ( \6334 , \6332 , \6333 );
nand \mul_7_15_g34874/U$1 ( \6335 , \4403 , \4585 );
nand \mul_7_15_g34729/U$1 ( \6336 , \6334 , \6335 );
not \mul_7_15_g34163/U$3 ( \6337 , \6336 );
not \mul_7_15_g34163/U$4 ( \6338 , \5361 );
or \mul_7_15_g34163/U$2 ( \6339 , \6337 , \6338 );
nand \mul_7_15_g34342/U$1 ( \6340 , \4055 , \6311 );
nand \mul_7_15_g34163/U$1 ( \6341 , \6339 , \6340 );
xor \mul_7_15_g34013/U$1 ( \6342 , \6210 , \6223 );
xor \mul_7_15_g33788/U$4 ( \6343 , \6341 , \6342 );
not \mul_7_15_g34514/U$2 ( \6344 , \6246 );
nand \mul_7_15_g34514/U$1 ( \6345 , \6344 , \4048 );
not \mul_7_15_g34318/U$3 ( \6346 , \5390 );
not \mul_7_15_g34802/U$3 ( \6347 , \4046 );
not \mul_7_15_g34802/U$4 ( \6348 , \6227 );
or \mul_7_15_g34802/U$2 ( \6349 , \6347 , \6348 );
not \mul_7_15_g35338/U$2 ( \6350 , \5270 );
nand \mul_7_15_g35338/U$1 ( \6351 , \6350 , \4256 );
nand \mul_7_15_g34802/U$1 ( \6352 , \6349 , \6351 );
not \mul_7_15_g34318/U$4 ( \6353 , \6352 );
or \mul_7_15_g34318/U$2 ( \6354 , \6346 , \6353 );
nand \mul_7_15_g34362/U$1 ( \6355 , \6231 , \5021 );
nand \mul_7_15_g34318/U$1 ( \6356 , \6354 , \6355 );
not \mul_7_15_g34317/U$1 ( \6357 , \6356 );
nand \mul_7_15_g34092/U$1 ( \6358 , \6345 , \6357 );
not \mul_7_15_g33964/U$3 ( \6359 , \6358 );
not \mul_7_15_g34770/U$3 ( \6360 , \4029 );
not \mul_7_15_g34770/U$4 ( \6361 , \5234 );
or \mul_7_15_g34770/U$2 ( \6362 , \6360 , \6361 );
nand \mul_7_15_g34879/U$1 ( \6363 , \4088 , \5339 );
nand \mul_7_15_g34770/U$1 ( \6364 , \6362 , \6363 );
not \mul_7_15_g34138/U$3 ( \6365 , \6364 );
not \mul_7_15_g34138/U$4 ( \6366 , \4085 );
or \mul_7_15_g34138/U$2 ( \6367 , \6365 , \6366 );
nand \mul_7_15_g34378/U$1 ( \6368 , \4331 , \6258 );
nand \mul_7_15_g34138/U$1 ( \6369 , \6367 , \6368 );
not \mul_7_15_g33964/U$4 ( \6370 , \6369 );
or \mul_7_15_g33964/U$2 ( \6371 , \6359 , \6370 );
not \mul_7_15_g34513/U$1 ( \6372 , \6345 );
nand \mul_7_15_g34094/U$1 ( \6373 , \6372 , \6356 );
nand \mul_7_15_g33964/U$1 ( \6374 , \6371 , \6373 );
and \mul_7_15_g33788/U$3 ( \6375 , \6343 , \6374 );
and \mul_7_15_g33788/U$5 ( \6376 , \6341 , \6342 );
or \mul_7_15_g33788/U$2 ( \6377 , \6375 , \6376 );
buf \mul_7_15_g33787/U$1 ( \6378 , \6377 );
xnor \g35401/U$1 ( \6379 , \6294 , \6303 );
xnor \mul_7_15_g35315/U$1 ( \6380 , \6379 , \6316 );
not \mul_7_15_g33888/U$1 ( \6381 , \6380 );
nor \mul_7_15_g33732/U$1 ( \6382 , \6378 , \6381 );
not \mul_7_15_g33615/U$4 ( \6383 , \6382 );
and \mul_7_15_g33615/U$2 ( \6384 , \6331 , \6383 );
and \mul_7_15_g33615/U$5 ( \6385 , \6378 , \6381 );
nor \mul_7_15_g33615/U$1 ( \6386 , \6384 , \6385 );
nand \mul_7_15_g33519/U$1 ( \6387 , \6327 , \6386 );
xor \mul_7_15_g33891/U$1 ( \6388 , \6240 , \6252 );
xor \mul_7_15_g33891/U$1_r1 ( \6389 , \6388 , \6268 );
not \mul_7_15_g34743/U$3 ( \6390 , \4023 );
not \mul_7_15_g34743/U$4 ( \6391 , \4069 );
or \mul_7_15_g34743/U$2 ( \6392 , \6390 , \6391 );
nand \mul_7_15_g34894/U$1 ( \6393 , \4407 , \5131 );
nand \mul_7_15_g34743/U$1 ( \6394 , \6392 , \6393 );
not \mul_7_15_g34173/U$3 ( \6395 , \6394 );
not \mul_7_15_g34173/U$4 ( \6396 , \4065 );
or \mul_7_15_g34173/U$2 ( \6397 , \6395 , \6396 );
nand \mul_7_15_g34360/U$1 ( \6398 , \4055 , \6336 );
nand \mul_7_15_g34173/U$1 ( \6399 , \6397 , \6398 );
not \g3/U$2 ( \6400 , \6399 );
not \mul_7_15_g34338/U$3 ( \6401 , \5019 );
not \mul_7_15_g34801/U$3 ( \6402 , \3958 );
not \mul_7_15_g34801/U$4 ( \6403 , \5874 );
or \mul_7_15_g34801/U$2 ( \6404 , \6402 , \6403 );
nand \mul_7_15_g34872/U$1 ( \6405 , \5873 , \4473 );
nand \mul_7_15_g34801/U$1 ( \6406 , \6404 , \6405 );
not \mul_7_15_g34338/U$4 ( \6407 , \6406 );
or \mul_7_15_g34338/U$2 ( \6408 , \6401 , \6407 );
nand \mul_7_15_g34430/U$1 ( \6409 , \6352 , \5021 );
nand \mul_7_15_g34338/U$1 ( \6410 , \6408 , \6409 );
nand \mul_7_15_g34812/U$1 ( \6411 , \4076 , \5388 );
and \mul_7_15_g34533/U$2 ( \6412 , \5749 , \6411 );
not \mul_7_15_g34565/U$3 ( \6413 , \4048 );
not \mul_7_15_g34565/U$4 ( \6414 , \3272 );
or \mul_7_15_g34565/U$2 ( \6415 , \6413 , \6414 );
nand \mul_7_15_g34565/U$1 ( \6416 , \6415 , \4088 );
nor \mul_7_15_g34533/U$1 ( \6417 , \6412 , \6416 );
nand \mul_7_15_g34098/U$1 ( \6418 , \6410 , \6417 );
nand \g3/U$1 ( \6419 , \6400 , \6418 );
not \g2/U$3 ( \6420 , \6419 );
not \mul_7_15_g34237/U$3 ( \6421 , \4662 );
not \mul_7_15_g34691/U$3 ( \6422 , \3963 );
not \mul_7_15_g34691/U$4 ( \6423 , \4666 );
or \mul_7_15_g34691/U$2 ( \6424 , \6422 , \6423 );
nand \mul_7_15_g34857/U$1 ( \6425 , \4665 , \4486 );
nand \mul_7_15_g34691/U$1 ( \6426 , \6424 , \6425 );
not \mul_7_15_g34237/U$4 ( \6427 , \6426 );
or \mul_7_15_g34237/U$2 ( \6428 , \6421 , \6427 );
nand \mul_7_15_g34388/U$1 ( \6429 , \5187 , \6214 );
nand \mul_7_15_g34237/U$1 ( \6430 , \6428 , \6429 );
not \g2/U$4 ( \6431 , \6430 );
or \g2/U$2 ( \6432 , \6420 , \6431 );
not \mul_7_15_g35309/U$2 ( \6433 , \6418 );
nand \mul_7_15_g35309/U$1 ( \6434 , \6433 , \6399 );
nand \g2/U$1 ( \6435 , \6432 , \6434 );
xor \g35393/U$1 ( \6436 , \6389 , \6435 );
xor \mul_7_15_g33788/U$1 ( \6437 , \6341 , \6342 );
xor \mul_7_15_g33788/U$1_r1 ( \6438 , \6437 , \6374 );
and \mul_7_15_g33685/U$2 ( \6439 , \6436 , \6438 );
not \mul_7_15_g33685/U$4 ( \6440 , \6436 );
not \mul_7_15_g33785/U$1 ( \6441 , \6438 );
and \mul_7_15_g33685/U$3 ( \6442 , \6440 , \6441 );
nor \mul_7_15_g33685/U$1 ( \6443 , \6439 , \6442 );
not \mul_7_15_g34081/U$3 ( \6444 , \6357 );
not \mul_7_15_g34512/U$1 ( \6445 , \6345 );
not \mul_7_15_g34081/U$4 ( \6446 , \6445 );
or \mul_7_15_g34081/U$2 ( \6447 , \6444 , \6446 );
or \mul_7_15_g34081/U$5 ( \6448 , \6372 , \6357 );
nand \mul_7_15_g34081/U$1 ( \6449 , \6447 , \6448 );
xor \mul_7_15_g33969/U$1 ( \6450 , \6449 , \6369 );
not \mul_7_15_g34808/U$3 ( \6451 , \5388 );
not \mul_7_15_g34808/U$4 ( \6452 , \4088 );
or \mul_7_15_g34808/U$2 ( \6453 , \6451 , \6452 );
nand \mul_7_15_g34946/U$1 ( \6454 , \4089 , \4048 );
nand \mul_7_15_g34808/U$1 ( \6455 , \6453 , \6454 );
and \mul_7_15_g34160/U$2 ( \6456 , \4086 , \6455 );
not \fopt35517/U$1 ( \6457 , \5241 );
and \mul_7_15_g34160/U$3 ( \6458 , \6457 , \6364 );
nor \mul_7_15_g34160/U$1 ( \6459 , \6456 , \6458 );
not \mul_7_15_g34159/U$1 ( \6460 , \6459 );
not \mul_7_15_g34005/U$3 ( \6461 , \6460 );
not \mul_7_15_g34782/U$3 ( \6462 , \4026 );
not \mul_7_15_g34782/U$4 ( \6463 , \4069 );
or \mul_7_15_g34782/U$2 ( \6464 , \6462 , \6463 );
nand \mul_7_15_g34926/U$1 ( \6465 , \5749 , \5344 );
nand \mul_7_15_g34782/U$1 ( \6466 , \6464 , \6465 );
and \mul_7_15_g34223/U$2 ( \6467 , \6466 , \4065 );
and \mul_7_15_g34223/U$3 ( \6468 , \4562 , \6394 );
nor \mul_7_15_g34223/U$1 ( \6469 , \6467 , \6468 );
not \mul_7_15_g34222/U$1 ( \6470 , \6469 );
not \mul_7_15_g34005/U$4 ( \6471 , \6470 );
or \mul_7_15_g34005/U$2 ( \6472 , \6461 , \6471 );
not \mul_7_15_g34018/U$3 ( \6473 , \6459 );
not \mul_7_15_g34018/U$4 ( \6474 , \6469 );
or \mul_7_15_g34018/U$2 ( \6475 , \6473 , \6474 );
not \mul_7_15_g34683/U$3 ( \6476 , \4019 );
not \mul_7_15_g34683/U$4 ( \6477 , \5178 );
or \mul_7_15_g34683/U$2 ( \6478 , \6476 , \6477 );
nand \mul_7_15_g34920/U$1 ( \6479 , \4665 , \4585 );
nand \mul_7_15_g34683/U$1 ( \6480 , \6478 , \6479 );
not \mul_7_15_g34230/U$3 ( \6481 , \6480 );
not \mul_7_15_g34230/U$4 ( \6482 , \4662 );
or \mul_7_15_g34230/U$2 ( \6483 , \6481 , \6482 );
nand \mul_7_15_g34498/U$1 ( \6484 , \5187 , \6426 );
nand \mul_7_15_g34230/U$1 ( \6485 , \6483 , \6484 );
nand \mul_7_15_g34018/U$1 ( \6486 , \6475 , \6485 );
nand \mul_7_15_g34005/U$1 ( \6487 , \6472 , \6486 );
xor \mul_7_15_g33684/U$4 ( \6488 , \6450 , \6487 );
xor \mul_7_15_g35316/U$1 ( \6489 , \6418 , \6399 );
xnor \mul_7_15_g35316/U$1_r1 ( \6490 , \6489 , \6430 );
and \mul_7_15_g33684/U$3 ( \6491 , \6488 , \6490 );
and \mul_7_15_g33684/U$5 ( \6492 , \6450 , \6487 );
or \mul_7_15_g33684/U$2 ( \6493 , \6491 , \6492 );
nand \mul_7_15_g33605/U$1 ( \6494 , \6443 , \6493 );
not \g35883/U$3 ( \6495 , \6494 );
xor \mul_7_15_g33684/U$1 ( \6496 , \6450 , \6487 );
xor \mul_7_15_g33684/U$1_r1 ( \6497 , \6496 , \6490 );
nor \mul_7_15_g34518/U$1 ( \6498 , \4103 , \5388 );
not \mul_7_15_g34790/U$3 ( \6499 , \3963 );
not \mul_7_15_g34790/U$4 ( \6500 , \5023 );
or \mul_7_15_g34790/U$2 ( \6501 , \6499 , \6500 );
not \mul_7_15_g35043/U$1 ( \6502 , \5576 );
nand \mul_7_15_g34880/U$1 ( \6503 , \6502 , \4486 );
nand \mul_7_15_g34790/U$1 ( \6504 , \6501 , \6503 );
not \mul_7_15_g34324/U$3 ( \6505 , \6504 );
not \mul_7_15_g34324/U$4 ( \6506 , \5020 );
or \mul_7_15_g34324/U$2 ( \6507 , \6505 , \6506 );
nand \mul_7_15_g34421/U$1 ( \6508 , \6406 , \5021 );
nand \mul_7_15_g34324/U$1 ( \6509 , \6507 , \6508 );
xor \mul_7_15_g33943/U$4 ( \6510 , \6498 , \6509 );
not \mul_7_15_g34228/U$3 ( \6511 , \4662 );
not \mul_7_15_g34754/U$3 ( \6512 , \4023 );
not \mul_7_15_g34754/U$4 ( \6513 , \4666 );
or \mul_7_15_g34754/U$2 ( \6514 , \6512 , \6513 );
not \mul_7_15_g35344/U$2 ( \6515 , \5178 );
nand \mul_7_15_g35344/U$1 ( \6516 , \6515 , \5131 );
nand \mul_7_15_g34754/U$1 ( \6517 , \6514 , \6516 );
not \mul_7_15_g34228/U$4 ( \6518 , \6517 );
or \mul_7_15_g34228/U$2 ( \6519 , \6511 , \6518 );
nand \mul_7_15_g34493/U$1 ( \6520 , \4672 , \6480 );
nand \mul_7_15_g34228/U$1 ( \6521 , \6519 , \6520 );
and \mul_7_15_g33943/U$3 ( \6522 , \6510 , \6521 );
and \mul_7_15_g33943/U$5 ( \6523 , \6498 , \6509 );
or \mul_7_15_g33943/U$2 ( \6524 , \6522 , \6523 );
xor \mul_7_15_g35326/U$1 ( \6525 , \6410 , \6417 );
or \mul_7_15_g35308/U$1 ( \6526 , \6524 , \6525 );
not \g35889/U$3 ( \6527 , \6526 );
not \mul_7_15_g34043/U$3 ( \6528 , \6470 );
not \mul_7_15_g34229/U$1 ( \6529 , \6485 );
not \mul_7_15_g34043/U$4 ( \6530 , \6529 );
or \mul_7_15_g34043/U$2 ( \6531 , \6528 , \6530 );
nand \mul_7_15_g34070/U$1 ( \6532 , \6485 , \6469 );
nand \mul_7_15_g34043/U$1 ( \6533 , \6531 , \6532 );
and \mul_7_15_g33984/U$2 ( \6534 , \6533 , \6460 );
not \mul_7_15_g33984/U$4 ( \6535 , \6533 );
and \mul_7_15_g33984/U$3 ( \6536 , \6535 , \6459 );
nor \mul_7_15_g33984/U$1 ( \6537 , \6534 , \6536 );
not \g35889/U$4 ( \6538 , \6537 );
or \g35889/U$2 ( \6539 , \6527 , \6538 );
nand \mul_7_15_g33874/U$1 ( \6540 , \6524 , \6525 );
nand \g35889/U$1 ( \6541 , \6539 , \6540 );
nand \mul_7_15_g33640/U$1 ( \6542 , \6497 , \6541 );
not \g35883/U$4 ( \6543 , \6542 );
or \g35883/U$2 ( \6544 , \6495 , \6543 );
or \g35998/U$1 ( \6545 , \6443 , \6493 );
nand \g35883/U$1 ( \6546 , \6544 , \6545 );
not \mul_7_15_g33725/U$3 ( \6547 , \6377 );
not \mul_7_15_g33725/U$4 ( \6548 , \6380 );
and \mul_7_15_g33725/U$2 ( \6549 , \6547 , \6548 );
and \mul_7_15_g33725/U$5 ( \6550 , \6377 , \6380 );
nor \mul_7_15_g33725/U$1 ( \6551 , \6549 , \6550 );
not \mul_7_15_g33679/U$1 ( \6552 , \6551 );
not \mul_7_15_g33625/U$3 ( \6553 , \6552 );
not \mul_7_15_g33625/U$4 ( \6554 , \6330 );
or \mul_7_15_g33625/U$2 ( \6555 , \6553 , \6554 );
nand \mul_7_15_g33629/U$1 ( \6556 , \6329 , \6551 );
nand \mul_7_15_g33625/U$1 ( \6557 , \6555 , \6556 );
not \mul_7_15_g33669/U$3 ( \6558 , \6389 );
not \mul_7_15_g33669/U$4 ( \6559 , \6438 );
or \mul_7_15_g33669/U$2 ( \6560 , \6558 , \6559 );
or \mul_7_15_g33690/U$2 ( \6561 , \6438 , \6389 );
nand \mul_7_15_g33690/U$1 ( \6562 , \6561 , \6435 );
nand \mul_7_15_g33669/U$1 ( \6563 , \6560 , \6562 );
nor \mul_7_15_g33554/U$1 ( \6564 , \6557 , \6563 );
or \mul_7_15_g33513/U$2 ( \6565 , \6546 , \6564 );
nand \mul_7_15_g33557/U$1 ( \6566 , \6557 , \6563 );
nand \mul_7_15_g33513/U$1 ( \6567 , \6565 , \6566 );
and \mul_7_15_g33467/U$2 ( \6568 , \6387 , \6567 );
nor \mul_7_15_g33522/U$1 ( \6569 , \6327 , \6386 );
nor \mul_7_15_g33467/U$1 ( \6570 , \6568 , \6569 );
buf \mul_7_15_g33553/U$1 ( \6571 , \6564 );
or \mul_7_15_g35286/U$1 ( \6572 , \6497 , \6541 );
nand \mul_7_15_g33584/U$1 ( \6573 , \6545 , \6572 );
nor \mul_7_15_g33520/U$1 ( \6574 , \6571 , \6573 );
xor \mul_7_15_g33769/U$1 ( \6575 , \6525 , \6524 );
xnor \mul_7_15_g33769/U$1_r1 ( \6576 , \6575 , \6537 );
xor \mul_7_15_g33943/U$1 ( \6577 , \6498 , \6509 );
xor \mul_7_15_g33943/U$1_r1 ( \6578 , \6577 , \6521 );
not \mul_7_15_g34777/U$3 ( \6579 , \4029 );
not \mul_7_15_g34777/U$4 ( \6580 , \4069 );
or \mul_7_15_g34777/U$2 ( \6581 , \6579 , \6580 );
nand \mul_7_15_g34876/U$1 ( \6582 , \4407 , \5339 );
nand \mul_7_15_g34777/U$1 ( \6583 , \6581 , \6582 );
not \mul_7_15_g34220/U$3 ( \6584 , \6583 );
not \mul_7_15_g34220/U$4 ( \6585 , \6162 );
or \mul_7_15_g34220/U$2 ( \6586 , \6584 , \6585 );
nand \mul_7_15_g34492/U$1 ( \6587 , \4055 , \6466 );
nand \mul_7_15_g34220/U$1 ( \6588 , \6586 , \6587 );
not \mul_7_15_g33990/U$2 ( \6589 , \6588 );
not \mul_7_15_g34562/U$3 ( \6590 , \5388 );
not \mul_7_15_g34562/U$4 ( \6591 , \4049 );
or \mul_7_15_g34562/U$2 ( \6592 , \6590 , \6591 );
nand \mul_7_15_g34562/U$1 ( \6593 , \6592 , \4665 );
nand \mul_7_15_g34815/U$1 ( \6594 , \1454 , \4048 );
nand \mul_7_15_g34540/U$1 ( \6595 , \6593 , \4070 , \6594 );
not \mul_7_15_g35328/U$2 ( \6596 , \6595 );
not \mul_7_15_g34336/U$3 ( \6597 , \5019 );
not \mul_7_15_g34794/U$3 ( \6598 , \4019 );
not \mul_7_15_g34794/U$4 ( \6599 , \5023 );
or \mul_7_15_g34794/U$2 ( \6600 , \6598 , \6599 );
nand \mul_7_15_g34883/U$1 ( \6601 , \6502 , \4585 );
nand \mul_7_15_g34794/U$1 ( \6602 , \6600 , \6601 );
not \mul_7_15_g34336/U$4 ( \6603 , \6602 );
or \mul_7_15_g34336/U$2 ( \6604 , \6597 , \6603 );
nand \mul_7_15_g34346/U$1 ( \6605 , \6504 , \5021 );
nand \mul_7_15_g34336/U$1 ( \6606 , \6604 , \6605 );
nand \mul_7_15_g35328/U$1 ( \6607 , \6596 , \6606 );
nand \mul_7_15_g33990/U$1 ( \6608 , \6589 , \6607 );
and \mul_7_15_g33840/U$2 ( \6609 , \6578 , \6608 );
not \mul_7_15_g33989/U$2 ( \6610 , \6588 );
nor \mul_7_15_g33989/U$1 ( \6611 , \6610 , \6607 );
nor \mul_7_15_g33840/U$1 ( \6612 , \6609 , \6611 );
nand \mul_7_15_g33661/U$1 ( \6613 , \6576 , \6612 );
not \mul_7_15_g33592/U$3 ( \6614 , \6613 );
not \mul_7_15_g33965/U$3 ( \6615 , \6588 );
not \mul_7_15_g33965/U$4 ( \6616 , \6607 );
and \mul_7_15_g33965/U$2 ( \6617 , \6615 , \6616 );
and \mul_7_15_g33965/U$5 ( \6618 , \6588 , \6607 );
nor \mul_7_15_g33965/U$1 ( \6619 , \6617 , \6618 );
xor \g35395/U$1 ( \6620 , \6578 , \6619 );
not \mul_7_15_g34084/U$3 ( \6621 , \6606 );
not \mul_7_15_g34084/U$4 ( \6622 , \6595 );
and \mul_7_15_g34084/U$2 ( \6623 , \6621 , \6622 );
and \mul_7_15_g34084/U$5 ( \6624 , \6606 , \6595 );
nor \mul_7_15_g34084/U$1 ( \6625 , \6623 , \6624 );
and \g35898/U$2 ( \6626 , \5178 , \4026 );
not \g35898/U$4 ( \6627 , \5178 );
and \g35898/U$3 ( \6628 , \6627 , \5344 );
or \g35898/U$1 ( \6629 , \6626 , \6628 );
not \mul_7_15_g34227/U$3 ( \6630 , \6629 );
not \mul_7_15_g34227/U$4 ( \6631 , \4662 );
or \mul_7_15_g34227/U$2 ( \6632 , \6630 , \6631 );
nand \mul_7_15_g34358/U$1 ( \6633 , \4672 , \6517 );
nand \mul_7_15_g34227/U$1 ( \6634 , \6632 , \6633 );
not \mul_7_15_g34226/U$1 ( \6635 , \6634 );
xor \mul_7_15_g33854/U$4 ( \6636 , \6625 , \6635 );
not \mul_7_15_g34162/U$3 ( \6637 , \4411 );
and \mul_7_15_g34804/U$2 ( \6638 , \5388 , \4070 );
not \mul_7_15_g34804/U$4 ( \6639 , \5388 );
and \mul_7_15_g34804/U$3 ( \6640 , \6639 , \4399 );
nor \mul_7_15_g34804/U$1 ( \6641 , \6638 , \6640 );
not \mul_7_15_g34162/U$4 ( \6642 , \6641 );
and \mul_7_15_g34162/U$2 ( \6643 , \6637 , \6642 );
not \mul_7_15_g35336/U$2 ( \6644 , \6583 );
nor \mul_7_15_g35336/U$1 ( \6645 , \6644 , \4056 );
nor \mul_7_15_g34162/U$1 ( \6646 , \6643 , \6645 );
and \mul_7_15_g33854/U$3 ( \6647 , \6636 , \6646 );
and \mul_7_15_g33854/U$5 ( \6648 , \6625 , \6635 );
or \mul_7_15_g33854/U$2 ( \6649 , \6647 , \6648 );
nand \mul_7_15_g33772/U$1 ( \6650 , \6620 , \6649 );
not \mul_7_15_g34787/U$3 ( \6651 , \4026 );
not \mul_7_15_g34787/U$4 ( \6652 , \5874 );
or \mul_7_15_g34787/U$2 ( \6653 , \6651 , \6652 );
nand \mul_7_15_g34843/U$1 ( \6654 , \5024 , \5344 );
nand \mul_7_15_g34787/U$1 ( \6655 , \6653 , \6654 );
not \mul_7_15_g34314/U$3 ( \6656 , \6655 );
not \mul_7_15_g34314/U$4 ( \6657 , \5020 );
or \mul_7_15_g34314/U$2 ( \6658 , \6656 , \6657 );
not \mul_7_15_g34786/U$3 ( \6659 , \4023 );
not \mul_7_15_g34786/U$4 ( \6660 , \5874 );
or \mul_7_15_g34786/U$2 ( \6661 , \6659 , \6660 );
nand \mul_7_15_g34902/U$1 ( \6662 , \5873 , \5131 );
nand \mul_7_15_g34786/U$1 ( \6663 , \6661 , \6662 );
nand \mul_7_15_g34350/U$1 ( \6664 , \6663 , \5021 );
nand \mul_7_15_g34314/U$1 ( \6665 , \6658 , \6664 );
not \mul_7_15_g34083/U$3 ( \6666 , \6665 );
not \g35896/U$2 ( \6667 , \5178 );
not \mul_7_15_g35346/U$2 ( \6668 , \4535 );
nand \mul_7_15_g35346/U$1 ( \6669 , \6668 , \4048 );
not \mul_7_15_g34561/U$3 ( \6670 , \5388 );
not \mul_7_15_g34561/U$4 ( \6671 , \4535 );
or \mul_7_15_g34561/U$2 ( \6672 , \6670 , \6671 );
nand \mul_7_15_g34561/U$1 ( \6673 , \6672 , \5873 );
nand \g35896/U$1 ( \6674 , \6667 , \6669 , \6673 );
not \mul_7_15_g34083/U$4 ( \6675 , \6674 );
and \mul_7_15_g34083/U$2 ( \6676 , \6666 , \6675 );
and \mul_7_15_g34083/U$5 ( \6677 , \6665 , \6674 );
nor \mul_7_15_g34083/U$1 ( \6678 , \6676 , \6677 );
not \mul_7_15_g34225/U$3 ( \6679 , \4663 );
and \mul_7_15_g34807/U$2 ( \6680 , \5388 , \4665 );
not \mul_7_15_g34807/U$4 ( \6681 , \5388 );
and \mul_7_15_g34807/U$3 ( \6682 , \6681 , \4666 );
nor \mul_7_15_g34807/U$1 ( \6683 , \6680 , \6682 );
not \mul_7_15_g34225/U$4 ( \6684 , \6683 );
and \mul_7_15_g34225/U$2 ( \6685 , \6679 , \6684 );
not \mul_7_15_g34732/U$3 ( \6686 , \4029 );
not \mul_7_15_g34732/U$4 ( \6687 , \4666 );
or \mul_7_15_g34732/U$2 ( \6688 , \6686 , \6687 );
not \mul_7_15_g35343/U$2 ( \6689 , \5178 );
nand \mul_7_15_g35343/U$1 ( \6690 , \6689 , \5339 );
nand \mul_7_15_g34732/U$1 ( \6691 , \6688 , \6690 );
and \mul_7_15_g35331/U$1 ( \6692 , \5187 , \6691 );
nor \mul_7_15_g34225/U$1 ( \6693 , \6685 , \6692 );
or \mul_7_15_g35310/U$1 ( \6694 , \6678 , \6693 );
not \mul_7_15_g34810/U$3 ( \6695 , \4048 );
not \mul_7_15_g34810/U$4 ( \6696 , \5874 );
or \mul_7_15_g34810/U$2 ( \6697 , \6695 , \6696 );
nand \mul_7_15_g34944/U$1 ( \6698 , \5024 , \5388 );
nand \mul_7_15_g34810/U$1 ( \6699 , \6697 , \6698 );
and \mul_7_15_g34315/U$2 ( \6700 , \5020 , \6699 );
not \mul_7_15_g34796/U$3 ( \6701 , \4029 );
not \mul_7_15_g34796/U$4 ( \6702 , \5874 );
or \mul_7_15_g34796/U$2 ( \6703 , \6701 , \6702 );
nand \mul_7_15_g34889/U$1 ( \6704 , \5873 , \5339 );
nand \mul_7_15_g34796/U$1 ( \6705 , \6703 , \6704 );
and \mul_7_15_g34315/U$3 ( \6706 , \6705 , \5021 );
nor \mul_7_15_g34315/U$1 ( \6707 , \6700 , \6706 );
nand \mul_7_15_g34836/U$1 ( \6708 , \5021 , \4048 );
nand \mul_7_15_g34560/U$1 ( \6709 , \5024 , \6708 );
nor \mul_7_15_g34090/U$1 ( \6710 , \6707 , \6709 );
not \g35892/U$3 ( \6711 , \6710 );
not \mul_7_15_g34319/U$3 ( \6712 , \5020 );
not \mul_7_15_g34319/U$4 ( \6713 , \6705 );
or \mul_7_15_g34319/U$2 ( \6714 , \6712 , \6713 );
nand \mul_7_15_g34487/U$1 ( \6715 , \6655 , \5021 );
nand \mul_7_15_g34319/U$1 ( \6716 , \6714 , \6715 );
not \mul_7_15_g34096/U$2 ( \6717 , \6716 );
nand \mul_7_15_g34511/U$1 ( \6718 , \5187 , \4048 );
nand \mul_7_15_g34096/U$1 ( \6719 , \6717 , \6718 );
not \g35892/U$4 ( \6720 , \6719 );
or \g35892/U$2 ( \6721 , \6711 , \6720 );
not \mul_7_15_g35325/U$2 ( \6722 , \6718 );
nand \mul_7_15_g35325/U$1 ( \6723 , \6722 , \6716 );
nand \g35892/U$1 ( \6724 , \6721 , \6723 );
nand \mul_7_15_g33988/U$1 ( \6725 , \6678 , \6693 );
nand \mul_7_15_g33860/U$1 ( \6726 , \6724 , \6725 );
nand \mul_7_15_g33839/U$1 ( \6727 , \6694 , \6726 );
not \g35888/U$3 ( \6728 , \6727 );
nand \mul_7_15_g34520/U$1 ( \6729 , \4055 , \4048 );
not \mul_7_15_g34793/U$1 ( \6730 , \6602 );
not \mul_7_15_g34331/U$3 ( \6731 , \6730 );
not \mul_7_15_g34331/U$4 ( \6732 , \5265 );
and \mul_7_15_g34331/U$2 ( \6733 , \6731 , \6732 );
and \mul_7_15_g34331/U$5 ( \6734 , \6663 , \5020 );
nor \mul_7_15_g34331/U$1 ( \6735 , \6733 , \6734 );
xor \mul_7_15_g33972/U$1 ( \6736 , \6729 , \6735 );
not \mul_7_15_g34247/U$3 ( \6737 , \6691 );
not \mul_7_15_g34247/U$4 ( \6738 , \4662 );
or \mul_7_15_g34247/U$2 ( \6739 , \6737 , \6738 );
nand \mul_7_15_g34340/U$1 ( \6740 , \5187 , \6629 );
nand \mul_7_15_g34247/U$1 ( \6741 , \6739 , \6740 );
xnor \mul_7_15_g33972/U$1_r1 ( \6742 , \6736 , \6741 );
not \mul_7_15_g35327/U$2 ( \6743 , \6674 );
nand \mul_7_15_g35327/U$1 ( \6744 , \6743 , \6665 );
nand \mul_7_15_g33859/U$1 ( \6745 , \6742 , \6744 );
not \g35888/U$4 ( \6746 , \6745 );
or \g35888/U$2 ( \6747 , \6728 , \6746 );
or \mul_7_15_g35307/U$1 ( \6748 , \6742 , \6744 );
nand \g35888/U$1 ( \6749 , \6747 , \6748 );
xor \mul_7_15_g33854/U$1 ( \6750 , \6625 , \6635 );
xor \mul_7_15_g33854/U$1_r1 ( \6751 , \6750 , \6646 );
not \mul_7_15_g34078/U$3 ( \6752 , \6729 );
not \mul_7_15_g34078/U$4 ( \6753 , \6735 );
or \mul_7_15_g34078/U$2 ( \6754 , \6752 , \6753 );
nand \mul_7_15_g34078/U$1 ( \6755 , \6754 , \6741 );
or \mul_7_15_g35321/U$1 ( \6756 , \6729 , \6735 );
and \mul_7_15_g35264/U$1 ( \6757 , \6755 , \6756 );
nand \mul_7_15_g33794/U$1 ( \6758 , \6751 , \6757 );
nand \mul_7_15_g33663/U$1 ( \6759 , \6650 , \6749 , \6758 );
nor \mul_7_15_g33797/U$1 ( \6760 , \6751 , \6757 );
nand \mul_7_15_g33731/U$1 ( \6761 , \6650 , \6760 );
or \mul_7_15_g35297/U$1 ( \6762 , \6620 , \6649 );
nand \mul_7_15_g33645/U$1 ( \6763 , \6759 , \6761 , \6762 );
not \mul_7_15_g33592/U$4 ( \6764 , \6763 );
or \mul_7_15_g33592/U$2 ( \6765 , \6614 , \6764 );
or \mul_7_15_g35289/U$1 ( \6766 , \6576 , \6612 );
nand \mul_7_15_g33592/U$1 ( \6767 , \6765 , \6766 );
nand \mul_7_15_g33486/U$1 ( \6768 , \6574 , \6767 , \6387 );
nand \mul_7_15_g33455/U$1 ( \6769 , \6570 , \6768 );
and \mul_7_15_g35285/U$2 ( \6770 , \6135 , \6189 );
not \mul_7_15_g35285/U$4 ( \6771 , \6135 );
and \mul_7_15_g35285/U$3 ( \6772 , \6771 , \6190 );
nor \mul_7_15_g35285/U$1 ( \6773 , \6770 , \6772 );
not \mul_7_15_g33581/U$3 ( \6774 , \6773 );
not \mul_7_15_g33581/U$4 ( \6775 , \6146 );
or \mul_7_15_g33581/U$2 ( \6776 , \6774 , \6775 );
or \mul_7_15_g33581/U$5 ( \6777 , \6773 , \6146 );
nand \mul_7_15_g33581/U$1 ( \6778 , \6776 , \6777 );
not \mul_7_15_g33546/U$1 ( \6779 , \6778 );
xor \mul_7_15_g33757/U$1 ( \6780 , \6065 , \6082 );
xor \mul_7_15_g33757/U$1_r1 ( \6781 , \6780 , \6115 );
xor \mul_7_15_g33711/U$4 ( \6782 , \6318 , \6322 );
and \mul_7_15_g33711/U$3 ( \6783 , \6782 , \6325 );
and \mul_7_15_g33711/U$5 ( \6784 , \6318 , \6322 );
or \mul_7_15_g33711/U$2 ( \6785 , \6783 , \6784 );
xor \mul_7_15_g33577/U$4 ( \6786 , \6781 , \6785 );
not \mul_7_15_g33824/U$3 ( \6787 , \6149 );
not \mul_7_15_g33824/U$4 ( \6788 , \6186 );
or \mul_7_15_g33824/U$2 ( \6789 , \6787 , \6788 );
nand \mul_7_15_g33831/U$1 ( \6790 , \6152 , \6187 );
nand \mul_7_15_g33824/U$1 ( \6791 , \6789 , \6790 );
and \mul_7_15_g33729/U$2 ( \6792 , \6791 , \6184 );
not \mul_7_15_g33729/U$4 ( \6793 , \6791 );
not \mul_7_15_g33808/U$1 ( \6794 , \6184 );
and \mul_7_15_g33729/U$3 ( \6795 , \6793 , \6794 );
nor \mul_7_15_g33729/U$1 ( \6796 , \6792 , \6795 );
and \mul_7_15_g33577/U$3 ( \6797 , \6786 , \6796 );
and \mul_7_15_g33577/U$5 ( \6798 , \6781 , \6785 );
or \mul_7_15_g33577/U$2 ( \6799 , \6797 , \6798 );
not \mul_7_15_g33576/U$1 ( \6800 , \6799 );
nand \mul_7_15_g33508/U$1 ( \6801 , \6779 , \6800 );
xor \mul_7_15_g33577/U$1 ( \6802 , \6781 , \6785 );
xor \mul_7_15_g33577/U$1_r1 ( \6803 , \6802 , \6796 );
not \mul_7_15_g33575/U$1 ( \6804 , \6803 );
or \g35885/U$2 ( \6805 , \6326 , \6288 );
buf \mul_7_15_g33807/U$1 ( \6806 , \6200 );
nand \g35885/U$1 ( \6807 , \6805 , \6806 );
nand \mul_7_15_g33658/U$1 ( \6808 , \6326 , \6288 );
nand \mul_7_15_g33616/U$1 ( \6809 , \6807 , \6808 );
not \mul_7_15_g33578/U$1 ( \6810 , \6809 );
nand \mul_7_15_g33537/U$1 ( \6811 , \6804 , \6810 );
and \mul_7_15_g33484/U$1 ( \6812 , \6801 , \6811 );
nand \mul_7_15_g35272/U$1 ( \6813 , \6198 , \6769 , \6812 );
not \mul_7_15_g33478/U$1 ( \6814 , \6126 );
not \mul_7_15_g33494/U$1 ( \6815 , \6023 );
nand \mul_7_15_g33446/U$1 ( \6816 , \6814 , \6815 );
not \mul_7_15_g33389/U$3 ( \6817 , \6816 );
not \mul_7_15_g33389/U$4 ( \6818 , \6197 );
or \mul_7_15_g33389/U$2 ( \6819 , \6817 , \6818 );
not \mul_7_15_g33477/U$1 ( \6820 , \6133 );
not \mul_7_15_g33547/U$1 ( \6821 , \6195 );
nand \mul_7_15_g33454/U$1 ( \6822 , \6820 , \6821 );
nand \mul_7_15_g33510/U$1 ( \6823 , \6778 , \6799 );
not \g35882/U$3 ( \6824 , \6823 );
nand \mul_7_15_g33535/U$1 ( \6825 , \6803 , \6809 );
not \g35882/U$4 ( \6826 , \6825 );
or \g35882/U$2 ( \6827 , \6824 , \6826 );
nand \g35882/U$1 ( \6828 , \6827 , \6801 );
nand \mul_7_15_g33405/U$1 ( \6829 , \6822 , \6828 , \6816 );
nand \mul_7_15_g33389/U$1 ( \6830 , \6819 , \6829 );
nand \mul_7_15_g33364/U$1 ( \6831 , \6813 , \6830 );
not \mul_7_15_g33435/U$3 ( \6832 , \5740 );
not \mul_7_15_g33496/U$3 ( \6833 , \5686 );
not \mul_7_15_g33496/U$4 ( \6834 , \5690 );
and \mul_7_15_g33496/U$2 ( \6835 , \6833 , \6834 );
and \mul_7_15_g33496/U$5 ( \6836 , \5686 , \5690 );
nor \mul_7_15_g33496/U$1 ( \6837 , \6835 , \6836 );
not \mul_7_15_g33435/U$4 ( \6838 , \6837 );
or \mul_7_15_g33435/U$2 ( \6839 , \6832 , \6838 );
or \mul_7_15_g33435/U$5 ( \6840 , \5740 , \6837 );
nand \mul_7_15_g33435/U$1 ( \6841 , \6839 , \6840 );
not \mul_7_15_g33410/U$1 ( \6842 , \6841 );
xor \mul_7_15_g35206/U$4 ( \6843 , \5954 , \5956 );
and \mul_7_15_g35206/U$3 ( \6844 , \6843 , \5959 );
and \mul_7_15_g35206/U$5 ( \6845 , \5954 , \5956 );
or \mul_7_15_g35206/U$2 ( \6846 , \6844 , \6845 );
not \mul_7_15_g33811/U$1 ( \6847 , \6009 );
nand \mul_7_15_g33776/U$1 ( \6848 , \6847 , \6006 );
not \mul_7_15_g33649/U$3 ( \6849 , \6848 );
not \mul_7_15_g33649/U$4 ( \6850 , \6001 );
or \mul_7_15_g33649/U$2 ( \6851 , \6849 , \6850 );
or \mul_7_15_g35295/U$1 ( \6852 , \6847 , \6006 );
nand \mul_7_15_g33649/U$1 ( \6853 , \6851 , \6852 );
xor \mul_7_15_g33476/U$4 ( \6854 , \6846 , \6853 );
xor \mul_7_15_g33569/U$1 ( \6855 , \5732 , \5734 );
xor \mul_7_15_g33569/U$1_r1 ( \6856 , \6855 , \5737 );
and \mul_7_15_g33476/U$3 ( \6857 , \6854 , \6856 );
and \mul_7_15_g33476/U$5 ( \6858 , \6846 , \6853 );
or \mul_7_15_g33476/U$2 ( \6859 , \6857 , \6858 );
not \mul_7_15_g33475/U$1 ( \6860 , \6859 );
nand \mul_7_15_g33384/U$1 ( \6861 , \6842 , \6860 );
xor \mul_7_15_g33476/U$1 ( \6862 , \6846 , \6853 );
xor \mul_7_15_g33476/U$1_r1 ( \6863 , \6862 , \6856 );
not \mul_7_15_g33474/U$1 ( \6864 , \6863 );
not \g36014/U$3 ( \6865 , \6018 );
not \g36014/U$4 ( \6866 , \5965 );
or \g36014/U$2 ( \6867 , \6865 , \6866 );
not \mul_7_15_g33745/U$1 ( \6868 , \5965 );
not \g36015/U$3 ( \6869 , \6868 );
not \g36015/U$4 ( \6870 , \6019 );
or \g36015/U$2 ( \6871 , \6869 , \6870 );
nand \g36015/U$1 ( \6872 , \6871 , \5922 );
nand \g36014/U$1 ( \6873 , \6867 , \6872 );
not \mul_7_15_g33495/U$1 ( \6874 , \6873 );
nand \mul_7_15_g33444/U$1 ( \6875 , \6864 , \6874 );
and \mul_7_15_g33362/U$1 ( \6876 , \6861 , \6875 );
nand \mul_7_15_g33328/U$1 ( \6877 , \5745 , \6831 , \6876 );
nand \mul_7_15_g33387/U$1 ( \6878 , \6841 , \6859 );
nand \mul_7_15_g33442/U$1 ( \6879 , \6863 , \6873 );
nand \mul_7_15_g33360/U$1 ( \6880 , \6878 , \6879 );
and \mul_7_15_g33343/U$1 ( \6881 , \6880 , \6861 );
nand \mul_7_15_g33320/U$1 ( \6882 , \6881 , \5745 );
buf \mul_7_15_g33396/U$1 ( \6883 , \5682 );
nor \mul_7_15_g33375/U$1 ( \6884 , \5684 , \5743 );
and \mul_7_15_g33341/U$2 ( \6885 , \6883 , \6884 );
nor \mul_7_15_g33398/U$1 ( \6886 , \5681 , \5563 );
nor \mul_7_15_g33341/U$1 ( \6887 , \6885 , \6886 );
nand \mul_7_15_g33312/U$1 ( \6888 , \6877 , \6882 , \6887 );
not \mul_7_15_g33302/U$4 ( \6889 , \6888 );
or \mul_7_15_g33302/U$2 ( \6890 , \5561 , \6889 );
or \mul_7_15_g35274/U$1 ( \6891 , \5206 , \5382 );
or \mul_7_15_g35273/U$1 ( \6892 , \5385 , \5509 );
nand \mul_7_15_g33346/U$1 ( \6893 , \6891 , \6892 );
not \mul_7_15_g33371/U$1 ( \6894 , \5383 );
nor \mul_7_15_g33319/U$1 ( \6895 , \5558 , \6894 );
and \mul_7_15_g33313/U$2 ( \6896 , \6893 , \6895 );
or \mul_7_15_g35271/U$1 ( \6897 , \5538 , \5542 );
not \mul_7_15_g33355/U$1 ( \6898 , \5557 );
or \mul_7_15_g33324/U$2 ( \6899 , \6897 , \6898 );
not \mul_7_15_g35275/U$2 ( \6900 , \5556 );
nand \mul_7_15_g35275/U$1 ( \6901 , \6900 , \5553 );
nand \mul_7_15_g33324/U$1 ( \6902 , \6899 , \6901 );
nor \mul_7_15_g33313/U$1 ( \6903 , \6896 , \6902 );
nand \mul_7_15_g33302/U$1 ( \6904 , \6890 , \6903 );
not \mul_7_15_g33290/U$4 ( \6905 , \6904 );
or \mul_7_15_g33290/U$2 ( \6906 , \4985 , \6905 );
not \mul_7_15_g33561/U$1 ( \6907 , \4960 );
not \mul_7_15_g33315/U$3 ( \6908 , \6907 );
not \mul_7_15_g33326/U$3 ( \6909 , \4927 );
nand \mul_7_15_g33414/U$1 ( \6910 , \4515 , \4692 );
not \mul_7_15_g33393/U$2 ( \6911 , \6910 );
nand \mul_7_15_g33393/U$1 ( \6912 , \6911 , \4766 );
nand \mul_7_15_g33458/U$1 ( \6913 , \4764 , \4698 );
nand \mul_7_15_g33460/U$1 ( \6914 , \4771 , \4832 );
nand \mul_7_15_g33526/U$1 ( \6915 , \4840 , \4883 );
and \mul_7_15_g33425/U$1 ( \6916 , \6913 , \6914 , \6915 );
and \mul_7_15_g33350/U$2 ( \6917 , \6912 , \6916 );
and \mul_7_15_g33424/U$2 ( \6918 , \4834 , \4885 );
not \fopt35509/U$1 ( \6919 , \6915 );
nor \mul_7_15_g33424/U$1 ( \6920 , \6918 , \6919 );
nor \mul_7_15_g33350/U$1 ( \6921 , \6917 , \6920 );
not \mul_7_15_g33326/U$4 ( \6922 , \6921 );
or \mul_7_15_g33326/U$2 ( \6923 , \6909 , \6922 );
or \mul_7_15_g35279/U$1 ( \6924 , \4920 , \4926 );
nand \mul_7_15_g33326/U$1 ( \6925 , \6923 , \6924 );
not \mul_7_15_g33315/U$4 ( \6926 , \6925 );
or \mul_7_15_g33315/U$2 ( \6927 , \6908 , \6926 );
nand \mul_7_15_g33558/U$1 ( \6928 , \4932 , \4959 );
nand \mul_7_15_g33315/U$1 ( \6929 , \6927 , \6928 );
not \fopt35588/U$1 ( \6930 , \4983 );
and \mul_7_15_g33299/U$2 ( \6931 , \6929 , \6930 );
and \mul_7_15_g33630/U$1 ( \6932 , \4964 , \4982 );
nor \mul_7_15_g33299/U$1 ( \6933 , \6931 , \6932 );
nand \mul_7_15_g33290/U$1 ( \6934 , \6906 , \6933 );
not \mul_7_15_g34658/U$1 ( \6935 , \4978 );
and \mul_7_15_g34293/U$2 ( \6936 , \4815 , \6935 );
and \mul_7_15_g34293/U$3 ( \6937 , \4859 , \4156 );
nor \mul_7_15_g34293/U$1 ( \6938 , \6936 , \6937 );
not \mul_7_15_g34033/U$3 ( \6939 , \6938 );
nand \mul_7_15_g34826/U$1 ( \6940 , \4156 , \4044 );
not \mul_7_15_g34033/U$4 ( \6941 , \6940 );
and \mul_7_15_g34033/U$2 ( \6942 , \6939 , \6941 );
and \mul_7_15_g34033/U$5 ( \6943 , \6938 , \6940 );
nor \mul_7_15_g34033/U$1 ( \6944 , \6942 , \6943 );
not \mul_7_15_g33843/U$3 ( \6945 , \6944 );
xor \mul_7_15_g33941/U$4 ( \6946 , \4972 , \4973 );
and \mul_7_15_g33941/U$3 ( \6947 , \6946 , \4980 );
and \mul_7_15_g33941/U$5 ( \6948 , \4972 , \4973 );
or \mul_7_15_g33941/U$2 ( \6949 , \6947 , \6948 );
not \mul_7_15_g33843/U$4 ( \6950 , \6949 );
or \mul_7_15_g33843/U$2 ( \6951 , \6945 , \6950 );
or \mul_7_15_g33843/U$5 ( \6952 , \6949 , \6944 );
nand \mul_7_15_g33843/U$1 ( \6953 , \6951 , \6952 );
not \mul_7_15_g33668/U$3 ( \6954 , \6953 );
xor \mul_7_15_g33743/U$4 ( \6955 , \4968 , \4969 );
and \mul_7_15_g33743/U$3 ( \6956 , \6955 , \4981 );
and \mul_7_15_g33743/U$5 ( \6957 , \4968 , \4969 );
or \mul_7_15_g33743/U$2 ( \6958 , \6956 , \6957 );
not \mul_7_15_g33668/U$4 ( \6959 , \6958 );
or \mul_7_15_g33668/U$2 ( \6960 , \6954 , \6959 );
or \mul_7_15_g33668/U$5 ( \6961 , \6958 , \6953 );
nand \mul_7_15_g33668/U$1 ( \6962 , \6960 , \6961 );
not \mul_7_15_g33667/U$1 ( \6963 , \6962 );
and \mul_7_15_g33280/U$2 ( \6964 , \6934 , \6963 );
not \mul_7_15_g33280/U$4 ( \6965 , \6934 );
and \mul_7_15_g33280/U$3 ( \6966 , \6965 , \6962 );
nor \mul_7_15_g33280/U$1 ( \6967 , \6964 , \6966 );
not \mul_7_15_g33337/U$1 ( \6968 , \4928 );
not \mul_7_15_g33288/U$3 ( \6969 , \6968 );
not \mul_7_15_g33288/U$4 ( \6970 , \6904 );
or \mul_7_15_g33288/U$2 ( \6971 , \6969 , \6970 );
not \mul_7_15_g33325/U$1 ( \6972 , \6925 );
nand \mul_7_15_g33288/U$1 ( \6973 , \6971 , \6972 );
nand \mul_7_15_g33528/U$1 ( \6974 , \6907 , \6928 );
not \mul_7_15_g33527/U$1 ( \6975 , \6974 );
and \mul_7_15_g33281/U$2 ( \6976 , \6973 , \6975 );
not \mul_7_15_g33281/U$4 ( \6977 , \6973 );
and \mul_7_15_g33281/U$3 ( \6978 , \6977 , \6974 );
nor \mul_7_15_g33281/U$1 ( \6979 , \6976 , \6978 );
and \mul_7_15_g35619/U$1 ( \6980 , \4836 , \4885 );
not \mul_7_15_g33292/U$3 ( \6981 , \6980 );
not \mul_7_15_g33292/U$4 ( \6982 , \6904 );
or \mul_7_15_g33292/U$2 ( \6983 , \6981 , \6982 );
not \mul_7_15_g33349/U$1 ( \6984 , \6921 );
nand \mul_7_15_g33292/U$1 ( \6985 , \6983 , \6984 );
nand \mul_7_15_g33500/U$1 ( \6986 , \6924 , \4927 );
not \mul_7_15_g33499/U$1 ( \6987 , \6986 );
and \mul_7_15_g33282/U$2 ( \6988 , \6985 , \6987 );
not \mul_7_15_g33282/U$4 ( \6989 , \6985 );
and \mul_7_15_g33282/U$3 ( \6990 , \6989 , \6986 );
nor \mul_7_15_g33282/U$1 ( \6991 , \6988 , \6990 );
not \mul_7_15_g33294/U$3 ( \6992 , \4836 );
not \mul_7_15_g33294/U$4 ( \6993 , \6904 );
or \mul_7_15_g33294/U$2 ( \6994 , \6992 , \6993 );
nand \mul_7_15_g33377/U$1 ( \6995 , \6912 , \6913 );
not \mul_7_15_g33462/U$1 ( \6996 , \4835 );
and \mul_7_15_g33340/U$2 ( \6997 , \6995 , \6996 );
not \mul_7_15_g33459/U$1 ( \6998 , \6914 );
nor \mul_7_15_g33340/U$1 ( \6999 , \6997 , \6998 );
nand \mul_7_15_g33294/U$1 ( \7000 , \6994 , \6999 );
not \g35846/U$2 ( \7001 , \6919 );
nand \g35846/U$1 ( \7002 , \7001 , \4885 );
not \mul_7_15_g33501/U$1 ( \7003 , \7002 );
and \mul_7_15_g33283/U$2 ( \7004 , \7000 , \7003 );
not \mul_7_15_g33283/U$4 ( \7005 , \7000 );
and \mul_7_15_g33283/U$3 ( \7006 , \7005 , \7002 );
nor \mul_7_15_g33283/U$1 ( \7007 , \7004 , \7006 );
not \mul_7_15_g33401/U$1 ( \7008 , \4767 );
not \mul_7_15_g33293/U$3 ( \7009 , \7008 );
not \mul_7_15_g33293/U$4 ( \7010 , \6904 );
or \mul_7_15_g33293/U$2 ( \7011 , \7009 , \7010 );
not \mul_7_15_g33376/U$1 ( \7012 , \6995 );
nand \mul_7_15_g33293/U$1 ( \7013 , \7011 , \7012 );
not \mul_7_15_g33437/U$2 ( \7014 , \6998 );
nand \mul_7_15_g33437/U$1 ( \7015 , \7014 , \4834 );
not \mul_7_15_g33436/U$1 ( \7016 , \7015 );
and \mul_7_15_g33284/U$2 ( \7017 , \7013 , \7016 );
not \mul_7_15_g33284/U$4 ( \7018 , \7013 );
and \mul_7_15_g33284/U$3 ( \7019 , \7018 , \7015 );
nor \mul_7_15_g33284/U$1 ( \7020 , \7017 , \7019 );
not \mul_7_15_g33291/U$3 ( \7021 , \4694 );
not \mul_7_15_g33291/U$4 ( \7022 , \6904 );
or \mul_7_15_g33291/U$2 ( \7023 , \7021 , \7022 );
nand \mul_7_15_g33291/U$1 ( \7024 , \7023 , \6910 );
nand \mul_7_15_g33439/U$1 ( \7025 , \6913 , \4766 );
not \mul_7_15_g33438/U$1 ( \7026 , \7025 );
and \mul_7_15_g33285/U$2 ( \7027 , \7024 , \7026 );
not \mul_7_15_g33285/U$4 ( \7028 , \7024 );
and \mul_7_15_g33285/U$3 ( \7029 , \7028 , \7025 );
nor \mul_7_15_g33285/U$1 ( \7030 , \7027 , \7029 );
not \mul_7_15_g33289/U$3 ( \7031 , \5543 );
not \mul_7_15_g33306/U$3 ( \7032 , \5511 );
not \mul_7_15_g33306/U$4 ( \7033 , \6888 );
or \mul_7_15_g33306/U$2 ( \7034 , \7032 , \7033 );
not \mul_7_15_g33369/U$1 ( \7035 , \6894 );
nand \mul_7_15_g33335/U$1 ( \7036 , \6893 , \7035 );
nand \mul_7_15_g33306/U$1 ( \7037 , \7034 , \7036 );
not \mul_7_15_g33289/U$4 ( \7038 , \7037 );
or \mul_7_15_g33289/U$2 ( \7039 , \7031 , \7038 );
nand \mul_7_15_g33289/U$1 ( \7040 , \7039 , \6897 );
nand \mul_7_15_g33334/U$1 ( \7041 , \6901 , \5557 );
not \mul_7_15_g33333/U$1 ( \7042 , \7041 );
and \mul_7_15_g33286/U$2 ( \7043 , \7040 , \7042 );
not \mul_7_15_g33286/U$4 ( \7044 , \7040 );
and \mul_7_15_g33286/U$3 ( \7045 , \7044 , \7041 );
nor \mul_7_15_g33286/U$1 ( \7046 , \7043 , \7045 );
not \mul_7_15_g35278/U$2 ( \7047 , \4927 );
nor \mul_7_15_g35278/U$1 ( \7048 , \7047 , \4960 );
and \mul_7_15_g33339/U$1 ( \7049 , \6980 , \7048 );
buf \fopt35661/U$1 ( \7050 , \6888 );
nand \mul_7_15_g33308/U$1 ( \7051 , \7049 , \7050 , \5560 );
not \mul_7_15_g33307/U$2 ( \7052 , \6903 );
nand \mul_7_15_g33307/U$1 ( \7053 , \7052 , \7049 );
not \mul_7_15_g33314/U$1 ( \7054 , \6929 );
nand \mul_7_15_g33298/U$1 ( \7055 , \7051 , \7053 , \7054 );
nor \mul_7_15_g33607/U$1 ( \7056 , \6932 , \4983 );
and \mul_7_15_g33287/U$2 ( \7057 , \7055 , \7056 );
not \mul_7_15_g33287/U$4 ( \7058 , \7055 );
not \mul_7_15_g33606/U$1 ( \7059 , \7056 );
and \mul_7_15_g33287/U$3 ( \7060 , \7058 , \7059 );
nor \mul_7_15_g33287/U$1 ( \7061 , \7057 , \7060 );
buf \mul_7_15_g33399/U$1 ( \7062 , \5510 );
not \mul_7_15_g33300/U$3 ( \7063 , \7062 );
not \mul_7_15_g33300/U$4 ( \7064 , \7050 );
or \mul_7_15_g33300/U$2 ( \7065 , \7063 , \7064 );
nand \mul_7_15_g33300/U$1 ( \7066 , \7065 , \6892 );
nand \mul_7_15_g33352/U$1 ( \7067 , \7035 , \6891 );
not \mul_7_15_g33351/U$1 ( \7068 , \7067 );
and \mul_7_15_g33297/U$2 ( \7069 , \7066 , \7068 );
not \mul_7_15_g33297/U$4 ( \7070 , \7066 );
and \mul_7_15_g33297/U$3 ( \7071 , \7070 , \7067 );
nor \mul_7_15_g33297/U$1 ( \7072 , \7069 , \7071 );
nand \mul_7_15_g33379/U$1 ( \7073 , \6892 , \7062 );
not \mul_7_15_g33378/U$1 ( \7074 , \7073 );
and \mul_7_15_g33303/U$2 ( \7075 , \7050 , \7074 );
not \mul_7_15_g33303/U$4 ( \7076 , \7050 );
and \mul_7_15_g33303/U$3 ( \7077 , \7076 , \7073 );
nor \mul_7_15_g33303/U$1 ( \7078 , \7075 , \7077 );
not \mul_7_15_g33380/U$2 ( \7079 , \6886 );
nand \mul_7_15_g33380/U$1 ( \7080 , \7079 , \6883 );
buf \mul_7_15_g33363/U$1 ( \7081 , \6831 );
not \mul_7_15_g33323/U$3 ( \7082 , \7081 );
not \mul_7_15_g33323/U$4 ( \7083 , \6876 );
or \mul_7_15_g33323/U$2 ( \7084 , \7082 , \7083 );
not \mul_7_15_g33342/U$1 ( \7085 , \6881 );
nand \mul_7_15_g33323/U$1 ( \7086 , \7084 , \7085 );
buf \mul_7_15_g33382/U$1 ( \7087 , \5744 );
and \mul_7_15_g33310/U$2 ( \7088 , \7086 , \7087 );
buf \mul_7_15_g33374/U$1 ( \7089 , \6884 );
nor \mul_7_15_g33310/U$1 ( \7090 , \7088 , \7089 );
and \mul_7_15_g33304/U$2 ( \7091 , \7080 , \7090 );
not \mul_7_15_g33304/U$4 ( \7092 , \7080 );
not \mul_7_15_g33309/U$1 ( \7093 , \7090 );
and \mul_7_15_g33304/U$3 ( \7094 , \7092 , \7093 );
nor \mul_7_15_g33304/U$1 ( \7095 , \7091 , \7094 );
not \mul_7_15_g33353/U$2 ( \7096 , \7087 );
nor \mul_7_15_g33353/U$1 ( \7097 , \7096 , \7089 );
and \mul_7_15_g33316/U$2 ( \7098 , \7097 , \7086 );
not \mul_7_15_g33316/U$4 ( \7099 , \7097 );
not \mul_7_15_g33322/U$1 ( \7100 , \7086 );
and \mul_7_15_g33316/U$3 ( \7101 , \7099 , \7100 );
nor \mul_7_15_g33316/U$1 ( \7102 , \7098 , \7101 );
not \mul_7_15_g33327/U$3 ( \7103 , \6875 );
not \mul_7_15_g33327/U$4 ( \7104 , \7081 );
or \mul_7_15_g33327/U$2 ( \7105 , \7103 , \7104 );
nand \mul_7_15_g33327/U$1 ( \7106 , \7105 , \6879 );
nand \mul_7_15_g35270/U$1 ( \7107 , \6878 , \6861 );
not \mul_7_15_g33344/U$1 ( \7108 , \7107 );
and \mul_7_15_g33317/U$2 ( \7109 , \7106 , \7108 );
not \mul_7_15_g33317/U$4 ( \7110 , \7106 );
and \mul_7_15_g33317/U$3 ( \7111 , \7110 , \7107 );
nor \mul_7_15_g33317/U$1 ( \7112 , \7109 , \7111 );
nand \mul_7_15_g33418/U$1 ( \7113 , \6875 , \6879 );
not \mul_7_15_g33417/U$1 ( \7114 , \7113 );
and \mul_7_15_g33329/U$2 ( \7115 , \7081 , \7114 );
not \mul_7_15_g33329/U$4 ( \7116 , \7081 );
and \mul_7_15_g33329/U$3 ( \7117 , \7116 , \7113 );
nor \mul_7_15_g33329/U$1 ( \7118 , \7115 , \7117 );
not \mul_7_15_g33403/U$3 ( \7119 , \6812 );
not \mul_7_15_g33403/U$4 ( \7120 , \6769 );
or \mul_7_15_g33403/U$2 ( \7121 , \7119 , \7120 );
nand \mul_7_15_g33403/U$1 ( \7122 , \7121 , \6828 );
buf \mul_7_15_g33448/U$1 ( \7123 , \6196 );
and \mul_7_15_g33365/U$2 ( \7124 , \7122 , \7123 );
not \mul_7_15_g33452/U$1 ( \7125 , \6822 );
nor \mul_7_15_g33365/U$1 ( \7126 , \7124 , \7125 );
nand \mul_7_15_g33416/U$1 ( \7127 , \6127 , \6816 );
and \mul_7_15_g33330/U$2 ( \7128 , \7126 , \7127 );
not \mul_7_15_g33330/U$4 ( \7129 , \7126 );
not \mul_7_15_g33415/U$1 ( \7130 , \7127 );
and \mul_7_15_g33330/U$3 ( \7131 , \7129 , \7130 );
nor \mul_7_15_g33330/U$1 ( \7132 , \7128 , \7131 );
nand \mul_7_15_g33420/U$1 ( \7133 , \6822 , \7123 );
not \mul_7_15_g33419/U$1 ( \7134 , \7133 );
and \mul_7_15_g33366/U$2 ( \7135 , \7122 , \7134 );
not \mul_7_15_g33366/U$4 ( \7136 , \7122 );
and \mul_7_15_g33366/U$3 ( \7137 , \7136 , \7133 );
nor \mul_7_15_g33366/U$1 ( \7138 , \7135 , \7137 );
and \mul_7_15_g33404/U$2 ( \7139 , \6769 , \6811 );
not \mul_7_15_g33533/U$1 ( \7140 , \6825 );
nor \mul_7_15_g33404/U$1 ( \7141 , \7139 , \7140 );
nand \mul_7_15_g35276/U$1 ( \7142 , \6823 , \6801 );
and \mul_7_15_g33367/U$2 ( \7143 , \7141 , \7142 );
not \mul_7_15_g33367/U$4 ( \7144 , \7141 );
not \mul_7_15_g33481/U$1 ( \7145 , \7142 );
and \mul_7_15_g33367/U$3 ( \7146 , \7144 , \7145 );
nor \mul_7_15_g33367/U$1 ( \7147 , \7143 , \7146 );
and \mul_7_15_g33394/U$1 ( \7148 , \6910 , \4694 );
nand \mul_7_15_g33504/U$1 ( \7149 , \6811 , \6825 );
not \mul_7_15_g33503/U$1 ( \7150 , \7149 );
and \mul_7_15_g33407/U$2 ( \7151 , \6769 , \7150 );
not \mul_7_15_g33407/U$4 ( \7152 , \6769 );
and \mul_7_15_g33407/U$3 ( \7153 , \7152 , \7149 );
nor \mul_7_15_g33407/U$1 ( \7154 , \7151 , \7153 );
not \mul_7_15_g33551/U$1 ( \7155 , \6571 );
not \mul_7_15_g33468/U$3 ( \7156 , \7155 );
not \mul_7_15_g33511/U$3 ( \7157 , \6767 );
not \mul_7_15_g33583/U$1 ( \7158 , \6573 );
not \mul_7_15_g33511/U$4 ( \7159 , \7158 );
or \mul_7_15_g33511/U$2 ( \7160 , \7157 , \7159 );
nand \mul_7_15_g33511/U$1 ( \7161 , \7160 , \6546 );
not \mul_7_15_g33468/U$4 ( \7162 , \7161 );
or \mul_7_15_g33468/U$2 ( \7163 , \7156 , \7162 );
nand \mul_7_15_g33468/U$1 ( \7164 , \7163 , \6566 );
not \mul_7_15_g35277/U$2 ( \7165 , \6569 );
nand \mul_7_15_g35277/U$1 ( \7166 , \7165 , \6387 );
not \mul_7_15_g33505/U$1 ( \7167 , \7166 );
and \mul_7_15_g33427/U$2 ( \7168 , \7164 , \7167 );
not \mul_7_15_g33427/U$4 ( \7169 , \7164 );
and \mul_7_15_g33427/U$3 ( \7170 , \7169 , \7166 );
nor \mul_7_15_g33427/U$1 ( \7171 , \7168 , \7170 );
not \mul_7_15_g33529/U$2 ( \7172 , \6571 );
nand \mul_7_15_g33529/U$1 ( \7173 , \7172 , \6566 );
not \mul_7_15_g33472/U$3 ( \7174 , \7173 );
not \mul_7_15_g33472/U$4 ( \7175 , \7161 );
or \mul_7_15_g33472/U$2 ( \7176 , \7174 , \7175 );
or \mul_7_15_g33472/U$5 ( \7177 , \7173 , \7161 );
nand \mul_7_15_g33472/U$1 ( \7178 , \7176 , \7177 );
not \mul_7_15_g33514/U$3 ( \7179 , \6572 );
not \mul_7_15_g33514/U$4 ( \7180 , \6767 );
or \mul_7_15_g33514/U$2 ( \7181 , \7179 , \7180 );
nand \mul_7_15_g33514/U$1 ( \7182 , \7181 , \6542 );
nand \mul_7_15_g33587/U$1 ( \7183 , \6545 , \6494 );
not \mul_7_15_g33586/U$1 ( \7184 , \7183 );
and \mul_7_15_g33473/U$2 ( \7185 , \7182 , \7184 );
not \mul_7_15_g33473/U$4 ( \7186 , \7182 );
and \mul_7_15_g33473/U$3 ( \7187 , \7186 , \7183 );
nor \mul_7_15_g33473/U$1 ( \7188 , \7185 , \7187 );
nand \mul_7_15_g33608/U$1 ( \7189 , \6542 , \6572 );
not \mul_7_15_g33515/U$3 ( \7190 , \7189 );
not \mul_7_15_g33515/U$4 ( \7191 , \6767 );
or \mul_7_15_g33515/U$2 ( \7192 , \7190 , \7191 );
or \mul_7_15_g33515/U$5 ( \7193 , \7189 , \6767 );
nand \mul_7_15_g33515/U$1 ( \7194 , \7192 , \7193 );
nand \mul_7_15_g33632/U$1 ( \7195 , \6766 , \6613 );
and \mul_7_15_g33647/U$2 ( \7196 , \6749 , \6758 );
nor \mul_7_15_g33647/U$1 ( \7197 , \7196 , \6760 );
nand \mul_7_15_g33734/U$1 ( \7198 , \6762 , \6650 );
nand \mul_7_15_g33834/U$1 ( \7199 , \6748 , \6745 );
nand \mul_7_15_g33955/U$1 ( \7200 , \6694 , \6725 );
nand \mul_7_15_g34077/U$1 ( \7201 , \6723 , \6719 );
and \mul_7_15_g34080/U$2 ( \7202 , \6707 , \6709 );
nor \mul_7_15_g34080/U$1 ( \7203 , \7202 , \6710 );
not \mul_7_15_g34835/U$1 ( \7204 , \6708 );
and \mul_7_15_g35348/U$1 ( \7205 , \6897 , \5543 );
xor \mul_7_15_g35268/U$1 ( \7206 , \7037 , \7205 );
xor \mul_7_15_g35282/U$1 ( \7207 , \7198 , \7197 );
not \mul_7_15_g35294/U$2 ( \7208 , \6760 );
nand \mul_7_15_g35294/U$1 ( \7209 , \7208 , \6758 );
xnor \mul_7_15_g35288/U$1 ( \7210 , \6749 , \7209 );
xnor \mul_7_15_g35298/U$1 ( \7211 , \6727 , \7199 );
xnor \mul_7_15_g35302/U$1 ( \7212 , \7200 , \6724 );
xnor \mul_7_15_g35311/U$1 ( \7213 , \6710 , \7201 );
not \mul_7_15_g35351/U$2 ( \7214 , \7195 );
xor \mul_7_15_g35351/U$1 ( \7215 , \6763 , \7214 );
xor \g35500/U$1 ( \7216 , \7148 , \6904 );
endmodule

