//
// Conformal-LEC Version 20.10-d005 (29-Apr-2020)
//
module top(RIdec64b8_720,RIbc62af0_23,RIbc62a78_22,RIbc62a00_21,RIbc62988_20,RIbc62910_19,RIbc62898_18,RIbc62820_17,RIbc627a8_16,
        RIbc62730_15,RIbc626b8_14,RIbc62640_13,RIdec37b8_688,RIfc8daa0_6634,RIdec0ab8_656,RIfc56348_6003,RIdebddb8_624,RIdebb0b8_592,RIdeb83b8_560,
        RIfc98798_6757,RIdeb29b8_496,RIfcbd098_7173,RIdeafcb8_464,RIfc8dc08_6635,RIdeacb80_432,RIdea6280_400,RIde9f980_368,RIfcd6868_7463,RIfc8ded8_6637,
        RIfc7dd80_6454,RIfc56618_6005,RIde92e10_306,RIde8f300_288,RIde8b160_268,RIde86fc0_248,RIde82ad8_227,RIfc8e040_6638,RIfcd96d0_7496,RIfca1e10_6864,
        RIfcbd200_7174,RIe16c5c0_2610,RIe16a298_2585,RIe168ab0_2568,RIe1664b8_2541,RIe1637b8_2509,RIee37f00_5095,RIe160ab8_2477,RIfc8ea18_6645,RIe15ddb8_2445,
        RIe1583b8_2381,RIe1556b8_2349,RIfe9f828_8159,RIe1529b8_2317,RIfe9f990_8160,RIe14fcb8_2285,RIfcbd368_7175,RIe14cfb8_2253,RIe14a2b8_2221,RIe1475b8_2189,
        RIfc8ee50_6648,RIfc45278_5809,RIfc98360_6754,RIfca2248_6867,RIe141d20_2126,RIe13f9f8_2101,RIdf3d900_2077,RIdf3b470_2051,RIfcd6ca0_7466,RIee2ff08_5004,
        RIfc8ece8_6647,RIee2dd48_4980,RIdf36718_1996,RIdf34120_1969,RIdf31f60_1945,RIfe9f6c0_8158,RIfcb4560_7074,RIfc45db8_5817,RIfc8e1a8_6639,RIfc7d678_6449,
        RIdf2aee0_1865,RIdf28ff0_1843,RIdf26e30_1819,RIdf25378_1800,RIfcb43f8_7073,RIfc8e748_6643,RIdf23488_1778,RIfcc2c00_7238,RIdf21e08_1762,RIdf20788_1746,
        RIdf1b760_1689,RIdf1a248_1674,RIdf18088_1650,RIdf15388_1618,RIdf12688_1586,RIdf0f988_1554,RIdf0cc88_1522,RIdf09f88_1490,RIdf07288_1458,RIdf04588_1426,
        RIdefeb88_1362,RIdefbe88_1330,RIdef9188_1298,RIdef6488_1266,RIdef3788_1234,RIdef0a88_1202,RIdeedd88_1170,RIdeeb088_1138,RIfc8efb8_6649,RIfc44e40_5806,
        RIfc57860_6018,RIfca23b0_6868,RIfe9faf8_8161,RIdee3900_1053,RIdee1740_1029,RIdedf6e8_1006,RIfcbd4d0_7176,RIee22678_4850,RIfc98090_6752,RIee21598_4838,
        RIfe9fc60_8162,RIded80c8_922,RIfe9fdc8_8163,RIded3be0_873,RIded18b8_848,RIdecebb8_816,RIdecbeb8_784,RIdec91b8_752,RIdeb56b8_528,RIde99080_336,
        RIe16f2c0_2642,RIe15b0b8_2413,RIe1448b8_2157,RIdf392b0_2027,RIdf2d910_1895,RIdf1e190_1719,RIdf01888_1394,RIdee8388_1106,RIdedd0f0_979,RIde7efc8_209,
        RIe19e750_3180,RIbc625c8_12,RIbc62550_11,RIbc624d8_10,RIbc62460_9,RIbc623e8_8,RIbc62370_7,RIbc622f8_6,RIbc62280_5,RIbc62208_4,
        RIbc62190_3,RIbc62118_2,RIe19ba50_3148,RIfc479d8_5837,RIe198d50_3116,RIfe9f558_8157,RIe196050_3084,RIe193350_3052,RIe190650_3020,RIe18ac50_2956,
        RIe187f50_2924,RIfc47870_5836,RIe185250_2892,RIf142ef8_5221,RIe182550_2860,RIe17f850_2828,RIe17cb50_2796,RIfcb5208_7083,RIfcbc6c0_7166,RIe177588_2735,
        RIe176610_2724,RIf13fdc0_5186,RIfe9f3f0_8156,RIfce40f8_7617,RIfc47708_5835,RIfc47438_5833,RIfca15a0_6858,RIfc99170_6764,RIe1745b8_2701,RIfc8cc90_6624,
        RIfc556a0_5994,RIfc7ee60_6466,RIfce8e50_7672,RIfe9f288_8155,RIe224aa8_4707,RIfc55808_5995,RIe221da8_4675,RIfcb50a0_7082,RIe21f0a8_4643,RIe2196a8_4579,
        RIe2169a8_4547,RIfcbc828_7167,RIe213ca8_4515,RIfc47000_5830,RIe210fa8_4483,RIfcbc990_7168,RIe20e2a8_4451,RIe20b5a8_4419,RIe2088a8_4387,RIfc46bc8_5827,
        RIfcd6598_7461,RIe2032e0_4326,RIe2016c0_4306,RIfc98ea0_6762,RIfc7eb90_6464,RIfce0318_7573,RIfcbcaf8_7169,RIfc8cf60_6626,RIfcb4dd0_7080,RIe1fd340_4258,
        RIe1fc260_4246,RIf15cf38_5517,RIfe9f120_8154,RIfc7ea28_6463,RIfc8d0c8_6627,RIfcbcc60_7170,RIfc98bd0_6760,RIfce2d48_7603,RIe1fb018_4233,RIfc55f10_6000,
        RIfc7e8c0_6462,RIfc8d230_6628,RIe1f6590_4180,RIfce58e0_7634,RIfc468f8_5825,RIfcc2ed0_7240,RIe1f4100_4154,RIfceedf0_7740,RIfc8d398_6629,RIfc8d500_6630,
        RIe1eef70_4096,RIe1ec810_4068,RIe1e9b10_4036,RIe1e6e10_4004,RIe1e4110_3972,RIe1e1410_3940,RIe1de710_3908,RIe1dba10_3876,RIe1d8d10_3844,RIe1d3310_3780,
        RIe1d0610_3748,RIe1cd910_3716,RIe1cac10_3684,RIe1c7f10_3652,RIe1c5210_3620,RIe1c2510_3588,RIe1bf810_3556,RIf14d0b0_5336,RIfe9efb8_8153,RIe1ba248_3495,
        RIe1b8088_3471,RIfec4dd0_8360,RIfec50a0_8362,RIe1b5ec8_3447,RIe1b46e0_3430,RIfcb4998_7077,RIfcb4c68_7079,RIfec5370_8364,RIfe9ee50_8152,RIfcbcdc8_7171,
        RIfc46358_5821,RIfec5208_8363,RIfec4f38_8361,RIe1a9b50_3308,RIe1a6e50_3276,RIe1a4150_3244,RIe1a1450_3212,RIe18d950_2988,RIe179e50_2764,RIe2277a8_4739,
        RIe21c3a8_4611,RIe205ba8_4355,RIe1ffc08_4287,RIe1f8fc0_4210,RIe1f1b08_4127,RIe1d6010_3812,RIe1bcb10_3524,RIe1af988_3375,RIe171fc0_2674,RIdec6080_717,
        RIdec3380_685,RIee204b8_4826,RIdec0680_653,RIfcd70d8_7469,RIdebd980_621,RIdebac80_589,RIdeb7f80_557,RIfcbe448_7187,RIdeb2580_493,RIfcb3480_7062,
        RIdeaf880_461,RIfc43928_5791,RIdeac1a8_429,RIdea58a8_397,RIde9efa8_365,RIfcd88c0_7486,RIee1c408_4780,RIfcc77f0_7292,RIfea04d0_8168,RIde92438_303,
        RIde8ec70_286,RIde8aad0_266,RIde86930_246,RIfca31c0_6878,RIfc59a20_6042,RIfcd1de0_7410,RIfc91448_6675,RIfc97280_6742,RIe16c188_2607,RIfc97118_6741,
        RIe168948_2567,RIe166080_2538,RIe163380_2506,RIee37ac8_5092,RIe160680_2474,RIfcd1c78_7409,RIe15d980_2442,RIe157f80_2378,RIe155280_2346,RIfc3f530_5746,
        RIe152580_2314,RIee35368_5064,RIe14f880_2282,RIfc7a3d8_6413,RIe14cb80_2250,RIe149e80_2218,RIe147180_2186,RIfc42b18_5781,RIfc7a270_6412,RIfc5a560_6050,
        RIfc96b78_6737,RIfea6fb0_8216,RIe13f5c0_2098,RIdf3d4c8_2074,RIdf3b038_2048,RIfce5bb0_7636,RIee2fc38_5002,RIfc91cb8_6681,RIee2d910_4977,RIdf362e0_1993,
        RIdf33e50_1967,RIdf31c90_1943,RIdf2fda0_1921,RIfc43658_5789,RIfc59e58_6045,RIfc96fb0_6740,RIfc7ac48_6419,RIfea0368_8167,RIdf28bb8_1840,RIdf26cc8_1818,
        RIdf25210_1799,RIfc91718_6677,RIfcb3318_7061,RIfc919e8_6679,RIfc91880_6678,RIfc430b8_5785,RIdf20350_1743,RIfc7a978_6417,RIdf19e10_1671,RIdf17c50_1647,
        RIdf14f50_1615,RIdf12250_1583,RIdf0f550_1551,RIdf0c850_1519,RIdf09b50_1487,RIdf06e50_1455,RIdf04150_1423,RIdefe750_1359,RIdefba50_1327,RIdef8d50_1295,
        RIdef6050_1263,RIdef3350_1231,RIdef0650_1199,RIdeed950_1167,RIdeeac50_1135,RIfcd1b10_7408,RIfc968a8_6735,RIfc91f88_6683,RIfcdfc10_7568,RIfea99e0_8246,
        RIdee3630_1051,RIdee1308_1026,RIdedf2b0_1003,RIfcc7d90_7296,RIfcd85f0_7484,RIfce3888_7611,RIfc5a830_6052,RIdeda3f0_947,RIfea9878_8245,RIded5f08_898,
        RIded37a8_870,RIded1480_845,RIdece780_813,RIdecba80_781,RIdec8d80_749,RIdeb5280_525,RIde986a8_333,RIe16ee88_2639,RIe15ac80_2410,RIe144480_2154,
        RIdf38e78_2024,RIdf2d4d8_1892,RIdf1dd58_1716,RIdf01450_1391,RIdee7f50_1103,RIdedccb8_976,RIde7e5f0_206,RIe19e318_3177,RIe19b618_3145,RIfc8f3f0_6652,
        RIe198918_3113,RIf144b18_5241,RIe195c18_3081,RIe192f18_3049,RIe190218_3017,RIe18a818_2953,RIe187b18_2921,RIf143d08_5231,RIe184e18_2889,RIfcb3cf0_7068,
        RIe182118_2857,RIe17f418_2825,RIe17c718_2793,RIfc448a0_5802,RIf141170_5200,RIfc7c9d0_6440,RIfea0098_8165,RIfc57e00_6022,RIf13f550_5180,RIfcd6e08_7467,
        RIee3d900_5159,RIfc8f6c0_6654,RIfce0048_7571,RIfca27e8_6871,RIe1742e8_2699,RIfc7c700_6438,RIfc8f990_6656,RIfce9828_7679,RIfc583a0_6026,RIf16cdc0_5698,
        RIe224670_4704,RIf16c118_5689,RIe221970_4672,RIfc58508_6027,RIe21ec70_4640,RIe219270_4576,RIe216570_4544,RIfc3ff08_5753,RIe213870_4512,RIf1696e8_5659,
        RIe210b70_4480,RIfc58940_6030,RIe20de70_4448,RIe20b170_4416,RIe208470_4384,RIfc8fc60_6658,RIfc97820_6746,RIe202ea8_4323,RIe201288_4303,RIfcc27c8_7235,
        RIfcdfee0_7570,RIfc44198_5797,RIfc58670_6028,RIf1608e0_5558,RIf15e9f0_5536,RIfe9ff30_8164,RIe1fc0f8_4245,RIfc7be90_6432,RIf15bb88_5503,RIfcd8cf8_7489,
        RIfcd8e60_7490,RIfca2d88_6875,RIfcbdea8_7183,RIfcb3a20_7066,RIe1fabe0_4230,RIfc90098_6661,RIfc90200_6662,RIfcd20b0_7412,RIe1f6158_4177,RIfc904d0_6664,
        RIfca2ef0_6876,RIfc97550_6744,RIe1f3e30_4152,RIfc59048_6035,RIfc907a0_6666,RIfc90638_6665,RIe1eeb38_4093,RIe1ec3d8_4065,RIe1e96d8_4033,RIe1e69d8_4001,
        RIe1e3cd8_3969,RIe1e0fd8_3937,RIe1de2d8_3905,RIe1db5d8_3873,RIe1d88d8_3841,RIe1d2ed8_3777,RIe1d01d8_3745,RIe1cd4d8_3713,RIe1ca7d8_3681,RIe1c7ad8_3649,
        RIe1c4dd8_3617,RIe1c20d8_3585,RIe1bf3d8_3553,RIfcc73b8_7289,RIfce3cc0_7614,RIe1b9e10_3492,RIe1b7c50_3468,RIfcd6f70_7468,RIf149e10_5300,RIe1b5a90_3444,
        RIfea0200_8166,RIfc90bd8_6669,RIfcdfd78_7569,RIe1b2ef8_3413,RIe1b15a8_3395,RIfc973e8_6743,RIfcc7520_7290,RIe1acdf0_3344,RIe1ab608_3327,RIe1a9718_3305,
        RIe1a6a18_3273,RIe1a3d18_3241,RIe1a1018_3209,RIe18d518_2985,RIe179a18_2761,RIe227370_4736,RIe21bf70_4608,RIe205770_4352,RIe1ff7d0_4284,RIe1f8b88_4207,
        RIe1f16d0_4124,RIe1d5bd8_3809,RIe1bc6d8_3521,RIe1af550_3372,RIe171b88_2671,RIdec5108_706,RIdec2408_674,RIfc93608_6699,RIdebf708_642,RIfc934a0_6698,
        RIdebca08_610,RIdeb9d08_578,RIdeb7008_546,RIfcdf7d8_7565,RIdeb1608_482,RIfc78218_6389,RIdeae908_450,RIfcc8498_7301,RIdea9d90_418,RIdea3490_386,
        RIde9cb90_354,RIee1cc78_4786,RIee1bb98_4774,RIee1b328_4768,RIee1aab8_4762,RIde909f8_295,RIde8d578_279,RIfea8ea0_8238,RIde85238_239,RIde813e0_220,
        RIfc938d8_6701,RIfce5e80_7638,RIfcbfd98_7205,RIfce8ce8_7671,RIe16b4e0_2598,RIfea8d38_8237,RIfea9f80_8250,RIe165108_2527,RIe162408_2495,RIfc779a8_6383,
        RIe15f708_2463,RIfe9dc08_8139,RIe15ca08_2431,RIe157008_2367,RIe154308_2335,RIfea7550_8220,RIe151608_2303,RIfcd6160_7458,RIe14e908_2271,RIfcd1408_7403,
        RIe14bc08_2239,RIe148f08_2207,RIe146208_2175,RIfceb718_7701,RIfcb19c8_7043,RIfc93e78_6705,RIfce7938_7657,RIe140da8_2115,RIdf3ecb0_2091,RIdf3c988_2066,
        RIfe9daa0_8138,RIfce8478_7665,RIfcdbf98_7525,RIfc776d8_6381,RIfc93fe0_6706,RIdf354d0_1983,RIdf33040_1957,RIdf30fe8_1934,RIdf2ee28_1910,RIee2ba20_4955,
        RIfc93ba8_6703,RIfc77de0_6386,RIee27ad8_4910,RIfe9d668_8135,RIfea8bd0_8236,RIdf26458_1812,RIfe9d7d0_8136,RIfcb1c98_7045,RIee26cc8_4900,RIdf22ab0_1771,
        RIfcc0068_7207,RIdf21598_1756,RIdf1f6a8_1734,RIdf1aef0_1683,RIfe9d938_8137,RIdf16cd8_1636,RIdf13fd8_1604,RIdf112d8_1572,RIdf0e5d8_1540,RIdf0b8d8_1508,
        RIdf08bd8_1476,RIdf05ed8_1444,RIdf031d8_1412,RIdefd7d8_1348,RIdefaad8_1316,RIdef7dd8_1284,RIdef50d8_1252,RIdef23d8_1220,RIdeef6d8_1188,RIdeec9d8_1156,
        RIdee9cd8_1124,RIfc942b0_6708,RIfcde6f8_7553,RIfcd1138_7401,RIfcde860_7554,RIdee4878_1064,RIdee2af0_1043,RIdee0a98_1020,RIdede8d8_996,RIfc5c9f0_6076,
        RIee22240_4847,RIfcc8768_7303,RIee21160_4835,RIded95e0_937,RIded7150_911,RIded5260_889,RIfea76b8_8221,RIded0508_834,RIdecd808_802,RIdecab08_770,
        RIdec7e08_738,RIdeb4308_514,RIde96290_322,RIe16df10_2628,RIe159d08_2399,RIe143508_2143,RIdf37f00_2013,RIdf2c560_1881,RIdf1cde0_1705,RIdf004d8_1380,
        RIdee6fd8_1092,RIdedbd40_965,RIde7c1d8_195,RIe19d3a0_3166,RIe19a6a0_3134,RIfcb2c10_7056,RIe1979a0_3102,RIfc923c0_6686,RIe194ca0_3070,RIe191fa0_3038,
        RIe18f2a0_3006,RIe1898a0_2942,RIe186ba0_2910,RIfc422a8_5775,RIe183ea0_2878,RIfcbecb8_7193,RIe1811a0_2846,RIe17e4a0_2814,RIe17b7a0_2782,RIf142250_5212,
        RIf140bd0_5196,RIfec43f8_8353,RIe175968_2715,RIfc79b68_6407,RIf13efb0_5176,RIfc92528_6687,RIfcb2aa8_7055,RIfcd8320_7482,RIfcea200_7686,RIfc79898_6405,
        RIe1734d8_2689,RIfcd7948_7475,RIfcd7678_7473,RIf16e170_5712,RIfc927f8_6689,RIfc92960_6690,RIe2236f8_4693,RIfc795c8_6403,RIe2209f8_4661,RIf16ad68_5675,
        RIe21dcf8_4629,RIe2182f8_4565,RIe2155f8_4533,RIfe9d398_8133,RIe2128f8_4501,RIfcdb9f8_7521,RIe20fbf8_4469,RIfc41d08_5771,RIe20cef8_4437,RIe20a1f8_4405,
        RIe2074f8_4373,RIfcd7510_7472,RIf166010_5620,RIfe9d230_8132,RIe2008b0_4296,RIf165098_5609,RIfc41ba0_5770,RIfc41a38_5769,RIfc92c30_6692,RIfc418d0_5768,
        RIfc79190_6400,RIe1fcad0_4252,RIfec4560_8354,RIfc79028_6399,RIfcbf258_7197,RIfcc1df0_7228,RIfcd81b8_7481,RIfc92d98_6693,RIfc5b4d8_6061,RIfcd77e0_7474,
        RIe1fa0a0_4222,RIf156188_5439,RIfe9d500_8134,RIf1546d0_5420,RIe1f5348_4167,RIfec4830_8356,RIfec46c8_8355,RIf1508f0_5376,RIe1f3020_4142,RIfce3180_7606,
        RIfce8fb8_7673,RIfcbf690_7200,RIe1edd28_4083,RIe1eb460_4054,RIe1e8760_4022,RIe1e5a60_3990,RIe1e2d60_3958,RIe1e0060_3926,RIe1dd360_3894,RIe1da660_3862,
        RIe1d7960_3830,RIe1d1f60_3766,RIe1cf260_3734,RIe1cc560_3702,RIe1c9860_3670,RIe1c6b60_3638,RIe1c3e60_3606,RIe1c1160_3574,RIe1be460_3542,RIfe9d0c8_8131,
        RIfe9cc90_8128,RIe1b9168_3483,RIe1b7110_3460,RIf14a3b0_5304,RIfe9cb28_8127,RIfe9cf60_8130,RIfe9c9c0_8126,RIfce2208_7595,RIfce9558_7677,RIfe9c858_8125,
        RIfe9cdf8_8129,RIf147110_5268,RIf146468_5259,RIe1ac2b0_3336,RIe1aaac8_3319,RIe1a87a0_3294,RIe1a5aa0_3262,RIe1a2da0_3230,RIe1a00a0_3198,RIe18c5a0_2974,
        RIe178aa0_2750,RIe2263f8_4725,RIe21aff8_4597,RIe2047f8_4341,RIe1fe858_4273,RIe1f7c10_4196,RIe1f0758_4113,RIe1d4c60_3798,RIe1bb760_3510,RIe1ae5d8_3361,
        RIe170c10_2660,RIdec4190_695,RIdec1490_663,RIfceaa70_7692,RIdebe790_631,RIfc954f8_6721,RIdebba90_599,RIdeb8d90_567,RIdeb6090_535,RIfcebb50_7704,
        RIdeb0690_471,RIee1e190_4801,RIdead990_439,RIfcdf0d0_7560,RIdea7978_407,RIdea1078_375,RIde9a778_343,RIee1c840_4783,RIfc957c8_6723,RIfcc8e70_7308,
        RIfc5e610_6096,RIfe9e8b0_8148,RIde8c1c8_273,RIde88028_253,RIde83b40_232,RIfcb0bb8_7033,RIfca4b10_6896,RIfc75d88_6363,RIfca4c78_6897,RIfc95390_6720,
        RIe16a9a0_2590,RIfcc8fd8_7309,RIe166e90_2548,RIe164190_2516,RIe161490_2484,RIfe9e748_8147,RIe15e790_2452,RIfc74f78_6353,RIe15ba90_2420,RIe156090_2356,
        RIe153390_2324,RIfc3ecc0_5740,RIe150690_2292,RIfce8b80_7670,RIe14d990_2260,RIfca6730_6916,RIe14ac90_2228,RIe147f90_2196,RIe145290_2164,RIfcee2b0_7732,
        RIfc5f2b8_6105,RIfc753b0_6356,RIfc74b40_6350,RIe140268_2107,RIdf3e170_2083,RIdf3be48_2058,RIdf39c88_2034,RIfcc1c88_7227,RIfcc1850_7224,RIfc965d8_6733,
        RIfc96038_6729,RIdf34828_1974,RIdf327d0_1951,RIdf301d8_1924,RIdf2e2e8_1902,RIfc5e778_6097,RIfcd0328_7391,RIfc757e8_6359,RIfcee6e8_7735,RIdf296f8_1848,
        RIdf273d0_1823,RIdf257b0_1803,RIdf23b90_1783,RIfc95d68_6727,RIfceda40_7726,RIfe9eb80_8150,RIfc75518_6357,RIfcd01c0_7390,RIdf1eb68_1726,RIfe9ece8_8151,
        RIfe9ea18_8149,RIdf15d60_1625,RIdf13060_1593,RIdf10360_1561,RIdf0d660_1529,RIdf0a960_1497,RIdf07c60_1465,RIdf04f60_1433,RIdf02260_1401,RIdefc860_1337,
        RIdef9b60_1305,RIdef6e60_1273,RIdef4160_1241,RIdef1460_1209,RIdeee760_1177,RIdeeba60_1145,RIdee8d60_1113,RIfc961a0_6730,RIfc96308_6731,RIfc5ee80_6102,
        RIfce6150_7640,RIdee42d8_1060,RIdee1e48_1034,RIdee00c0_1013,RIdeddac8_986,RIfc96470_6732,RIfc75248_6355,RIfc74ca8_6351,RIfcb0618_7029,RIded8938_928,
        RIded6610_903,RIded4450_879,RIded2290_855,RIdecf590_823,RIdecc890_791,RIdec9b90_759,RIdec6e90_727,RIdeb3390_503,RIde93e78_311,RIe16cf98_2617,
        RIe158d90_2388,RIe142590_2132,RIdf36f88_2002,RIdf2b5e8_1870,RIdf1be68_1694,RIdeff560_1369,RIdee6060_1081,RIdedadc8_954,RIde79dc0_184,RIe19c428_3155,
        RIe199728_3123,RIfe9e310_8144,RIe196a28_3091,RIfcc04a0_7210,RIe193d28_3059,RIe191028_3027,RIe18e328_2995,RIe188928_2931,RIe185c28_2899,RIfce1830_7588,
        RIe182f28_2867,RIfe9e478_8145,RIe180228_2835,RIe17d528_2803,RIe17a828_2771,RIf141878_5205,RIfcb12c0_7038,RIfc94418_6709,RIe174f90_2708,RIfc77408_6379,
        RIf13ea10_5172,RIfcdc100_7526,RIfc94580_6710,RIfc946e8_6711,RIfced338_7721,RIfce5fe8_7639,RIe172998_2681,RIfcdc268_7527,RIfcddff0_7548,RIfcc0608_7211,
        RIfce7230_7652,RIfc40340_5756,RIe222780_4682,RIfcdd618_7541,RIe21fa80_4650,RIfcd0b98_7397,RIe21cd80_4618,RIe217380_4554,RIe214680_4522,RIfec4998_8357,
        RIe211980_4490,RIf168608_5647,RIe20ec80_4458,RIfcc0770_7212,RIe20bf80_4426,RIe209280_4394,RIe206580_4362,RIfce2370_7596,RIfcee580_7734,RIfec4c68_8359,
        RIfec4b00_8358,RIfc949b8_6713,RIfcebcb8_7705,RIf162938_5581,RIf1612b8_5565,RIfccd088_7355,RIfcc08d8_7213,RIfe9e040_8142,RIfe9e1a8_8143,RIfcead40_7694,
        RIf15ad78_5493,RIfc94c88_6715,RIfccc3e0_7346,RIfc765f8_6369,RIfc94df0_6716,RIfcc0a40_7214,RIe1f9998_4217,RIfcc8d08_7307,RIfce8748_7667,RIfceb2e0_7698,
        RIe1f4970_4160,RIf152510_5396,RIf1512c8_5383,RIfcb0ff0_7036,RIe1f24e0_4134,RIfc761c0_6366,RIfc950c0_6718,RIfcc0e78_7217,RIe1ed1e8_4075,RIe1ea4e8_4043,
        RIe1e77e8_4011,RIe1e4ae8_3979,RIe1e1de8_3947,RIe1df0e8_3915,RIe1dc3e8_3883,RIe1d96e8_3851,RIe1d69e8_3819,RIe1d0fe8_3755,RIe1ce2e8_3723,RIe1cb5e8_3691,
        RIe1c88e8_3659,RIe1c5be8_3627,RIe1c2ee8_3595,RIe1c01e8_3563,RIe1bd4e8_3531,RIf14bfd0_5324,RIf14ac20_5310,RIfe9ded8_8141,RIe1b65d0_3452,RIfcecd98_7717,
        RIfc76490_6368,RIe1b4c80_3434,RIe1b38d0_3420,RIfcc0fe0_7218,RIfceaea8_7695,RIe1b1f80_3402,RIe1b0360_3382,RIfcd0760_7394,RIf145ec8_5255,RIfe9e5e0_8146,
        RIfe9dd70_8140,RIe1a7828_3283,RIe1a4b28_3251,RIe1a1e28_3219,RIe19f128_3187,RIe18b628_2963,RIe177b28_2739,RIe225480_4714,RIe21a080_4586,RIe203880_4330,
        RIe1fd8e0_4262,RIe1f6c98_4185,RIe1ef7e0_4102,RIe1d3ce8_3787,RIe1ba7e8_3499,RIe1ad660_3350,RIe16fc98_2649,RIdec6788_722,RIdec3a88_690,RIee20788_4828,
        RIdec0d88_658,RIee1f810_4817,RIdebe088_626,RIdebb388_594,RIdeb8688_562,RIfc9b1c8_6787,RIdeb2c88_498,RIfce1f38_7593,RIdeaff88_466,RIfc892e8_6583,
        RIdead210_434,RIdea6910_402,RIdea0010_370,RIee1d650_4793,RIee1c570_4781,RIee1b5f8_4770,RIee1aef0_4765,RIfe99888_8091,RIfe99450_8088,RIfe99720_8090,
        RIfe995b8_8089,RIde83168_229,RIfcc43e8_7255,RIfcd5a58_7453,RIfc89450_6584,RIfcc5798_7269,RIe16c890_2612,RIe16a568_2587,RIe168d80_2570,RIe166788_2543,
        RIe163a88_2511,RIfc83618_6517,RIe160d88_2479,RIee36718_5078,RIe15e088_2447,RIe158688_2383,RIe155988_2351,RIfc3f800_5748,RIe152c88_2319,RIfc895b8_6585,
        RIe14ff88_2287,RIfc51cf8_5953,RIe14d288_2255,RIe14a588_2223,RIe147888_2191,RIee34990_5057,RIee338b0_5045,RIfc831e0_6514,RIfcd3b68_7431,RIe141ff0_2128,
        RIe13fcc8_2103,RIdf3dbd0_2079,RIdf3b740_2053,RIfcb6f90_7104,RIee301d8_5006,RIfcba938_7145,RIee2e018_4982,RIdf369e8_1998,RIdf343f0_1971,RIdf32230_1947,
        RIfe99e28_8095,RIfc83078_6513,RIfcb6e28_7103,RIfc9ad90_6784,RIfcbad70_7148,RIdf2b1b0_1867,RIdf292c0_1845,RIfe99b58_8093,RIfe999f0_8092,RIfc9ac28_6783,
        RIfc4a9a8_5871,RIdf23758_1780,RIfc82da8_6511,RIdf220d8_1764,RIdf20a58_1748,RIdf1ba30_1691,RIfe99cc0_8094,RIdf18358_1652,RIdf15658_1620,RIdf12958_1588,
        RIdf0fc58_1556,RIdf0cf58_1524,RIdf0a258_1492,RIdf07558_1460,RIdf04858_1428,RIdefee58_1364,RIdefc158_1332,RIdef9458_1300,RIdef6758_1268,RIdef3a58_1236,
        RIdef0d58_1204,RIdeee058_1172,RIdeeb358_1140,RIee25918_4886,RIee24b08_4876,RIfc52568_5959,RIfc826a0_6506,RIdee5958_1076,RIdee3bd0_1055,RIfe99f90_8096,
        RIdedf9b8_1008,RIfce4800_7622,RIfc89b58_6589,RIfc9f3e0_6834,RIfc82538_6505,RIdeda828_950,RIded8398_924,RIfeabe70_8272,RIded3eb0_875,RIded1b88_850,
        RIdecee88_818,RIdecc188_786,RIdec9488_754,RIdeb5988_530,RIde99710_338,RIe16f590_2644,RIe15b388_2415,RIe144b88_2159,RIdf39580_2029,RIdf2dbe0_1897,
        RIdf1e460_1721,RIdf01b58_1396,RIdee8658_1108,RIdedd3c0_981,RIde7f658_211,RIe19ea20_3182,RIe19bd20_3150,RIf145928_5251,RIe199020_3118,RIfe98910_8080,
        RIe196320_3086,RIe193620_3054,RIe190920_3022,RIe18af20_2958,RIe188220_2926,RIf143e70_5232,RIe185520_2894,RIfc95c00_6726,RIe182820_2862,RIe17fb20_2830,
        RIe17ce20_2798,RIf142520_5214,RIf141440_5202,RIe1776f0_2736,RIfeab8d0_8268,RIfcc5bd0_7272,RIfc62dc8_6147,RIee3e710_5169,RIfc9cb18_6805,RIee3c820_5147,
        RIee3b470_5133,RIee3a390_5121,RIe174888_2703,RIf170498_5737,RIfc68660_6210,RIf16e878_5717,RIfc6ea38_6281,RIfe98d48_8083,RIe224d78_4709,RIf16c280_5690,
        RIe222078_4677,RIf16b308_5679,RIe21f378_4645,RIe219978_4581,RIe216c78_4549,RIf16a390_5668,RIe213f78_4517,RIf169b20_5662,RIe211278_4485,RIf1681d0_5644,
        RIe20e578_4453,RIe20b878_4421,RIe208b78_4389,RIfcd4ae0_7442,RIfc61478_6129,RIfeab060_8262,RIe201990_4308,RIfc70ec8_6307,RIfc70928_6303,RIfcec528_7711,
        RIfcbe880_7190,RIf160d18_5561,RIf15ee28_5539,RIfe98be0_8082,RIfe98eb0_8084,RIf15d0a0_5518,RIf15bcf0_5504,RIfcd4540_7438,RIf159e00_5482,RIf1592c0_5474,
        RIf158078_5461,RIfca3a30_6884,RIfea7988_8223,RIf156728_5443,RIf155be8_5435,RIf154b08_5423,RIfe98a78_8081,RIf1538c0_5410,RIf1520d8_5393,RIf150e90_5380,
        RIe1f43d0_4156,RIf14fdb0_5368,RIfcd2380_7414,RIf14e2f8_5349,RIe1ef240_4098,RIe1ecae0_4070,RIe1e9de0_4038,RIe1e70e0_4006,RIe1e43e0_3974,RIe1e16e0_3942,
        RIe1de9e0_3910,RIe1dbce0_3878,RIe1d8fe0_3846,RIe1d35e0_3782,RIe1d08e0_3750,RIe1cdbe0_3718,RIe1caee0_3686,RIe1c81e0_3654,RIe1c54e0_3622,RIe1c27e0_3590,
        RIe1bfae0_3558,RIfc44b70_5804,RIf14bd00_5322,RIfe992e8_8087,RIfe987a8_8079,RIf14a950_5308,RIf149f78_5301,RIfe99180_8086,RIfe98640_8078,RIf149438_5293,
        RIfcec7f8_7713,RIfe984d8_8077,RIe1b1b48_3399,RIfc4b650_5880,RIfcda918_7509,RIfe98370_8076,RIfe99018_8085,RIe1a9e20_3310,RIe1a7120_3278,RIe1a4420_3246,
        RIe1a1720_3214,RIe18dc20_2990,RIe17a120_2766,RIe227a78_4741,RIe21c678_4613,RIe205e78_4357,RIe1ffed8_4289,RIe1f9290_4212,RIe1f1dd8_4129,RIe1d62e0_3814,
        RIe1bcde0_3526,RIe1afc58_3377,RIe172290_2676,RIdec6620_721,RIdec3920_689,RIfc49328_5855,RIdec0c20_657,RIfc80eb8_6489,RIdebdf20_625,RIdebb220_593,
        RIdeb8520_561,RIfc80648_6483,RIdeb2b20_497,RIfc8b340_6606,RIdeafe20_465,RIfc491c0_5854,RIdeacec8_433,RIdea65c8_401,RIde9fcc8_369,RIfcd9c70_7500,
        RIfe98208_8075,RIfce4698_7621,RIfe980a0_8074,RIde93158_307,RIde8f648_289,RIde8b4a8_269,RIde87308_249,RIde82e20_228,RIfcbba18_7157,RIfc48d88_5851,
        RIfc99f80_6774,RIfc8b4a8_6607,RIe16c728_2611,RIe16a400_2586,RIe168c18_2569,RIe166620_2542,RIe163920_2510,RIee38068_5096,RIe160c20_2478,RIfc48248_5843,
        RIe15df20_2446,RIe158520_2382,RIe155820_2350,RIfcbbe50_7160,RIe152b20_2318,RIfc47e10_5840,RIe14fe20_2286,RIfca0e98_6853,RIe14d120_2254,RIe14a420_2222,
        RIe147720_2190,RIfc8be80_6614,RIfc7fb08_6475,RIfc480e0_5842,RIfc99878_6769,RIe141e88_2127,RIe13fb60_2102,RIdf3da68_2078,RIdf3b5d8_2052,RIfe97f38_8073,
        RIee30070_5005,RIee2eb58_4990,RIee2deb0_4981,RIdf36880_1997,RIdf34288_1970,RIdf320c8_1946,RIfe97dd0_8072,RIfcc3740_7246,RIfc48ab8_5849,RIfce05e8_7575,
        RIfc80210_6480,RIdf2b048_1866,RIdf29158_1844,RIdf26f98_1820,RIdf254e0_1801,RIfc8bbb0_6612,RIfc48950_5848,RIdf235f0_1779,RIfc8bd18_6613,RIdf21f70_1763,
        RIdf208f0_1747,RIdf1b8c8_1690,RIdf1a3b0_1675,RIdf181f0_1651,RIdf154f0_1619,RIdf127f0_1587,RIdf0faf0_1555,RIdf0cdf0_1523,RIdf0a0f0_1491,RIdf073f0_1459,
        RIdf046f0_1427,RIdefecf0_1363,RIdefbff0_1331,RIdef92f0_1299,RIdef65f0_1267,RIdef38f0_1235,RIdef0bf0_1203,RIdeedef0_1171,RIdeeb1f0_1139,RIfcbc120_7162,
        RIfcd9838_7497,RIfc99710_6768,RIfca1168_6855,RIdee57f0_1075,RIdee3a68_1054,RIdee18a8_1030,RIdedf850_1007,RIfc549f8_5985,RIfcb5370_7084,RIfce43c8_7619,
        RIfce0480_7574,RIdeda6c0_949,RIded8230_923,RIded6070_899,RIded3d48_874,RIded1a20_849,RIdeced20_817,RIdecc020_785,RIdec9320_753,RIdeb5820_529,
        RIde993c8_337,RIe16f428_2643,RIe15b220_2414,RIe144a20_2158,RIdf39418_2028,RIdf2da78_1896,RIdf1e2f8_1720,RIdf019f0_1395,RIdee84f0_1107,RIdedd258_980,
        RIde7f310_210,RIe19e8b8_3181,RIe19bbb8_3149,RIfe976c8_8067,RIe198eb8_3117,RIf144c80_5242,RIe1961b8_3085,RIe1934b8_3053,RIe1907b8_3021,RIe18adb8_2957,
        RIe1880b8_2925,RIfe97560_8066,RIe1853b8_2893,RIfcc3fb0_7252,RIe1826b8_2861,RIe17f9b8_2829,RIe17ccb8_2797,RIfcd3730_7428,RIf1412d8_5201,RIfcc4118_7253,
        RIfe97830_8068,RIfc4a6d8_5869,RIf13f6b8_5181,RIfc9f980_6838,RIfc9fae8_6839,RIfcc3e48_7251,RIfc89e28_6591,RIfc89cc0_6590,RIe174720_2702,RIfc4a408_5867,
        RIfce27a8_7599,RIfc530a8_5967,RIfcd5d28_7455,RIf16cf28_5699,RIe224c10_4708,RIfc53210_5968,RIe221f10_4676,RIf16b1a0_5678,RIe21f210_4644,RIe219810_4580,
        RIe216b10_4548,RIfc401d8_5755,RIe213e10_4516,RIf1699b8_5661,RIe211110_4484,RIfc81cc8_6499,RIe20e410_4452,RIe20b710_4420,RIe208a10_4388,RIfc8a0f8_6593,
        RIfcb6720_7098,RIe203448_4327,RIe201828_4307,RIfc53378_5969,RIfc8a3c8_6595,RIfcb65b8_7097,RIfc49fd0_5864,RIf160bb0_5560,RIf15ecc0_5538,RIe1fd4a8_4259,
        RIfe97b00_8070,RIfc8a530_6596,RIfe97c68_8071,RIfc8a800_6598,RIfc8a698_6597,RIfc9a7f0_6780,RIfc81890_6496,RIfcd5e90_7456,RIe1fb180_4234,RIfc49e68_5863,
        RIfc81728_6495,RIfcbb1a8_7151,RIe1f66f8_4181,RIfcd3460_7426,RIfcb62e8_7095,RIfc9a520_6778,RIe1f4268_4155,RIfc49d00_5862,RIfcd9dd8_7501,RIfcbb310_7152,
        RIe1ef0d8_4097,RIe1ec978_4069,RIe1e9c78_4037,RIe1e6f78_4005,RIe1e4278_3973,RIe1e1578_3941,RIe1de878_3909,RIe1dbb78_3877,RIe1d8e78_3845,RIe1d3478_3781,
        RIe1d0778_3749,RIe1cda78_3717,RIe1cad78_3685,RIe1c8078_3653,RIe1c5378_3621,RIe1c2678_3589,RIe1bf978_3557,RIfc49a30_5860,RIfcb6018_7093,RIe1ba3b0_3496,
        RIe1b81f0_3472,RIfce0a20_7578,RIfcbb5e0_7154,RIe1b6030_3448,RIfe97998_8069,RIfce5610_7632,RIfcc3a10_7248,RIe1b3330_3416,RIe1b19e0_3398,RIfc495f8_5857,
        RIfc81188_6491,RIe1ad228_3347,RIe1aba40_3330,RIe1a9cb8_3309,RIe1a6fb8_3277,RIe1a42b8_3245,RIe1a15b8_3213,RIe18dab8_2989,RIe179fb8_2765,RIe227910_4740,
        RIe21c510_4612,RIe205d10_4356,RIe1ffd70_4288,RIe1f9128_4211,RIe1f1c70_4128,RIe1d6178_3813,RIe1bcc78_3525,RIe1afaf0_3376,RIe172128_2675,RIdec6a58_724,
        RIdec3d58_692,RIfc723e0_6322,RIdec1058_660,RIfc59fc0_6046,RIdebe358_628,RIdebb658_596,RIdeb8958_564,RIfcb96f0_7132,RIdeb2f58_500,RIfce1c68_7591,
        RIdeb0258_468,RIfc9b498_6789,RIdead558_436,RIdea6fa0_404,RIdea06a0_372,RIfc81458_6493,RIfc83780_6518,RIfc4e620_5914,RIfcd3e38_7433,RIde937e8_309,
        RIde8f990_290,RIde8bb38_271,RIde87650_250,RIde834b0_230,RIfc42c80_5782,RIfc65960_6178,RIfc6c710_6256,RIee392b0_5109,RIe16cb60_2614,RIe16a6d0_2588,
        RIe169050_2572,RIe166a58_2545,RIe163d58_2513,RIfec3cf0_8348,RIe161058_2481,RIfcd54b8_7449,RIe15e358_2449,RIe158958_2385,RIe155c58_2353,RIfe9ba48_8115,
        RIe152f58_2321,RIfec4128_8351,RIe150258_2289,RIfcb9b28_7135,RIe14d558_2257,RIe14a858_2225,RIe147b58_2193,RIfcdb2f0_7516,RIfc553d0_5992,RIfc9a0e8_6775,
        RIfcbd908_7179,RIe1422c0_2130,RIe13ff98_2105,RIdf3dea0_2081,RIdf3ba10_2055,RIfc87128_6559,RIee304a8_5008,RIfcc51f8_7265,RIee2e2e8_4984,RIdf36cb8_2000,
        RIfec3fc0_8350,RIdf32500_1949,RIfec3e58_8349,RIee2c830_4965,RIee2ad78_4946,RIee296f8_4930,RIee284b0_4917,RIfe9b8e0_8114,RIfe9b610_8112,RIfe9b778_8113,
        RIfe9b4a8_8111,RIfcb7c38_7113,RIfc86b88_6555,RIdf238c0_1781,RIfc75ab8_6361,RIdf22240_1765,RIfeaa3b8_8253,RIdf1bb98_1692,RIdf1a680_1677,RIdf18628_1654,
        RIdf15928_1622,RIdf12c28_1590,RIdf0ff28_1558,RIdf0d228_1526,RIdf0a528_1494,RIdf07828_1462,RIdf04b28_1430,RIdeff128_1366,RIdefc428_1334,RIdef9728_1302,
        RIdef6a28_1270,RIdef3d28_1238,RIdef1028_1206,RIdeee328_1174,RIdeeb628_1142,RIee25a80_4887,RIee24c70_4877,RIfcddd20_7546,RIfccc110_7344,RIdee5c28_1078,
        RIdee3ea0_1057,RIdee1b78_1032,RIdedfc88_1010,RIfc6a6b8_6233,RIee227e0_4851,RIfc88be0_6578,RIee21868_4840,RIdedaaf8_952,RIded8668_926,RIded6340_901,
        RIded4180_877,RIded1e58_852,RIdecf158_820,RIdecc458_788,RIdec9758_756,RIdeb5c58_532,RIde99da0_340,RIe16f860_2646,RIe15b658_2417,RIe144e58_2161,
        RIdf39850_2031,RIdf2deb0_1899,RIdf1e730_1723,RIdf01e28_1398,RIdee8928_1110,RIdedd690_983,RIde7fce8_213,RIe19ecf0_3184,RIe19bff0_3152,RIf145a90_5252,
        RIe1992f0_3120,RIf144de8_5243,RIe1965f0_3088,RIe1938f0_3056,RIe190bf0_3024,RIe18b1f0_2960,RIe1884f0_2928,RIfc72980_6326,RIe1857f0_2896,RIf143060_5222,
        RIe182af0_2864,RIe17fdf0_2832,RIe17d0f0_2800,RIf142688_5215,RIf141710_5204,RIe177858_2737,RIe176778_2725,RIfcea638_7689,RIfca54e8_6903,RIee3e878_5170,
        RIee3dbd0_5161,RIee3c988_5148,RIee3b5d8_5134,RIee3a4f8_5122,RIe174b58_2705,RIf170600_5738,RIfc76fd0_6376,RIf16e9e0_5718,RIfced608_7723,RIf16d090_5700,
        RIe225048_4711,RIf16c550_5692,RIe222348_4679,RIf16b470_5680,RIe21f648_4647,RIe219c48_4583,RIe216f48_4551,RIf16a4f8_5669,RIe214248_4519,RIf169df0_5664,
        RIe211548_4487,RIf1684a0_5646,RIe20e848_4455,RIe20bb48_4423,RIe208e48_4391,RIf1673c0_5634,RIf166448_5623,RIfe9c6f0_8124,RIfe9c150_8120,RIf1654d0_5612,
        RIfcc4550_7256,RIf1635e0_5590,RIf162500_5578,RIf160fe8_5563,RIf15f0f8_5541,RIfe9bfe8_8119,RIfe9c588_8123,RIf15d208_5519,RIf15bfc0_5506,RIfc4d540_5902,
        RIfc9c848_6803,RIfec4290_8352,RIfe9c2b8_8121,RIfcc01d0_7208,RIe1fb2e8_4235,RIfe9c420_8122,RIfca3e68_6887,RIf154c70_5424,RIe1f69c8_4183,RIf153a28_5411,
        RIf152240_5394,RIf150ff8_5381,RIe1f46a0_4158,RIfca6028_6911,RIfc43bf8_5793,RIf14e460_5350,RIe1ef3a8_4099,RIe1ecdb0_4072,RIe1ea0b0_4040,RIe1e73b0_4008,
        RIe1e46b0_3976,RIe1e19b0_3944,RIe1decb0_3912,RIe1dbfb0_3880,RIe1d92b0_3848,RIe1d38b0_3784,RIe1d0bb0_3752,RIe1cdeb0_3720,RIe1cb1b0_3688,RIe1c84b0_3656,
        RIe1c57b0_3624,RIe1c2ab0_3592,RIe1bfdb0_3560,RIfc4d6a8_5903,RIf14be68_5323,RIe1ba680_3498,RIfe9be80_8118,RIfc86e58_6557,RIfcd46a8_7439,RIe1b6300_3450,
        RIfe9bd18_8117,RIf1495a0_5294,RIf1481f0_5280,RIe1b3600_3418,RIe1b1e18_3401,RIfc69470_6220,RIfcbfac8_7203,RIfe9bbb0_8116,RIe1abd10_3332,RIe1aa0f0_3312,
        RIe1a73f0_3280,RIe1a46f0_3248,RIe1a19f0_3216,RIe18def0_2992,RIe17a3f0_2768,RIe227d48_4743,RIe21c948_4615,RIe206148_4359,RIe2001a8_4291,RIe1f9560_4214,
        RIe1f20a8_4131,RIe1d65b0_3816,RIe1bd0b0_3528,RIe1aff28_3379,RIe172560_2678,RIdec68f0_723,RIdec3bf0_691,RIee208f0_4829,RIdec0ef0_659,RIfc7ce08_6443,
        RIdebe1f0_627,RIdebb4f0_595,RIdeb87f0_563,RIfc9b8d0_6792,RIdeb2df0_499,RIfcc6710_7280,RIdeb00f0_467,RIfc5ff60_6114,RIdead3f0_435,RIdea6c58_403,
        RIdea0358_371,RIfce5070_7628,RIee1c6d8_4782,RIfce70c8_7651,RIee1b058_4766,RIde934a0_308,RIfe9b1d8_8109,RIde8b7f0_270,RIfe9b340_8110,RIfc6b798_6245,
        RIfcb2238_7049,RIfcd3a00_7430,RIfcdb020_7514,RIfc511b8_5945,RIe16c9f8_2613,RIfcb27d8_7053,RIe168ee8_2571,RIe1668f0_2544,RIe163bf0_2512,RIee381d0_5097,
        RIe160ef0_2480,RIfcdfaa8_7567,RIe15e1f0_2448,RIe1587f0_2384,RIe155af0_2352,RIfc3f968_5749,RIe152df0_2320,RIfcd5080_7446,RIe1500f0_2288,RIfc84b30_6532,
        RIe14d3f0_2256,RIe14a6f0_2224,RIe1479f0_2192,RIfcea098_7685,RIfc92f00_6694,RIfc54890_5984,RIfcdcc40_7534,RIe142158_2129,RIe13fe30_2104,RIdf3dd38_2080,
        RIdf3b8a8_2054,RIfc57590_6016,RIee30340_5007,RIfcd0490_7392,RIee2e180_4983,RIdf36b50_1999,RIdf34558_1972,RIdf32398_1948,RIfe9b070_8108,RIfcb1860_7042,
        RIfca1b40_6862,RIfc5c018_6069,RIfe9ada0_8106,RIdf2b318_1868,RIdf29428_1846,RIdf27100_1821,RIfe9af08_8107,RIfc5e1d8_6093,RIfcdcda8_7535,RIfcac400_6982,
        RIfc691a0_6218,RIfcaad80_6966,RIdf20bc0_1749,RIfc61b80_6134,RIdf1a518_1676,RIdf184c0_1653,RIdf157c0_1621,RIdf12ac0_1589,RIdf0fdc0_1557,RIdf0d0c0_1525,
        RIdf0a3c0_1493,RIdf076c0_1461,RIdf049c0_1429,RIdefefc0_1365,RIdefc2c0_1333,RIdef95c0_1301,RIdef68c0_1269,RIdef3bc0_1237,RIdef0ec0_1205,RIdeee1c0_1173,
        RIdeeb4c0_1141,RIfc69b78_6225,RIfc6b900_6246,RIfc4d270_5900,RIfced770_7724,RIdee5ac0_1077,RIdee3d38_1056,RIdee1a10_1031,RIdedfb20_1009,RIfc7ff40_6478,
        RIfca4408_6891,RIfcb5640_7086,RIee21700_4839,RIdeda990_951,RIded8500_925,RIded61d8_900,RIded4018_876,RIded1cf0_851,RIdeceff0_819,RIdecc2f0_787,
        RIdec95f0_755,RIdeb5af0_531,RIde99a58_339,RIe16f6f8_2645,RIe15b4f0_2416,RIe144cf0_2160,RIdf396e8_2030,RIdf2dd48_1898,RIdf1e5c8_1722,RIdf01cc0_1397,
        RIdee87c0_1109,RIdedd528_982,RIde7f9a0_212,RIe19eb88_3183,RIe19be88_3151,RIfe9a698_8101,RIe199188_3119,RIfe9a530_8100,RIe196488_3087,RIe193788_3055,
        RIe190a88_3023,RIe18b088_2959,RIe188388_2927,RIfe9a800_8102,RIe185688_2895,RIfc8d938_6633,RIe182988_2863,RIe17fc88_2831,RIe17cf88_2799,RIfe9a3c8_8099,
        RIf1415a8_5203,RIfe9a260_8098,RIfe9a0f8_8097,RIfcb9150_7128,RIf13f820_5182,RIfc9fc50_6840,RIfce5340_7630,RIfc5cb58_6077,RIfc576f8_6017,RIfc780b0_6388,
        RIe1749f0_2704,RIfc7adb0_6420,RIfc7c2c8_6435,RIfcb2d78_7057,RIfc7e758_6461,RIfe9aad0_8104,RIe224ee0_4710,RIf16c3e8_5691,RIe2221e0_4678,RIfcd3898_7429,
        RIe21f4e0_4646,RIe219ae0_4582,RIe216de0_4550,RIfc880a0_6570,RIe2140e0_4518,RIf169c88_5663,RIe2113e0_4486,RIf168338_5645,RIe20e6e0_4454,RIe20b9e0_4422,
        RIe208ce0_4390,RIfce4c38_7625,RIfc9c6e0_6802,RIe2035b0_4328,RIe201af8_4309,RIfc500d8_5933,RIfc85c10_6544,RIfce81a8_7663,RIfce9c60_7682,RIf160e80_5562,
        RIf15ef90_5540,RIfe9a968_8103,RIfe9ac38_8105,RIfca8d28_6943,RIf15be58_5505,RIfcedba8_7727,RIfc6a988_6235,RIfc71cd8_6317,RIfccb198_7333,RIfcaa3a8_6959,
        RIfec3b88_8347,RIfc4c730_5892,RIfc6d688_6267,RIfca8e90_6944,RIe1f6860_4182,RIfc64e20_6170,RIfcaee30_7012,RIfccee10_7376,RIe1f4538_4157,RIfc63ea8_6159,
        RIfcaecc8_7011,RIfcae458_7005,RIfeab1c8_8263,RIe1ecc48_4071,RIe1e9f48_4039,RIe1e7248_4007,RIe1e4548_3975,RIe1e1848_3943,RIe1deb48_3911,RIe1dbe48_3879,
        RIe1d9148_3847,RIe1d3748_3783,RIe1d0a48_3751,RIe1cdd48_3719,RIe1cb048_3687,RIe1c8348_3655,RIe1c5648_3623,RIe1c2948_3591,RIe1bfc48_3559,RIfcc70e8_7287,
        RIfca7ae0_6930,RIe1ba518_3497,RIe1b8358_3473,RIfc598b8_6041,RIfcc2228_7231,RIe1b6198_3449,RIe1b4848_3431,RIfc82f10_6512,RIfc55970_5996,RIe1b3498_3417,
        RIe1b1cb0_3400,RIfcb7698_7109,RIfc4b4e8_5879,RIe1ad390_3348,RIe1abba8_3331,RIe1a9f88_3311,RIe1a7288_3279,RIe1a4588_3247,RIe1a1888_3215,RIe18dd88_2991,
        RIe17a288_2767,RIe227be0_4742,RIe21c7e0_4614,RIe205fe0_4358,RIe200040_4290,RIe1f93f8_4213,RIe1f1f40_4130,RIe1d6448_3815,RIe1bcf48_3527,RIe1afdc0_3378,
        RIe1723f8_2677,RIdec6d28_726,RIdec4028_694,RIee20bc0_4831,RIdec1328_662,RIfcbaed8_7149,RIdebe628_630,RIdebb928_598,RIdeb8c28_566,RIfc412b8_5767,
        RIdeb3228_502,RIfc9ea08_6827,RIdeb0528_470,RIee1e028_4800,RIdead828_438,RIdea7630_406,RIdea0d30_374,RIfcbac08_7147,RIfc55538_5993,RIfcba668_7143,
        RIfc4af48_5875,RIfe912f0_7996,RIfe91458_7997,RIde8be80_272,RIde87ce0_252,RIfc85238_6537,RIfc88640_6574,RIfcda210_7504,RIfcd5788_7451,RIee39418_5110,
        RIe16ce30_2616,RIfc884d8_6573,RIe169320_2574,RIe166d28_2547,RIe164028_2515,RIfe90918_7989,RIe161328_2483,RIee36880_5079,RIe15e628_2451,RIe158c28_2387,
        RIe155f28_2355,RIfe91188_7995,RIe153228_2323,RIfe91020_7994,RIe150528_2291,RIfcda378_7505,RIe14d828_2259,RIe14ab28_2227,RIe147e28_2195,RIfe90eb8_7993,
        RIfe90d50_7992,RIfcb99c0_7134,RIfc9c2a8_6799,RIfe90be8_7991,RIfe90a80_7990,RIdf3e008_2082,RIdf3bce0_2057,RIfcec690_7712,RIee30778_5010,RIfc87dd0_6568,
        RIee2e5b8_4986,RIdf36e20_2001,RIdf346c0_1973,RIdf32668_1950,RIdf30070_1923,RIee2c998_4966,RIee2aee0_4947,RIee299c8_4932,RIee28618_4918,RIfe90378_7985,
        RIfe907b0_7988,RIfe904e0_7986,RIfe90648_7987,RIfc9d928_6815,RIfc86048_6547,RIfcb92b8_7129,RIfc4ee90_5920,RIfc86a20_6554,RIdf20e90_1751,RIfcb8fe8_7127,
        RIdf1a950_1679,RIdf188f8_1656,RIdf15bf8_1624,RIdf12ef8_1592,RIdf101f8_1560,RIdf0d4f8_1528,RIdf0a7f8_1496,RIdf07af8_1464,RIdf04df8_1432,RIdeff3f8_1368,
        RIdefc6f8_1336,RIdef99f8_1304,RIdef6cf8_1272,RIdef3ff8_1240,RIdef12f8_1208,RIdeee5f8_1176,RIdeeb8f8_1144,RIfc857d8_6541,RIee24dd8_4878,RIfc4ff70_5932,
        RIfc50240_5934,RIdee5ef8_1080,RIdee4170_1059,RIfe915c0_7998,RIdedff58_1012,RIfcd4810_7440,RIee22948_4852,RIfce1560_7586,RIee219d0_4841,RIdedac60_953,
        RIfe91728_7999,RIded64a8_902,RIfe91890_8000,RIded2128_854,RIdecf428_822,RIdecc728_790,RIdec9a28_758,RIdeb5f28_534,RIde9a430_342,RIe16fb30_2648,
        RIe15b928_2419,RIe145128_2163,RIdf39b20_2033,RIdf2e180_1901,RIdf1ea00_1725,RIdf020f8_1400,RIdee8bf8_1112,RIdedd960_985,RIde80378_215,RIe19efc0_3186,
        RIe19c2c0_3154,RIf145d60_5254,RIe1995c0_3122,RIfc637a0_6154,RIe1968c0_3090,RIe193bc0_3058,RIe190ec0_3026,RIe18b4c0_2962,RIe1887c0_2930,RIfc62af8_6145,
        RIe185ac0_2898,RIfe8fc70_7980,RIe182dc0_2866,RIe1800c0_2834,RIe17d3c0_2802,RIfe90210_7984,RIfe8ff40_7982,RIfc72f20_6330,RIe176a48_2727,RIfcaf6a0_7018,
        RIfc61040_6126,RIf13e8a8_5171,RIfe900a8_7983,RIee3caf0_5149,RIee3b740_5135,RIee3a660_5123,RIe174e28_2707,RIf170768_5739,RIfc5fdf8_6113,RIf16eb48_5719,
        RIfcaaab0_6964,RIf16d1f8_5701,RIe225318_4713,RIf16c6b8_5693,RIe222618_4681,RIf16b5d8_5681,RIe21f918_4649,RIe219f18_4585,RIe217218_4553,RIfca62f8_6913,
        RIe214518_4521,RIfcc9578_7313,RIe211818_4489,RIfca5a88_6907,RIe20eb18_4457,RIe20be18_4425,RIe209118_4393,RIf167690_5636,RIf166718_5625,RIfe8f9a0_7978,
        RIfe8f838_7977,RIf165638_5613,RIf164990_5604,RIf1638b0_5592,RIf1627d0_5580,RIf161150_5564,RIf15f260_5542,RIe1fd778_4261,RIe1fc530_4248,RIf15d4d8_5521,
        RIf15c290_5508,RIfca20e0_6866,RIf159f68_5483,RIf159428_5475,RIf1581e0_5462,RIfc5ebb0_6100,RIfe8fdd8_7981,RIfc69e48_6227,RIfc5e8e0_6098,RIf154f40_5426,
        RIe1f6b30_4184,RIf153b90_5412,RIf1523a8_5395,RIfce88b0_7668,RIfe8fb08_7979,RIfcebe20_7706,RIfcb1158_7037,RIf14e730_5352,RIe1ef678_4101,RIe1ed080_4074,
        RIe1ea380_4042,RIe1e7680_4010,RIe1e4980_3978,RIe1e1c80_3946,RIe1def80_3914,RIe1dc280_3882,RIe1d9580_3850,RIe1d3b80_3786,RIe1d0e80_3754,RIe1ce180_3722,
        RIe1cb480_3690,RIe1c8780_3658,RIe1c5a80_3626,RIe1c2d80_3594,RIe1c0080_3562,RIfcc8ba0_7306,RIfc5d698_6085,RIfec35e8_8343,RIfeabd08_8271,RIfc5cf90_6080,
        RIfc5ce28_6079,RIfec31b0_8340,RIe1b4b18_3433,RIf149708_5295,RIf148358_5281,RIe1b3768_3419,RIfec3480_8342,RIfc483b0_5844,RIfc80be8_6487,RIe1ad4f8_3349,
        RIfec3318_8341,RIe1aa3c0_3314,RIe1a76c0_3282,RIe1a49c0_3250,RIe1a1cc0_3218,RIe18e1c0_2994,RIe17a6c0_2770,RIe228018_4745,RIe21cc18_4617,RIe206418_4361,
        RIe200478_4293,RIe1f9830_4216,RIe1f2378_4133,RIe1d6880_3818,RIe1bd380_3530,RIe1b01f8_3381,RIe172830_2680,RIdec6bc0_725,RIdec3ec0_693,RIee20a58_4830,
        RIdec11c0_661,RIee1f978_4818,RIdebe4c0_629,RIdebb7c0_597,RIdeb8ac0_565,RIee1efa0_4811,RIdeb30c0_501,RIfcb04b0_7028,RIdeb03c0_469,RIfc5e4a8_6095,
        RIdead6c0_437,RIdea72e8_405,RIdea09e8_373,RIfcb2508_7051,RIfcd16d8_7405,RIfc5d800_6086,RIfc63d40_6158,RIde93b30_310,RIfea7820_8222,RIfea73e8_8219,
        RIde87998_251,RIde837f8_231,RIfc7bd28_6431,RIfcc7ef8_7297,RIfc7a108_6411,RIfc7a6a8_6415,RIe16ccc8_2615,RIe16a838_2589,RIe1691b8_2573,RIe166bc0_2546,
        RIe163ec0_2514,RIee38338_5098,RIe1611c0_2482,RIfc54b60_5986,RIe15e4c0_2450,RIe158ac0_2386,RIe155dc0_2354,RIee35a70_5069,RIe1530c0_2322,RIee357a0_5067,
        RIe1503c0_2290,RIfc9fdb8_6841,RIe14d6c0_2258,RIe14a9c0_2226,RIe147cc0_2194,RIee34af8_5058,RIee33a18_5046,RIee327d0_5033,RIfcbcf30_7172,RIe142428_2131,
        RIe140100_2106,RIfea7280_8218,RIdf3bb78_2056,RIfc731f0_6332,RIee30610_5009,RIfcbe010_7184,RIee2e450_4985,RIfec2ee0_8338,RIfec3048_8339,RIfec2c10_8336,
        RIfec2d78_8337,RIfcb46c8_7075,RIfcb4830_7076,RIee29860_4931,RIfcb88e0_7122,RIdf2b480_1869,RIdf29590_1847,RIdf27268_1822,RIdf25648_1802,RIfcc9de8_7319,
        RIfc53648_5971,RIdf23a28_1782,RIfc823d0_6504,RIdf223a8_1766,RIdf20d28_1750,RIdf1bd00_1693,RIdf1a7e8_1678,RIdf18790_1655,RIdf15a90_1623,RIdf12d90_1591,
        RIdf10090_1559,RIdf0d390_1527,RIdf0a690_1495,RIdf07990_1463,RIdf04c90_1431,RIdeff290_1367,RIdefc590_1335,RIdef9890_1303,RIdef6b90_1271,RIdef3e90_1239,
        RIdef1190_1207,RIdeee490_1175,RIdeeb790_1143,RIee25be8_4888,RIfc6af28_6239,RIee23fc8_4868,RIfccf680_7382,RIdee5d90_1079,RIdee4008_1058,RIdee1ce0_1033,
        RIdedfdf0_1011,RIfc6b090_6240,RIfc534e0_5970,RIfca5920_6906,RIfc66770_6188,RIfe8f6d0_7976,RIded87d0_927,RIfe8f568_7975,RIded42e8_878,RIded1fc0_853,
        RIdecf2c0_821,RIdecc5c0_789,RIdec98c0_757,RIdeb5dc0_533,RIde9a0e8_341,RIe16f9c8_2647,RIe15b7c0_2418,RIe144fc0_2162,RIdf399b8_2032,RIdf2e018_1900,
        RIdf1e898_1724,RIdf01f90_1399,RIdee8a90_1111,RIdedd7f8_984,RIde80030_214,RIe19ee58_3185,RIe19c158_3153,RIf145bf8_5253,RIe199458_3121,RIfe8f298_7973,
        RIe196758_3089,RIe193a58_3057,RIe190d58_3025,RIe18b358_2961,RIe188658_2929,RIfe8f130_7972,RIe185958_2897,RIfc9f278_6833,RIe182c58_2865,RIe17ff58_2833,
        RIe17d258_2801,RIf1427f0_5216,RIfe8efc8_7971,RIe1779c0_2738,RIe1768e0_2726,RIfc81e30_6500,RIfc9ff20_6842,RIfca0088_6843,RIfc81b60_6498,RIfce5778_7633,
        RIfce08b8_7577,RIfc815c0_6494,RIe174cc0_2706,RIfca04c0_6846,RIfc53eb8_5977,RIfcc65a8_7279,RIfc80d50_6488,RIfc804e0_6482,RIe2251b0_4712,RIfc80378_6481,
        RIe2224b0_4680,RIfcb5910_7088,RIe21f7b0_4648,RIe219db0_4584,RIe2170b0_4552,RIfca01f0_6844,RIe2143b0_4520,RIfc82c40_6510,RIe2116b0_4488,RIfc7f6d0_6472,
        RIe20e9b0_4456,RIe20bcb0_4424,RIe208fb0_4392,RIf167528_5635,RIf1665b0_5624,RIe203718_4329,RIe201c60_4310,RIfc9da90_6816,RIfcc5360_7266,RIf163748_5591,
        RIf162668_5579,RIfc7e320_6458,RIfc87998_6565,RIe1fd610_4260,RIe1fc3c8_4247,RIf15d370_5520,RIf15c128_5507,RIfcc5d38_7273,RIfce7d70_7660,RIfc4bd58_5885,
        RIfc55c40_5998,RIfca2ab8_6873,RIe1fb450_4236,RIf156890_5444,RIfcd5ff8_7457,RIf154dd8_5425,RIfec2aa8_8335,RIfcb4b00_7078,RIfcd9400_7494,RIf151160_5382,
        RIe1f4808_4159,RIfc44738_5801,RIfc90908_6667,RIf14e5c8_5351,RIe1ef510_4100,RIe1ecf18_4073,RIe1ea218_4041,RIe1e7518_4009,RIe1e4818_3977,RIe1e1b18_3945,
        RIe1dee18_3913,RIe1dc118_3881,RIe1d9418_3849,RIe1d3a18_3785,RIe1d0d18_3753,RIe1ce018_3721,RIe1cb318_3689,RIe1c8618_3657,RIe1c5918_3625,RIe1c2c18_3593,
        RIe1bff18_3561,RIf14d218_5337,RIfe8ee60_7970,RIfea8090_8228,RIe1b84c0_3474,RIf14aab8_5309,RIfc6c170_6252,RIe1b6468_3451,RIe1b49b0_3432,RIfcafad8_7021,
        RIfcaa948_6963,RIfe8ecf8_7969,RIfe8f400_7974,RIfc67f58_6205,RIfca8ff8_6945,RIfe8eb90_7968,RIe1abe78_3333,RIe1aa258_3313,RIe1a7558_3281,RIe1a4858_3249,
        RIe1a1b58_3217,RIe18e058_2993,RIe17a558_2769,RIe227eb0_4744,RIe21cab0_4616,RIe2062b0_4360,RIe200310_4292,RIe1f96c8_4215,RIe1f2210_4132,RIe1d6718_3817,
        RIe1bd218_3529,RIe1b0090_3380,RIe1726c8_2679,RIdec4460_697,RIdec1760_665,RIee1fae0_4819,RIdebea60_633,RIee1f108_4812,RIdebbd60_601,RIdeb9060_569,
        RIdeb6360_537,RIee1eb68_4808,RIdeb0960_473,RIee1e460_4803,RIdeadc60_441,RIee1d7b8_4794,RIdea8008_409,RIdea1708_377,RIde9ae08_345,RIfe957d8_8045,
        RIfe95508_8043,RIfe95670_8044,RIee1a7e8_4760,RIfe95aa8_8047,RIfe95238_8041,RIfe95940_8046,RIfe953a0_8042,RIee1a0e0_4755,RIee19ca8_4752,RIee19870_4749,
        RIee19438_4746,RIee38ba8_5104,RIfe95c10_8048,RIee384a0_5099,RIfea9440_8242,RIe164460_2518,RIe161760_2486,RIfe942c0_8030,RIe15ea60_2454,RIfe94158_8029,
        RIe15bd60_2422,RIe156360_2358,RIe153660_2326,RIfe94428_8031,RIe150960_2294,RIfe94590_8032,RIe14dc60_2262,RIfc5c2e8_6071,RIe14af60_2230,RIe148260_2198,
        RIe145560_2166,RIee33ce8_5048,RIee32aa0_5035,RIee31858_5022,RIfc5d530_6084,RIe140538_2109,RIdf3e2d8_2084,RIdf3c118_2060,RIdf39df0_2035,RIfcdd780_7542,
        RIee2ee28_4992,RIfcc88d0_7304,RIee2cc68_4968,RIdf34990_1975,RIdf32aa0_1953,RIdf304a8_1926,RIdf2e5b8_1904,RIee2b1b0_4949,RIfe946f8_8033,RIfcb2940_7054,
        RIee273d0_4905,RIfe949c8_8035,RIdf27538_1824,RIfe94b30_8036,RIfe94860_8034,RIee26f98_4902,RIee269f8_4898,RIee26728_4896,RIee26458_4894,RIee26188_4892,
        RIfe94c98_8037,RIee25d50_4889,RIfea9170_8240,RIdf16030_1627,RIdf13330_1595,RIdf10630_1563,RIdf0d930_1531,RIdf0ac30_1499,RIdf07f30_1467,RIdf05230_1435,
        RIdf02530_1403,RIdefcb30_1339,RIdef9e30_1307,RIdef7130_1275,RIdef4430_1243,RIdef1730_1211,RIdeeea30_1179,RIdeebd30_1147,RIdee9030_1115,RIee250a8_4880,
        RIee24298_4870,RIee23758_4862,RIee22d80_4855,RIfe950d0_8040,RIfe94f68_8039,RIfe94e00_8038,RIdeddd98_988,RIee22ab0_4853,RIee21e08_4844,RIfca46d8_6893,
        RIfc5dad0_6088,RIfeaa250_8252,RIfe96048_8051,RIfe95d78_8049,RIfe95ee0_8050,RIdecf860_825,RIdeccb60_793,RIdec9e60_761,RIdec7160_729,RIdeb3660_505,
        RIde94508_313,RIe16d268_2619,RIe159060_2390,RIe142860_2134,RIdf37258_2004,RIdf2b8b8_1872,RIdf1c138_1696,RIdeff830_1371,RIdee6330_1083,RIdedb098_956,
        RIde7a450_186,RIe19c6f8_3157,RIe1999f8_3125,RIf1450b8_5245,RIe196cf8_3093,RIf143fd8_5233,RIe193ff8_3061,RIe1912f8_3029,RIe18e5f8_2997,RIe188bf8_2933,
        RIe185ef8_2901,RIfe973f8_8065,RIe1831f8_2869,RIf142958_5217,RIe1804f8_2837,RIe17d7f8_2805,RIe17aaf8_2773,RIf141b48_5207,RIfc542f0_5980,RIfc800a8_6479,
        RIe175260_2710,RIfca0bc8_6851,RIfc48680_5846,RIee3dea0_5163,RIfcc6878_7281,RIee3ba10_5137,RIee3a930_5125,RIfe97290_8064,RIe172b00_2682,RIf16f958_5729,
        RIf16ee18_5721,RIf16da68_5707,RIf16d360_5702,RIfe96e58_8061,RIe222a50_4684,RIfe96cf0_8060,RIe21fd50_4652,RIf16a660_5670,RIe21d050_4620,RIe217650_4556,
        RIe214950_4524,RIf169f58_5665,RIe211c50_4492,RIf168770_5648,RIe20ef50_4460,RIf1677f8_5637,RIe20c250_4428,RIe209550_4396,RIe206850_4364,RIf166880_5626,
        RIf1657a0_5614,RIe201dc8_4311,RIe2005e0_4294,RIfe96b88_8059,RIf163b80_5594,RIf162c08_5583,RIf161420_5566,RIf15f530_5544,RIf15d7a8_5523,RIfe968b8_8057,
        RIfe96a20_8058,RIfcb3fc0_7070,RIfc7cf70_6444,RIfc579c8_6019,RIf159590_5476,RIf1584b0_5464,RIf157268_5451,RIf1569f8_5445,RIfe965e8_8055,RIf155d50_5436,
        RIf155210_5428,RIf153e60_5414,RIfe96750_8056,RIf1527e0_5398,RIf151430_5384,RIfcd2650_7416,RIe1f2648_4135,RIf14f108_5359,RIfc7f298_6469,RIf14d4e8_5339,
        RIe1ed350_4076,RIe1ea7b8_4045,RIe1e7ab8_4013,RIe1e4db8_3981,RIe1e20b8_3949,RIe1df3b8_3917,RIe1dc6b8_3885,RIe1d99b8_3853,RIe1d6cb8_3821,RIe1d12b8_3757,
        RIe1ce5b8_3725,RIe1cb8b8_3693,RIe1c8bb8_3661,RIe1c5eb8_3629,RIe1c31b8_3597,RIe1c04b8_3565,RIe1bd7b8_3533,RIf14c138_5325,RIf14ad88_5311,RIe1b8790_3476,
        RIfe96480_8054,RIf14a0e0_5302,RIf149870_5296,RIfe97128_8063,RIfe96318_8053,RIf148628_5283,RIfc58d78_6033,RIe1b20e8_3403,RIe1b04c8_3383,RIf146cd8_5265,
        RIfc591b0_6036,RIfe961b0_8052,RIfe96fc0_8062,RIe1a7af8_3285,RIe1a4df8_3253,RIe1a20f8_3221,RIe19f3f8_3189,RIe18b8f8_2965,RIe177df8_2741,RIe225750_4716,
        RIe21a350_4588,RIe203b50_4332,RIe1fdbb0_4264,RIe1f6f68_4187,RIe1efab0_4104,RIe1d3fb8_3789,RIe1baab8_3501,RIe1ad930_3352,RIe16ff68_2651,RIdec42f8_696,
        RIdec15f8_664,RIfcc6cb0_7284,RIdebe8f8_632,RIfe93780_8022,RIdebbbf8_600,RIdeb8ef8_568,RIdeb61f8_536,RIee1ea00_4807,RIdeb07f8_472,RIee1e2f8_4802,
        RIdeadaf8_440,RIfc5d3c8_6083,RIdea7cc0_408,RIdea13c0_376,RIde9aac0_344,RIfc58238_6025,RIfcc3b78_7249,RIfc7d0d8_6445,RIfc59750_6040,RIfe93a50_8024,
        RIfe938e8_8023,RIde88370_254,RIde83e88_233,RIfc5f420_6106,RIfc976b8_6745,RIfc90a70_6668,RIfc60500_6118,RIee38a40_5103,RIe16ab08_2591,RIe169488_2575,
        RIe166ff8_2549,RIe1642f8_2517,RIe1615f8_2485,RIee369e8_5080,RIe15e8f8_2453,RIee35bd8_5070,RIe15bbf8_2421,RIe1561f8_2357,RIe1534f8_2325,RIfc3ee28_5741,
        RIe1507f8_2293,RIfce6c90_7648,RIe14daf8_2261,RIfcca7c0_7326,RIe14adf8_2229,RIe1480f8_2197,RIe1453f8_2165,RIee33b80_5047,RIee32938_5034,RIee316f0_5021,
        RIee30bb0_5013,RIe1403d0_2108,RIfe93618_8021,RIdf3bfb0_2059,RIfe934b0_8020,RIfcd0d00_7398,RIee2ecc0_4991,RIee2e720_4987,RIee2cb00_4967,RIfe93bb8_8025,
        RIdf32938_1952,RIdf30340_1925,RIdf2e450_1903,RIee2b048_4948,RIee29b30_4933,RIfc67148_6195,RIfc6fb18_6293,RIdf29860_1849,RIfe931e0_8018,RIfe93348_8019,
        RIfe93078_8017,RIfc672b0_6196,RIfca8788_6939,RIdf22510_1767,RIfcea7a0_7690,RIdf20ff8_1752,RIdf1ecd0_1727,RIdf1aab8_1680,RIfea7c58_8225,RIdf15ec8_1626,
        RIdf131c8_1594,RIdf104c8_1562,RIdf0d7c8_1530,RIdf0aac8_1498,RIdf07dc8_1466,RIdf050c8_1434,RIdf023c8_1402,RIdefc9c8_1338,RIdef9cc8_1306,RIdef6fc8_1274,
        RIdef42c8_1242,RIdef15c8_1210,RIdeee8c8_1178,RIdeebbc8_1146,RIdee8ec8_1114,RIee24f40_4879,RIee24130_4869,RIee235f0_4861,RIee22c18_4854,RIfe93d20_8026,
        RIdee1fb0_1035,RIdee0228_1014,RIdeddc30_987,RIfc684f8_6209,RIee21ca0_4843,RIfc68390_6208,RIee20d28_4832,RIded8aa0_929,RIfe93ff0_8028,RIded45b8_880,
        RIfe93e88_8027,RIdecf6f8_824,RIdecc9f8_792,RIdec9cf8_760,RIdec6ff8_728,RIdeb34f8_504,RIde941c0_312,RIe16d100_2618,RIe158ef8_2389,RIe1426f8_2133,
        RIdf370f0_2003,RIdf2b750_1871,RIdf1bfd0_1695,RIdeff6c8_1370,RIdee61c8_1082,RIdedaf30_955,RIde7a108_185,RIe19c590_3156,RIe199890_3124,RIf144f50_5244,
        RIe196b90_3092,RIfc76058_6365,RIe193e90_3060,RIe191190_3028,RIe18e490_2996,RIe188a90_2932,RIe185d90_2900,RIfccd8f8_7361,RIe183090_2868,RIfc76e68_6375,
        RIe180390_2836,RIe17d690_2804,RIe17a990_2772,RIf1419e0_5206,RIf140630_5192,RIe176bb0_2728,RIe1750f8_2709,RIfcd1840_7406,RIfc5f6f0_6108,RIee3dd38_5162,
        RIee3cc58_5150,RIee3b8a8_5136,RIee3a7c8_5124,RIee39580_5111,RIfea9008_8239,RIf16f7f0_5728,RIf16ecb0_5720,RIf16d900_5706,RIfc78ec0_6398,RIfcc8060_7298,
        RIe2228e8_4683,RIfc5a3f8_6049,RIe21fbe8_4651,RIfc74000_6342,RIe21cee8_4619,RIe2174e8_4555,RIe2147e8_4523,RIfca2c20_6874,RIe211ae8_4491,RIfca2950_6872,
        RIe20ede8_4459,RIfcc24f8_7233,RIe20c0e8_4427,RIe2093e8_4395,RIe2066e8_4363,RIfc45110_5808,RIfcc6f80_7286,RIfe92f10_8016,RIfe92970_8012,RIf164af8_5605,
        RIf163a18_5593,RIf162aa0_5582,RIfe92ad8_8013,RIf15f3c8_5543,RIf15d640_5522,RIfe92808_8011,RIfe92c40_8014,RIfe926a0_8010,RIfe92da8_8015,RIfe92538_8009,
        RIfcb5a78_7089,RIf158348_5463,RIf157100_5450,RIfc53be8_5975,RIfec38b8_8345,RIfcc5ea0_7274,RIf1550a8_5427,RIf153cf8_5413,RIfec3a20_8346,RIf152678_5397,
        RIfec3750_8344,RIf14ff18_5369,RIfe923d0_8008,RIf14efa0_5358,RIf14e898_5353,RIf14d380_5338,RIfe92268_8007,RIe1ea650_4044,RIe1e7950_4012,RIe1e4c50_3980,
        RIe1e1f50_3948,RIe1df250_3916,RIe1dc550_3884,RIe1d9850_3852,RIe1d6b50_3820,RIe1d1150_3756,RIe1ce450_3724,RIe1cb750_3692,RIe1c8a50_3660,RIe1c5d50_3628,
        RIe1c3050_3596,RIe1c0350_3564,RIe1bd650_3532,RIfcda4e0_7506,RIfc9d220_6810,RIe1b8628_3475,RIe1b6738_3453,RIfc4f2c8_5923,RIfce16c8_7587,RIfe91cc8_8003,
        RIfe91e30_8004,RIf1484c0_5282,RIf147548_5271,RIfe91f98_8005,RIfe91b60_8002,RIf146b70_5264,RIfc9f548_6835,RIfe92100_8006,RIfe919f8_8001,RIe1a7990_3284,
        RIe1a4c90_3252,RIe1a1f90_3220,RIe19f290_3188,RIe18b790_2964,RIe177c90_2740,RIe2255e8_4715,RIe21a1e8_4587,RIe2039e8_4331,RIe1fda48_4263,RIe1f6e00_4186,
        RIe1ef948_4103,RIe1d3e50_3788,RIe1ba950_3500,RIe1ad7c8_3351,RIe16fe00_2650,RIdec4730_699,RIdec1a30_667,RIfce3f90_7616,RIdebed30_635,RIfcc3308_7243,
        RIdebc030_603,RIdeb9330_571,RIdeb6630_539,RIfc8c588_6619,RIdeb0c30_475,RIfc5a998_6053,RIdeadf30_443,RIfc99b48_6771,RIdea8698_411,RIdea1d98_379,
        RIde9b498_347,RIfc78bf0_6396,RIfcbc558_7165,RIfca12d0_6856,RIfca3fd0_6888,RIfec2670_8332,RIfec2508_8331,RIde88a00_256,RIde84518_235,RIfcc35d8_7245,
        RIfcb57a8_7087,RIfc5a290_6048,RIfca3058_6877,RIee38e78_5106,RIfec27d8_8333,RIfca3328_6879,RIe1672c8_2551,RIe164730_2520,RIe161a30_2488,RIee36cb8_5082,
        RIe15ed30_2456,RIfcc7250_7288,RIe15c030_2424,RIe156630_2360,RIe153930_2328,RIfcc7688_7291,RIe150c30_2296,RIfc8af08_6603,RIe14df30_2264,RIfc9a250_6776,
        RIe14b230_2232,RIe148530_2200,RIe145830_2168,RIfc9aac0_6782,RIfc56bb8_6009,RIfca1ca8_6863,RIfcec960_7714,RIe1406a0_2110,RIdf3e440_2085,RIdf3c280_2061,
        RIdf39f58_2036,RIfc9a958_6781,RIee2f0f8_4994,RIfcdb458_7517,RIee2cf38_4970,RIdf34c60_1977,RIfec2940_8334,RIdf30778_1928,RIdf2e888_1906,RIee2b480_4951,
        RIfec23a0_8330,RIee288e8_4920,RIfec2238_8329,RIdf29b30_1851,RIdf27808_1826,RIdf25a80_1805,RIdf23e60_1785,RIfc55100_5990,RIfcd9f40_7502,RIfc54f98_5989,
        RIfc54cc8_5987,RIfc4b218_5877,RIdf1efa0_1729,RIfcc69e0_7282,RIdf18bc8_1658,RIdf16300_1629,RIdf13600_1597,RIdf10900_1565,RIdf0dc00_1533,RIdf0af00_1501,
        RIdf08200_1469,RIdf05500_1437,RIdf02800_1405,RIdefce00_1341,RIdefa100_1309,RIdef7400_1277,RIdef4700_1245,RIdef1a00_1213,RIdeeed00_1181,RIdeec000_1149,
        RIdee9300_1117,RIfce4ad0_7624,RIfc9e8a0_6826,RIfcc46b8_7257,RIfcd4108_7435,RIdee4440_1061,RIdee2280_1037,RIdee0390_1015,RIdede068_990,RIfcda0a8_7503,
        RIfce54a8_7631,RIfca0790_6848,RIfc50ee8_5943,RIded8d70_931,RIded68e0_905,RIded4888_882,RIded2560_857,RIdecfb30_827,RIdecce30_795,RIdeca130_763,
        RIdec7430_731,RIdeb3930_507,RIde94b98_315,RIe16d538_2621,RIe159330_2392,RIe142b30_2136,RIdf37528_2006,RIdf2bb88_1874,RIdf1c408_1698,RIdeffb00_1373,
        RIdee6600_1085,RIdedb368_958,RIde7aae0_188,RIe19c9c8_3159,RIe199cc8_3127,RIfe8ea28_7967,RIe196fc8_3095,RIfec20d0_8328,RIe1942c8_3063,RIe1915c8_3031,
        RIe18e8c8_2999,RIe188ec8_2935,RIe1861c8_2903,RIfc68228_6207,RIe1834c8_2871,RIfccb5d0_7336,RIe1807c8_2839,RIe17dac8_2807,RIe17adc8_2775,RIf141e18_5209,
        RIf140900_5194,RIf140090_5188,RIe1753c8_2711,RIf13f988_5183,RIf13ece0_5174,RIee3e170_5165,RIee3cf28_5152,RIee3bce0_5139,RIee3ac00_5127,RIee39850_5113,
        RIe172dd0_2684,RIf16fc28_5731,RIf16f0e8_5723,RIf16dd38_5709,RIfce9120_7674,RIfc404a8_5757,RIe222d20_4686,RIf16b8a8_5683,RIe220020_4654,RIf16a930_5672,
        RIe21d320_4622,RIe217920_4558,RIe214c20_4526,RIfc5b910_6064,RIe211f20_4494,RIfe8e8c0_7966,RIe20f220_4462,RIfe8e758_7965,RIe20c520_4430,RIe209820_4398,
        RIe206b20_4366,RIf166b50_5628,RIf165a70_5616,RIfe8dd80_7958,RIfe8dab0_7956,RIf164c60_5606,RIf163e50_5596,RIf162ed8_5585,RIf1616f0_5568,RIf15f800_5546,
        RIf15da78_5525,RIfe8d948_7955,RIfe8dc18_7957,RIf15c560_5510,RIf15b048_5495,RIfc62828_6143,RIf159860_5478,RIf158780_5466,RIf157538_5453,RIfca6e38_6921,
        RIe1f9b00_4218,RIfc61e50_6136,RIfc61748_6131,RIf154130_5416,RIe1f4ad8_4161,RIf152ab0_5400,RIf151700_5386,RIf1501e8_5371,RIe1f27b0_4136,RIfc60ed8_6125,
        RIfc7b620_6426,RIf14d7b8_5341,RIe1ed4b8_4077,RIe1eaa88_4047,RIe1e7d88_4015,RIe1e5088_3983,RIe1e2388_3951,RIe1df688_3919,RIe1dc988_3887,RIe1d9c88_3855,
        RIe1d6f88_3823,RIe1d1588_3759,RIe1ce888_3727,RIe1cbb88_3695,RIe1c8e88_3663,RIe1c6188_3631,RIe1c3488_3599,RIe1c0788_3567,RIe1bda88_3535,RIfca4de0_6898,
        RIfc5ea48_6099,RIe1b8a60_3478,RIe1b6a08_3455,RIfcbd638_7177,RIfc44fa8_5807,RIfe8e5f0_7964,RIfe8e1b8_7961,RIf1488f8_5285,RIf147818_5273,RIfe8e050_7960,
        RIfe8e488_7963,RIf146e40_5266,RIf146030_5256,RIfe8dee8_7959,RIfe8e320_7962,RIe1a7dc8_3287,RIe1a50c8_3255,RIe1a23c8_3223,RIe19f6c8_3191,RIe18bbc8_2967,
        RIe1780c8_2743,RIe225a20_4718,RIe21a620_4590,RIe203e20_4334,RIe1fde80_4266,RIe1f7238_4189,RIe1efd80_4106,RIe1d4288_3791,RIe1bad88_3503,RIe1adc00_3354,
        RIe170238_2653,RIdec45c8_698,RIdec18c8_666,RIfce85e0_7666,RIdebebc8_634,RIfcb8bb0_7124,RIdebbec8_602,RIdeb91c8_570,RIdeb64c8_538,RIfc85d78_6545,
        RIdeb0ac8_474,RIfc85aa8_6543,RIdeaddc8_442,RIfc4d3d8_5901,RIdea8350_410,RIdea1a50_378,RIde9b150_346,RIfc85ee0_6546,RIfc9c9b0_6804,RIfce13f8_7585,
        RIfcb8778_7121,RIfe8d510_7952,RIfe8d3a8_7951,RIde886b8_255,RIde841d0_234,RIde806c0_216,RIfcb8070_7116,RIfce1128_7583,RIfc9c140_6798,RIee38d10_5105,
        RIe16ac70_2592,RIfc850d0_6536,RIe167160_2550,RIe1645c8_2519,RIe1618c8_2487,RIee36b50_5081,RIe15ebc8_2455,RIee35d40_5071,RIe15bec8_2423,RIe1564c8_2359,
        RIe1537c8_2327,RIfc3ef90_5742,RIe150ac8_2295,RIfe8d7e0_7954,RIe14ddc8_2263,RIfce0fc0_7582,RIe14b0c8_2231,RIe1483c8_2199,RIe1456c8_2167,RIee33e50_5049,
        RIee32c08_5036,RIee319c0_5023,RIee30d18_5014,RIfe8cf70_7948,RIfe8ce08_7947,RIfe8d240_7950,RIfe8d0d8_7949,RIfce9dc8_7683,RIee2ef90_4993,RIfce51d8_7629,
        RIee2cdd0_4969,RIdf34af8_1976,RIfe8d678_7953,RIdf30610_1927,RIdf2e720_1905,RIee2b318_4950,RIee29c98_4934,RIee28780_4919,RIee27538_4906,RIdf299c8_1850,
        RIdf276a0_1825,RIdf25918_1804,RIdf23cf8_1784,RIfc83ff0_6524,RIfcb73c8_7107,RIfc51320_5946,RIfcdaa80_7510,RIfc83d20_6522,RIdf1ee38_1728,RIfc51b90_5952,
        RIdf18a60_1657,RIdf16198_1628,RIdf13498_1596,RIdf10798_1564,RIdf0da98_1532,RIdf0ad98_1500,RIdf08098_1468,RIdf05398_1436,RIdf02698_1404,RIdefcc98_1340,
        RIdef9f98_1308,RIdef7298_1276,RIdef4598_1244,RIdef1898_1212,RIdeeeb98_1180,RIdeebe98_1148,RIdee9198_1116,RIee25210_4881,RIee24400_4871,RIee238c0_4863,
        RIee22ee8_4856,RIfe8cca0_7946,RIdee2118_1036,RIfe8cb38_7945,RIdeddf00_989,RIfcc5a68_7271,RIee21f70_4845,RIfcb6cc0_7102,RIee20e90_4833,RIded8c08_930,
        RIded6778_904,RIded4720_881,RIded23f8_856,RIdecf9c8_826,RIdecccc8_794,RIdec9fc8_762,RIdec72c8_730,RIdeb37c8_506,RIde94850_314,RIe16d3d0_2620,
        RIe1591c8_2391,RIe1429c8_2135,RIdf373c0_2005,RIdf2ba20_1873,RIdf1c2a0_1697,RIdeff998_1372,RIdee6498_1084,RIdedb200_957,RIde7a798_187,RIe19c860_3158,
        RIe199b60_3126,RIf145220_5246,RIe196e60_3094,RIf144140_5234,RIe194160_3062,RIe191460_3030,RIe18e760_2998,RIe188d60_2934,RIe186060_2902,RIf1431c8_5223,
        RIe183360_2870,RIf142ac0_5218,RIe180660_2838,RIe17d960_2806,RIe17ac60_2774,RIf141cb0_5208,RIf140798_5193,RIf13ff28_5187,RIfe8be90_7936,RIfceb880_7702,
        RIf13eb78_5173,RIee3e008_5164,RIee3cdc0_5151,RIee3bb78_5138,RIee3aa98_5126,RIee396e8_5112,RIe172c68_2683,RIf16fac0_5730,RIf16ef80_5722,RIf16dbd0_5708,
        RIfcc4af0_7260,RIf16c820_5694,RIe222bb8_4685,RIf16b740_5682,RIe21feb8_4653,RIf16a7c8_5671,RIe21d1b8_4621,RIe2177b8_4557,RIe214ab8_4525,RIfe8c430_7940,
        RIe211db8_4493,RIf1688d8_5649,RIe20f0b8_4461,RIf167960_5638,RIe20c3b8_4429,RIe2096b8_4397,RIe2069b8_4365,RIf1669e8_5627,RIf165908_5615,RIfe8c9d0_7944,
        RIfe8c700_7942,RIfc9c578_6801,RIf163ce8_5595,RIf162d70_5584,RIf161588_5567,RIf15f698_5545,RIf15d910_5524,RIfe8c598_7941,RIfe8c868_7943,RIf15c3f8_5509,
        RIf15aee0_5494,RIf15a0d0_5484,RIf1596f8_5477,RIf158618_5465,RIf1573d0_5452,RIf156b60_5446,RIfec1f68_8327,RIf155eb8_5437,RIf155378_5429,RIf153fc8_5415,
        RIfe8bff8_7937,RIf152948_5399,RIf151598_5385,RIf150080_5370,RIfe8c2c8_7939,RIf14f270_5360,RIfc503a8_5935,RIf14d650_5340,RIfe8c160_7938,RIe1ea920_4046,
        RIe1e7c20_4014,RIe1e4f20_3982,RIe1e2220_3950,RIe1df520_3918,RIe1dc820_3886,RIe1d9b20_3854,RIe1d6e20_3822,RIe1d1420_3758,RIe1ce720_3726,RIe1cba20_3694,
        RIe1c8d20_3662,RIe1c6020_3630,RIe1c3320_3598,RIe1c0620_3566,RIe1bd920_3534,RIf14c2a0_5326,RIf14aef0_5312,RIe1b88f8_3477,RIe1b68a0_3454,RIfcd4db0_7444,
        RIfc4ebc0_5918,RIfec1e00_8326,RIfe8bd28_7935,RIf148790_5284,RIf1476b0_5272,RIfe8ba58_7933,RIfec1b30_8324,RIfc4e788_5915,RIfcb8e80_7126,RIfe8bbc0_7934,
        RIfec1c98_8325,RIe1a7c60_3286,RIe1a4f60_3254,RIe1a2260_3222,RIe19f560_3190,RIe18ba60_2966,RIe177f60_2742,RIe2258b8_4717,RIe21a4b8_4589,RIe203cb8_4333,
        RIe1fdd18_4265,RIe1f70d0_4188,RIe1efc18_4105,RIe1d4120_3790,RIe1bac20_3502,RIe1ada98_3353,RIe1700d0_2652,RIdec4a00_701,RIdec1d00_669,RIfcad7b0_6996,
        RIdebf000_637,RIfc64cb8_6169,RIdebc300_605,RIdeb9600_573,RIdeb6900_541,RIfc6f9b0_6292,RIdeb0f00_477,RIfc657f8_6177,RIdeae200_445,RIfce69c0_7646,
        RIdea8d28_413,RIdea2428_381,RIde9bb28_349,RIfc6fc80_6294,RIee1b760_4771,RIfca8080_6934,RIfe8b8f0_7932,RIde90020_292,RIde8c510_274,RIde89090_258,
        RIde84ba8_237,RIfc65ac8_6179,RIfcad210_6992,RIfcce168_7367,RIfcce2d0_7368,RIfc51488_5947,RIe16af40_2594,RIfc65c30_6180,RIe167598_2553,RIe164a00_2522,
        RIe161d00_2490,RIfc66e78_6193,RIe15f000_2458,RIfc6e498_6277,RIe15c300_2426,RIe156900_2362,RIe153c00_2330,RIfc6e330_6276,RIe150f00_2298,RIfccda60_7362,
        RIe14e200_2266,RIfc6e1c8_6275,RIe14b500_2234,RIe148800_2202,RIe145b00_2170,RIee33fb8_5050,RIee32d70_5037,RIee31c90_5025,RIee30fe8_5016,RIfea8630_8232,
        RIdf3e5a8_2086,RIdf3c550_2063,RIfea8798_8233,RIfc6e060_6274,RIfcac6d0_6984,RIfc56078_6001,RIfc6e600_6278,RIdf34dc8_1978,RIdf32d70_1955,RIfea84c8_8231,
        RIdf2eb58_1908,RIee2b750_4953,RIfc6ee70_6284,RIfc6efd8_6285,RIee27808_4908,RIfe8b788_7931,RIdf27ad8_1828,RIdf25d50_1807,RIdf24130_1787,RIfc66608_6187,
        RIfccde98_7365,RIfc66a40_6190,RIfc668d8_6189,RIfcacf40_6990,RIfeaaef8_8261,RIfc6e8d0_6280,RIdf18d30_1659,RIdf165d0_1631,RIdf138d0_1599,RIdf10bd0_1567,
        RIdf0ded0_1535,RIdf0b1d0_1503,RIdf084d0_1471,RIdf057d0_1439,RIdf02ad0_1407,RIdefd0d0_1343,RIdefa3d0_1311,RIdef76d0_1279,RIdef49d0_1247,RIdef1cd0_1215,
        RIdeeefd0_1183,RIdeec2d0_1151,RIdee95d0_1119,RIfc6dc28_6271,RIfc67c88_6203,RIfccb300_7334,RIfccd4c0_7358,RIfea81f8_8229,RIfea8360_8230,RIdee04f8_1016,
        RIdede338_992,RIfc6def8_6273,RIfcac130_6980,RIfc67b20_6202,RIfc67df0_6204,RIded9040_933,RIded6a48_906,RIded4b58_884,RIded26c8_858,RIdecfe00_829,
        RIdecd100_797,RIdeca400_765,RIdec7700_733,RIdeb3c00_509,RIde95228_317,RIe16d808_2623,RIe159600_2394,RIe142e00_2138,RIdf377f8_2008,RIdf2be58_1876,
        RIdf1c6d8_1700,RIdeffdd0_1375,RIdee68d0_1087,RIdedb638_960,RIde7b170_190,RIe19cc98_3161,RIe199f98_3129,RIfc73088_6331,RIe197298_3097,RIf1442a8_5235,
        RIe194598_3065,RIe191898_3033,RIe18eb98_3001,RIe189198_2937,RIe186498_2905,RIfc72278_6321,RIe183798_2873,RIfc61ce8_6135,RIe180a98_2841,RIe17dd98_2809,
        RIe17b098_2777,RIfcaf268_7015,RIfca6a00_6918,RIfcc9b18_7317,RIe175530_2712,RIfc72818_6325,RIfc726b0_6324,RIfccf7e8_7383,RIfc72548_6323,RIee3be48_5140,
        RIee3ad68_5128,RIfc71fa8_6319,RIe1730a0_2686,RIfcaef98_7013,RIfccf518_7381,RIfc71e40_6318,RIfc62120_6138,RIfe8b350_7928,RIe222ff0_4688,RIfcc9f50_7320,
        RIe2202f0_4656,RIfc4a570_5868,RIe21d5f0_4624,RIe217bf0_4560,RIe214ef0_4528,RIfccf3b0_7380,RIe2121f0_4496,RIf168ba8_5651,RIe20f4f0_4464,RIfc71300_6310,
        RIe20c7f0_4432,RIe209af0_4400,RIe206df0_4368,RIfc718a0_6314,RIfc71a08_6315,RIe202098_4313,RIfe8b1e8_7927,RIfc715d0_6312,RIfce6588_7643,RIfc62c60_6146,
        RIf161858_5569,RIf15fad0_5548,RIf15dbe0_5526,RIe1fc698_4249,RIfe8b4b8_7929,RIfcae5c0_7006,RIfc63098_6149,RIfc63200_6150,RIfc71198_6309,RIf158a50_5468,
        RIf1576a0_5454,RIfcdc808_7531,RIfe8b620_7930,RIfc634d0_6152,RIfcceb40_7374,RIf154400_5418,RIe1f4da8_4163,RIf152c18_5401,RIf151868_5387,RIfc4d108_5899,
        RIe1f2a80_4138,RIfc70a90_6304,RIfc63bd8_6157,RIfca7810_6928,RIe1ed788_4079,RIe1ead58_4049,RIe1e8058_4017,RIe1e5358_3985,RIe1e2658_3953,RIe1df958_3921,
        RIe1dcc58_3889,RIe1d9f58_3857,RIe1d7258_3825,RIe1d1858_3761,RIe1ceb58_3729,RIe1cbe58_3697,RIe1c9158_3665,RIe1c6458_3633,RIe1c3758_3601,RIe1c0a58_3569,
        RIe1bdd58_3537,RIf14c408_5327,RIf14b1c0_5314,RIe1b8d30_3480,RIe1b6cd8_3457,RIfc707c0_6302,RIfca7c48_6931,RIe1b4de8_3435,RIe1b3a38_3421,RIfc70220_6298,
        RIfcce870_7372,RIe1b23b8_3405,RIe1b0630_3384,RIfc645b0_6164,RIfc700b8_6297,RIfeaac28_8259,RIe1aa690_3316,RIe1a8098_3289,RIe1a5398_3257,RIe1a2698_3225,
        RIe19f998_3193,RIe18be98_2969,RIe178398_2745,RIe225cf0_4720,RIe21a8f0_4592,RIe2040f0_4336,RIe1fe150_4268,RIe1f7508_4191,RIe1f0050_4108,RIe1d4558_3793,
        RIe1bb058_3505,RIe1aded0_3356,RIe170508_2655,RIdec4898_700,RIdec1b98_668,RIfc661d0_6184,RIdebee98_636,RIfce6b28_7647,RIdebc198_604,RIdeb9498_572,
        RIdeb6798_540,RIfc40d18_5763,RIdeb0d98_476,RIfcad648_6995,RIdeae098_444,RIfcaa510_6960,RIdea89e0_412,RIdea20e0_380,RIde9b7e0_348,RIfcab320_6970,
        RIfca8350_6936,RIfc6f6e0_6290,RIfcaa240_6958,RIde8fcd8_291,RIfe8aae0_7922,RIde88d48_257,RIde84860_236,RIde80a08_217,RIfc64718_6165,RIfcae020_7002,
        RIfcadeb8_7001,RIee38fe0_5107,RIe16add8_2593,RIe1695f0_2576,RIe167430_2552,RIe164898_2521,RIe161b98_2489,RIfe8a3d8_7917,RIe15ee98_2457,RIfe8a270_7916,
        RIe15c198_2425,RIe156798_2361,RIe153a98_2329,RIfc3f0f8_5743,RIe150d98_2297,RIfcab050_6968,RIe14e098_2265,RIfcca658_7325,RIe14b398_2233,RIe148698_2201,
        RIe145998_2169,RIfe8a810_7920,RIfe8a6a8_7919,RIee31b28_5024,RIee30e80_5015,RIe140808_2111,RIfe8a540_7918,RIdf3c3e8_2062,RIdf3a0c0_2037,RIfc6b1f8_6241,
        RIee2f260_4995,RIfc70d60_6306,RIee2d0a0_4971,RIfe8a978_7921,RIdf32c08_1954,RIdf308e0_1929,RIdf2e9f0_1907,RIee2b5e8_4952,RIee29e00_4935,RIee28a50_4921,
        RIee276a0_4907,RIdf29c98_1852,RIdf27970_1827,RIdf25be8_1806,RIdf23fc8_1786,RIfc6aaf0_6236,RIfc6ac58_6237,RIdf22678_1768,RIfcdd4b0_7540,RIdf21160_1753,
        RIdf1f108_1730,RIdf1ac20_1681,RIfeaa7f0_8256,RIdf16468_1630,RIdf13768_1598,RIdf10a68_1566,RIdf0dd68_1534,RIdf0b068_1502,RIdf08368_1470,RIdf05668_1438,
        RIdf02968_1406,RIdefcf68_1342,RIdefa268_1310,RIdef7568_1278,RIdef4868_1246,RIdef1b68_1214,RIdeeee68_1182,RIdeec168_1150,RIdee9468_1118,RIee25378_4882,
        RIee24568_4872,RIee23a28_4864,RIee23050_4857,RIfe8adb0_7924,RIdee23e8_1038,RIfe8ac48_7923,RIdede1d0_991,RIfca5650_6904,RIee220d8_4846,RIfceeb20_7738,
        RIee20ff8_4834,RIded8ed8_932,RIfe8af18_7925,RIded49f0_883,RIfe8b080_7926,RIdecfc98_828,RIdeccf98_796,RIdeca298_764,RIdec7598_732,RIdeb3a98_508,
        RIde94ee0_316,RIe16d6a0_2622,RIe159498_2393,RIe142c98_2137,RIdf37690_2007,RIdf2bcf0_1875,RIdf1c570_1699,RIdeffc68_1374,RIdee6768_1086,RIdedb4d0_959,
        RIde7ae28_189,RIe19cb30_3160,RIe199e30_3128,RIf145388_5247,RIe197130_3096,RIfe8a108_7915,RIe194430_3064,RIe191730_3032,RIe18ea30_3000,RIe189030_2936,
        RIe186330_2904,RIfc6c878_6257,RIe183630_2872,RIfcabcf8_6977,RIe180930_2840,RIe17dc30_2808,RIe17af30_2776,RIfcccc50_7352,RIfcccdb8_7353,RIe176d18_2729,
        RIfea7af0_8224,RIfe89fa0_7914,RIfe89e38_7913,RIfcdd078_7537,RIfccb738_7337,RIfca9868_6951,RIfcabb90_6976,RIfca99d0_6952,RIe172f38_2685,RIf16fd90_5732,
        RIf16f250_5724,RIfc6c440_6254,RIfcaba28_6975,RIfc40610_5758,RIe222e88_4687,RIfc5d260_6082,RIe220188_4655,RIfcab758_6973,RIe21d488_4623,RIe217a88_4559,
        RIe214d88_4527,RIfe892f8_7905,RIe212088_4495,RIf168a40_5650,RIe20f388_4463,RIf167ac8_5639,RIe20c688_4431,RIe209988_4399,RIe206c88_4367,RIfc6c2d8_6253,
        RIfceec88_7739,RIe201f30_4312,RIe200748_4295,RIf164dc8_5607,RIf163fb8_5597,RIf163040_5586,RIfe895c8_7907,RIf15f968_5547,RIfe89898_7909,RIfe89460_7906,
        RIe1fb5b8_4237,RIf15c6c8_5511,RIfe89730_7908,RIf15a238_5485,RIf1599c8_5479,RIf1588e8_5467,RIfe89cd0_7912,RIfc5ba78_6065,RIe1f9c68_4219,RIfc5bd48_6067,
        RIf1554e0_5430,RIf154298_5417,RIe1f4c40_4162,RIfe89b68_7911,RIfe89a00_7910,RIf150350_5372,RIe1f2918_4137,RIf14f3d8_5361,RIfccc818_7349,RIf14d920_5342,
        RIe1ed620_4078,RIe1eabf0_4048,RIe1e7ef0_4016,RIe1e51f0_3984,RIe1e24f0_3952,RIe1df7f0_3920,RIe1dcaf0_3888,RIe1d9df0_3856,RIe1d70f0_3824,RIe1d16f0_3760,
        RIe1ce9f0_3728,RIe1cbcf0_3696,RIe1c8ff0_3664,RIe1c62f0_3632,RIe1c35f0_3600,RIe1c08f0_3568,RIe1bdbf0_3536,RIfc680c0_6206,RIf14b058_5313,RIe1b8bc8_3479,
        RIe1b6b70_3456,RIfcac298_6981,RIf1499d8_5297,RIfe89190_7904,RIfec19c8_8323,RIf148a60_5286,RIfccdd30_7364,RIe1b2250_3404,RIfec1860_8322,RIfc6e768_6279,
        RIfc54728_5983,RIe1abfe0_3334,RIe1aa528_3315,RIe1a7f30_3288,RIe1a5230_3256,RIe1a2530_3224,RIe19f830_3192,RIe18bd30_2968,RIe178230_2744,RIe225b88_4719,
        RIe21a788_4591,RIe203f88_4335,RIe1fdfe8_4267,RIe1f73a0_4190,RIe1efee8_4107,RIe1d43f0_3792,RIe1baef0_3504,RIe1add68_3355,RIe1703a0_2654,RIdec4cd0_703,
        RIdec1fd0_671,RIfc7b4b8_6425,RIdebf2d0_639,RIfc7b1e8_6423,RIdebc5d0_607,RIdeb98d0_575,RIdeb6bd0_543,RIfe83358_7837,RIdeb11d0_479,RIee1e5c8_4804,
        RIdeae4d0_447,RIfc437c0_5790,RIdea93b8_415,RIdea2ab8_383,RIde9c1b8_351,RIfc90ea8_6671,RIfc7af18_6421,RIfe83088_7835,RIee1a950_4761,RIde906b0_294,
        RIde8cba0_276,RIfe82f20_7834,RIfe82db8_7833,RIee1a248_4756,RIfe831f0_7836,RIfcc2390_7232,RIee195a0_4747,RIfcbe718_7189,RIfea9e18_8249,RIfc43220_5786,
        RIe167868_2555,RIe164cd0_2524,RIe161fd0_2492,RIee36f88_5084,RIe15f2d0_2460,RIee35ea8_5072,RIe15c5d0_2428,RIe156bd0_2364,RIe153ed0_2332,RIfe83628_7839,
        RIe1511d0_2300,RIfebfda8_8303,RIe14e4d0_2268,RIfebfc40_8302,RIe14b7d0_2236,RIe148ad0_2204,RIe145dd0_2172,RIee34120_5051,RIee32ed8_5038,RIee31df8_5026,
        RIfcc1f58_7229,RIe140ad8_2113,RIdf3e878_2088,RIfe834c0_7838,RIdf3a390_2039,RIfc5a6c8_6051,RIfc91e20_6682,RIee2e888_4988,RIfc96a10_6736,RIdf35098_1980,
        RIfeab600_8266,RIdf30bb0_1931,RIfeab768_8267,RIfcbe9e8_7191,RIfc79fa0_6410,RIfc96740_6734,RIfc92258_6685,RIfea7118_8217,RIfea95a8_8243,RIdf26020_1809,
        RIdf24400_1789,RIfc79a00_6406,RIfc5add0_6056,RIfce5d18_7637,RIfc92690_6688,RIfce3018_7605,RIdf1f270_1731,RIfc79730_6404,RIdf19000_1661,RIdf168a0_1633,
        RIdf13ba0_1601,RIdf10ea0_1569,RIdf0e1a0_1537,RIdf0b4a0_1505,RIdf087a0_1473,RIdf05aa0_1441,RIdf02da0_1409,RIdefd3a0_1345,RIdefa6a0_1313,RIdef79a0_1281,
        RIdef4ca0_1249,RIdef1fa0_1217,RIdeef2a0_1185,RIdeec5a0_1153,RIdee98a0_1121,RIfc5b7a8_6063,RIfc5b640_6062,RIfc931d0_6696,RIfcecac8_7715,RIdee4710_1063,
        RIdee26b8_1040,RIdee07c8_1018,RIdede4a0_993,RIfcbf0f0_7196,RIfcbf528_7199,RIfc792f8_6401,RIfc93068_6695,RIded91a8_934,RIded6d18_908,RIded4e28_886,
        RIded2998_860,RIded00d0_831,RIdecd3d0_799,RIdeca6d0_767,RIdec79d0_735,RIdeb3ed0_511,RIde958b8_319,RIe16dad8_2625,RIe1598d0_2396,RIe1430d0_2140,
        RIdf37ac8_2010,RIdf2c128_1878,RIdf1c9a8_1702,RIdf000a0_1377,RIdee6ba0_1089,RIdedb908_962,RIde7b800_192,RIe19cf68_3163,RIe19a268_3131,RIfc8d7d0_6632,
        RIe197568_3099,RIfc561e0_6002,RIe194868_3067,RIe191b68_3035,RIe18ee68_3003,RIe189468_2939,RIe186768_2907,RIf143330_5224,RIe183a68_2875,RIfc7d948_6451,
        RIe180d68_2843,RIe17e068_2811,RIe17b368_2779,RIfc564b0_6004,RIfcd6700_7462,RIfc461f0_5820,RIe175698_2713,RIfc46088_5819,RIfc45f20_5818,RIfc7dc18_6453,
        RIfcd69d0_7464,RIfc98630_6756,RIfcc2a98_7237,RIfc7d510_6448,RIe173208_2687,RIfc8e478_6641,RIfc45ae8_5815,RIfc8e8b0_6644,RIfc45980_5814,RIfe82ae8_7831,
        RIe2232c0_4690,RIf16ba10_5684,RIe2205c0_4658,RIfcd24e8_7415,RIe21d8c0_4626,RIe217ec0_4562,RIe2151c0_4530,RIfebf268_8295,RIe2124c0_4498,RIf168d10_5652,
        RIe20f7c0_4466,RIfc7d240_6446,RIe20cac0_4434,RIe209dc0_4402,RIe2070c0_4370,RIf166e20_5630,RIfebf6a0_8298,RIfebf808_8299,RIfebf538_8297,RIfc8eb80_6646,
        RIf164120_5598,RIfc453e0_5810,RIf161b28_5571,RIf15fc38_5549,RIf15dd48_5527,RIe1fc968_4251,RIe1fb888_4239,RIfebf3d0_8296,RIf15b318_5497,RIfca2518_6869,
        RIfc8f120_6650,RIfebfad8_8301,RIfebf970_8300,RIfc7cca0_6442,RIe1f9dd0_4220,RIfe82c50_7832,RIf155648_5431,RIfc8f288_6651,RIe1f4f10_4164,RIf152d80_5402,
        RIfc8f828_6655,RIfcb3b88_7067,RIe1f2d50_4140,RIfc445d0_5800,RIfc8faf8_6657,RIf14da88_5343,RIe1eda58_4081,RIe1eb028_4051,RIe1e8328_4019,RIe1e5628_3987,
        RIe1e2928_3955,RIe1dfc28_3923,RIe1dcf28_3891,RIe1da228_3859,RIe1d7528_3827,RIe1d1b28_3763,RIe1cee28_3731,RIe1cc128_3699,RIe1c9428_3667,RIe1c6728_3635,
        RIe1c3a28_3603,RIe1c0d28_3571,RIe1be028_3539,RIfc7bff8_6433,RIfc44030_5796,RIe1b9000_3482,RIe1b6fa8_3459,RIfcbdd40_7182,RIfc8ff30_6660,RIe1b50b8_3437,
        RIe1b3d08_3423,RIfcbe178_7185,RIfc43d60_5794,RIe1b2520_3406,RIe1b0798_3385,RIfcdb5c0_7518,RIfc7ba58_6429,RIe1ac148_3335,RIe1aa960_3318,RIe1a8368_3291,
        RIe1a5668_3259,RIe1a2968_3227,RIe19fc68_3195,RIe18c168_2971,RIe178668_2747,RIe225fc0_4722,RIe21abc0_4594,RIe2043c0_4338,RIe1fe420_4270,RIe1f77d8_4193,
        RIe1f0320_4110,RIe1d4828_3795,RIe1bb328_3507,RIe1ae1a0_3358,RIe1707d8_2657,RIdec4b68_702,RIdec1e68_670,RIfc5df08_6091,RIdebf168_638,RIfce6df8_7649,
        RIdebc468_606,RIdeb9768_574,RIdeb6a68_542,RIfc75ef0_6364,RIdeb1068_478,RIfcc12b0_7220,RIdeae368_446,RIfc5e340_6094,RIdea9070_414,RIdea2770_382,
        RIde9be70_350,RIfced4a0_7722,RIfcc1418_7221,RIfc95930_6724,RIfcec0f0_7708,RIde90368_293,RIde8c858_275,RIde893d8_259,RIde84ef0_238,RIde80d50_218,
        RIfc95a98_6725,RIfced068_7719,RIfced1d0_7720,RIfcedfe0_7730,RIe16b0a8_2595,RIe169758_2577,RIe167700_2554,RIe164b68_2523,RIe161e68_2491,RIee36e20_5083,
        RIe15f168_2459,RIfc426e0_5778,RIe15c468_2427,RIe156a68_2363,RIe153d68_2331,RIfe82818_7829,RIe151068_2299,RIee34c60_5059,RIe14e368_2267,RIfc5f9c0_6110,
        RIe14b668_2235,RIe148968_2203,RIe145c68_2171,RIfccfef0_7388,RIfca57b8_6905,RIfc600c8_6115,RIfcafda8_7023,RIe140970_2112,RIdf3e710_2087,RIdf3c6b8_2064,
        RIdf3a228_2038,RIfc5fc90_6112,RIee2f3c8_4996,RIfc742d0_6344,RIee2d208_4972,RIdf34f30_1979,RIfebf100_8294,RIdf30a48_1930,RIdf2ecc0_1909,RIfcb08e8_7031,
        RIfcee418_7733,RIfc95ed0_6728,RIfcdef68_7559,RIdf29e00_1853,RIdf27c40_1829,RIdf25eb8_1808,RIdf24298_1788,RIfc5ed18_6101,RIfcee850_7736,RIdf227e0_1769,
        RIfc5efe8_6103,RIdf212c8_1754,RIfeaa520_8254,RIdf1ad88_1682,RIdf18e98_1660,RIdf16738_1632,RIdf13a38_1600,RIdf10d38_1568,RIdf0e038_1536,RIdf0b338_1504,
        RIdf08638_1472,RIdf05938_1440,RIdf02c38_1408,RIdefd238_1344,RIdefa538_1312,RIdef7838_1280,RIdef4b38_1248,RIdef1e38_1216,RIdeef138_1184,RIdeec438_1152,
        RIdee9738_1120,RIfcc96e0_7314,RIfccfd88_7387,RIfc60aa0_6122,RIfca5ec0_6910,RIdee45a8_1062,RIdee2550_1039,RIdee0660_1017,RIfe826b0_7828,RIfcdeb30_7556,
        RIfc73bc8_6339,RIfca5bf0_6908,RIfc73a60_6338,RIfe82980_7830,RIded6bb0_907,RIded4cc0_885,RIded2830_859,RIdecff68_830,RIdecd268_798,RIdeca568_766,
        RIdec7868_734,RIdeb3d68_510,RIde95570_318,RIe16d970_2624,RIe159768_2395,RIe142f68_2139,RIdf37960_2009,RIdf2bfc0_1877,RIdf1c840_1701,RIdefff38_1376,
        RIdee6a38_1088,RIdedb7a0_961,RIde7b4b8_191,RIe19ce00_3162,RIe19a100_3130,RIfce96c0_7678,RIe197400_3098,RIf144410_5236,RIe194700_3066,RIe191a00_3034,
        RIe18ed00_3002,RIe189300_2938,RIe186600_2906,RIfebee30_8292,RIe183900_2874,RIfcdbcc8_7523,RIe180c00_2842,RIe17df00_2810,RIe17b200_2778,RIf141f80_5210,
        RIfce7398_7653,RIfcb1e00_7046,RIfe82548_7827,RIfca42a0_6890,RIfcbff00_7206,RIfcaaee8_6967,RIee3d090_5153,RIfc5c180_6070,RIfce35b8_7609,RIee399b8_5114,
        RIfea8a68_8235,RIf16fef8_5733,RIfebecc8_8291,RIfc5c450_6072,RIfce9288_7675,RIfc40778_5759,RIe223158_4689,RIfce77d0_7656,RIe220458_4657,RIfce24d8_7597,
        RIe21d758_4625,RIe217d58_4561,RIe215058_4529,RIfce8a18_7669,RIe212358_4497,RIfce1998_7589,RIe20f658_4465,RIfc77840_6382,RIe20c958_4433,RIe209c58_4401,
        RIe206f58_4369,RIf166cb8_5629,RIf165bd8_5617,RIfe81fa8_7823,RIfe81e40_7822,RIfc5c888_6075,RIfceb178_7697,RIf1631a8_5587,RIf1619c0_5570,RIfccf248_7379,
        RIfc77570_6380,RIe1fc800_4250,RIe1fb720_4238,RIf15c830_5512,RIf15b1b0_5496,RIfcd0fd0_7400,RIfccc6b0_7348,RIf158bb8_5469,RIf157808_5455,RIfc5d0f8_6081,
        RIfebef98_8293,RIfcc8a38_7305,RIfcd7ab0_7476,RIfcb1428_7039,RIfeaa0e8_8251,RIfccc548_7347,RIfce3450_7608,RIf1504b8_5373,RIe1f2be8_4139,RIf14f540_5362,
        RIfc772a0_6378,RIfcec258_7709,RIe1ed8f0_4080,RIe1eaec0_4050,RIe1e81c0_4018,RIe1e54c0_3986,RIe1e27c0_3954,RIe1dfac0_3922,RIe1dcdc0_3890,RIe1da0c0_3858,
        RIe1d73c0_3826,RIe1d19c0_3762,RIe1cecc0_3730,RIe1cbfc0_3698,RIe1c92c0_3666,RIe1c65c0_3634,RIe1c38c0_3602,RIe1c0bc0_3570,RIe1bdec0_3538,RIf14c570_5328,
        RIf14b328_5315,RIe1b8e98_3481,RIe1b6e40_3458,RIfc76760_6370,RIfc94b20_6714,RIe1b4f50_3436,RIe1b3ba0_3422,RIfcec3c0_7710,RIfceb010_7696,RIfe823e0_7826,
        RIfe82110_7824,RIfcdd8e8_7543,RIfcc0ba8_7215,RIfe82278_7825,RIe1aa7f8_3317,RIe1a8200_3290,RIe1a5500_3258,RIe1a2800_3226,RIe19fb00_3194,RIe18c000_2970,
        RIe178500_2746,RIe225e58_4721,RIe21aa58_4593,RIe204258_4337,RIe1fe2b8_4269,RIe1f7670_4192,RIe1f01b8_4109,RIe1d46c0_3794,RIe1bb1c0_3506,RIe1ae038_3357,
        RIe170670_2656,RIdec4fa0_705,RIdec22a0_673,RIee1fdb0_4821,RIdebf5a0_641,RIee1f270_4813,RIdebc8a0_609,RIdeb9ba0_577,RIdeb6ea0_545,RIee1ecd0_4809,
        RIdeb14a0_481,RIee1e730_4805,RIdeae7a0_449,RIee1d920_4795,RIdea9a48_417,RIdea3148_385,RIde9c848_353,RIee1cb10_4785,RIee1ba30_4773,RIee1b1c0_4767,
        RIfec04b0_8308,RIfe850e0_7858,RIde8d230_278,RIfea9cb0_8248,RIfe84f78_7857,RIee1a3b0_4757,RIfe853b0_7860,RIee199d8_4750,RIfe85248_7859,RIee39148_5108,
        RIe16b378_2597,RIee38608_5100,RIe167b38_2557,RIe164fa0_2526,RIe1622a0_2494,RIfe85950_7864,RIe15f5a0_2462,RIee36010_5073,RIe15c8a0_2430,RIe156ea0_2366,
        RIe1541a0_2334,RIfe85c20_7866,RIe1514a0_2302,RIee34dc8_5060,RIe14e7a0_2270,RIfc861b0_6548,RIe14baa0_2238,RIe148da0_2206,RIe1460a0_2174,RIee343f0_5053,
        RIfe85518_7861,RIfe857e8_7863,RIfe85680_7862,RIe140c40_2114,RIdf3eb48_2090,RIdf3c820_2065,RIdf3a660_2041,RIfc9d4f0_6812,RIee2f698_4998,RIfc52298_5957,
        RIee2d4d8_4974,RIdf35368_1982,RIdf32ed8_1956,RIdf30e80_1933,RIfe85ab8_7865,RIee2b8b8_4954,RIee29f68_4936,RIee28bb8_4922,RIee27970_4909,RIdf2a0d0_1855,
        RIfe84e10_7856,RIdf262f0_1811,RIfe84ca8_7855,RIee27100_4903,RIee26b60_4899,RIfcd32f8_7425,RIee265c0_4895,RIfc9e300_6822,RIdf1f540_1733,RIee25eb8_4890,
        RIfe84b40_7854,RIdf16b70_1635,RIdf13e70_1603,RIdf11170_1571,RIdf0e470_1539,RIdf0b770_1507,RIdf08a70_1475,RIdf05d70_1443,RIdf03070_1411,RIdefd670_1347,
        RIdefa970_1315,RIdef7c70_1283,RIdef4f70_1251,RIdef2270_1219,RIdeef570_1187,RIdeec870_1155,RIdee9b70_1123,RIfec0348_8307,RIfcb54d8_7085,RIee23cf8_4866,
        RIfc54e30_5988,RIfec0078_8305,RIdee2988_1042,RIfec01e0_8306,RIdede770_995,RIfcd7ee8_7479,RIfcd43d8_7437,RIfc88eb0_6580,RIfc9e5d0_6824,RIded9478_936,
        RIded6fe8_910,RIded50f8_888,RIfeab330_8264,RIded03a0_833,RIdecd6a0_801,RIdeca9a0_769,RIdec7ca0_737,RIdeb41a0_513,RIde95f48_321,RIe16dda8_2627,
        RIe159ba0_2398,RIe1433a0_2142,RIdf37d98_2012,RIdf2c3f8_1880,RIdf1cc78_1704,RIdf00370_1379,RIdee6e70_1091,RIdedbbd8_964,RIde7be90_194,RIe19d238_3165,
        RIe19a538_3133,RIf145658_5249,RIe197838_3101,RIf1446e0_5238,RIe194b38_3069,RIe191e38_3037,RIe18f138_3005,RIe189738_2941,RIe186a38_2909,RIf143600_5226,
        RIe183d38_2877,RIf142c28_5219,RIe181038_2845,RIe17e338_2813,RIe17b638_2781,RIf1420e8_5211,RIf140a68_5195,RIf1401f8_5189,RIfebff10_8304,RIf13faf0_5184,
        RIf13ee48_5175,RIee3e2d8_5166,RIee3d1f8_5154,RIee3c118_5142,RIee3b038_5130,RIee39c88_5116,RIfe838f8_7841,RIf1701c8_5735,RIfc5ab00_6054,RIf16e008_5711,
        RIfcb0e88_7035,RIf16caf0_5696,RIe223590_4692,RIf16bce0_5686,RIe220890_4660,RIf16ac00_5674,RIe21db90_4628,RIe218190_4564,RIe215490_4532,RIf16a228_5667,
        RIe212790_4500,RIf168fe0_5654,RIe20fa90_4468,RIf167d98_5641,RIe20cd90_4436,RIe20a090_4404,RIe207390_4372,RIf1670f0_5632,RIf165ea8_5619,RIe202200_4314,
        RIfe83e98_7845,RIf164f30_5608,RIf1643f0_5600,RIfce8310_7664,RIf161df8_5573,RIf15ff08_5551,RIf15e018_5529,RIfe83d30_7844,RIfe84000_7846,RIf15cb00_5514,
        RIf15b5e8_5499,RIf15a508_5487,RIfc887a8_6575,RIf158d20_5470,RIf157970_5456,RIf156cc8_5447,RIfe84438_7849,RIf156020_5438,RIfc51fc8_5955,RIf154568_5419,
        RIe1f51e0_4166,RIf153050_5404,RIf1519d0_5388,RIf150788_5375,RIfe842d0_7848,RIf14f810_5364,RIf14eb68_5355,RIf14dd58_5345,RIfe84168_7847,RIe1eb2f8_4053,
        RIe1e85f8_4021,RIe1e58f8_3989,RIe1e2bf8_3957,RIe1dfef8_3925,RIe1dd1f8_3893,RIe1da4f8_3861,RIe1d77f8_3829,RIe1d1df8_3765,RIe1cf0f8_3733,RIe1cc3f8_3701,
        RIe1c96f8_3669,RIe1c69f8_3637,RIe1c3cf8_3605,RIe1c0ff8_3573,RIe1be2f8_3541,RIf14c840_5330,RIf14b5f8_5317,RIfe83a60_7842,RIfe849d8_7853,RIfc74168_6343,
        RIf149b40_5298,RIfe83bc8_7843,RIfe84708_7851,RIf148d30_5288,RIf147ae8_5275,RIfe84870_7852,RIe1b0900_3386,RIf146fa8_5267,RIf146300_5258,RIfe845a0_7850,
        RIfe83790_7840,RIe1a8638_3293,RIe1a5938_3261,RIe1a2c38_3229,RIe19ff38_3197,RIe18c438_2973,RIe178938_2749,RIe226290_4724,RIe21ae90_4596,RIe204690_4340,
        RIe1fe6f0_4272,RIe1f7aa8_4195,RIe1f05f0_4112,RIe1d4af8_3797,RIe1bb5f8_3509,RIe1ae470_3360,RIe170aa8_2659,RIdec4e38_704,RIdec2138_672,RIee1fc48_4820,
        RIdebf438_640,RIfc49490_5856,RIdebc738_608,RIdeb9a38_576,RIdeb6d38_544,RIfc48ef0_5852,RIdeb1338_480,RIfcd9b08_7499,RIdeae638_448,RIfc8b610_6608,
        RIdea9700_416,RIdea2e00_384,RIde9c500_352,RIee1c9a8_4784,RIee1b8c8_4772,RIfc80918_6485,RIfcdad50_7512,RIfe86e68_7879,RIde8cee8_277,RIfe86d00_7878,
        RIfec0d20_8314,RIde81098_219,RIfc8b8e0_6610,RIfcd2d58_7421,RIfce4530_7620,RIfc8ba48_6611,RIe16b210_2596,RIe1698c0_2578,RIe1679d0_2556,RIe164e38_2525,
        RIe162138_2493,RIee370f0_5085,RIe15f438_2461,RIfc999e0_6770,RIe15c738_2429,RIe156d38_2365,RIe154038_2333,RIfc3f260_5744,RIe151338_2301,RIfc48518_5845,
        RIe14e638_2269,RIfc99e18_6773,RIe14b938_2237,RIe148c38_2205,RIe145f38_2173,RIee34288_5052,RIee33040_5039,RIee31f60_5027,RIfcd99a0_7498,RIfe86b98_7877,
        RIdf3e9e0_2089,RIfe86a30_7876,RIdf3a4f8_2040,RIfcc3470_7244,RIee2f530_4997,RIfc7fdd8_6477,RIee2d370_4973,RIdf35200_1981,RIfec0ff0_8316,RIdf30d18_1932,
        RIfec0e88_8315,RIfcd2a88_7419,RIfc8c858_6621,RIfc47ca8_5839,RIfcd6430_7460,RIdf29f68_1854,RIdf27da8_1830,RIdf26188_1810,RIdf24568_1790,RIfc8cb28_6623,
        RIfcdb188_7515,RIdf22948_1770,RIfc475a0_5834,RIdf21430_1755,RIdf1f3d8_1732,RIfec0bb8_8313,RIfe868c8_7875,RIdf16a08_1634,RIdf13d08_1602,RIdf11008_1570,
        RIdf0e308_1538,RIdf0b608_1506,RIdf08908_1474,RIdf05c08_1442,RIdf02f08_1410,RIdefd508_1346,RIdefa808_1314,RIdef7b08_1282,RIdef4e08_1250,RIdef2108_1218,
        RIdeef408_1186,RIdeec708_1154,RIdee9a08_1122,RIee254e0_4883,RIee246d0_4873,RIee23b90_4865,RIee231b8_4858,RIfe86fd0_7880,RIdee2820_1041,RIdee0930_1019,
        RIdede608_994,RIfc55da8_5999,RIfc98a68_6759,RIfcc3038_7241,RIfc464c0_5822,RIded9310_935,RIded6e80_909,RIded4f90_887,RIded2b00_861,RIded0238_832,
        RIdecd538_800,RIdeca838_768,RIdec7b38_736,RIdeb4038_512,RIde95c00_320,RIe16dc40_2626,RIe159a38_2397,RIe143238_2141,RIdf37c30_2011,RIdf2c290_1879,
        RIdf1cb10_1703,RIdf00208_1378,RIdee6d08_1090,RIdedba70_963,RIde7bb48_193,RIe19d0d0_3164,RIe19a3d0_3132,RIf1454f0_5248,RIe1976d0_3100,RIf144578_5237,
        RIe1949d0_3068,RIe191cd0_3036,RIe18efd0_3004,RIe1895d0_2940,RIe1868d0_2908,RIf143498_5225,RIe183bd0_2876,RIfc51758_5949,RIe180ed0_2844,RIe17e1d0_2812,
        RIe17b4d0_2780,RIfc9b060_6786,RIfc9ee40_6830,RIe176e80_2730,RIe175800_2714,RIfcb70f8_7105,RIfce0cf0_7580,RIfcc4280_7254,RIfcba7d0_7144,RIee3bfb0_5141,
        RIee3aed0_5129,RIee39b20_5115,RIe173370_2688,RIf170060_5734,RIf16f3b8_5725,RIf16dea0_5710,RIf16d4c8_5703,RIf16c988_5695,RIe223428_4691,RIf16bb78_5685,
        RIe220728_4659,RIf16aa98_5673,RIe21da28_4627,RIe218028_4563,RIe215328_4531,RIf16a0c0_5666,RIe212628_4499,RIf168e78_5653,RIe20f928_4467,RIf167c30_5640,
        RIe20cc28_4435,RIe209f28_4403,RIe207228_4371,RIf166f88_5631,RIf165d40_5618,RIfec0618_8309,RIfe86760_7874,RIfc52b08_5963,RIf164288_5599,RIf163310_5588,
        RIf161c90_5572,RIf15fda0_5550,RIf15deb0_5528,RIfe865f8_7873,RIfe85d88_7867,RIf15c998_5513,RIf15b480_5498,RIf15a3a0_5486,RIf159b30_5480,RIfc83348_6515,
        RIfc4ade0_5874,RIfc89720_6586,RIe1f9f38_4221,RIfc4ac78_5873,RIfc9f110_6832,RIfc4ab10_5872,RIe1f5078_4165,RIf152ee8_5403,RIfc899f0_6588,RIf150620_5374,
        RIe1f2eb8_4141,RIf14f6a8_5363,RIf14ea00_5354,RIf14dbf0_5344,RIe1edbc0_4082,RIe1eb190_4052,RIe1e8490_4020,RIe1e5790_3988,RIe1e2a90_3956,RIe1dfd90_3924,
        RIe1dd090_3892,RIe1da390_3860,RIe1d7690_3828,RIe1d1c90_3764,RIe1cef90_3732,RIe1cc290_3700,RIe1c9590_3668,RIe1c6890_3636,RIe1c3b90_3604,RIe1c0e90_3572,
        RIe1be190_3540,RIf14c6d8_5329,RIf14b490_5316,RIfe85ef0_7868,RIfe86490_7872,RIf14a248_5303,RIfc819f8_6497,RIfec0a50_8312,RIfe861c0_7870,RIf148bc8_5287,
        RIf147980_5274,RIfe86328_7871,RIfec0780_8310,RIfcbb478_7153,RIf146198_5257,RIfe86058_7869,RIfec08e8_8311,RIe1a84d0_3292,RIe1a57d0_3260,RIe1a2ad0_3228,
        RIe19fdd0_3196,RIe18c2d0_2972,RIe1787d0_2748,RIe226128_4723,RIe21ad28_4595,RIe204528_4339,RIe1fe588_4271,RIe1f7940_4194,RIe1f0488_4111,RIe1d4990_3796,
        RIe1bb490_3508,RIe1ae308_3359,RIe170940_2658,RIdec53d8_708,RIdec26d8_676,RIee20080_4823,RIdebf9d8_644,RIee1f3d8_4814,RIdebccd8_612,RIdeb9fd8_580,
        RIdeb72d8_548,RIee1ee38_4810,RIdeb18d8_484,RIee1e898_4806,RIdeaebd8_452,RIee1da88_4796,RIdeaa420_420,RIdea3b20_388,RIde9d220_356,RIee1cde0_4787,
        RIee1bd00_4775,RIee1b490_4769,RIfcd8a28_7487,RIde91088_297,RIde8d8c0_280,RIfe7dac0_7774,RIfe7d958_7773,RIee1a518_4758,RIee19e10_4753,RIee19b40_4751,
        RIfc768c8_6371,RIfcd05f8_7393,RIfe7dd90_7776,RIee38770_5101,RIfe7dc28_7775,RIe1653d8_2529,RIe1626d8_2497,RIee373c0_5087,RIe15f9d8_2465,RIee362e0_5075,
        RIe15ccd8_2433,RIe1572d8_2369,RIe1545d8_2337,RIfe7def8_7777,RIe1518d8_2305,RIfebdeb8_8281,RIe14ebd8_2273,RIfc649e8_6167,RIe14bed8_2241,RIe1491d8_2209,
        RIe1464d8_2177,RIfe7d7f0_7772,RIfe7d688_7771,RIee32230_5029,RIfceb9e8_7703,RIfebdd50_8280,RIfe7d520_7770,RIfebdbe8_8279,RIfe7d3b8_7769,RIfc734c0_6334,
        RIee2f968_5000,RIfccfab8_7385,RIee2d7a8_4976,RIdf357a0_1985,RIdf33310_1959,RIdf312b8_1936,RIdf2f0f8_1912,RIee2bcf0_4957,RIee2a238_4938,RIee28e88_4924,
        RIee27c40_4911,RIfe7ce18_7765,RIfe7ccb0_7764,RIfe7cf80_7766,RIfe7cb48_7763,RIee27268_4904,RIee26e30_4901,RIee26890_4897,RIfcaa0d8_6957,RIee262f0_4893,
        RIfe7d250_7768,RIee26020_4891,RIfe7d0e8_7767,RIdf16fa8_1638,RIdf142a8_1606,RIdf115a8_1574,RIdf0e8a8_1542,RIdf0bba8_1510,RIdf08ea8_1478,RIdf061a8_1446,
        RIdf034a8_1414,RIdefdaa8_1350,RIdefada8_1318,RIdef80a8_1286,RIdef53a8_1254,RIdef26a8_1222,RIdeef9a8_1190,RIdeecca8_1158,RIdee9fa8_1126,RIee25648_4884,
        RIee249a0_4875,RIfebe020_8282,RIee23488_4860,RIfebe2f0_8284,RIfebe188_8283,RIfe7e1c8_7779,RIfe7e060_7778,RIfcbf7f8_7201,RIfc7aae0_6418,RIfc787b8_6393,
        RIfc618b0_6132,RIded98b0_939,RIded72b8_912,RIded5530_891,RIded2dd0_863,RIded07d8_836,RIdecdad8_804,RIdecadd8_772,RIdec80d8_740,RIdeb45d8_516,
        RIde96920_324,RIe16e1e0_2630,RIe159fd8_2401,RIe1437d8_2145,RIdf381d0_2015,RIdf2c830_1883,RIdf1d0b0_1707,RIdf007a8_1382,RIdee72a8_1094,RIdedc010_967,
        RIde7c868_197,RIe19d670_3168,RIe19a970_3136,RIfe7b630_7748,RIe197c70_3104,RIfe7b4c8_7747,RIe194f70_3072,RIe192270_3040,RIe18f570_3008,RIe189b70_2944,
        RIe186e70_2912,RIfe7b360_7746,RIe184170_2880,RIfe7b1f8_7745,RIe181470_2848,RIe17e770_2816,RIe17ba70_2784,RIf1423b8_5213,RIf140ea0_5198,RIf140360_5190,
        RIfe7b798_7749,RIf13fc58_5185,RIf13f280_5178,RIfc79460_6402,RIee3d4c8_5156,RIfe7b090_7744,RIfe7af28_7743,RIee39df0_5117,RIe1737a8_2691,RIfe7adc0_7742,
        RIfe7ac58_7741,RIf16e440_5714,RIfcb20d0_7048,RIfe7bd38_7753,RIe2239c8_4695,RIf16be48_5687,RIe220cc8_4663,RIf16aed0_5676,RIe21dfc8_4631,RIe2185c8_4567,
        RIe2158c8_4535,RIfebd7b0_8276,RIe212bc8_4503,RIfebd648_8275,RIe20fec8_4471,RIfe7b900_7750,RIe20d1c8_4439,RIe20a4c8_4407,RIe2077c8_4375,RIf167258_5633,
        RIf166178_5621,RIe2024d0_4316,RIfe7bbd0_7752,RIf165368_5611,RIf1646c0_5602,RIfcd0a30_7396,RIf1620c8_5575,RIf1601d8_5553,RIf15e2e8_5531,RIfe7ba68_7751,
        RIfe7bea0_7754,RIf15cdd0_5516,RIf15b8b8_5501,RIf15a7d8_5489,RIfca4840_6894,RIf158ff0_5472,RIf157c40_5458,RIf156f98_5449,RIfe7c170_7756,RIf156458_5441,
        RIf155918_5433,RIf1549a0_5422,RIe1f54b0_4168,RIfe7c008_7755,RIf151b38_5389,RIf150bc0_5378,RIe1f32f0_4144,RIf14fae0_5366,RIf14ee38_5357,RIf14e028_5347,
        RIe1edff8_4085,RIe1eb730_4056,RIe1e8a30_4024,RIe1e5d30_3992,RIe1e3030_3960,RIe1e0330_3928,RIe1dd630_3896,RIe1da930_3864,RIe1d7c30_3832,RIe1d2230_3768,
        RIe1cf530_3736,RIe1cc830_3704,RIe1c9b30_3672,RIe1c6e30_3640,RIe1c4130_3608,RIe1c1430_3576,RIe1be730_3544,RIf14cb10_5332,RIf14b8c8_5319,RIfebda80_8278,
        RIfe7c878_7761,RIf14a680_5306,RIfe7c2d8_7757,RIfe7c9e0_7762,RIfe7c440_7758,RIf149000_5290,RIf147db8_5277,RIe1b2688_3407,RIfebd918_8277,RIfe7c5a8_7759,
        RIf146738_5261,RIfe7c710_7760,RIe1aad98_3321,RIe1a8a70_3296,RIe1a5d70_3264,RIe1a3070_3232,RIe1a0370_3200,RIe18c870_2976,RIe178d70_2752,RIe2266c8_4727,
        RIe21b2c8_4599,RIe204ac8_4343,RIe1feb28_4275,RIe1f7ee0_4198,RIe1f0a28_4115,RIe1d4f30_3800,RIe1bba30_3512,RIe1ae8a8_3363,RIe170ee0_2662,RIdec5270_707,
        RIdec2570_675,RIee1ff18_4822,RIdebf870_643,RIfe7f848_7795,RIdebcb70_611,RIdeb9e70_579,RIdeb7170_547,RIfe7fc80_7798,RIdeb1770_483,RIfca5d58_6909,
        RIdeaea70_451,RIfcaf808_7019,RIdeaa0d8_419,RIdea37d8_387,RIde9ced8_355,RIfcdc3d0_7528,RIfcce438_7369,RIfcb0a50_7032,RIfc75680_6358,RIde90d40_296,
        RIfe7f9b0_7796,RIde89720_260,RIde85580_240,RIde81728_221,RIfc52f40_5966,RIfc82100_6502,RIfca7108_6923,RIfe7fb18_7797,RIe16b648_2599,RIe169a28_2579,
        RIe167ca0_2558,RIe165270_2528,RIe162570_2496,RIee37258_5086,RIe15f870_2464,RIee36178_5074,RIe15cb70_2432,RIe157170_2368,RIe154470_2336,RIfc86fc0_6558,
        RIe151770_2304,RIfc4eff8_5921,RIe14ea70_2272,RIfce1290_7584,RIe14bd70_2240,RIe149070_2208,RIe146370_2176,RIee34558_5054,RIee331a8_5040,RIee320c8_5028,
        RIee31150_5017,RIfe800b8_7801,RIfe7ff50_7800,RIdf3caf0_2067,RIfe7fde8_7799,RIfcc8330_7300,RIee2f800_4999,RIfca0d30_6852,RIee2d640_4975,RIdf35638_1984,
        RIdf331a8_1958,RIdf31150_1935,RIdf2ef90_1911,RIee2bb88_4956,RIee2a0d0_4937,RIee28d20_4923,RIfe7f578_7793,RIdf2a238_1856,RIdf27f10_1831,RIfe7f6e0_7794,
        RIdf246d0_1791,RIfcce9d8_7373,RIfc63638_6153,RIdf22c18_1772,RIfc62990_6144,RIdf21700_1757,RIdf1f810_1735,RIfeaa958_8257,RIdf19168_1662,RIdf16e40_1637,
        RIdf14140_1605,RIdf11440_1573,RIdf0e740_1541,RIdf0ba40_1509,RIdf08d40_1477,RIdf06040_1445,RIdf03340_1413,RIdefd940_1349,RIdefac40_1317,RIdef7f40_1285,
        RIdef5240_1253,RIdef2540_1221,RIdeef840_1189,RIdeecb40_1157,RIdee9e40_1125,RIfcb7800_7110,RIee24838_4874,RIfc4cb68_5895,RIee23320_4859,RIfe80388_7803,
        RIdee2c58_1044,RIfe80220_7802,RIdedea40_997,RIfc98900_6758,RIee223a8_4848,RIfcc8600_7302,RIee212c8_4836,RIded9748_938,RIfe804f0_7804,RIded53c8_890,
        RIded2c68_862,RIded0670_835,RIdecd970_803,RIdecac70_771,RIdec7f70_739,RIdeb4470_515,RIde965d8_323,RIe16e078_2629,RIe159e70_2400,RIe143670_2144,
        RIdf38068_2014,RIdf2c6c8_1882,RIdf1cf48_1706,RIdf00640_1381,RIdee7140_1093,RIdedbea8_966,RIde7c520_196,RIe19d508_3167,RIe19a808_3135,RIfe7ee70_7788,
        RIe197b08_3103,RIfe7efd8_7789,RIe194e08_3071,RIe192108_3039,RIe18f408_3007,RIe189a08_2943,RIe186d08_2911,RIf143768_5227,RIe184008_2879,RIfc4bbf0_5884,
        RIe181308_2847,RIe17e608_2815,RIe17b908_2783,RIfe7f410_7792,RIf140d38_5197,RIe176fe8_2731,RIe175ad0_2716,RIfe7f2a8_7791,RIf13f118_5177,RIee3e440_5167,
        RIee3d360_5155,RIee3c280_5143,RIee3b1a0_5131,RIfe7f140_7790,RIe173640_2690,RIf170330_5736,RIf16f520_5726,RIf16e2d8_5713,RIf16d630_5704,RIfe7ea38_7785,
        RIe223860_4694,RIfc9c410_6800,RIe220b60_4662,RIfcb8340_7118,RIe21de60_4630,RIe218460_4566,RIe215760_4534,RIfc9cc80_6806,RIe212a60_4502,RIfc4ddb0_5908,
        RIe20fd60_4470,RIfc873f8_6561,RIe20d060_4438,RIe20a360_4406,RIe207660_4374,RIfc86750_6552,RIfc4e4b8_5913,RIe202368_4315,RIe200a18_4297,RIf165200_5610,
        RIf164558_5601,RIf163478_5589,RIf161f60_5574,RIf160070_5552,RIf15e180_5530,RIe1fcc38_4253,RIe1fb9f0_4240,RIf15cc68_5515,RIf15b750_5500,RIf15a670_5488,
        RIf159c98_5481,RIf158e88_5471,RIf157ad8_5457,RIf156e30_5448,RIfe7e768_7783,RIf1562f0_5440,RIf1557b0_5432,RIf154838_5421,RIfe7e8d0_7784,RIf1531b8_5405,
        RIfc52400_5958,RIf150a58_5377,RIe1f3188_4143,RIf14f978_5365,RIf14ecd0_5356,RIf14dec0_5346,RIe1ede90_4084,RIe1eb5c8_4055,RIe1e88c8_4023,RIe1e5bc8_3991,
        RIe1e2ec8_3959,RIe1e01c8_3927,RIe1dd4c8_3895,RIe1da7c8_3863,RIe1d7ac8_3831,RIe1d20c8_3767,RIe1cf3c8_3735,RIe1cc6c8_3703,RIe1c99c8_3671,RIe1c6cc8_3639,
        RIe1c3fc8_3607,RIe1c12c8_3575,RIe1be5c8_3543,RIf14c9a8_5331,RIf14b760_5318,RIfe7ed08_7787,RIfe7e600_7782,RIf14a518_5305,RIfca1f78_6865,RIfe7eba0_7786,
        RIfe7e498_7781,RIf148e98_5289,RIf147c50_5276,RIfe7e330_7780,RIe1b0a68_3387,RIf147278_5269,RIf1465d0_5260,RIe1ac418_3337,RIe1aac30_3320,RIe1a8908_3295,
        RIe1a5c08_3263,RIe1a2f08_3231,RIe1a0208_3199,RIe18c708_2975,RIe178c08_2751,RIe226560_4726,RIe21b160_4598,RIe204960_4342,RIe1fe9c0_4274,RIe1f7d78_4197,
        RIe1f08c0_4114,RIe1d4dc8_3799,RIe1bb8c8_3511,RIe1ae740_3362,RIe170d78_2661,RIdec56a8_710,RIdec29a8_678,RIfc54020_5978,RIdebfca8_646,RIee1f540_4815,
        RIdebcfa8_614,RIdeba2a8_582,RIdeb75a8_550,RIfc4fe08_5931,RIdeb1ba8_486,RIfc6b630_6244,RIdeaeea8_454,RIfc6a118_6229,RIdeaaab0_422,RIdea41b0_390,
        RIde9d8b0_358,RIfc69ce0_6226,RIee1be68_4776,RIfc653c0_6174,RIee1ac20_4763,RIde91718_299,RIde8df50_282,RIde89db0_262,RIde85c10_242,RIde81db8_223,
        RIfca76a8_6927,RIfcca4f0_7324,RIfc4ce38_5897,RIfc6b360_6242,RIe16b918_2601,RIe169cf8_2581,RIe167f70_2560,RIe1656a8_2531,RIe1629a8_2499,RIee37690_5089,
        RIe15fca8_2467,RIfce93f0_7676,RIe15cfa8_2435,RIe1575a8_2371,RIe1548a8_2339,RIee35908_5068,RIe151ba8_2307,RIee34f30_5061,RIe14eea8_2275,RIfce32e8_7607,
        RIe14c1a8_2243,RIe1494a8_2211,RIe1467a8_2179,RIfcde2c0_7550,RIfc687c8_6211,RIfca9160_6946,RIfcb1590_7040,RIe141078_2117,RIdf3ef80_2093,RIdf3cdc0_2069,
        RIfebeb60_8290,RIfc64448_6163,RIee2fad0_5001,RIfca7978_6929,RIfc676e8_6199,RIdf35a70_1987,RIdf335e0_1961,RIdf31420_1937,RIdf2f3c8_1914,RIfccef78_7377,
        RIfca6fa0_6922,RIfc62558_6141,RIfc61fb8_6137,RIfe81b70_7820,RIdf281e0_1833,RIfe81cd8_7821,RIdf249a0_1793,RIfc44300_5798,RIfcafc40_7022,RIdf22ee8_1774,
        RIfcaac18_6965,RIdf219d0_1759,RIdf1fae0_1737,RIdf1b1c0_1685,RIdf19438_1664,RIdf17278_1640,RIdf14578_1608,RIdf11878_1576,RIdf0eb78_1544,RIdf0be78_1512,
        RIdf09178_1480,RIdf06478_1448,RIdf03778_1416,RIdefdd78_1352,RIdefb078_1320,RIdef8378_1288,RIdef5678_1256,RIdef2978_1224,RIdeefc78_1192,RIdeecf78_1160,
        RIdeea278_1128,RIfc611a8_6127,RIfc61a18_6133,RIfca65c8_6915,RIfca6b68_6919,RIdee4b48_1066,RIdee2dc0_1045,RIdee0c00_1021,RIdedeba8_998,RIfc626c0_6142,
        RIfc738f8_6337,RIfcb31b0_7060,RIee21430_4837,RIded9a18_940,RIded7588_914,RIded5698_892,RIded30a0_865,RIded0aa8_838,RIdecdda8_806,RIdecb0a8_774,
        RIdec83a8_742,RIdeb48a8_518,RIde96fb0_326,RIe16e4b0_2632,RIe15a2a8_2403,RIe143aa8_2147,RIdf384a0_2017,RIdf2cb00_1885,RIdf1d380_1709,RIdf00a78_1384,
        RIdee7578_1096,RIdedc2e0_969,RIde7cef8_199,RIe19d940_3170,RIe19ac40_3138,RIfc64880_6166,RIe197f40_3106,RIf144848_5239,RIe195240_3074,RIe192540_3042,
        RIe18f840_3010,RIe189e40_2946,RIe187140_2914,RIf143a38_5229,RIe184440_2882,RIfc6f140_6286,RIe181740_2850,RIe17ea40_2818,RIe17bd40_2786,RIfc64f88_6171,
        RIf141008_5199,RIe177150_2732,RIfe81738_7817,RIfccabf8_7329,RIf13f3e8_5179,RIfca81e8_6935,RIee3d630_5157,RIfc66068_6183,RIfc6ed08_6283,RIfcdde88_7547,
        RIe173a78_2693,RIfc66338_6185,RIfc6eba0_6282,RIfc664a0_6186,RIfcacdd8_6989,RIfe81468_7815,RIe223c98_4697,RIfc66d10_6192,RIe220f98_4665,RIf16b038_5677,
        RIe21e298_4633,RIe218898_4569,RIe215b98_4537,RIfc3fc38_5751,RIe212e98_4505,RIfc67850_6200,RIe210198_4473,RIf167f00_5642,RIe20d498_4441,RIe20a798_4409,
        RIe207a98_4377,RIfcacb08_6987,RIfcac9a0_6986,RIfea8900_8234,RIfe818a0_7818,RIfca8a58_6941,RIfccad60_7330,RIfcac838_6985,RIfc67418_6197,RIf160340_5554,
        RIf15e450_5532,RIfe81a08_7819,RIfe81300_7814,RIfc6dac0_6270,RIf15ba20_5502,RIfc6d958_6269,RIfc6d7f0_6268,RIfc587d8_6029,RIfc6cf80_6262,RIfc6d3b8_6265,
        RIfe815d0_7816,RIfc6d520_6266,RIfcabe60_6978,RIfc6d0e8_6263,RIe1f5780_4170,RIfc6c5a8_6255,RIfc68d68_6215,RIfc68c00_6214,RIe1f3458_4145,RIfc68a98_6213,
        RIfccb8a0_7338,RIfca9b38_6953,RIe1ee160_4086,RIe1eba00_4058,RIe1e8d00_4026,RIe1e6000_3994,RIe1e3300_3962,RIe1e0600_3930,RIe1dd900_3898,RIe1dac00_3866,
        RIe1d7f00_3834,RIe1d2500_3770,RIe1cf800_3738,RIe1ccb00_3706,RIe1c9e00_3674,RIe1c7100_3642,RIe1c4400_3610,RIe1c1700_3578,RIe1bea00_3546,RIfc6bbd0_6248,
        RIfcdd348_7539,RIe1b9438_3485,RIe1b73e0_3462,RIfcab5f0_6972,RIfccbb70_7340,RIe1b5220_3438,RIe1b3e70_3424,RIfc6c9e0_6258,RIfcab488_6971,RIfea7dc0_8226,
        RIe1b0bd0_3388,RIfc6ce18_6261,RIfcabfc8_6979,RIe1ac580_3338,RIe1aaf00_3322,RIe1a8d40_3298,RIe1a6040_3266,RIe1a3340_3234,RIe1a0640_3202,RIe18cb40_2978,
        RIe179040_2754,RIe226998_4729,RIe21b598_4601,RIe204d98_4345,RIe1fedf8_4277,RIe1f81b0_4200,RIe1f0cf8_4117,RIe1d5200_3802,RIe1bbd00_3514,RIe1aeb78_3365,
        RIe1711b0_2664,RIdec5540_709,RIdec2840_677,RIfcc4dc0_7262,RIdebfb40_645,RIfc9d7c0_6814,RIdebce40_613,RIdeba140_581,RIdeb7440_549,RIfc4d978_5905,
        RIdeb1a40_485,RIfc9dbf8_6817,RIdeaed40_453,RIfcb8610_7120,RIdeaa768_421,RIdea3e68_389,RIde9d568_357,RIfc50678_5937,RIfc507e0_5938,RIfc9dec8_6819,
        RIfc853a0_6538,RIde913d0_298,RIde8dc08_281,RIde89a68_261,RIde858c8_241,RIde81a70_222,RIfc84860_6530,RIfc50948_5939,RIfc84c98_6533,RIfcb7da0_7114,
        RIe16b7b0_2600,RIe169b90_2580,RIe167e08_2559,RIe165540_2530,RIe162840_2498,RIee37528_5088,RIe15fb40_2466,RIfcb5be0_7090,RIe15ce40_2434,RIe157440_2370,
        RIe154740_2338,RIfcd35c8_7427,RIe151a40_2306,RIfc53a80_5974,RIe14ed40_2274,RIfcc6170_7276,RIe14c040_2242,RIe149340_2210,RIe146640_2178,RIfc7f130_6468,
        RIee33310_5041,RIfcb4f38_7081,RIfc47f78_5841,RIe140f10_2116,RIdf3ee18_2092,RIdf3cc58_2068,RIdf3a7c8_2042,RIfc7fc70_6476,RIfcd27b8_7417,RIfca1000_6854,
        RIfcc6b48_7283,RIdf35908_1986,RIdf33478_1960,RIfebe9f8_8289,RIdf2f260_1913,RIfcb7968_7111,RIee2a3a0_4939,RIfc51050_5944,RIfcd3fa0_7434,RIdf2a3a0_1857,
        RIdf28078_1832,RIfe81198_7813,RIdf24838_1792,RIfc84428_6527,RIfce7ed8_7661,RIdf22d80_1773,RIfc515f0_5948,RIdf21868_1758,RIdf1f978_1736,RIdf1b058_1684,
        RIdf192d0_1663,RIdf17110_1639,RIdf14410_1607,RIdf11710_1575,RIdf0ea10_1543,RIdf0bd10_1511,RIdf09010_1479,RIdf06310_1447,RIdf03610_1415,RIdefdc10_1351,
        RIdefaf10_1319,RIdef8210_1287,RIdef5510_1255,RIdef2810_1223,RIdeefb10_1191,RIdeece10_1159,RIdeea110_1127,RIfc7e1b8_6457,RIfca19d8_6861,RIfc7dab0_6452,
        RIfc7e488_6459,RIdee49e0_1065,RIfe80d60_7810,RIfeabba0_8270,RIfe80bf8_7809,RIfcb3750_7064,RIfce9f30_7684,RIfc7e5f0_6460,RIfc56a50_6008,RIfe81030_7812,
        RIded7420_913,RIfe80ec8_7811,RIded2f38_864,RIded0940_837,RIdecdc40_805,RIdecaf40_773,RIdec8240_741,RIdeb4740_517,RIde96c68_325,RIe16e348_2631,
        RIe15a140_2402,RIe143940_2146,RIdf38338_2016,RIdf2c998_1884,RIdf1d218_1708,RIdf00910_1383,RIdee7410_1095,RIdedc178_968,RIde7cbb0_198,RIe19d7d8_3169,
        RIe19aad8_3137,RIfcc2d68_7239,RIe197dd8_3105,RIfc5c5b8_6073,RIe1950d8_3073,RIe1923d8_3041,RIe18f6d8_3009,RIe189cd8_2945,RIe186fd8_2913,RIf1438d0_5228,
        RIe1842d8_2881,RIfc5b370_6060,RIe1815d8_2849,RIe17e8d8_2817,RIe17bbd8_2785,RIfcbb748_7155,RIfc59480_6038,RIfcbbce8_7159,RIe175c38_2717,RIfcdb890_7520,
        RIfc59b88_6043,RIfc8ada0_6602,RIfcb5eb0_7092,RIfc57c98_6021,RIfc57158_6013,RIfc58aa8_6031,RIe173910_2692,RIfcc62d8_7277,RIfc8a968_6599,RIfc57428_6015,
        RIfc56d20_6010,RIfc408e0_5760,RIe223b30_4696,RIfc82970_6508,RIe220e30_4664,RIfcecc30_7716,RIe21e130_4632,RIe218730_4568,RIe215a30_4536,RIfc3fad0_5750,
        RIe212d30_4504,RIf169148_5655,RIe210030_4472,RIfc545c0_5982,RIe20d330_4440,RIe20a630_4408,RIe207930_4376,RIfc88d48_6579,RIfc4bec0_5886,RIe202638_4317,
        RIe200b80_4298,RIfc88910_6576,RIfc4c190_5888,RIfc4c2f8_5889,RIfcba398_7141,RIfcd4270_7436,RIfcba0c8_7139,RIe1fcda0_4254,RIe1fbb58_4241,RIfc53d50_5976,
        RIfc9b768_6791,RIfc537b0_5972,RIfc4c5c8_5891,RIfc9e468_6823,RIf157da8_5459,RIfcb9f60_7138,RIe1fa208_4223,RIfc849c8_6531,RIfc529a0_5962,RIfc9f6b0_6836,
        RIe1f5618_4169,RIf153320_5406,RIfcc4988_7259,RIf150d28_5379,RIfebe458_8285,RIfc87f38_6569,RIfcb7f08_7115,RIf14e190_5348,RIfe80658_7805,RIe1eb898_4057,
        RIe1e8b98_4025,RIe1e5e98_3993,RIe1e3198_3961,RIe1e0498_3929,RIe1dd798_3897,RIe1daa98_3865,RIe1d7d98_3833,RIe1d2398_3769,RIe1cf698_3737,RIe1cc998_3705,
        RIe1c9c98_3673,RIe1c6f98_3641,RIe1c4298_3609,RIe1c1598_3577,RIe1be898_3545,RIf14cc78_5333,RIf14ba30_5320,RIe1b92d0_3484,RIe1b7278_3461,RIf14a7e8_5307,
        RIf149ca8_5299,RIfebe5c0_8286,RIfe807c0_7806,RIfc50510_5936,RIfce4f08_7627,RIfe80a90_7808,RIfebe890_8288,RIfc9cde8_6807,RIfc87560_6562,RIfe80928_7807,
        RIfebe728_8287,RIe1a8bd8_3297,RIe1a5ed8_3265,RIe1a31d8_3233,RIe1a04d8_3201,RIe18c9d8_2977,RIe178ed8_2753,RIe226830_4728,RIe21b430_4600,RIe204c30_4344,
        RIe1fec90_4276,RIe1f8048_4199,RIe1f0b90_4116,RIe1d5098_3801,RIe1bbb98_3513,RIe1aea10_3364,RIe171048_2663,RIdec5978_712,RIdec2c78_680,RIfc8aad0_6600,
        RIdebff78_648,RIfc8ac38_6601,RIdebd278_616,RIdeba578_584,RIdeb7878_552,RIfc40e80_5764,RIdeb1e78_488,RIfcdaeb8_7513,RIdeaf178_456,RIee1dbf0_4797,
        RIdeab140_424,RIdea4840_392,RIde9df40_360,RIfc8b070_6604,RIfcc38a8_7247,RIfc807b0_6484,RIfcbb8b0_7156,RIde91a60_300,RIde8e298_283,RIde8a440_264,
        RIde862a0_244,RIde82100_224,RIfcbbb80_7158,RIfc8c150_6616,RIfcbbfb8_7161,RIfc54458_5981,RIe16bbe8_2603,RIfc8c2b8_6617,RIe168240_2562,RIe165978_2533,
        RIe162c78_2501,RIee37960_5091,RIe15ff78_2469,RIfcd6b38_7465,RIe15d278_2437,RIe157878_2373,RIe154b78_2341,RIfc8e5e0_6642,RIe151e78_2309,RIfcb4290_7072,
        RIe14f178_2277,RIfc56ff0_6012,RIe14c478_2245,RIe149778_2213,RIe146a78_2181,RIee346c0_5055,RIee335e0_5043,RIee32398_5030,RIee31420_5019,RIe141348_2119,
        RIe13f020_2094,RIfec16f8_8321,RIdf3a930_2043,RIfce3e28_7615,RIfc56780_6006,RIfcb4128_7071,RIfce2eb0_7604,RIdf35d40_1989,RIfe88218_7893,RIdf316f0_1939,
        RIdf2f698_1916,RIfc7f9a0_6474,RIfce4260_7618,RIfcd62c8_7459,RIfce9990_7680,RIdf2a670_1859,RIdf284b0_1835,RIdf26728_1814,RIdf24c70_1795,RIfc7ecf8_6465,
        RIfcc31a0_7242,RIfc99008_6763,RIfc46e98_5829,RIfce2a78_7601,RIdf1fdb0_1739,RIfcc6e18_7285,RIdf19708_1666,RIdf17548_1642,RIdf14848_1610,RIdf11b48_1578,
        RIdf0ee48_1546,RIdf0c148_1514,RIdf09448_1482,RIdf06748_1450,RIdf03a48_1418,RIdefe048_1354,RIdefb348_1322,RIdef8648_1290,RIdef5948_1258,RIdef2c48_1226,
        RIdeeff48_1194,RIdeed248_1162,RIdeea548_1130,RIfcd9130_7492,RIfc7cb38_6441,RIfc97af0_6748,RIfcb3e58_7069,RIdee4e18_1068,RIdee3090_1047,RIdee0ed0_1023,
        RIfe88380_7894,RIfc97dc0_6750,RIfcc2930_7236,RIfcd9298_7493,RIfc7c868_6439,RIded9ce8_942,RIded76f0_915,RIded5968_894,RIded3370_867,RIded0d78_840,
        RIdece078_808,RIdecb378_776,RIdec8678_744,RIdeb4b78_520,RIde97640_328,RIe16e780_2634,RIe15a578_2405,RIe143d78_2149,RIdf38770_2019,RIdf2cdd0_1887,
        RIdf1d650_1711,RIdf00d48_1386,RIdee7848_1098,RIdedc5b0_971,RIde7d588_201,RIe19dc10_3172,RIe19af10_3140,RIfec1590_8320,RIe198210_3108,RIfec1428_8319,
        RIe195510_3076,RIe192810_3044,RIe18fb10_3012,RIe18a110_2948,RIe187410_2916,RIfec12c0_8318,RIe184710_2884,RIfc88370_6572,RIe181a10_2852,RIe17ed10_2820,
        RIe17c010_2788,RIfc6ccb0_6260,RIfc5f858_6109,RIfca88f0_6940,RIe175f08_2719,RIfc81020_6490,RIfcc6008_7275,RIfc4ea58_5917,RIfc42140_5774,RIfca3b98_6885,
        RIfc5ac68_6055,RIfc984c8_6755,RIe173d48_2695,RIfc9b330_6788,RIf16f688_5727,RIfc42410_5776,RIfc5f588_6107,RIfe880b0_7892,RIe223f68_4699,RIf16bfb0_5688,
        RIe221268_4667,RIfc86cf0_6556,RIe21e568_4635,RIe218b68_4571,RIe215e68_4539,RIfe87de0_7890,RIe213168_4507,RIf1692b0_5656,RIe210468_4475,RIfcdf670_7564,
        RIe20d768_4443,RIe20aa68_4411,RIe207d68_4379,RIfca6460_6914,RIf1662e0_5622,RIe202908_4319,RIfe87b10_7888,RIfc58c10_6032,RIfc50ab0_5940,RIfccd790_7360,
        RIfccd1f0_7356,RIf160610_5556,RIf15e720_5534,RIfe87c78_7889,RIfe87f48_7891,RIfce7668_7655,RIfc86480_6550,RIfcd2218_7413,RIfcb01e0_7026,RIfc47b40_5838,
        RIfc84158_6525,RIfc4b920_5882,RIe1fa4d8_4225,RIfc4ba88_5883,RIfcb7530_7108,RIfcd58f0_7452,RIe1f5a50_4172,RIf153488_5407,RIf151ca0_5390,RIfc51e60_5954,
        RIe1f3728_4147,RIfc9aef8_6785,RIfcbaaa0_7146,RIfc52130_5956,RIe1ee430_4088,RIe1ebcd0_4060,RIe1e8fd0_4028,RIe1e62d0_3996,RIe1e35d0_3964,RIe1e08d0_3932,
        RIe1ddbd0_3900,RIe1daed0_3868,RIe1d81d0_3836,RIe1d27d0_3772,RIe1cfad0_3740,RIe1ccdd0_3708,RIe1ca0d0_3676,RIe1c73d0_3644,RIe1c46d0_3612,RIe1c19d0_3580,
        RIe1becd0_3548,RIfce0b88_7579,RIfc82808_6507,RIe1b9708_3487,RIe1b76b0_3464,RIfcd5bc0_7454,RIfcb69f0_7100,RIe1b54f0_3440,RIe1b4140_3426,RIfc89f90_6592,
        RIfce9af8_7681,RIe1b2958_3409,RIe1b0ea0_3390,RIfc4a138_5865,RIfc8a260_6594,RIe1ac850_3340,RIe1ab1d0_3324,RIe1a9010_3300,RIe1a6310_3268,RIe1a3610_3236,
        RIe1a0910_3204,RIe18ce10_2980,RIe179310_2756,RIe226c68_4731,RIe21b868_4603,RIe205068_4347,RIe1ff0c8_4279,RIe1f8480_4202,RIe1f0fc8_4119,RIe1d54d0_3804,
        RIe1bbfd0_3516,RIe1aee48_3367,RIe171480_2666,RIdec5810_711,RIdec2b10_679,RIfce6f60_7650,RIdebfe10_647,RIfc95228_6719,RIdebd110_615,RIdeba410_583,
        RIdeb7710_551,RIfe879a8_7887,RIdeb1d10_487,RIfcc16e8_7223,RIdeaf010_455,RIfca4f48_6899,RIdeaadf8_423,RIdea44f8_391,RIde9dbf8_359,RIee1cf48_4788,
        RIee1bfd0_4777,RIfc95660_6722,RIfcee148_7731,RIfe87840_7886,RIfe876d8_7885,RIde8a0f8_263,RIde85f58_243,RIfcb0780_7030,RIfcee9b8_7737,RIfc5f150_6104,
        RIfcdee00_7558,RIfcd8050_7480,RIe16ba80_2602,RIfca5380_6902,RIe1680d8_2561,RIe165810_2532,RIe162b10_2500,RIee377f8_5090,RIe15fe10_2468,RIee36448_5076,
        RIe15d110_2436,RIe157710_2372,RIe154a10_2340,RIfc3f3c8_5745,RIe151d10_2308,RIfcde9c8_7555,RIe14f010_2276,RIfc4a2a0_5866,RIe14c310_2244,RIe149610_2212,
        RIe146910_2180,RIfc62288_6139,RIee33478_5042,RIfc71b70_6316,RIee312b8_5018,RIe1411e0_2118,RIfe87570_7884,RIdf3cf28_2070,RIfe87408_7883,RIfcc99b0_7316,
        RIfccf0e0_7378,RIfcaeb60_7010,RIfcca220_7322,RIdf35bd8_1988,RIdf33748_1962,RIdf31588_1938,RIdf2f530_1915,RIee2be58_4958,RIee2a508_4940,RIee28ff0_4925,
        RIee27da8_4912,RIdf2a508_1858,RIdf28348_1834,RIdf265c0_1813,RIdf24b08_1794,RIfc74708_6347,RIfc42578_5777,RIfc43388_5787,RIfc745a0_6346,RIfcb0078_7025,
        RIdf1fc48_1738,RIfcaff10_7024,RIdf195a0_1665,RIdf173e0_1641,RIdf146e0_1609,RIdf119e0_1577,RIdf0ece0_1545,RIdf0bfe0_1513,RIdf092e0_1481,RIdf065e0_1449,
        RIdf038e0_1417,RIdefdee0_1353,RIdefb1e0_1321,RIdef84e0_1289,RIdef57e0_1257,RIdef2ae0_1225,RIdeefde0_1193,RIdeed0e0_1161,RIdeea3e0_1129,RIee257b0_4885,
        RIfca73d8_6925,RIee23e60_4867,RIfce66f0_7644,RIdee4cb0_1067,RIdee2f28_1046,RIdee0d68_1022,RIdeded10_999,RIfcca388_7323,RIfce6858_7645,RIfcceca8_7375,
        RIfcdc970_7532,RIded9b80_941,RIfeaaac0_8258,RIded5800_893,RIded3208_866,RIded0c10_839,RIdecdf10_807,RIdecb210_775,RIdec8510_743,RIdeb4a10_519,
        RIde972f8_327,RIe16e618_2633,RIe15a410_2404,RIe143c10_2148,RIdf38608_2018,RIdf2cc68_1886,RIdf1d4e8_1710,RIdf00be0_1385,RIdee76e0_1097,RIdedc448_970,
        RIde7d240_200,RIe19daa8_3171,RIe19ada8_3139,RIf1457c0_5250,RIe1980a8_3107,RIf1449b0_5240,RIe1953a8_3075,RIe1926a8_3043,RIe18f9a8_3011,RIe189fa8_2947,
        RIe1872a8_2915,RIf143ba0_5230,RIe1845a8_2883,RIfc912e0_6674,RIe1818a8_2851,RIe17eba8_2819,RIe17bea8_2787,RIfc915b0_6676,RIfcbe5b0_7188,RIfce3b58_7613,
        RIe175da0_2718,RIfceb448_7699,RIfcc7958_7293,RIfc42de8_5783,RIfc96e48_6739,RIfc7a810_6416,RIfc96ce0_6738,RIfcc7ac0_7294,RIe173be0_2694,RIfce39f0_7612,
        RIfc7a540_6414,RIfc91b50_6680,RIfc429b0_5780,RIfea9710_8244,RIe223e00_4698,RIfcd8488_7483,RIe221100_4666,RIfc920f0_6684,RIe21e400_4634,RIe218a00_4570,
        RIe215d00_4538,RIfc79e38_6409,RIe213000_4506,RIfcbee20_7194,RIe210300_4474,RIf168068_5643,RIe20d600_4442,RIe20a900_4410,RIe207c00_4378,RIfc5af38_6057,
        RIfcd73a8_7471,RIe2027a0_4318,RIe200ce8_4299,RIfcb2670_7052,RIfcdf940_7566,RIfc5b208_6059,RIfcbf3c0_7198,RIf1604a8_5555,RIf15e5b8_5533,RIfe872a0_7882,
        RIfe87138_7881,RIfc78920_6394,RIfec1158_8317,RIfc93338_6697,RIfcea368_7687,RIfcb23a0_7050,RIfc5bbe0_6066,RIfcede78_7729,RIe1fa370_4224,RIfcd4c48_7443,
        RIfce1dd0_7592,RIfcbf960_7202,RIe1f58e8_4171,RIfcbfc30_7204,RIfc78380_6390,RIfc93770_6700,RIe1f35c0_4146,RIfcb1f68_7047,RIfce1b00_7590,RIfc93a40_6702,
        RIe1ee2c8_4087,RIe1ebb68_4059,RIe1e8e68_4027,RIe1e6168_3995,RIe1e3468_3963,RIe1e0768_3931,RIe1dda68_3899,RIe1dad68_3867,RIe1d8068_3835,RIe1d2668_3771,
        RIe1cf968_3739,RIe1ccc68_3707,RIe1c9f68_3675,RIe1c7268_3643,RIe1c4568_3611,RIe1c1868_3579,RIe1beb68_3547,RIfcdec98_7557,RIfc94148_6707,RIe1b95a0_3486,
        RIe1b7548_3463,RIfcd12a0_7402,RIfceabd8_7693,RIe1b5388_3439,RIe1b3fd8_3425,RIfc94850_6712,RIfcd7c18_7477,RIe1b27f0_3408,RIe1b0d38_3389,RIfc76a30_6372,
        RIfce2640_7598,RIe1ac6e8_3339,RIe1ab068_3323,RIe1a8ea8_3299,RIe1a61a8_3267,RIe1a34a8_3235,RIe1a07a8_3203,RIe18cca8_2979,RIe1791a8_2755,RIe226b00_4730,
        RIe21b700_4602,RIe204f00_4346,RIe1fef60_4278,RIe1f8318_4201,RIe1f0e60_4118,RIe1d5368_3803,RIe1bbe68_3515,RIe1aece0_3366,RIe171318_2665,RIdec5c48_714,
        RIdec2f48_682,RIfc7c160_6434,RIdec0248_650,RIfcb38b8_7065,RIdebd548_618,RIdeba848_586,RIdeb7b48_554,RIfce7c08_7659,RIdeb2148_490,RIfce7aa0_7658,
        RIdeaf448_458,RIfca38c8_6883,RIdeab7d0_426,RIdea4ed0_394,RIde9e5d0_362,RIfc41e70_5772,RIfc5b0a0_6058,RIfcdbb60_7522,RIfc78650_6392,RIfea92d8_8241,
        RIde8e5e0_284,RIfea0d40_8174,RIfea0bd8_8173,RIfcdf508_7563,RIfcb1b30_7044,RIfc5ccc0_6078,RIfcb16f8_7041,RIfc77b10_6384,RIe16beb8_2605,RIe169e60_2582,
        RIe168510_2564,RIe165c48_2535,RIe162f48_2503,RIfc4f9d0_5928,RIe160248_2471,RIfc4e8f0_5916,RIe15d548_2439,RIe157b48_2375,RIe154e48_2343,RIfc4e1e8_5911,
        RIe152148_2311,RIfc868b8_6553,RIe14f448_2279,RIfc865e8_6551,RIe14c748_2247,RIe149a48_2215,RIe146d48_2183,RIfc9eb70_6828,RIfc9ecd8_6829,RIfcc5630_7268,
        RIfc83bb8_6521,RIe141618_2121,RIfea0ea8_8175,RIdf3d1f8_2072,RIdf3ac00_2045,RIee308e0_5011,RIfcd3cd0_7432,RIfc84e00_6534,RIfc834b0_6516,RIdf36010_1991,
        RIdf33a18_1964,RIdf31858_1940,RIdf2f968_1918,RIee2c128_4960,RIee2a7d8_4942,RIee292c0_4927,RIee28078_4914,RIdf2a940_1861,RIdf28780_1837,RIfea0a70_8172,
        RIfea0908_8171,RIfcd4f18_7445,RIfca0628_6847,RIdf23050_1775,RIfcd3190_7424,RIdf21b38_1760,RIdf20080_1741,RIdf1b328_1686,RIdf199d8_1668,RIdf17818_1644,
        RIdf14b18_1612,RIdf11e18_1580,RIdf0f118_1548,RIdf0c418_1516,RIdf09718_1484,RIdf06a18_1452,RIdf03d18_1420,RIdefe318_1356,RIdefb618_1324,RIdef8918_1292,
        RIdef5c18_1260,RIdef2f18_1228,RIdef0218_1196,RIdeed518_1164,RIdeea818_1132,RIfcdf3a0_7562,RIfca5218_6901,RIfcdc538_7529,RIfcdc6a0_7530,RIdee50e8_1070,
        RIdee3360_1049,RIfea07a0_8170,RIdedefe0_1001,RIfcb0d20_7034,RIfcd4978_7441,RIfca49a8_6895,RIfca1708_6859,RIded9fb8_944,RIded79c0_917,RIded5ad0_895,
        RIfeab498_8265,RIded1048_842,RIdece348_810,RIdecb648_778,RIdec8948_746,RIdeb4e48_522,RIde97cd0_330,RIe16ea50_2636,RIe15a848_2407,RIe144048_2151,
        RIdf38a40_2021,RIdf2d0a0_1889,RIdf1d920_1713,RIdf01018_1388,RIdee7b18_1100,RIdedc880_973,RIde7dc18_203,RIe19dee0_3174,RIe19b1e0_3142,RIfc67580_6198,
        RIe1984e0_3110,RIfccb030_7332,RIe1957e0_3078,RIe192ae0_3046,RIe18fde0_3014,RIe18a3e0_2950,RIe1876e0_2918,RIfc6a550_6232,RIe1849e0_2886,RIfcaa7e0_6962,
        RIe181ce0_2854,RIe17efe0_2822,RIe17c2e0_2790,RIfc65d98_6181,RIfc65690_6176,RIe1772b8_2733,RIfea0638_8169,RIfcca928_7327,RIfc607d0_6120,RIfc65258_6173,
        RIee3d798_5158,RIee3c3e8_5144,RIfca9430_6948,RIee39f58_5118,RIe174018_2697,RIfcecf00_7718,RIfc650f0_6172,RIf16e5a8_5715,RIfc43a90_5792,RIfc65528_6175,
        RIe224238_4701,RIfca9f70_6956,RIe221538_4669,RIfc6b4c8_6243,RIe21e838_4637,RIe218e38_4573,RIe216138_4541,RIfc3fda0_5752,RIe213438_4509,RIfc61310_6128,
        RIe210738_4477,RIfc60c08_6123,RIe20da38_4445,RIe20ad38_4413,RIe208038_4381,RIfc66ba8_6191,RIfccbcd8_7341,RIe202bd8_4321,RIe200fb8_4301,RIfcadbe8_6999,
        RIfccbe40_7342,RIfca7540_6926,RIfc6a3e8_6231,RIfca6898_6917,RIfc73358_6333,RIe1fd070_4256,RIe1fbe28_4243,RIfcc2660_7234,RIfc44468_5799,RIf15a940_5490,
        RIfca7270_6924,RIfc5e070_6092,RIfc5dda0_6090,RIfc7e050_6456,RIe1fa7a8_4227,RIfc5d968_6087,RIfcd9568_7495,RIfc8d668_6631,RIe1f5d20_4174,RIfca4138_6889,
        RIfc8cdf8_6625,RIfcc7c28_7295,RIe1f39f8_4149,RIfc99440_6766,RIfcbc3f0_7164,RIfc5a128_6047,RIe1ee700_4090,RIe1ebfa0_4062,RIe1e92a0_4030,RIe1e65a0_3998,
        RIe1e38a0_3966,RIe1e0ba0_3934,RIe1ddea0_3902,RIe1db1a0_3870,RIe1d84a0_3838,RIe1d2aa0_3774,RIe1cfda0_3742,RIe1cd0a0_3710,RIe1ca3a0_3678,RIe1c76a0_3646,
        RIe1c49a0_3614,RIe1c1ca0_3582,RIe1befa0_3550,RIf14cde0_5334,RIf14bb98_5321,RIe1b99d8_3489,RIe1b7980_3466,RIfc4c460_5890,RIfc9e738_6825,RIe1b5658_3441,
        RIfec54d8_8365,RIf149168_5291,RIf147f20_5278,RIe1b2ac0_3410,RIe1b1170_3392,RIf1473e0_5270,RIf1468a0_5262,RIe1acb20_3342,RIe1ab338_3325,RIe1a92e0_3302,
        RIe1a65e0_3270,RIe1a38e0_3238,RIe1a0be0_3206,RIe18d0e0_2982,RIe1795e0_2758,RIe226f38_4733,RIe21bb38_4605,RIe205338_4349,RIe1ff398_4281,RIe1f8750_4204,
        RIe1f1298_4121,RIe1d57a0_3806,RIe1bc2a0_3518,RIe1af118_3369,RIe171750_2668,RIdec5ae0_713,RIdec2de0_681,RIfc82268_6503,RIdec00e0_649,RIfcb8d18_7125,
        RIdebd3e0_617,RIdeba6e0_585,RIdeb79e0_553,RIfcb9858_7133,RIdeb1fe0_489,RIfc9efa8_6831,RIdeaf2e0_457,RIfce0750_7576,RIdeab488_425,RIdea4b88_393,
        RIde9e288_361,RIee1d0b0_4789,RIee1c138_4778,RIfcd0e68_7399,RIfc76d00_6374,RIfe89028_7903,RIfe88d58_7901,RIfe88ec0_7902,RIfe88bf0_7900,RIfcda7b0_7508,
        RIfc4d810_5904,RIfc52dd8_5965,RIfcde590_7552,RIfc4f868_5927,RIe16bd50_2604,RIfc68930_6212,RIe1683a8_2563,RIe165ae0_2534,RIe162de0_2502,RIfe88a88_7899,
        RIe1600e0_2470,RIfcc9140_7310,RIe15d3e0_2438,RIe1579e0_2374,RIe154ce0_2342,RIfc698a8_6223,RIe151fe0_2310,RIee35098_5062,RIe14f2e0_2278,RIfcc0338_7209,
        RIe14c5e0_2246,RIe1498e0_2214,RIe146be0_2182,RIfc88208_6571,RIfc85670_6540,RIfc81f98_6501,RIfcc4f28_7263,RIe1414b0_2120,RIe13f188_2095,RIdf3d090_2071,
        RIdf3aa98_2044,RIfcd2920_7418,RIfc7d7e0_6450,RIfc49760_5858,RIfce5a48_7635,RIdf35ea8_1990,RIdf338b0_1963,RIfe88920_7898,RIdf2f800_1917,RIee2bfc0_4959,
        RIee2a670_4941,RIee29158_4926,RIee27f10_4913,RIdf2a7d8_1860,RIdf28618_1836,RIdf26890_1815,RIdf24dd8_1796,RIfcad918_6997,RIfc69fb0_6228,RIfc63368_6151,
        RIfc623f0_6140,RIfc60938_6121,RIdf1ff18_1740,RIfcba500_7142,RIdf19870_1667,RIdf176b0_1643,RIdf149b0_1611,RIdf11cb0_1579,RIdf0efb0_1547,RIdf0c2b0_1515,
        RIdf095b0_1483,RIdf068b0_1451,RIdf03bb0_1419,RIdefe1b0_1355,RIdefb4b0_1323,RIdef87b0_1291,RIdef5ab0_1259,RIdef2db0_1227,RIdef00b0_1195,RIdeed3b0_1163,
        RIdeea6b0_1131,RIfcc9848_7315,RIfc69a10_6224,RIfcacc70_6988,RIfccbfa8_7343,RIdee4f80_1069,RIdee31f8_1048,RIdee1038_1024,RIdedee78_1000,RIfc84590_6528,
        RIfc9bba0_6794,RIee21b38_4842,RIfc47168_5831,RIded9e50_943,RIded7858_916,RIfe887b8_7897,RIded34d8_868,RIded0ee0_841,RIdece1e0_809,RIdecb4e0_777,
        RIdec87e0_745,RIdeb4ce0_521,RIde97988_329,RIe16e8e8_2635,RIe15a6e0_2406,RIe143ee0_2150,RIdf388d8_2020,RIdf2cf38_1888,RIdf1d7b8_1712,RIdf00eb0_1387,
        RIdee79b0_1099,RIdedc718_972,RIde7d8d0_202,RIe19dd78_3173,RIe19b078_3141,RIfca1438_6857,RIe198378_3109,RIfca35f8_6881,RIe195678_3077,RIe192978_3045,
        RIe18fc78_3013,RIe18a278_2949,RIe187578_2917,RIfcba230_7140,RIe184878_2885,RIf142d90_5220,RIe181b78_2853,RIe17ee78_2821,RIe17c178_2789,RIfc9be70_6796,
        RIfc9bd08_6795,RIfc4ccd0_5896,RIe176070_2720,RIfc87c68_6567,RIfc87b00_6566,RIfcc4c58_7261,RIfc4fca0_5930,RIfc4f598_5925,RIfc876c8_6563,RIfc4dae0_5906,
        RIe173eb0_2696,RIfcb9420_7130,RIfc4e080_5910,RIfc4e350_5912,RIfc9d388_6811,RIfc40a48_5761,RIe2240d0_4700,RIfc85508_6539,RIe2213d0_4668,RIfc9ba38_6793,
        RIe21e6d0_4636,RIe218cd0_4572,RIe215fd0_4540,RIfc52c70_5964,RIe2132d0_4508,RIfca3760_6882,RIe2105d0_4476,RIfc97988_6747,RIe20d8d0_4444,RIe20abd0_4412,
        RIe207ed0_4380,RIfceb5b0_7700,RIfcddbb8_7545,RIe202a70_4320,RIe200e50_4300,RIfc73d30_6340,RIfcaf100_7014,RIfc71468_6311,RIfcdcad8_7533,RIfcdda50_7544,
        RIfca8620_6938,RIe1fcf08_4255,RIe1fbcc0_4242,RIfc6c008_6251,RIfcdd1e0_7538,RIfca9700_6950,RIfca92c8_6947,RIfcce5a0_7370,RIfc6ba68_6247,RIfc6f410_6288,
        RIe1fa640_4226,RIfcce000_7366,RIfc53918_5973,RIfcce708_7371,RIe1f5bb8_4173,RIf1535f0_5408,RIf151e08_5391,RIfc72db8_6329,RIe1f3890_4148,RIf14fc48_5367,
        RIfc72c50_6328,RIfc73e98_6341,RIe1ee598_4089,RIe1ebe38_4061,RIe1e9138_4029,RIe1e6438_3997,RIe1e3738_3965,RIe1e0a38_3933,RIe1ddd38_3901,RIe1db038_3869,
        RIe1d8338_3837,RIe1d2938_3773,RIe1cfc38_3741,RIe1ccf38_3709,RIe1ca238_3677,RIe1c7538_3645,RIe1c4838_3613,RIe1c1b38_3581,RIe1bee38_3549,RIfcb8a48_7123,
        RIfcb84a8_7119,RIe1b9870_3488,RIe1b7818_3465,RIfc85940_6542,RIfc9e198_6821,RIfeac140_8274,RIe1b42a8_3427,RIfc518c0_5950,RIfc838e8_6519,RIfe884e8_7895,
        RIe1b1008_3391,RIfcc5900_7270,RIfc82ad8_6509,RIe1ac9b8_3341,RIfe88650_7896,RIe1a9178_3301,RIe1a6478_3269,RIe1a3778_3237,RIe1a0a78_3205,RIe18cf78_2981,
        RIe179478_2757,RIe226dd0_4732,RIe21b9d0_4604,RIe2051d0_4348,RIe1ff230_4280,RIe1f85e8_4203,RIe1f1130_4120,RIe1d5638_3805,RIe1bc138_3517,RIe1aefb0_3368,
        RIe1715e8_2667,RIdec5f18_716,RIdec3218_684,RIee20350_4825,RIdec0518_652,RIee1f6a8_4816,RIdebd818_620,RIdebab18_588,RIdeb7e18_556,RIfce4da0_7626,
        RIdeb2418_492,RIfcea908_7691,RIdeaf718_460,RIfce20a0_7594,RIdeabe60_428,RIdea5560_396,RIde9ec60_364,RIfce6420_7642,RIee1c2a0_4779,RIfc75950_6360,
        RIee1ad88_4764,RIde920f0_302,RIfea4148_8211,RIfeaa688_8255,RIfea3fe0_8210,RIde82790_226,RIfc6f848_6291,RIfc5dc38_6089,RIfc76b98_6373,RIfcae2f0_7004,
        RIe16c020_2606,RIe16a130_2584,RIe1687e0_2566,RIe165f18_2537,RIe163218_2505,RIfcadd50_7000,RIe160518_2473,RIfc55268_5991,RIe15d818_2441,RIe157e18_2377,
        RIe155118_2345,RIfc45548_5811,RIe152418_2313,RIfc498c8_5859,RIe14f718_2281,RIfcbda70_7180,RIe14ca18_2249,RIe149d18_2217,RIe147018_2185,RIee34828_5056,
        RIee33748_5044,RIee32668_5032,RIee31588_5020,RIe1418e8_2123,RIe13f458_2097,RIdf3d360_2073,RIdf3aed0_2047,RIfc526d0_5960,RIfc42848_5779,RIfcae9f8_7009,
        RIfcb7260_7106,RIfea42b0_8212,RIdf33ce8_1966,RIdf31b28_1942,RIdf2fc38_1920,RIee2c3f8_4962,RIfc4cfa0_5898,RIfc572c0_6014,RIfc4f430_5924,RIfea3e78_8209,
        RIdf28a50_1839,RIdf26b60_1817,RIdf250a8_1798,RIfc9b600_6790,RIfcb9df8_7137,RIdf23320_1777,RIfc86318_6549,RIfeabfd8_8273,RIdf201e8_1742,RIdf1b5f8_1688,
        RIdf19ca8_1670,RIdf17ae8_1646,RIdf14de8_1614,RIdf120e8_1582,RIdf0f3e8_1550,RIdf0c6e8_1518,RIdf099e8_1486,RIdf06ce8_1454,RIdf03fe8_1422,RIdefe5e8_1358,
        RIdefb8e8_1326,RIdef8be8_1294,RIdef5ee8_1262,RIdef31e8_1230,RIdef04e8_1198,RIdeed7e8_1166,RIdeeaae8_1134,RIfc89018_6581,RIfcc54c8_7267,RIfc89180_6582,
        RIfc4b380_5878,RIdee53b8_1072,RIdee34c8_1050,RIfea3d10_8208,RIdedf148_1002,RIfcae188_7003,RIfc4b0b0_5876,RIfc74870_6348,RIfce4968_7623,RIdeda288_946,
        RIded7c90_919,RIded5da0_897,RIded3640_869,RIded1318_844,RIdece618_812,RIdecb918_780,RIdec8c18_748,RIdeb5118_524,RIde98360_332,RIe16ed20_2638,
        RIe15ab18_2409,RIe144318_2153,RIdf38d10_2023,RIdf2d370_1891,RIdf1dbf0_1715,RIdf012e8_1390,RIdee7de8_1102,RIdedcb50_975,RIde7e2a8_205,RIe19e1b0_3176,
        RIe19b4b0_3144,RIfc9cf50_6808,RIe1987b0_3112,RIfc87290_6560,RIe195ab0_3080,RIe192db0_3048,RIe1900b0_3016,RIe18a6b0_2952,RIe1879b0_2920,RIfc842c0_6526,
        RIe184cb0_2888,RIfc83a50_6520,RIe181fb0_2856,RIe17f2b0_2824,RIe17c5b0_2792,RIfc9d0b8_6809,RIfc9e030_6820,RIe177420_2734,RIe176340_2722,RIfc4f700_5926,
        RIfcc4820_7258,RIfc4fb38_5929,RIfce8040_7662,RIee3c6b8_5146,RIee3b308_5132,RIfc812f0_6492,RIe174180_2698,RIfcd3028_7423,RIfc7f400_6470,RIfc46a60_5826,
        RIfc472d0_5832,RIf16cc58_5697,RIe224508_4703,RIfc7d3a8_6447,RIe221808_4671,RIfc97c58_6749,RIe21eb08_4639,RIe219108_4575,RIe216408_4543,RIfcdbe30_7524,
        RIe213708_4511,RIf169580_5658,RIe210a08_4479,RIfca4570_6892,RIe20dd08_4447,RIe20b008_4415,RIe208308_4383,RIfc7b080_6422,RIfc59cf0_6044,RIfea9b48_8247,
        RIfea4418_8213,RIfc79cd0_6408,RIfcd19a8_7407,RIfcc81c8_7299,RIf162230_5576,RIf160778_5557,RIf15e888_5535,RIfea4580_8214,RIfea46e8_8215,RIfc77f48_6387,
        RIfc41fd8_5773,RIf15aaa8_5491,RIfc7c430_6436,RIf159158_5473,RIf157f10_5460,RIfcae890_7008,RIe1faa78_4229,RIfc4a840_5870,RIfc4ed28_5919,RIfce0e58_7581,
        RIe1f5ff0_4176,RIf153758_5409,RIf151f70_5392,RIfccb468_7335,RIe1f3cc8_4151,RIfc68ed0_6216,RIfc6d250_6264,RIfca9ca0_6954,RIe1ee9d0_4092,RIe1ec270_4064,
        RIe1e9570_4032,RIe1e6870_4000,RIe1e3b70_3968,RIe1e0e70_3936,RIe1de170_3904,RIe1db470_3872,RIe1d8770_3840,RIe1d2d70_3776,RIe1d0070_3744,RIe1cd370_3712,
        RIe1ca670_3680,RIe1c7970_3648,RIe1c4c70_3616,RIe1c1f70_3584,RIe1bf270_3552,RIfc784e8_6391,RIfcbef88_7195,RIe1b9ca8_3491,RIe1b7ae8_3467,RIfcc20c0_7230,
        RIfca6190_6912,RIe1b5928_3443,RIe1b4410_3428,RIfcb81d8_7117,RIfcc5090_7264,RIe1b2d90_3412,RIe1b1440_3394,RIfcd5350_7448,RIfcb9588_7131,RIe1acc88_3343,
        RIe1ab4a0_3326,RIe1a95b0_3304,RIe1a68b0_3272,RIe1a3bb0_3240,RIe1a0eb0_3208,RIe18d3b0_2984,RIe1798b0_2760,RIe227208_4735,RIe21be08_4607,RIe205608_4351,
        RIe1ff668_4283,RIe1f8a20_4206,RIe1f1568_4123,RIe1d5a70_3808,RIe1bc570_3520,RIe1af3e8_3371,RIe171a20_2670,RIdec5db0_715,RIdec30b0_683,RIee201e8_4824,
        RIdec03b0_651,RIfcaf538_7017,RIdebd6b0_619,RIdeba9b0_587,RIdeb7cb0_555,RIfc40fe8_5765,RIdeb22b0_491,RIfcd08c8_7395,RIdeaf5b0_459,RIee1dd58_4798,
        RIdeabb18_427,RIdea5218_395,RIde9e918_363,RIee1d218_4790,RIfcedd10_7728,RIfce62b8_7641,RIfcc92a8_7311,RIde91da8_301,RIde8e928_285,RIde8a788_265,
        RIde865e8_245,RIde82448_225,RIfea1448_8179,RIfc750e0_6354,RIfcc19b8_7225,RIfced8d8_7725,RIfec5eb0_8372,RIe169fc8_2583,RIe168678_2565,RIe165db0_2536,
        RIe1630b0_2504,RIfccfc20_7386,RIe1603b0_2472,RIee365b0_5077,RIe15d6b0_2440,RIe157cb0_2376,RIe154fb0_2344,RIfea1718_8181,RIe1522b0_2312,RIee35200_5063,
        RIe14f5b0_2280,RIfcb0348_7027,RIe14c8b0_2248,RIe149bb0_2216,RIe146eb0_2184,RIfc73790_6336,RIfcdf238_7561,RIee32500_5031,RIfc94f58_6717,RIe141780_2122,
        RIe13f2f0_2096,RIfec5be0_8370,RIdf3ad68_2046,RIfea15b0_8180,RIfc5fb28_6111,RIfcae728_7007,RIfc74438_6345,RIdf36178_1992,RIdf33b80_1965,RIdf319c0_1941,
        RIdf2fad0_1919,RIee2c290_4961,RIee2a940_4943,RIfc70658_6301,RIfc704f0_6300,RIdf2aaa8_1862,RIdf288e8_1838,RIdf269f8_1816,RIdf24f40_1797,RIfc64b50_6168,
        RIfccaa90_7328,RIdf231b8_1776,RIfcad4e0_6994,RIdf21ca0_1761,RIfeaad90_8260,RIdf1b490_1687,RIdf19b40_1669,RIdf17980_1645,RIdf14c80_1613,RIdf11f80_1581,
        RIdf0f280_1549,RIdf0c580_1517,RIdf09880_1485,RIdf06b80_1453,RIdf03e80_1421,RIdefe480_1357,RIdefb780_1325,RIdef8a80_1293,RIdef5d80_1261,RIdef3080_1229,
        RIdef0380_1197,RIdeed680_1165,RIdeea980_1133,RIfc595e8_6039,RIfcac568_6983,RIfcccf20_7354,RIfccd358_7357,RIdee5250_1071,RIfea7f28_8227,RIdee11a0_1025,
        RIfea12e0_8178,RIfc679b8_6201,RIee22510_4849,RIfc6dd90_6272,RIfc6cb48_6259,RIdeda120_945,RIded7b28_918,RIded5c38_896,RIfec5d48_8371,RIded11b0_843,
        RIdece4b0_811,RIdecb7b0_779,RIdec8ab0_747,RIdeb4fb0_523,RIde98018_331,RIe16ebb8_2637,RIe15a9b0_2408,RIe1441b0_2152,RIdf38ba8_2022,RIdf2d208_1890,
        RIdf1da88_1714,RIdf01180_1389,RIdee7c80_1101,RIdedc9e8_974,RIde7df60_204,RIe19e048_3175,RIe19b348_3143,RIfcc3ce0_7250,RIe198648_3111,RIfc7efc8_6467,
        RIe195948_3079,RIe192c48_3047,RIe18ff48_3015,RIe18a548_2951,RIe187848_2919,RIfc46790_5824,RIe184b48_2887,RIfc98d38_6761,RIe181e48_2855,RIe17f148_2823,
        RIe17c448_2791,RIfcb5d48_7091,RIfc995a8_6767,RIfc9a3b8_6777,RIe1761d8_2721,RIfc54188_5979,RIfcd2bf0_7420,RIfc8b778_6609,RIfc7dee8_6455,RIee3c550_5145,
        RIfc8c420_6618,RIee3a0c0_5119,RIfeaba38_8269,RIfc46628_5823,RIfcbc288_7163,RIf16e710_5716,RIfc8fdc8_6659,RIfc48c20_5850,RIe2243a0_4702,RIfca0358_6845,
        RIe2216a0_4670,RIfc9a688_6779,RIe21e9a0_4638,RIe218fa0_4574,RIe2162a0_4542,RIfc456b0_5812,RIe2135a0_4510,RIf169418_5657,RIe2108a0_4478,RIfc8bfe8_6615,
        RIe20dba0_4446,RIe20aea0_4414,RIe2081a0_4382,RIfc8c9c0_6622,RIfc7f568_6471,RIe202d40_4322,RIe201120_4302,RIfce2910_7600,RIfc487e8_5847,RIfc46d30_5828,
        RIfc992d8_6765,RIfca2680_6870,RIfc44a08_5803,RIe1fd1d8_4257,RIe1fbf90_4244,RIfc580d0_6024,RIfcbdbd8_7181,RIfc8dd70_6636,RIfce01b0_7572,RIfc7bbc0_6430,
        RIfc90368_6663,RIfc7b8f0_6428,RIe1fa910_4228,RIfcd8b90_7488,RIfc43ec8_5795,RIfc7b788_6427,RIe1f5e88_4175,RIfc7b350_6424,RIfc90d40_6670,RIfca3490_6880,
        RIe1f3b60_4150,RIfc91010_6672,RIfcdb728_7519,RIfcd8758_7485,RIe1ee868_4091,RIe1ec108_4063,RIe1e9408_4031,RIe1e6708_3999,RIe1e3a08_3967,RIe1e0d08_3935,
        RIe1de008_3903,RIe1db308_3871,RIe1d8608_3839,RIe1d2c08_3775,RIe1cff08_3743,RIe1cd208_3711,RIe1ca508_3679,RIe1c7808_3647,RIe1c4b08_3615,RIe1c1e08_3583,
        RIe1bf108_3551,RIf14cf48_5335,RIfc78d58_6397,RIe1b9b40_3490,RIfec5910_8368,RIfc78a88_6395,RIfcd51e8_7447,RIe1b57c0_3442,RIfea1010_8176,RIf1492d0_5292,
        RIfec5a78_8369,RIe1b2c28_3411,RIe1b12d8_3393,RIfec5640_8366,RIf146a08_5263,RIfec57a8_8367,RIfea1178_8177,RIe1a9448_3303,RIe1a6748_3271,RIe1a3a48_3239,
        RIe1a0d48_3207,RIe18d248_2983,RIe179748_2759,RIe2270a0_4734,RIe21bca0_4606,RIe2054a0_4350,RIe1ff500_4282,RIe1f88b8_4205,RIe1f1400_4122,RIe1d5908_3807,
        RIe1bc408_3519,RIe1af280_3370,RIe1718b8_2669,RIdec6350_719,RIdec3650_687,RIfcaf3d0_7016,RIdec0950_655,RIfc6a280_6230,RIdebdc50_623,RIdebaf50_591,
        RIdeb8250_559,RIfc42f50_5784,RIdeb2850_495,RIfc981f8_6753,RIdeafb50_463,RIfc8c6f0_6620,RIdeac838_431,RIdea5f38_399,RIde9f638_367,RIee1d4e8_4792,
        RIfcda648_7507,RIfcc6440_7278,RIfcd5620_7450,RIde92ac8_305,RIfea34a0_8202,RIfea31d0_8200,RIfea3338_8201,RIfcb6b58_7101,RIfcb6888_7099,RIfc9dd60_6818,
        RIee19708_4748,RIfc50c18_5941,RIe16c458_2609,RIfc80a80_6486,RIfec62e8_8375,RIe166350_2540,RIe163650_2508,RIee37d98_5094,RIe160950_2476,RIfcaa678_6961,
        RIe15dc50_2444,RIe158250_2380,RIe155550_2348,RIfea3ba8_8207,RIe152850_2316,RIee35638_5066,RIe14fb50_2284,RIfc62f30_6148,RIe14ce50_2252,RIe14a150_2220,
        RIe147450_2188,RIfc97f28_6751,RIfc89888_6587,RIfc8f558_6653,RIfc52838_5961,RIe141bb8_2125,RIe13f890_2100,RIdf3d798_2076,RIdf3b308_2050,RIee30a48_5012,
        RIfc568e8_6007,RIee2e9f0_4989,RIee2dbe0_4979,RIdf365b0_1995,RIfea38d8_8205,RIfea3a40_8206,RIdf2ff08_1922,RIee2c6c8_4964,RIee2ac10_4945,RIee29590_4929,
        RIee28348_4916,RIdf2ad78_1864,RIdf28e88_1842,RIfea3608_8203,RIfea3770_8204,RIfcc0d10_7216,RIfc75c20_6362,RIfca50b0_6900,RIfc74e10_6352,RIfcc9410_7312,
        RIdf20620_1745,RIfc73628_6335,RIdf1a0e0_1673,RIdf17f20_1649,RIdf15220_1617,RIdf12520_1585,RIdf0f820_1553,RIdf0cb20_1521,RIdf09e20_1489,RIdf07120_1457,
        RIdf04420_1425,RIdefea20_1361,RIdefbd20_1329,RIdef9020_1297,RIdef6320_1265,RIdef3620_1233,RIdef0920_1201,RIdeedc20_1169,RIdeeaf20_1137,RIfcab8c0_6974,
        RIfc7c598_6437,RIfc5beb0_6068,RIfc58ee0_6034,RIdee5688_1074,RIdee3798_1052,RIdee15d8_1028,RIdedf580_1005,RIfcb3048_7059,RIfc72ae8_6327,RIfca3d00_6886,
        RIfcb6450_7096,RIdeda558_948,RIded7f60_921,RIfea3068_8199,RIded3a78_872,RIded1750_847,RIdecea50_815,RIdecbd50_783,RIdec9050_751,RIdeb5550_527,
        RIde98d38_335,RIe16f158_2641,RIe15af50_2412,RIe144750_2156,RIdf39148_2026,RIdf2d7a8_1894,RIdf1e028_1718,RIdf01720_1393,RIdee8220_1105,RIdedcf88_978,
        RIde7ec80_208,RIe19e5e8_3179,RIe19b8e8_3147,RIfca84b8_6937,RIe198be8_3115,RIfc846f8_6529,RIe195ee8_3083,RIe1931e8_3051,RIe1904e8_3019,RIe18aae8_2955,
        RIe187de8_2923,RIfce2be0_7602,RIe1850e8_2891,RIfc8e310_6640,RIe1823e8_2859,RIe17f6e8_2827,RIe17c9e8_2795,RIfcd1570_7404,RIfccc278_7345,RIf1404c8_5191,
        RIfea2d98_8197,RIfcc1b20_7226,RIfc60398_6117,RIee3e5a8_5168,RIee3da68_5160,RIfc642e0_6162,RIfca7f18_6933,RIee3a228_5120,RIfec6180_8374,RIfca9598_6949,
        RIfc5c720_6074,RIfc6bea0_6250,RIfccaec8_7331,RIfc44cd8_5805,RIe224940_4706,RIfcb6180_7094,RIe221c40_4674,RIfc55ad8_5997,RIe21ef40_4642,RIe219540_4578,
        RIe216840_4546,RIfc4dc48_5907,RIe213b40_4514,RIfcdcf10_7536,RIe210e40_4482,RIfcab1b8_6969,RIe20e140_4450,RIe20b440_4418,RIe208740_4386,RIfce3720_7610,
        RIfc64178_6161,RIe203178_4325,RIe201558_4305,RIfcd2ec0_7422,RIf164828_5603,RIfc7f838_6473,RIf162398_5577,RIfcc9c80_7318,RIfca8bc0_6942,RIfea2ac8_8195,
        RIfea2c30_8196,RIfc59318_6037,RIfc4f160_5922,RIf15ac10_5492,RIfcebf88_7707,RIfcbb040_7150,RIfca1870_6860,RIfc93d10_6704,RIe1faeb0_4232,RIf1565c0_5442,
        RIf155a80_5434,RIfc45c50_5816,RIe1f6428_4179,RIfccdbc8_7363,RIfcccae8_7351,RIfca6cd0_6920,RIfec6018_8373,RIfc64010_6160,RIfc434f0_5788,RIfc4c028_5887,
        RIe1eee08_4095,RIe1ec6a8_4067,RIe1e99a8_4035,RIe1e6ca8_4003,RIe1e3fa8_3971,RIe1e12a8_3939,RIe1de5a8_3907,RIe1db8a8_3875,RIe1d8ba8_3843,RIe1d31a8_3779,
        RIe1d04a8_3747,RIe1cd7a8_3715,RIe1caaa8_3683,RIe1c7da8_3651,RIe1c50a8_3619,RIe1c23a8_3587,RIe1bf6a8_3555,RIfc63908_6155,RIfc6bd38_6249,RIe1ba0e0_3494,
        RIe1b7f20_3470,RIfc66fe0_6194,RIfc92ac8_6691,RIe1b5d60_3446,RIfea2f00_8198,RIfc9bfd8_6797,RIfc50d80_5942,RIe1b31c8_3415,RIe1b1878_3397,RIfc4df18_5909,
        RIfc9d658_6813,RIe1ad0c0_3346,RIe1ab8d8_3329,RIe1a99e8_3307,RIe1a6ce8_3275,RIe1a3fe8_3243,RIe1a12e8_3211,RIe18d7e8_2987,RIe179ce8_2763,RIe227640_4738,
        RIe21c240_4610,RIe205a40_4354,RIe1ffaa0_4286,RIe1f8e58_4209,RIe1f19a0_4126,RIe1d5ea8_3811,RIe1bc9a8_3523,RIe1af820_3374,RIe171e58_2673,RIdec61e8_718,
        RIdec34e8_686,RIee20620_4827,RIdec07e8_654,RIfc4b7b8_5881,RIdebdae8_622,RIdebade8_590,RIdeb80e8_558,RIfc41150_5766,RIdeb26e8_494,RIfc87830_6564,
        RIdeaf9e8_462,RIee1dec0_4799,RIdeac4f0_430,RIdea5bf0_398,RIde9f2f0_366,RIee1d380_4791,RIfc77c78_6385,RIfc84f68_6535,RIfc6ff50_6296,RIde92780_304,
        RIde8efb8_287,RIde8ae18_267,RIde86c78_247,RIee1a680_4759,RIee19f78_4754,RIfcd7240_7470,RIfcbeb50_7192,RIfc76328_6367,RIe16c2f0_2608,RIee388d8_5102,
        RIfea20f0_8188,RIe1661e8_2539,RIe1634e8_2507,RIee37c30_5093,RIe1607e8_2475,RIfce7500_7654,RIe15dae8_2443,RIe1580e8_2379,RIe1553e8_2347,RIfc3f698_5747,
        RIe1526e8_2315,RIee354d0_5065,RIe14f9e8_2283,RIfc83e88_6523,RIe14cce8_2251,RIe149fe8_2219,RIe1472e8_2187,RIfcea4d0_7688,RIfcb7ad0_7112,RIfc695d8_6221,
        RIfc51a28_5951,RIe141a50_2124,RIe13f728_2099,RIdf3d630_2075,RIdf3b1a0_2049,RIfca9e08_6955,RIee2fda0_5003,RIfc88a78_6577,RIee2da78_4978,RIdf36448_1994,
        RIdf33fb8_1968,RIdf31df8_1944,RIfea2258_8189,RIee2c560_4963,RIee2aaa8_4944,RIee29428_4928,RIee281e0_4915,RIdf2ac10_1863,RIdf28d20_1841,RIfea27f8_8193,
        RIfea2960_8194,RIfcdabe8_7511,RIfca08f8_6849,RIfc8b1d8_6605,RIfc49058_5853,RIfca0a60_6850,RIdf204b8_1744,RIfc99cb0_6772,RIdf19f78_1672,RIdf17db8_1648,
        RIdf150b8_1616,RIdf123b8_1584,RIdf0f6b8_1552,RIdf0c9b8_1520,RIdf09cb8_1488,RIdf06fb8_1456,RIdf042b8_1424,RIdefe8b8_1360,RIdefbbb8_1328,RIdef8eb8_1296,
        RIdef61b8_1264,RIdef34b8_1232,RIdef07b8_1200,RIdeedab8_1168,RIdeeadb8_1136,RIfcd1f48_7411,RIfc57f68_6023,RIfcbe2e0_7186,RIfcd8fc8_7491,RIdee5520_1073,
        RIfea2690_8192,RIdee1470_1027,RIdedf418_1004,RIfc57b30_6020,RIfcb35e8_7063,RIfcbd7a0_7178,RIfc91178_6673,RIfea2528_8191,RIded7df8_920,RIfea23c0_8190,
        RIded3910_871,RIded15e8_846,RIdece8e8_814,RIdecbbe8_782,RIdec8ee8_750,RIdeb53e8_526,RIde989f0_334,RIe16eff0_2640,RIe15ade8_2411,RIe1445e8_2155,
        RIdf38fe0_2025,RIdf2d640_1893,RIdf1dec0_1717,RIdf015b8_1392,RIdee80b8_1104,RIdedce20_977,RIde7e938_207,RIe19e480_3178,RIe19b780_3146,RIfccc980_7350,
        RIe198a80_3114,RIfcc1148_7219,RIe195d80_3082,RIe193080_3050,RIe190380_3018,RIe18a980_2954,RIe187c80_2922,RIfcb2ee0_7058,RIe184f80_2890,RIfc615e0_6130,
        RIe182280_2858,RIe17f580_2826,RIe17c880_2794,RIfc69038_6217,RIfc4c898_5893,RIfc6f2a8_6287,RIe1764a8_2723,RIfcad0a8_6991,RIfc6adc0_6238,RIfc70388_6299,
        RIfea1b50_8184,RIfea1f88_8187,RIfc56e88_6011,RIfea1cb8_8185,RIe174450_2700,RIfc60d70_6124,RIfc6a820_6234,RIfea1e20_8186,RIf16d798_5705,RIfc40bb0_5762,
        RIe2247d8_4705,RIfc77138_6377,RIe221ad8_4673,RIfcd7d80_7478,RIe21edd8_4641,RIe2193d8_4577,RIe2166d8_4545,RIfc40070_5754,RIe2139d8_4513,RIf169850_5660,
        RIe210cd8_4481,RIfcc1580_7222,RIe20dfd8_4449,RIe20b2d8_4417,RIe2085d8_4385,RIfcd0058_7389,RIfc749d8_6349,RIe203010_4324,RIe2013f0_4304,RIfc60230_6116,
        RIfc60668_6119,RIfcaf970_7020,RIfc45818_5813,RIf160a48_5559,RIf15eb58_5537,RIfea1880_8182,RIfea19e8_8183,RIfc72110_6320,RIfc49b98_5861,RIfcca0b8_7321,
        RIfc71738_6313,RIfc4ca00_5894,RIfc71030_6308,RIfcde428_7551,RIe1fad48_4231,RIfc70bf8_6305,RIfc63a70_6156,RIfca7db0_6932,RIe1f62c0_4178,RIfcada80_6998,
        RIfc6fde8_6295,RIfc6f578_6289,RIe1f3f98_4153,RIfcde158_7549,RIfcad378_6993,RIfc65f00_6182,RIe1eeca0_4094,RIe1ec540_4066,RIe1e9840_4034,RIe1e6b40_4002,
        RIe1e3e40_3970,RIe1e1140_3938,RIe1de440_3906,RIe1db740_3874,RIe1d8a40_3842,RIe1d3040_3778,RIe1d0340_3746,RIe1cd640_3714,RIe1ca940_3682,RIe1c7c40_3650,
        RIe1c4f40_3618,RIe1c2240_3586,RIe1bf540_3554,RIfc69308_6219,RIfccba08_7339,RIe1b9f78_3493,RIe1b7db8_3469,RIfccd628_7359,RIfc69740_6222,RIe1b5bf8_3445,
        RIe1b4578_3429,RIfccf950_7384,RIf148088_5279,RIe1b3060_3414,RIe1b1710_3396,RIfc9f818_6837,RIfcb9c90_7136,RIe1acf58_3345,RIe1ab770_3328,RIe1a9880_3306,
        RIe1a6b80_3274,RIe1a3e80_3242,RIe1a1180_3210,RIe18d680_2986,RIe179b80_2762,RIe2274d8_4737,RIe21c0d8_4609,RIe2058d8_4353,RIe1ff938_4285,RIe1f8cf0_4208,
        RIe1f1838_4125,RIe1d5d40_3810,RIe1bc840_3522,RIe1af6b8_3373,RIe171cf0_2672,R_58_102f1b78,R_59_be1fc68,R_5a_10279198,R_5b_102299e8,R_5c_101d0448,
        R_5d_f7f82f0,R_5e_be21600,R_5f_f7fa5b8,R_60_1027d530,R_61_10205ae8,R_62_10283510,R_63_f82b578,R_64_ace4e68,R_65_f8204e0,R_66_1027a0b0,
        R_67_1022dc30,R_68_102478a8,R_69_10286f78,R_6a_f7edd80,R_6b_101c3628,R_6c_f7fbe00,R_6d_f7ce9f8,R_6e_f7c8830,R_6f_101ffc68,R_70_f7d4000,
        R_71_acee958,R_72_94046c0,R_73_101ee420,R_74_102eb268,R_75_b320c50,R_76_ad80a90,R_77_1027fd48,R_78_f7ce4b8,R_79_ad77048,R_7a_102a6ae0,
        R_7b_f7e4c78,R_7c_e2a6ce0,R_7d_101e86e0,R_7e_e2a9cc8,R_7f_10292be0,R_80_b33cde8,R_81_101e2908,R_82_102e9780,R_83_f8157a0,R_84_f819358,
        R_85_ace8b70,R_86_be142b0,R_87_f81b770,R_88_b330278,R_89_f7fe9f8,R_8a_101cf488,R_8b_f8225c0,R_8c_101d4738,R_8d_101c4000,R_8e_101fe960,
        R_8f_102a0330,R_90_f7f4bd0,R_91_1023e5a8,R_92_10248da8,R_93_be2c938,R_94_f7f5458,R_95_f7c6808,R_96_be316a8,R_97_e2a0328,R_98_be2d850,
        R_99_10217db0,R_9a_f7ec340,R_9b_be23ec0,R_9c_101d4540,R_9d_f800828,R_9e_102970c8,R_9f_10221de0,R_a0_ad8d568,R_a1_be4eb58,R_a2_f7c5500,
        R_a3_ad88f30,R_a4_f82f088,R_a5_f7dcbc8,R_a6_10292940,R_a7_be138d8,R_a8_acee418,R_a9_ad84450,R_aa_be10838,R_ab_be31fd8,R_ac_acdaef0,
        R_ad_acea908,R_ae_101f8830,R_af_f7dec98,R_b0_101e2c50,R_b1_f801b30,R_b2_be16e00,R_b3_102e3cf0,R_b4_10291788);
input RIdec64b8_720,RIbc62af0_23,RIbc62a78_22,RIbc62a00_21,RIbc62988_20,RIbc62910_19,RIbc62898_18,RIbc62820_17,RIbc627a8_16,
        RIbc62730_15,RIbc626b8_14,RIbc62640_13,RIdec37b8_688,RIfc8daa0_6634,RIdec0ab8_656,RIfc56348_6003,RIdebddb8_624,RIdebb0b8_592,RIdeb83b8_560,
        RIfc98798_6757,RIdeb29b8_496,RIfcbd098_7173,RIdeafcb8_464,RIfc8dc08_6635,RIdeacb80_432,RIdea6280_400,RIde9f980_368,RIfcd6868_7463,RIfc8ded8_6637,
        RIfc7dd80_6454,RIfc56618_6005,RIde92e10_306,RIde8f300_288,RIde8b160_268,RIde86fc0_248,RIde82ad8_227,RIfc8e040_6638,RIfcd96d0_7496,RIfca1e10_6864,
        RIfcbd200_7174,RIe16c5c0_2610,RIe16a298_2585,RIe168ab0_2568,RIe1664b8_2541,RIe1637b8_2509,RIee37f00_5095,RIe160ab8_2477,RIfc8ea18_6645,RIe15ddb8_2445,
        RIe1583b8_2381,RIe1556b8_2349,RIfe9f828_8159,RIe1529b8_2317,RIfe9f990_8160,RIe14fcb8_2285,RIfcbd368_7175,RIe14cfb8_2253,RIe14a2b8_2221,RIe1475b8_2189,
        RIfc8ee50_6648,RIfc45278_5809,RIfc98360_6754,RIfca2248_6867,RIe141d20_2126,RIe13f9f8_2101,RIdf3d900_2077,RIdf3b470_2051,RIfcd6ca0_7466,RIee2ff08_5004,
        RIfc8ece8_6647,RIee2dd48_4980,RIdf36718_1996,RIdf34120_1969,RIdf31f60_1945,RIfe9f6c0_8158,RIfcb4560_7074,RIfc45db8_5817,RIfc8e1a8_6639,RIfc7d678_6449,
        RIdf2aee0_1865,RIdf28ff0_1843,RIdf26e30_1819,RIdf25378_1800,RIfcb43f8_7073,RIfc8e748_6643,RIdf23488_1778,RIfcc2c00_7238,RIdf21e08_1762,RIdf20788_1746,
        RIdf1b760_1689,RIdf1a248_1674,RIdf18088_1650,RIdf15388_1618,RIdf12688_1586,RIdf0f988_1554,RIdf0cc88_1522,RIdf09f88_1490,RIdf07288_1458,RIdf04588_1426,
        RIdefeb88_1362,RIdefbe88_1330,RIdef9188_1298,RIdef6488_1266,RIdef3788_1234,RIdef0a88_1202,RIdeedd88_1170,RIdeeb088_1138,RIfc8efb8_6649,RIfc44e40_5806,
        RIfc57860_6018,RIfca23b0_6868,RIfe9faf8_8161,RIdee3900_1053,RIdee1740_1029,RIdedf6e8_1006,RIfcbd4d0_7176,RIee22678_4850,RIfc98090_6752,RIee21598_4838,
        RIfe9fc60_8162,RIded80c8_922,RIfe9fdc8_8163,RIded3be0_873,RIded18b8_848,RIdecebb8_816,RIdecbeb8_784,RIdec91b8_752,RIdeb56b8_528,RIde99080_336,
        RIe16f2c0_2642,RIe15b0b8_2413,RIe1448b8_2157,RIdf392b0_2027,RIdf2d910_1895,RIdf1e190_1719,RIdf01888_1394,RIdee8388_1106,RIdedd0f0_979,RIde7efc8_209,
        RIe19e750_3180,RIbc625c8_12,RIbc62550_11,RIbc624d8_10,RIbc62460_9,RIbc623e8_8,RIbc62370_7,RIbc622f8_6,RIbc62280_5,RIbc62208_4,
        RIbc62190_3,RIbc62118_2,RIe19ba50_3148,RIfc479d8_5837,RIe198d50_3116,RIfe9f558_8157,RIe196050_3084,RIe193350_3052,RIe190650_3020,RIe18ac50_2956,
        RIe187f50_2924,RIfc47870_5836,RIe185250_2892,RIf142ef8_5221,RIe182550_2860,RIe17f850_2828,RIe17cb50_2796,RIfcb5208_7083,RIfcbc6c0_7166,RIe177588_2735,
        RIe176610_2724,RIf13fdc0_5186,RIfe9f3f0_8156,RIfce40f8_7617,RIfc47708_5835,RIfc47438_5833,RIfca15a0_6858,RIfc99170_6764,RIe1745b8_2701,RIfc8cc90_6624,
        RIfc556a0_5994,RIfc7ee60_6466,RIfce8e50_7672,RIfe9f288_8155,RIe224aa8_4707,RIfc55808_5995,RIe221da8_4675,RIfcb50a0_7082,RIe21f0a8_4643,RIe2196a8_4579,
        RIe2169a8_4547,RIfcbc828_7167,RIe213ca8_4515,RIfc47000_5830,RIe210fa8_4483,RIfcbc990_7168,RIe20e2a8_4451,RIe20b5a8_4419,RIe2088a8_4387,RIfc46bc8_5827,
        RIfcd6598_7461,RIe2032e0_4326,RIe2016c0_4306,RIfc98ea0_6762,RIfc7eb90_6464,RIfce0318_7573,RIfcbcaf8_7169,RIfc8cf60_6626,RIfcb4dd0_7080,RIe1fd340_4258,
        RIe1fc260_4246,RIf15cf38_5517,RIfe9f120_8154,RIfc7ea28_6463,RIfc8d0c8_6627,RIfcbcc60_7170,RIfc98bd0_6760,RIfce2d48_7603,RIe1fb018_4233,RIfc55f10_6000,
        RIfc7e8c0_6462,RIfc8d230_6628,RIe1f6590_4180,RIfce58e0_7634,RIfc468f8_5825,RIfcc2ed0_7240,RIe1f4100_4154,RIfceedf0_7740,RIfc8d398_6629,RIfc8d500_6630,
        RIe1eef70_4096,RIe1ec810_4068,RIe1e9b10_4036,RIe1e6e10_4004,RIe1e4110_3972,RIe1e1410_3940,RIe1de710_3908,RIe1dba10_3876,RIe1d8d10_3844,RIe1d3310_3780,
        RIe1d0610_3748,RIe1cd910_3716,RIe1cac10_3684,RIe1c7f10_3652,RIe1c5210_3620,RIe1c2510_3588,RIe1bf810_3556,RIf14d0b0_5336,RIfe9efb8_8153,RIe1ba248_3495,
        RIe1b8088_3471,RIfec4dd0_8360,RIfec50a0_8362,RIe1b5ec8_3447,RIe1b46e0_3430,RIfcb4998_7077,RIfcb4c68_7079,RIfec5370_8364,RIfe9ee50_8152,RIfcbcdc8_7171,
        RIfc46358_5821,RIfec5208_8363,RIfec4f38_8361,RIe1a9b50_3308,RIe1a6e50_3276,RIe1a4150_3244,RIe1a1450_3212,RIe18d950_2988,RIe179e50_2764,RIe2277a8_4739,
        RIe21c3a8_4611,RIe205ba8_4355,RIe1ffc08_4287,RIe1f8fc0_4210,RIe1f1b08_4127,RIe1d6010_3812,RIe1bcb10_3524,RIe1af988_3375,RIe171fc0_2674,RIdec6080_717,
        RIdec3380_685,RIee204b8_4826,RIdec0680_653,RIfcd70d8_7469,RIdebd980_621,RIdebac80_589,RIdeb7f80_557,RIfcbe448_7187,RIdeb2580_493,RIfcb3480_7062,
        RIdeaf880_461,RIfc43928_5791,RIdeac1a8_429,RIdea58a8_397,RIde9efa8_365,RIfcd88c0_7486,RIee1c408_4780,RIfcc77f0_7292,RIfea04d0_8168,RIde92438_303,
        RIde8ec70_286,RIde8aad0_266,RIde86930_246,RIfca31c0_6878,RIfc59a20_6042,RIfcd1de0_7410,RIfc91448_6675,RIfc97280_6742,RIe16c188_2607,RIfc97118_6741,
        RIe168948_2567,RIe166080_2538,RIe163380_2506,RIee37ac8_5092,RIe160680_2474,RIfcd1c78_7409,RIe15d980_2442,RIe157f80_2378,RIe155280_2346,RIfc3f530_5746,
        RIe152580_2314,RIee35368_5064,RIe14f880_2282,RIfc7a3d8_6413,RIe14cb80_2250,RIe149e80_2218,RIe147180_2186,RIfc42b18_5781,RIfc7a270_6412,RIfc5a560_6050,
        RIfc96b78_6737,RIfea6fb0_8216,RIe13f5c0_2098,RIdf3d4c8_2074,RIdf3b038_2048,RIfce5bb0_7636,RIee2fc38_5002,RIfc91cb8_6681,RIee2d910_4977,RIdf362e0_1993,
        RIdf33e50_1967,RIdf31c90_1943,RIdf2fda0_1921,RIfc43658_5789,RIfc59e58_6045,RIfc96fb0_6740,RIfc7ac48_6419,RIfea0368_8167,RIdf28bb8_1840,RIdf26cc8_1818,
        RIdf25210_1799,RIfc91718_6677,RIfcb3318_7061,RIfc919e8_6679,RIfc91880_6678,RIfc430b8_5785,RIdf20350_1743,RIfc7a978_6417,RIdf19e10_1671,RIdf17c50_1647,
        RIdf14f50_1615,RIdf12250_1583,RIdf0f550_1551,RIdf0c850_1519,RIdf09b50_1487,RIdf06e50_1455,RIdf04150_1423,RIdefe750_1359,RIdefba50_1327,RIdef8d50_1295,
        RIdef6050_1263,RIdef3350_1231,RIdef0650_1199,RIdeed950_1167,RIdeeac50_1135,RIfcd1b10_7408,RIfc968a8_6735,RIfc91f88_6683,RIfcdfc10_7568,RIfea99e0_8246,
        RIdee3630_1051,RIdee1308_1026,RIdedf2b0_1003,RIfcc7d90_7296,RIfcd85f0_7484,RIfce3888_7611,RIfc5a830_6052,RIdeda3f0_947,RIfea9878_8245,RIded5f08_898,
        RIded37a8_870,RIded1480_845,RIdece780_813,RIdecba80_781,RIdec8d80_749,RIdeb5280_525,RIde986a8_333,RIe16ee88_2639,RIe15ac80_2410,RIe144480_2154,
        RIdf38e78_2024,RIdf2d4d8_1892,RIdf1dd58_1716,RIdf01450_1391,RIdee7f50_1103,RIdedccb8_976,RIde7e5f0_206,RIe19e318_3177,RIe19b618_3145,RIfc8f3f0_6652,
        RIe198918_3113,RIf144b18_5241,RIe195c18_3081,RIe192f18_3049,RIe190218_3017,RIe18a818_2953,RIe187b18_2921,RIf143d08_5231,RIe184e18_2889,RIfcb3cf0_7068,
        RIe182118_2857,RIe17f418_2825,RIe17c718_2793,RIfc448a0_5802,RIf141170_5200,RIfc7c9d0_6440,RIfea0098_8165,RIfc57e00_6022,RIf13f550_5180,RIfcd6e08_7467,
        RIee3d900_5159,RIfc8f6c0_6654,RIfce0048_7571,RIfca27e8_6871,RIe1742e8_2699,RIfc7c700_6438,RIfc8f990_6656,RIfce9828_7679,RIfc583a0_6026,RIf16cdc0_5698,
        RIe224670_4704,RIf16c118_5689,RIe221970_4672,RIfc58508_6027,RIe21ec70_4640,RIe219270_4576,RIe216570_4544,RIfc3ff08_5753,RIe213870_4512,RIf1696e8_5659,
        RIe210b70_4480,RIfc58940_6030,RIe20de70_4448,RIe20b170_4416,RIe208470_4384,RIfc8fc60_6658,RIfc97820_6746,RIe202ea8_4323,RIe201288_4303,RIfcc27c8_7235,
        RIfcdfee0_7570,RIfc44198_5797,RIfc58670_6028,RIf1608e0_5558,RIf15e9f0_5536,RIfe9ff30_8164,RIe1fc0f8_4245,RIfc7be90_6432,RIf15bb88_5503,RIfcd8cf8_7489,
        RIfcd8e60_7490,RIfca2d88_6875,RIfcbdea8_7183,RIfcb3a20_7066,RIe1fabe0_4230,RIfc90098_6661,RIfc90200_6662,RIfcd20b0_7412,RIe1f6158_4177,RIfc904d0_6664,
        RIfca2ef0_6876,RIfc97550_6744,RIe1f3e30_4152,RIfc59048_6035,RIfc907a0_6666,RIfc90638_6665,RIe1eeb38_4093,RIe1ec3d8_4065,RIe1e96d8_4033,RIe1e69d8_4001,
        RIe1e3cd8_3969,RIe1e0fd8_3937,RIe1de2d8_3905,RIe1db5d8_3873,RIe1d88d8_3841,RIe1d2ed8_3777,RIe1d01d8_3745,RIe1cd4d8_3713,RIe1ca7d8_3681,RIe1c7ad8_3649,
        RIe1c4dd8_3617,RIe1c20d8_3585,RIe1bf3d8_3553,RIfcc73b8_7289,RIfce3cc0_7614,RIe1b9e10_3492,RIe1b7c50_3468,RIfcd6f70_7468,RIf149e10_5300,RIe1b5a90_3444,
        RIfea0200_8166,RIfc90bd8_6669,RIfcdfd78_7569,RIe1b2ef8_3413,RIe1b15a8_3395,RIfc973e8_6743,RIfcc7520_7290,RIe1acdf0_3344,RIe1ab608_3327,RIe1a9718_3305,
        RIe1a6a18_3273,RIe1a3d18_3241,RIe1a1018_3209,RIe18d518_2985,RIe179a18_2761,RIe227370_4736,RIe21bf70_4608,RIe205770_4352,RIe1ff7d0_4284,RIe1f8b88_4207,
        RIe1f16d0_4124,RIe1d5bd8_3809,RIe1bc6d8_3521,RIe1af550_3372,RIe171b88_2671,RIdec5108_706,RIdec2408_674,RIfc93608_6699,RIdebf708_642,RIfc934a0_6698,
        RIdebca08_610,RIdeb9d08_578,RIdeb7008_546,RIfcdf7d8_7565,RIdeb1608_482,RIfc78218_6389,RIdeae908_450,RIfcc8498_7301,RIdea9d90_418,RIdea3490_386,
        RIde9cb90_354,RIee1cc78_4786,RIee1bb98_4774,RIee1b328_4768,RIee1aab8_4762,RIde909f8_295,RIde8d578_279,RIfea8ea0_8238,RIde85238_239,RIde813e0_220,
        RIfc938d8_6701,RIfce5e80_7638,RIfcbfd98_7205,RIfce8ce8_7671,RIe16b4e0_2598,RIfea8d38_8237,RIfea9f80_8250,RIe165108_2527,RIe162408_2495,RIfc779a8_6383,
        RIe15f708_2463,RIfe9dc08_8139,RIe15ca08_2431,RIe157008_2367,RIe154308_2335,RIfea7550_8220,RIe151608_2303,RIfcd6160_7458,RIe14e908_2271,RIfcd1408_7403,
        RIe14bc08_2239,RIe148f08_2207,RIe146208_2175,RIfceb718_7701,RIfcb19c8_7043,RIfc93e78_6705,RIfce7938_7657,RIe140da8_2115,RIdf3ecb0_2091,RIdf3c988_2066,
        RIfe9daa0_8138,RIfce8478_7665,RIfcdbf98_7525,RIfc776d8_6381,RIfc93fe0_6706,RIdf354d0_1983,RIdf33040_1957,RIdf30fe8_1934,RIdf2ee28_1910,RIee2ba20_4955,
        RIfc93ba8_6703,RIfc77de0_6386,RIee27ad8_4910,RIfe9d668_8135,RIfea8bd0_8236,RIdf26458_1812,RIfe9d7d0_8136,RIfcb1c98_7045,RIee26cc8_4900,RIdf22ab0_1771,
        RIfcc0068_7207,RIdf21598_1756,RIdf1f6a8_1734,RIdf1aef0_1683,RIfe9d938_8137,RIdf16cd8_1636,RIdf13fd8_1604,RIdf112d8_1572,RIdf0e5d8_1540,RIdf0b8d8_1508,
        RIdf08bd8_1476,RIdf05ed8_1444,RIdf031d8_1412,RIdefd7d8_1348,RIdefaad8_1316,RIdef7dd8_1284,RIdef50d8_1252,RIdef23d8_1220,RIdeef6d8_1188,RIdeec9d8_1156,
        RIdee9cd8_1124,RIfc942b0_6708,RIfcde6f8_7553,RIfcd1138_7401,RIfcde860_7554,RIdee4878_1064,RIdee2af0_1043,RIdee0a98_1020,RIdede8d8_996,RIfc5c9f0_6076,
        RIee22240_4847,RIfcc8768_7303,RIee21160_4835,RIded95e0_937,RIded7150_911,RIded5260_889,RIfea76b8_8221,RIded0508_834,RIdecd808_802,RIdecab08_770,
        RIdec7e08_738,RIdeb4308_514,RIde96290_322,RIe16df10_2628,RIe159d08_2399,RIe143508_2143,RIdf37f00_2013,RIdf2c560_1881,RIdf1cde0_1705,RIdf004d8_1380,
        RIdee6fd8_1092,RIdedbd40_965,RIde7c1d8_195,RIe19d3a0_3166,RIe19a6a0_3134,RIfcb2c10_7056,RIe1979a0_3102,RIfc923c0_6686,RIe194ca0_3070,RIe191fa0_3038,
        RIe18f2a0_3006,RIe1898a0_2942,RIe186ba0_2910,RIfc422a8_5775,RIe183ea0_2878,RIfcbecb8_7193,RIe1811a0_2846,RIe17e4a0_2814,RIe17b7a0_2782,RIf142250_5212,
        RIf140bd0_5196,RIfec43f8_8353,RIe175968_2715,RIfc79b68_6407,RIf13efb0_5176,RIfc92528_6687,RIfcb2aa8_7055,RIfcd8320_7482,RIfcea200_7686,RIfc79898_6405,
        RIe1734d8_2689,RIfcd7948_7475,RIfcd7678_7473,RIf16e170_5712,RIfc927f8_6689,RIfc92960_6690,RIe2236f8_4693,RIfc795c8_6403,RIe2209f8_4661,RIf16ad68_5675,
        RIe21dcf8_4629,RIe2182f8_4565,RIe2155f8_4533,RIfe9d398_8133,RIe2128f8_4501,RIfcdb9f8_7521,RIe20fbf8_4469,RIfc41d08_5771,RIe20cef8_4437,RIe20a1f8_4405,
        RIe2074f8_4373,RIfcd7510_7472,RIf166010_5620,RIfe9d230_8132,RIe2008b0_4296,RIf165098_5609,RIfc41ba0_5770,RIfc41a38_5769,RIfc92c30_6692,RIfc418d0_5768,
        RIfc79190_6400,RIe1fcad0_4252,RIfec4560_8354,RIfc79028_6399,RIfcbf258_7197,RIfcc1df0_7228,RIfcd81b8_7481,RIfc92d98_6693,RIfc5b4d8_6061,RIfcd77e0_7474,
        RIe1fa0a0_4222,RIf156188_5439,RIfe9d500_8134,RIf1546d0_5420,RIe1f5348_4167,RIfec4830_8356,RIfec46c8_8355,RIf1508f0_5376,RIe1f3020_4142,RIfce3180_7606,
        RIfce8fb8_7673,RIfcbf690_7200,RIe1edd28_4083,RIe1eb460_4054,RIe1e8760_4022,RIe1e5a60_3990,RIe1e2d60_3958,RIe1e0060_3926,RIe1dd360_3894,RIe1da660_3862,
        RIe1d7960_3830,RIe1d1f60_3766,RIe1cf260_3734,RIe1cc560_3702,RIe1c9860_3670,RIe1c6b60_3638,RIe1c3e60_3606,RIe1c1160_3574,RIe1be460_3542,RIfe9d0c8_8131,
        RIfe9cc90_8128,RIe1b9168_3483,RIe1b7110_3460,RIf14a3b0_5304,RIfe9cb28_8127,RIfe9cf60_8130,RIfe9c9c0_8126,RIfce2208_7595,RIfce9558_7677,RIfe9c858_8125,
        RIfe9cdf8_8129,RIf147110_5268,RIf146468_5259,RIe1ac2b0_3336,RIe1aaac8_3319,RIe1a87a0_3294,RIe1a5aa0_3262,RIe1a2da0_3230,RIe1a00a0_3198,RIe18c5a0_2974,
        RIe178aa0_2750,RIe2263f8_4725,RIe21aff8_4597,RIe2047f8_4341,RIe1fe858_4273,RIe1f7c10_4196,RIe1f0758_4113,RIe1d4c60_3798,RIe1bb760_3510,RIe1ae5d8_3361,
        RIe170c10_2660,RIdec4190_695,RIdec1490_663,RIfceaa70_7692,RIdebe790_631,RIfc954f8_6721,RIdebba90_599,RIdeb8d90_567,RIdeb6090_535,RIfcebb50_7704,
        RIdeb0690_471,RIee1e190_4801,RIdead990_439,RIfcdf0d0_7560,RIdea7978_407,RIdea1078_375,RIde9a778_343,RIee1c840_4783,RIfc957c8_6723,RIfcc8e70_7308,
        RIfc5e610_6096,RIfe9e8b0_8148,RIde8c1c8_273,RIde88028_253,RIde83b40_232,RIfcb0bb8_7033,RIfca4b10_6896,RIfc75d88_6363,RIfca4c78_6897,RIfc95390_6720,
        RIe16a9a0_2590,RIfcc8fd8_7309,RIe166e90_2548,RIe164190_2516,RIe161490_2484,RIfe9e748_8147,RIe15e790_2452,RIfc74f78_6353,RIe15ba90_2420,RIe156090_2356,
        RIe153390_2324,RIfc3ecc0_5740,RIe150690_2292,RIfce8b80_7670,RIe14d990_2260,RIfca6730_6916,RIe14ac90_2228,RIe147f90_2196,RIe145290_2164,RIfcee2b0_7732,
        RIfc5f2b8_6105,RIfc753b0_6356,RIfc74b40_6350,RIe140268_2107,RIdf3e170_2083,RIdf3be48_2058,RIdf39c88_2034,RIfcc1c88_7227,RIfcc1850_7224,RIfc965d8_6733,
        RIfc96038_6729,RIdf34828_1974,RIdf327d0_1951,RIdf301d8_1924,RIdf2e2e8_1902,RIfc5e778_6097,RIfcd0328_7391,RIfc757e8_6359,RIfcee6e8_7735,RIdf296f8_1848,
        RIdf273d0_1823,RIdf257b0_1803,RIdf23b90_1783,RIfc95d68_6727,RIfceda40_7726,RIfe9eb80_8150,RIfc75518_6357,RIfcd01c0_7390,RIdf1eb68_1726,RIfe9ece8_8151,
        RIfe9ea18_8149,RIdf15d60_1625,RIdf13060_1593,RIdf10360_1561,RIdf0d660_1529,RIdf0a960_1497,RIdf07c60_1465,RIdf04f60_1433,RIdf02260_1401,RIdefc860_1337,
        RIdef9b60_1305,RIdef6e60_1273,RIdef4160_1241,RIdef1460_1209,RIdeee760_1177,RIdeeba60_1145,RIdee8d60_1113,RIfc961a0_6730,RIfc96308_6731,RIfc5ee80_6102,
        RIfce6150_7640,RIdee42d8_1060,RIdee1e48_1034,RIdee00c0_1013,RIdeddac8_986,RIfc96470_6732,RIfc75248_6355,RIfc74ca8_6351,RIfcb0618_7029,RIded8938_928,
        RIded6610_903,RIded4450_879,RIded2290_855,RIdecf590_823,RIdecc890_791,RIdec9b90_759,RIdec6e90_727,RIdeb3390_503,RIde93e78_311,RIe16cf98_2617,
        RIe158d90_2388,RIe142590_2132,RIdf36f88_2002,RIdf2b5e8_1870,RIdf1be68_1694,RIdeff560_1369,RIdee6060_1081,RIdedadc8_954,RIde79dc0_184,RIe19c428_3155,
        RIe199728_3123,RIfe9e310_8144,RIe196a28_3091,RIfcc04a0_7210,RIe193d28_3059,RIe191028_3027,RIe18e328_2995,RIe188928_2931,RIe185c28_2899,RIfce1830_7588,
        RIe182f28_2867,RIfe9e478_8145,RIe180228_2835,RIe17d528_2803,RIe17a828_2771,RIf141878_5205,RIfcb12c0_7038,RIfc94418_6709,RIe174f90_2708,RIfc77408_6379,
        RIf13ea10_5172,RIfcdc100_7526,RIfc94580_6710,RIfc946e8_6711,RIfced338_7721,RIfce5fe8_7639,RIe172998_2681,RIfcdc268_7527,RIfcddff0_7548,RIfcc0608_7211,
        RIfce7230_7652,RIfc40340_5756,RIe222780_4682,RIfcdd618_7541,RIe21fa80_4650,RIfcd0b98_7397,RIe21cd80_4618,RIe217380_4554,RIe214680_4522,RIfec4998_8357,
        RIe211980_4490,RIf168608_5647,RIe20ec80_4458,RIfcc0770_7212,RIe20bf80_4426,RIe209280_4394,RIe206580_4362,RIfce2370_7596,RIfcee580_7734,RIfec4c68_8359,
        RIfec4b00_8358,RIfc949b8_6713,RIfcebcb8_7705,RIf162938_5581,RIf1612b8_5565,RIfccd088_7355,RIfcc08d8_7213,RIfe9e040_8142,RIfe9e1a8_8143,RIfcead40_7694,
        RIf15ad78_5493,RIfc94c88_6715,RIfccc3e0_7346,RIfc765f8_6369,RIfc94df0_6716,RIfcc0a40_7214,RIe1f9998_4217,RIfcc8d08_7307,RIfce8748_7667,RIfceb2e0_7698,
        RIe1f4970_4160,RIf152510_5396,RIf1512c8_5383,RIfcb0ff0_7036,RIe1f24e0_4134,RIfc761c0_6366,RIfc950c0_6718,RIfcc0e78_7217,RIe1ed1e8_4075,RIe1ea4e8_4043,
        RIe1e77e8_4011,RIe1e4ae8_3979,RIe1e1de8_3947,RIe1df0e8_3915,RIe1dc3e8_3883,RIe1d96e8_3851,RIe1d69e8_3819,RIe1d0fe8_3755,RIe1ce2e8_3723,RIe1cb5e8_3691,
        RIe1c88e8_3659,RIe1c5be8_3627,RIe1c2ee8_3595,RIe1c01e8_3563,RIe1bd4e8_3531,RIf14bfd0_5324,RIf14ac20_5310,RIfe9ded8_8141,RIe1b65d0_3452,RIfcecd98_7717,
        RIfc76490_6368,RIe1b4c80_3434,RIe1b38d0_3420,RIfcc0fe0_7218,RIfceaea8_7695,RIe1b1f80_3402,RIe1b0360_3382,RIfcd0760_7394,RIf145ec8_5255,RIfe9e5e0_8146,
        RIfe9dd70_8140,RIe1a7828_3283,RIe1a4b28_3251,RIe1a1e28_3219,RIe19f128_3187,RIe18b628_2963,RIe177b28_2739,RIe225480_4714,RIe21a080_4586,RIe203880_4330,
        RIe1fd8e0_4262,RIe1f6c98_4185,RIe1ef7e0_4102,RIe1d3ce8_3787,RIe1ba7e8_3499,RIe1ad660_3350,RIe16fc98_2649,RIdec6788_722,RIdec3a88_690,RIee20788_4828,
        RIdec0d88_658,RIee1f810_4817,RIdebe088_626,RIdebb388_594,RIdeb8688_562,RIfc9b1c8_6787,RIdeb2c88_498,RIfce1f38_7593,RIdeaff88_466,RIfc892e8_6583,
        RIdead210_434,RIdea6910_402,RIdea0010_370,RIee1d650_4793,RIee1c570_4781,RIee1b5f8_4770,RIee1aef0_4765,RIfe99888_8091,RIfe99450_8088,RIfe99720_8090,
        RIfe995b8_8089,RIde83168_229,RIfcc43e8_7255,RIfcd5a58_7453,RIfc89450_6584,RIfcc5798_7269,RIe16c890_2612,RIe16a568_2587,RIe168d80_2570,RIe166788_2543,
        RIe163a88_2511,RIfc83618_6517,RIe160d88_2479,RIee36718_5078,RIe15e088_2447,RIe158688_2383,RIe155988_2351,RIfc3f800_5748,RIe152c88_2319,RIfc895b8_6585,
        RIe14ff88_2287,RIfc51cf8_5953,RIe14d288_2255,RIe14a588_2223,RIe147888_2191,RIee34990_5057,RIee338b0_5045,RIfc831e0_6514,RIfcd3b68_7431,RIe141ff0_2128,
        RIe13fcc8_2103,RIdf3dbd0_2079,RIdf3b740_2053,RIfcb6f90_7104,RIee301d8_5006,RIfcba938_7145,RIee2e018_4982,RIdf369e8_1998,RIdf343f0_1971,RIdf32230_1947,
        RIfe99e28_8095,RIfc83078_6513,RIfcb6e28_7103,RIfc9ad90_6784,RIfcbad70_7148,RIdf2b1b0_1867,RIdf292c0_1845,RIfe99b58_8093,RIfe999f0_8092,RIfc9ac28_6783,
        RIfc4a9a8_5871,RIdf23758_1780,RIfc82da8_6511,RIdf220d8_1764,RIdf20a58_1748,RIdf1ba30_1691,RIfe99cc0_8094,RIdf18358_1652,RIdf15658_1620,RIdf12958_1588,
        RIdf0fc58_1556,RIdf0cf58_1524,RIdf0a258_1492,RIdf07558_1460,RIdf04858_1428,RIdefee58_1364,RIdefc158_1332,RIdef9458_1300,RIdef6758_1268,RIdef3a58_1236,
        RIdef0d58_1204,RIdeee058_1172,RIdeeb358_1140,RIee25918_4886,RIee24b08_4876,RIfc52568_5959,RIfc826a0_6506,RIdee5958_1076,RIdee3bd0_1055,RIfe99f90_8096,
        RIdedf9b8_1008,RIfce4800_7622,RIfc89b58_6589,RIfc9f3e0_6834,RIfc82538_6505,RIdeda828_950,RIded8398_924,RIfeabe70_8272,RIded3eb0_875,RIded1b88_850,
        RIdecee88_818,RIdecc188_786,RIdec9488_754,RIdeb5988_530,RIde99710_338,RIe16f590_2644,RIe15b388_2415,RIe144b88_2159,RIdf39580_2029,RIdf2dbe0_1897,
        RIdf1e460_1721,RIdf01b58_1396,RIdee8658_1108,RIdedd3c0_981,RIde7f658_211,RIe19ea20_3182,RIe19bd20_3150,RIf145928_5251,RIe199020_3118,RIfe98910_8080,
        RIe196320_3086,RIe193620_3054,RIe190920_3022,RIe18af20_2958,RIe188220_2926,RIf143e70_5232,RIe185520_2894,RIfc95c00_6726,RIe182820_2862,RIe17fb20_2830,
        RIe17ce20_2798,RIf142520_5214,RIf141440_5202,RIe1776f0_2736,RIfeab8d0_8268,RIfcc5bd0_7272,RIfc62dc8_6147,RIee3e710_5169,RIfc9cb18_6805,RIee3c820_5147,
        RIee3b470_5133,RIee3a390_5121,RIe174888_2703,RIf170498_5737,RIfc68660_6210,RIf16e878_5717,RIfc6ea38_6281,RIfe98d48_8083,RIe224d78_4709,RIf16c280_5690,
        RIe222078_4677,RIf16b308_5679,RIe21f378_4645,RIe219978_4581,RIe216c78_4549,RIf16a390_5668,RIe213f78_4517,RIf169b20_5662,RIe211278_4485,RIf1681d0_5644,
        RIe20e578_4453,RIe20b878_4421,RIe208b78_4389,RIfcd4ae0_7442,RIfc61478_6129,RIfeab060_8262,RIe201990_4308,RIfc70ec8_6307,RIfc70928_6303,RIfcec528_7711,
        RIfcbe880_7190,RIf160d18_5561,RIf15ee28_5539,RIfe98be0_8082,RIfe98eb0_8084,RIf15d0a0_5518,RIf15bcf0_5504,RIfcd4540_7438,RIf159e00_5482,RIf1592c0_5474,
        RIf158078_5461,RIfca3a30_6884,RIfea7988_8223,RIf156728_5443,RIf155be8_5435,RIf154b08_5423,RIfe98a78_8081,RIf1538c0_5410,RIf1520d8_5393,RIf150e90_5380,
        RIe1f43d0_4156,RIf14fdb0_5368,RIfcd2380_7414,RIf14e2f8_5349,RIe1ef240_4098,RIe1ecae0_4070,RIe1e9de0_4038,RIe1e70e0_4006,RIe1e43e0_3974,RIe1e16e0_3942,
        RIe1de9e0_3910,RIe1dbce0_3878,RIe1d8fe0_3846,RIe1d35e0_3782,RIe1d08e0_3750,RIe1cdbe0_3718,RIe1caee0_3686,RIe1c81e0_3654,RIe1c54e0_3622,RIe1c27e0_3590,
        RIe1bfae0_3558,RIfc44b70_5804,RIf14bd00_5322,RIfe992e8_8087,RIfe987a8_8079,RIf14a950_5308,RIf149f78_5301,RIfe99180_8086,RIfe98640_8078,RIf149438_5293,
        RIfcec7f8_7713,RIfe984d8_8077,RIe1b1b48_3399,RIfc4b650_5880,RIfcda918_7509,RIfe98370_8076,RIfe99018_8085,RIe1a9e20_3310,RIe1a7120_3278,RIe1a4420_3246,
        RIe1a1720_3214,RIe18dc20_2990,RIe17a120_2766,RIe227a78_4741,RIe21c678_4613,RIe205e78_4357,RIe1ffed8_4289,RIe1f9290_4212,RIe1f1dd8_4129,RIe1d62e0_3814,
        RIe1bcde0_3526,RIe1afc58_3377,RIe172290_2676,RIdec6620_721,RIdec3920_689,RIfc49328_5855,RIdec0c20_657,RIfc80eb8_6489,RIdebdf20_625,RIdebb220_593,
        RIdeb8520_561,RIfc80648_6483,RIdeb2b20_497,RIfc8b340_6606,RIdeafe20_465,RIfc491c0_5854,RIdeacec8_433,RIdea65c8_401,RIde9fcc8_369,RIfcd9c70_7500,
        RIfe98208_8075,RIfce4698_7621,RIfe980a0_8074,RIde93158_307,RIde8f648_289,RIde8b4a8_269,RIde87308_249,RIde82e20_228,RIfcbba18_7157,RIfc48d88_5851,
        RIfc99f80_6774,RIfc8b4a8_6607,RIe16c728_2611,RIe16a400_2586,RIe168c18_2569,RIe166620_2542,RIe163920_2510,RIee38068_5096,RIe160c20_2478,RIfc48248_5843,
        RIe15df20_2446,RIe158520_2382,RIe155820_2350,RIfcbbe50_7160,RIe152b20_2318,RIfc47e10_5840,RIe14fe20_2286,RIfca0e98_6853,RIe14d120_2254,RIe14a420_2222,
        RIe147720_2190,RIfc8be80_6614,RIfc7fb08_6475,RIfc480e0_5842,RIfc99878_6769,RIe141e88_2127,RIe13fb60_2102,RIdf3da68_2078,RIdf3b5d8_2052,RIfe97f38_8073,
        RIee30070_5005,RIee2eb58_4990,RIee2deb0_4981,RIdf36880_1997,RIdf34288_1970,RIdf320c8_1946,RIfe97dd0_8072,RIfcc3740_7246,RIfc48ab8_5849,RIfce05e8_7575,
        RIfc80210_6480,RIdf2b048_1866,RIdf29158_1844,RIdf26f98_1820,RIdf254e0_1801,RIfc8bbb0_6612,RIfc48950_5848,RIdf235f0_1779,RIfc8bd18_6613,RIdf21f70_1763,
        RIdf208f0_1747,RIdf1b8c8_1690,RIdf1a3b0_1675,RIdf181f0_1651,RIdf154f0_1619,RIdf127f0_1587,RIdf0faf0_1555,RIdf0cdf0_1523,RIdf0a0f0_1491,RIdf073f0_1459,
        RIdf046f0_1427,RIdefecf0_1363,RIdefbff0_1331,RIdef92f0_1299,RIdef65f0_1267,RIdef38f0_1235,RIdef0bf0_1203,RIdeedef0_1171,RIdeeb1f0_1139,RIfcbc120_7162,
        RIfcd9838_7497,RIfc99710_6768,RIfca1168_6855,RIdee57f0_1075,RIdee3a68_1054,RIdee18a8_1030,RIdedf850_1007,RIfc549f8_5985,RIfcb5370_7084,RIfce43c8_7619,
        RIfce0480_7574,RIdeda6c0_949,RIded8230_923,RIded6070_899,RIded3d48_874,RIded1a20_849,RIdeced20_817,RIdecc020_785,RIdec9320_753,RIdeb5820_529,
        RIde993c8_337,RIe16f428_2643,RIe15b220_2414,RIe144a20_2158,RIdf39418_2028,RIdf2da78_1896,RIdf1e2f8_1720,RIdf019f0_1395,RIdee84f0_1107,RIdedd258_980,
        RIde7f310_210,RIe19e8b8_3181,RIe19bbb8_3149,RIfe976c8_8067,RIe198eb8_3117,RIf144c80_5242,RIe1961b8_3085,RIe1934b8_3053,RIe1907b8_3021,RIe18adb8_2957,
        RIe1880b8_2925,RIfe97560_8066,RIe1853b8_2893,RIfcc3fb0_7252,RIe1826b8_2861,RIe17f9b8_2829,RIe17ccb8_2797,RIfcd3730_7428,RIf1412d8_5201,RIfcc4118_7253,
        RIfe97830_8068,RIfc4a6d8_5869,RIf13f6b8_5181,RIfc9f980_6838,RIfc9fae8_6839,RIfcc3e48_7251,RIfc89e28_6591,RIfc89cc0_6590,RIe174720_2702,RIfc4a408_5867,
        RIfce27a8_7599,RIfc530a8_5967,RIfcd5d28_7455,RIf16cf28_5699,RIe224c10_4708,RIfc53210_5968,RIe221f10_4676,RIf16b1a0_5678,RIe21f210_4644,RIe219810_4580,
        RIe216b10_4548,RIfc401d8_5755,RIe213e10_4516,RIf1699b8_5661,RIe211110_4484,RIfc81cc8_6499,RIe20e410_4452,RIe20b710_4420,RIe208a10_4388,RIfc8a0f8_6593,
        RIfcb6720_7098,RIe203448_4327,RIe201828_4307,RIfc53378_5969,RIfc8a3c8_6595,RIfcb65b8_7097,RIfc49fd0_5864,RIf160bb0_5560,RIf15ecc0_5538,RIe1fd4a8_4259,
        RIfe97b00_8070,RIfc8a530_6596,RIfe97c68_8071,RIfc8a800_6598,RIfc8a698_6597,RIfc9a7f0_6780,RIfc81890_6496,RIfcd5e90_7456,RIe1fb180_4234,RIfc49e68_5863,
        RIfc81728_6495,RIfcbb1a8_7151,RIe1f66f8_4181,RIfcd3460_7426,RIfcb62e8_7095,RIfc9a520_6778,RIe1f4268_4155,RIfc49d00_5862,RIfcd9dd8_7501,RIfcbb310_7152,
        RIe1ef0d8_4097,RIe1ec978_4069,RIe1e9c78_4037,RIe1e6f78_4005,RIe1e4278_3973,RIe1e1578_3941,RIe1de878_3909,RIe1dbb78_3877,RIe1d8e78_3845,RIe1d3478_3781,
        RIe1d0778_3749,RIe1cda78_3717,RIe1cad78_3685,RIe1c8078_3653,RIe1c5378_3621,RIe1c2678_3589,RIe1bf978_3557,RIfc49a30_5860,RIfcb6018_7093,RIe1ba3b0_3496,
        RIe1b81f0_3472,RIfce0a20_7578,RIfcbb5e0_7154,RIe1b6030_3448,RIfe97998_8069,RIfce5610_7632,RIfcc3a10_7248,RIe1b3330_3416,RIe1b19e0_3398,RIfc495f8_5857,
        RIfc81188_6491,RIe1ad228_3347,RIe1aba40_3330,RIe1a9cb8_3309,RIe1a6fb8_3277,RIe1a42b8_3245,RIe1a15b8_3213,RIe18dab8_2989,RIe179fb8_2765,RIe227910_4740,
        RIe21c510_4612,RIe205d10_4356,RIe1ffd70_4288,RIe1f9128_4211,RIe1f1c70_4128,RIe1d6178_3813,RIe1bcc78_3525,RIe1afaf0_3376,RIe172128_2675,RIdec6a58_724,
        RIdec3d58_692,RIfc723e0_6322,RIdec1058_660,RIfc59fc0_6046,RIdebe358_628,RIdebb658_596,RIdeb8958_564,RIfcb96f0_7132,RIdeb2f58_500,RIfce1c68_7591,
        RIdeb0258_468,RIfc9b498_6789,RIdead558_436,RIdea6fa0_404,RIdea06a0_372,RIfc81458_6493,RIfc83780_6518,RIfc4e620_5914,RIfcd3e38_7433,RIde937e8_309,
        RIde8f990_290,RIde8bb38_271,RIde87650_250,RIde834b0_230,RIfc42c80_5782,RIfc65960_6178,RIfc6c710_6256,RIee392b0_5109,RIe16cb60_2614,RIe16a6d0_2588,
        RIe169050_2572,RIe166a58_2545,RIe163d58_2513,RIfec3cf0_8348,RIe161058_2481,RIfcd54b8_7449,RIe15e358_2449,RIe158958_2385,RIe155c58_2353,RIfe9ba48_8115,
        RIe152f58_2321,RIfec4128_8351,RIe150258_2289,RIfcb9b28_7135,RIe14d558_2257,RIe14a858_2225,RIe147b58_2193,RIfcdb2f0_7516,RIfc553d0_5992,RIfc9a0e8_6775,
        RIfcbd908_7179,RIe1422c0_2130,RIe13ff98_2105,RIdf3dea0_2081,RIdf3ba10_2055,RIfc87128_6559,RIee304a8_5008,RIfcc51f8_7265,RIee2e2e8_4984,RIdf36cb8_2000,
        RIfec3fc0_8350,RIdf32500_1949,RIfec3e58_8349,RIee2c830_4965,RIee2ad78_4946,RIee296f8_4930,RIee284b0_4917,RIfe9b8e0_8114,RIfe9b610_8112,RIfe9b778_8113,
        RIfe9b4a8_8111,RIfcb7c38_7113,RIfc86b88_6555,RIdf238c0_1781,RIfc75ab8_6361,RIdf22240_1765,RIfeaa3b8_8253,RIdf1bb98_1692,RIdf1a680_1677,RIdf18628_1654,
        RIdf15928_1622,RIdf12c28_1590,RIdf0ff28_1558,RIdf0d228_1526,RIdf0a528_1494,RIdf07828_1462,RIdf04b28_1430,RIdeff128_1366,RIdefc428_1334,RIdef9728_1302,
        RIdef6a28_1270,RIdef3d28_1238,RIdef1028_1206,RIdeee328_1174,RIdeeb628_1142,RIee25a80_4887,RIee24c70_4877,RIfcddd20_7546,RIfccc110_7344,RIdee5c28_1078,
        RIdee3ea0_1057,RIdee1b78_1032,RIdedfc88_1010,RIfc6a6b8_6233,RIee227e0_4851,RIfc88be0_6578,RIee21868_4840,RIdedaaf8_952,RIded8668_926,RIded6340_901,
        RIded4180_877,RIded1e58_852,RIdecf158_820,RIdecc458_788,RIdec9758_756,RIdeb5c58_532,RIde99da0_340,RIe16f860_2646,RIe15b658_2417,RIe144e58_2161,
        RIdf39850_2031,RIdf2deb0_1899,RIdf1e730_1723,RIdf01e28_1398,RIdee8928_1110,RIdedd690_983,RIde7fce8_213,RIe19ecf0_3184,RIe19bff0_3152,RIf145a90_5252,
        RIe1992f0_3120,RIf144de8_5243,RIe1965f0_3088,RIe1938f0_3056,RIe190bf0_3024,RIe18b1f0_2960,RIe1884f0_2928,RIfc72980_6326,RIe1857f0_2896,RIf143060_5222,
        RIe182af0_2864,RIe17fdf0_2832,RIe17d0f0_2800,RIf142688_5215,RIf141710_5204,RIe177858_2737,RIe176778_2725,RIfcea638_7689,RIfca54e8_6903,RIee3e878_5170,
        RIee3dbd0_5161,RIee3c988_5148,RIee3b5d8_5134,RIee3a4f8_5122,RIe174b58_2705,RIf170600_5738,RIfc76fd0_6376,RIf16e9e0_5718,RIfced608_7723,RIf16d090_5700,
        RIe225048_4711,RIf16c550_5692,RIe222348_4679,RIf16b470_5680,RIe21f648_4647,RIe219c48_4583,RIe216f48_4551,RIf16a4f8_5669,RIe214248_4519,RIf169df0_5664,
        RIe211548_4487,RIf1684a0_5646,RIe20e848_4455,RIe20bb48_4423,RIe208e48_4391,RIf1673c0_5634,RIf166448_5623,RIfe9c6f0_8124,RIfe9c150_8120,RIf1654d0_5612,
        RIfcc4550_7256,RIf1635e0_5590,RIf162500_5578,RIf160fe8_5563,RIf15f0f8_5541,RIfe9bfe8_8119,RIfe9c588_8123,RIf15d208_5519,RIf15bfc0_5506,RIfc4d540_5902,
        RIfc9c848_6803,RIfec4290_8352,RIfe9c2b8_8121,RIfcc01d0_7208,RIe1fb2e8_4235,RIfe9c420_8122,RIfca3e68_6887,RIf154c70_5424,RIe1f69c8_4183,RIf153a28_5411,
        RIf152240_5394,RIf150ff8_5381,RIe1f46a0_4158,RIfca6028_6911,RIfc43bf8_5793,RIf14e460_5350,RIe1ef3a8_4099,RIe1ecdb0_4072,RIe1ea0b0_4040,RIe1e73b0_4008,
        RIe1e46b0_3976,RIe1e19b0_3944,RIe1decb0_3912,RIe1dbfb0_3880,RIe1d92b0_3848,RIe1d38b0_3784,RIe1d0bb0_3752,RIe1cdeb0_3720,RIe1cb1b0_3688,RIe1c84b0_3656,
        RIe1c57b0_3624,RIe1c2ab0_3592,RIe1bfdb0_3560,RIfc4d6a8_5903,RIf14be68_5323,RIe1ba680_3498,RIfe9be80_8118,RIfc86e58_6557,RIfcd46a8_7439,RIe1b6300_3450,
        RIfe9bd18_8117,RIf1495a0_5294,RIf1481f0_5280,RIe1b3600_3418,RIe1b1e18_3401,RIfc69470_6220,RIfcbfac8_7203,RIfe9bbb0_8116,RIe1abd10_3332,RIe1aa0f0_3312,
        RIe1a73f0_3280,RIe1a46f0_3248,RIe1a19f0_3216,RIe18def0_2992,RIe17a3f0_2768,RIe227d48_4743,RIe21c948_4615,RIe206148_4359,RIe2001a8_4291,RIe1f9560_4214,
        RIe1f20a8_4131,RIe1d65b0_3816,RIe1bd0b0_3528,RIe1aff28_3379,RIe172560_2678,RIdec68f0_723,RIdec3bf0_691,RIee208f0_4829,RIdec0ef0_659,RIfc7ce08_6443,
        RIdebe1f0_627,RIdebb4f0_595,RIdeb87f0_563,RIfc9b8d0_6792,RIdeb2df0_499,RIfcc6710_7280,RIdeb00f0_467,RIfc5ff60_6114,RIdead3f0_435,RIdea6c58_403,
        RIdea0358_371,RIfce5070_7628,RIee1c6d8_4782,RIfce70c8_7651,RIee1b058_4766,RIde934a0_308,RIfe9b1d8_8109,RIde8b7f0_270,RIfe9b340_8110,RIfc6b798_6245,
        RIfcb2238_7049,RIfcd3a00_7430,RIfcdb020_7514,RIfc511b8_5945,RIe16c9f8_2613,RIfcb27d8_7053,RIe168ee8_2571,RIe1668f0_2544,RIe163bf0_2512,RIee381d0_5097,
        RIe160ef0_2480,RIfcdfaa8_7567,RIe15e1f0_2448,RIe1587f0_2384,RIe155af0_2352,RIfc3f968_5749,RIe152df0_2320,RIfcd5080_7446,RIe1500f0_2288,RIfc84b30_6532,
        RIe14d3f0_2256,RIe14a6f0_2224,RIe1479f0_2192,RIfcea098_7685,RIfc92f00_6694,RIfc54890_5984,RIfcdcc40_7534,RIe142158_2129,RIe13fe30_2104,RIdf3dd38_2080,
        RIdf3b8a8_2054,RIfc57590_6016,RIee30340_5007,RIfcd0490_7392,RIee2e180_4983,RIdf36b50_1999,RIdf34558_1972,RIdf32398_1948,RIfe9b070_8108,RIfcb1860_7042,
        RIfca1b40_6862,RIfc5c018_6069,RIfe9ada0_8106,RIdf2b318_1868,RIdf29428_1846,RIdf27100_1821,RIfe9af08_8107,RIfc5e1d8_6093,RIfcdcda8_7535,RIfcac400_6982,
        RIfc691a0_6218,RIfcaad80_6966,RIdf20bc0_1749,RIfc61b80_6134,RIdf1a518_1676,RIdf184c0_1653,RIdf157c0_1621,RIdf12ac0_1589,RIdf0fdc0_1557,RIdf0d0c0_1525,
        RIdf0a3c0_1493,RIdf076c0_1461,RIdf049c0_1429,RIdefefc0_1365,RIdefc2c0_1333,RIdef95c0_1301,RIdef68c0_1269,RIdef3bc0_1237,RIdef0ec0_1205,RIdeee1c0_1173,
        RIdeeb4c0_1141,RIfc69b78_6225,RIfc6b900_6246,RIfc4d270_5900,RIfced770_7724,RIdee5ac0_1077,RIdee3d38_1056,RIdee1a10_1031,RIdedfb20_1009,RIfc7ff40_6478,
        RIfca4408_6891,RIfcb5640_7086,RIee21700_4839,RIdeda990_951,RIded8500_925,RIded61d8_900,RIded4018_876,RIded1cf0_851,RIdeceff0_819,RIdecc2f0_787,
        RIdec95f0_755,RIdeb5af0_531,RIde99a58_339,RIe16f6f8_2645,RIe15b4f0_2416,RIe144cf0_2160,RIdf396e8_2030,RIdf2dd48_1898,RIdf1e5c8_1722,RIdf01cc0_1397,
        RIdee87c0_1109,RIdedd528_982,RIde7f9a0_212,RIe19eb88_3183,RIe19be88_3151,RIfe9a698_8101,RIe199188_3119,RIfe9a530_8100,RIe196488_3087,RIe193788_3055,
        RIe190a88_3023,RIe18b088_2959,RIe188388_2927,RIfe9a800_8102,RIe185688_2895,RIfc8d938_6633,RIe182988_2863,RIe17fc88_2831,RIe17cf88_2799,RIfe9a3c8_8099,
        RIf1415a8_5203,RIfe9a260_8098,RIfe9a0f8_8097,RIfcb9150_7128,RIf13f820_5182,RIfc9fc50_6840,RIfce5340_7630,RIfc5cb58_6077,RIfc576f8_6017,RIfc780b0_6388,
        RIe1749f0_2704,RIfc7adb0_6420,RIfc7c2c8_6435,RIfcb2d78_7057,RIfc7e758_6461,RIfe9aad0_8104,RIe224ee0_4710,RIf16c3e8_5691,RIe2221e0_4678,RIfcd3898_7429,
        RIe21f4e0_4646,RIe219ae0_4582,RIe216de0_4550,RIfc880a0_6570,RIe2140e0_4518,RIf169c88_5663,RIe2113e0_4486,RIf168338_5645,RIe20e6e0_4454,RIe20b9e0_4422,
        RIe208ce0_4390,RIfce4c38_7625,RIfc9c6e0_6802,RIe2035b0_4328,RIe201af8_4309,RIfc500d8_5933,RIfc85c10_6544,RIfce81a8_7663,RIfce9c60_7682,RIf160e80_5562,
        RIf15ef90_5540,RIfe9a968_8103,RIfe9ac38_8105,RIfca8d28_6943,RIf15be58_5505,RIfcedba8_7727,RIfc6a988_6235,RIfc71cd8_6317,RIfccb198_7333,RIfcaa3a8_6959,
        RIfec3b88_8347,RIfc4c730_5892,RIfc6d688_6267,RIfca8e90_6944,RIe1f6860_4182,RIfc64e20_6170,RIfcaee30_7012,RIfccee10_7376,RIe1f4538_4157,RIfc63ea8_6159,
        RIfcaecc8_7011,RIfcae458_7005,RIfeab1c8_8263,RIe1ecc48_4071,RIe1e9f48_4039,RIe1e7248_4007,RIe1e4548_3975,RIe1e1848_3943,RIe1deb48_3911,RIe1dbe48_3879,
        RIe1d9148_3847,RIe1d3748_3783,RIe1d0a48_3751,RIe1cdd48_3719,RIe1cb048_3687,RIe1c8348_3655,RIe1c5648_3623,RIe1c2948_3591,RIe1bfc48_3559,RIfcc70e8_7287,
        RIfca7ae0_6930,RIe1ba518_3497,RIe1b8358_3473,RIfc598b8_6041,RIfcc2228_7231,RIe1b6198_3449,RIe1b4848_3431,RIfc82f10_6512,RIfc55970_5996,RIe1b3498_3417,
        RIe1b1cb0_3400,RIfcb7698_7109,RIfc4b4e8_5879,RIe1ad390_3348,RIe1abba8_3331,RIe1a9f88_3311,RIe1a7288_3279,RIe1a4588_3247,RIe1a1888_3215,RIe18dd88_2991,
        RIe17a288_2767,RIe227be0_4742,RIe21c7e0_4614,RIe205fe0_4358,RIe200040_4290,RIe1f93f8_4213,RIe1f1f40_4130,RIe1d6448_3815,RIe1bcf48_3527,RIe1afdc0_3378,
        RIe1723f8_2677,RIdec6d28_726,RIdec4028_694,RIee20bc0_4831,RIdec1328_662,RIfcbaed8_7149,RIdebe628_630,RIdebb928_598,RIdeb8c28_566,RIfc412b8_5767,
        RIdeb3228_502,RIfc9ea08_6827,RIdeb0528_470,RIee1e028_4800,RIdead828_438,RIdea7630_406,RIdea0d30_374,RIfcbac08_7147,RIfc55538_5993,RIfcba668_7143,
        RIfc4af48_5875,RIfe912f0_7996,RIfe91458_7997,RIde8be80_272,RIde87ce0_252,RIfc85238_6537,RIfc88640_6574,RIfcda210_7504,RIfcd5788_7451,RIee39418_5110,
        RIe16ce30_2616,RIfc884d8_6573,RIe169320_2574,RIe166d28_2547,RIe164028_2515,RIfe90918_7989,RIe161328_2483,RIee36880_5079,RIe15e628_2451,RIe158c28_2387,
        RIe155f28_2355,RIfe91188_7995,RIe153228_2323,RIfe91020_7994,RIe150528_2291,RIfcda378_7505,RIe14d828_2259,RIe14ab28_2227,RIe147e28_2195,RIfe90eb8_7993,
        RIfe90d50_7992,RIfcb99c0_7134,RIfc9c2a8_6799,RIfe90be8_7991,RIfe90a80_7990,RIdf3e008_2082,RIdf3bce0_2057,RIfcec690_7712,RIee30778_5010,RIfc87dd0_6568,
        RIee2e5b8_4986,RIdf36e20_2001,RIdf346c0_1973,RIdf32668_1950,RIdf30070_1923,RIee2c998_4966,RIee2aee0_4947,RIee299c8_4932,RIee28618_4918,RIfe90378_7985,
        RIfe907b0_7988,RIfe904e0_7986,RIfe90648_7987,RIfc9d928_6815,RIfc86048_6547,RIfcb92b8_7129,RIfc4ee90_5920,RIfc86a20_6554,RIdf20e90_1751,RIfcb8fe8_7127,
        RIdf1a950_1679,RIdf188f8_1656,RIdf15bf8_1624,RIdf12ef8_1592,RIdf101f8_1560,RIdf0d4f8_1528,RIdf0a7f8_1496,RIdf07af8_1464,RIdf04df8_1432,RIdeff3f8_1368,
        RIdefc6f8_1336,RIdef99f8_1304,RIdef6cf8_1272,RIdef3ff8_1240,RIdef12f8_1208,RIdeee5f8_1176,RIdeeb8f8_1144,RIfc857d8_6541,RIee24dd8_4878,RIfc4ff70_5932,
        RIfc50240_5934,RIdee5ef8_1080,RIdee4170_1059,RIfe915c0_7998,RIdedff58_1012,RIfcd4810_7440,RIee22948_4852,RIfce1560_7586,RIee219d0_4841,RIdedac60_953,
        RIfe91728_7999,RIded64a8_902,RIfe91890_8000,RIded2128_854,RIdecf428_822,RIdecc728_790,RIdec9a28_758,RIdeb5f28_534,RIde9a430_342,RIe16fb30_2648,
        RIe15b928_2419,RIe145128_2163,RIdf39b20_2033,RIdf2e180_1901,RIdf1ea00_1725,RIdf020f8_1400,RIdee8bf8_1112,RIdedd960_985,RIde80378_215,RIe19efc0_3186,
        RIe19c2c0_3154,RIf145d60_5254,RIe1995c0_3122,RIfc637a0_6154,RIe1968c0_3090,RIe193bc0_3058,RIe190ec0_3026,RIe18b4c0_2962,RIe1887c0_2930,RIfc62af8_6145,
        RIe185ac0_2898,RIfe8fc70_7980,RIe182dc0_2866,RIe1800c0_2834,RIe17d3c0_2802,RIfe90210_7984,RIfe8ff40_7982,RIfc72f20_6330,RIe176a48_2727,RIfcaf6a0_7018,
        RIfc61040_6126,RIf13e8a8_5171,RIfe900a8_7983,RIee3caf0_5149,RIee3b740_5135,RIee3a660_5123,RIe174e28_2707,RIf170768_5739,RIfc5fdf8_6113,RIf16eb48_5719,
        RIfcaaab0_6964,RIf16d1f8_5701,RIe225318_4713,RIf16c6b8_5693,RIe222618_4681,RIf16b5d8_5681,RIe21f918_4649,RIe219f18_4585,RIe217218_4553,RIfca62f8_6913,
        RIe214518_4521,RIfcc9578_7313,RIe211818_4489,RIfca5a88_6907,RIe20eb18_4457,RIe20be18_4425,RIe209118_4393,RIf167690_5636,RIf166718_5625,RIfe8f9a0_7978,
        RIfe8f838_7977,RIf165638_5613,RIf164990_5604,RIf1638b0_5592,RIf1627d0_5580,RIf161150_5564,RIf15f260_5542,RIe1fd778_4261,RIe1fc530_4248,RIf15d4d8_5521,
        RIf15c290_5508,RIfca20e0_6866,RIf159f68_5483,RIf159428_5475,RIf1581e0_5462,RIfc5ebb0_6100,RIfe8fdd8_7981,RIfc69e48_6227,RIfc5e8e0_6098,RIf154f40_5426,
        RIe1f6b30_4184,RIf153b90_5412,RIf1523a8_5395,RIfce88b0_7668,RIfe8fb08_7979,RIfcebe20_7706,RIfcb1158_7037,RIf14e730_5352,RIe1ef678_4101,RIe1ed080_4074,
        RIe1ea380_4042,RIe1e7680_4010,RIe1e4980_3978,RIe1e1c80_3946,RIe1def80_3914,RIe1dc280_3882,RIe1d9580_3850,RIe1d3b80_3786,RIe1d0e80_3754,RIe1ce180_3722,
        RIe1cb480_3690,RIe1c8780_3658,RIe1c5a80_3626,RIe1c2d80_3594,RIe1c0080_3562,RIfcc8ba0_7306,RIfc5d698_6085,RIfec35e8_8343,RIfeabd08_8271,RIfc5cf90_6080,
        RIfc5ce28_6079,RIfec31b0_8340,RIe1b4b18_3433,RIf149708_5295,RIf148358_5281,RIe1b3768_3419,RIfec3480_8342,RIfc483b0_5844,RIfc80be8_6487,RIe1ad4f8_3349,
        RIfec3318_8341,RIe1aa3c0_3314,RIe1a76c0_3282,RIe1a49c0_3250,RIe1a1cc0_3218,RIe18e1c0_2994,RIe17a6c0_2770,RIe228018_4745,RIe21cc18_4617,RIe206418_4361,
        RIe200478_4293,RIe1f9830_4216,RIe1f2378_4133,RIe1d6880_3818,RIe1bd380_3530,RIe1b01f8_3381,RIe172830_2680,RIdec6bc0_725,RIdec3ec0_693,RIee20a58_4830,
        RIdec11c0_661,RIee1f978_4818,RIdebe4c0_629,RIdebb7c0_597,RIdeb8ac0_565,RIee1efa0_4811,RIdeb30c0_501,RIfcb04b0_7028,RIdeb03c0_469,RIfc5e4a8_6095,
        RIdead6c0_437,RIdea72e8_405,RIdea09e8_373,RIfcb2508_7051,RIfcd16d8_7405,RIfc5d800_6086,RIfc63d40_6158,RIde93b30_310,RIfea7820_8222,RIfea73e8_8219,
        RIde87998_251,RIde837f8_231,RIfc7bd28_6431,RIfcc7ef8_7297,RIfc7a108_6411,RIfc7a6a8_6415,RIe16ccc8_2615,RIe16a838_2589,RIe1691b8_2573,RIe166bc0_2546,
        RIe163ec0_2514,RIee38338_5098,RIe1611c0_2482,RIfc54b60_5986,RIe15e4c0_2450,RIe158ac0_2386,RIe155dc0_2354,RIee35a70_5069,RIe1530c0_2322,RIee357a0_5067,
        RIe1503c0_2290,RIfc9fdb8_6841,RIe14d6c0_2258,RIe14a9c0_2226,RIe147cc0_2194,RIee34af8_5058,RIee33a18_5046,RIee327d0_5033,RIfcbcf30_7172,RIe142428_2131,
        RIe140100_2106,RIfea7280_8218,RIdf3bb78_2056,RIfc731f0_6332,RIee30610_5009,RIfcbe010_7184,RIee2e450_4985,RIfec2ee0_8338,RIfec3048_8339,RIfec2c10_8336,
        RIfec2d78_8337,RIfcb46c8_7075,RIfcb4830_7076,RIee29860_4931,RIfcb88e0_7122,RIdf2b480_1869,RIdf29590_1847,RIdf27268_1822,RIdf25648_1802,RIfcc9de8_7319,
        RIfc53648_5971,RIdf23a28_1782,RIfc823d0_6504,RIdf223a8_1766,RIdf20d28_1750,RIdf1bd00_1693,RIdf1a7e8_1678,RIdf18790_1655,RIdf15a90_1623,RIdf12d90_1591,
        RIdf10090_1559,RIdf0d390_1527,RIdf0a690_1495,RIdf07990_1463,RIdf04c90_1431,RIdeff290_1367,RIdefc590_1335,RIdef9890_1303,RIdef6b90_1271,RIdef3e90_1239,
        RIdef1190_1207,RIdeee490_1175,RIdeeb790_1143,RIee25be8_4888,RIfc6af28_6239,RIee23fc8_4868,RIfccf680_7382,RIdee5d90_1079,RIdee4008_1058,RIdee1ce0_1033,
        RIdedfdf0_1011,RIfc6b090_6240,RIfc534e0_5970,RIfca5920_6906,RIfc66770_6188,RIfe8f6d0_7976,RIded87d0_927,RIfe8f568_7975,RIded42e8_878,RIded1fc0_853,
        RIdecf2c0_821,RIdecc5c0_789,RIdec98c0_757,RIdeb5dc0_533,RIde9a0e8_341,RIe16f9c8_2647,RIe15b7c0_2418,RIe144fc0_2162,RIdf399b8_2032,RIdf2e018_1900,
        RIdf1e898_1724,RIdf01f90_1399,RIdee8a90_1111,RIdedd7f8_984,RIde80030_214,RIe19ee58_3185,RIe19c158_3153,RIf145bf8_5253,RIe199458_3121,RIfe8f298_7973,
        RIe196758_3089,RIe193a58_3057,RIe190d58_3025,RIe18b358_2961,RIe188658_2929,RIfe8f130_7972,RIe185958_2897,RIfc9f278_6833,RIe182c58_2865,RIe17ff58_2833,
        RIe17d258_2801,RIf1427f0_5216,RIfe8efc8_7971,RIe1779c0_2738,RIe1768e0_2726,RIfc81e30_6500,RIfc9ff20_6842,RIfca0088_6843,RIfc81b60_6498,RIfce5778_7633,
        RIfce08b8_7577,RIfc815c0_6494,RIe174cc0_2706,RIfca04c0_6846,RIfc53eb8_5977,RIfcc65a8_7279,RIfc80d50_6488,RIfc804e0_6482,RIe2251b0_4712,RIfc80378_6481,
        RIe2224b0_4680,RIfcb5910_7088,RIe21f7b0_4648,RIe219db0_4584,RIe2170b0_4552,RIfca01f0_6844,RIe2143b0_4520,RIfc82c40_6510,RIe2116b0_4488,RIfc7f6d0_6472,
        RIe20e9b0_4456,RIe20bcb0_4424,RIe208fb0_4392,RIf167528_5635,RIf1665b0_5624,RIe203718_4329,RIe201c60_4310,RIfc9da90_6816,RIfcc5360_7266,RIf163748_5591,
        RIf162668_5579,RIfc7e320_6458,RIfc87998_6565,RIe1fd610_4260,RIe1fc3c8_4247,RIf15d370_5520,RIf15c128_5507,RIfcc5d38_7273,RIfce7d70_7660,RIfc4bd58_5885,
        RIfc55c40_5998,RIfca2ab8_6873,RIe1fb450_4236,RIf156890_5444,RIfcd5ff8_7457,RIf154dd8_5425,RIfec2aa8_8335,RIfcb4b00_7078,RIfcd9400_7494,RIf151160_5382,
        RIe1f4808_4159,RIfc44738_5801,RIfc90908_6667,RIf14e5c8_5351,RIe1ef510_4100,RIe1ecf18_4073,RIe1ea218_4041,RIe1e7518_4009,RIe1e4818_3977,RIe1e1b18_3945,
        RIe1dee18_3913,RIe1dc118_3881,RIe1d9418_3849,RIe1d3a18_3785,RIe1d0d18_3753,RIe1ce018_3721,RIe1cb318_3689,RIe1c8618_3657,RIe1c5918_3625,RIe1c2c18_3593,
        RIe1bff18_3561,RIf14d218_5337,RIfe8ee60_7970,RIfea8090_8228,RIe1b84c0_3474,RIf14aab8_5309,RIfc6c170_6252,RIe1b6468_3451,RIe1b49b0_3432,RIfcafad8_7021,
        RIfcaa948_6963,RIfe8ecf8_7969,RIfe8f400_7974,RIfc67f58_6205,RIfca8ff8_6945,RIfe8eb90_7968,RIe1abe78_3333,RIe1aa258_3313,RIe1a7558_3281,RIe1a4858_3249,
        RIe1a1b58_3217,RIe18e058_2993,RIe17a558_2769,RIe227eb0_4744,RIe21cab0_4616,RIe2062b0_4360,RIe200310_4292,RIe1f96c8_4215,RIe1f2210_4132,RIe1d6718_3817,
        RIe1bd218_3529,RIe1b0090_3380,RIe1726c8_2679,RIdec4460_697,RIdec1760_665,RIee1fae0_4819,RIdebea60_633,RIee1f108_4812,RIdebbd60_601,RIdeb9060_569,
        RIdeb6360_537,RIee1eb68_4808,RIdeb0960_473,RIee1e460_4803,RIdeadc60_441,RIee1d7b8_4794,RIdea8008_409,RIdea1708_377,RIde9ae08_345,RIfe957d8_8045,
        RIfe95508_8043,RIfe95670_8044,RIee1a7e8_4760,RIfe95aa8_8047,RIfe95238_8041,RIfe95940_8046,RIfe953a0_8042,RIee1a0e0_4755,RIee19ca8_4752,RIee19870_4749,
        RIee19438_4746,RIee38ba8_5104,RIfe95c10_8048,RIee384a0_5099,RIfea9440_8242,RIe164460_2518,RIe161760_2486,RIfe942c0_8030,RIe15ea60_2454,RIfe94158_8029,
        RIe15bd60_2422,RIe156360_2358,RIe153660_2326,RIfe94428_8031,RIe150960_2294,RIfe94590_8032,RIe14dc60_2262,RIfc5c2e8_6071,RIe14af60_2230,RIe148260_2198,
        RIe145560_2166,RIee33ce8_5048,RIee32aa0_5035,RIee31858_5022,RIfc5d530_6084,RIe140538_2109,RIdf3e2d8_2084,RIdf3c118_2060,RIdf39df0_2035,RIfcdd780_7542,
        RIee2ee28_4992,RIfcc88d0_7304,RIee2cc68_4968,RIdf34990_1975,RIdf32aa0_1953,RIdf304a8_1926,RIdf2e5b8_1904,RIee2b1b0_4949,RIfe946f8_8033,RIfcb2940_7054,
        RIee273d0_4905,RIfe949c8_8035,RIdf27538_1824,RIfe94b30_8036,RIfe94860_8034,RIee26f98_4902,RIee269f8_4898,RIee26728_4896,RIee26458_4894,RIee26188_4892,
        RIfe94c98_8037,RIee25d50_4889,RIfea9170_8240,RIdf16030_1627,RIdf13330_1595,RIdf10630_1563,RIdf0d930_1531,RIdf0ac30_1499,RIdf07f30_1467,RIdf05230_1435,
        RIdf02530_1403,RIdefcb30_1339,RIdef9e30_1307,RIdef7130_1275,RIdef4430_1243,RIdef1730_1211,RIdeeea30_1179,RIdeebd30_1147,RIdee9030_1115,RIee250a8_4880,
        RIee24298_4870,RIee23758_4862,RIee22d80_4855,RIfe950d0_8040,RIfe94f68_8039,RIfe94e00_8038,RIdeddd98_988,RIee22ab0_4853,RIee21e08_4844,RIfca46d8_6893,
        RIfc5dad0_6088,RIfeaa250_8252,RIfe96048_8051,RIfe95d78_8049,RIfe95ee0_8050,RIdecf860_825,RIdeccb60_793,RIdec9e60_761,RIdec7160_729,RIdeb3660_505,
        RIde94508_313,RIe16d268_2619,RIe159060_2390,RIe142860_2134,RIdf37258_2004,RIdf2b8b8_1872,RIdf1c138_1696,RIdeff830_1371,RIdee6330_1083,RIdedb098_956,
        RIde7a450_186,RIe19c6f8_3157,RIe1999f8_3125,RIf1450b8_5245,RIe196cf8_3093,RIf143fd8_5233,RIe193ff8_3061,RIe1912f8_3029,RIe18e5f8_2997,RIe188bf8_2933,
        RIe185ef8_2901,RIfe973f8_8065,RIe1831f8_2869,RIf142958_5217,RIe1804f8_2837,RIe17d7f8_2805,RIe17aaf8_2773,RIf141b48_5207,RIfc542f0_5980,RIfc800a8_6479,
        RIe175260_2710,RIfca0bc8_6851,RIfc48680_5846,RIee3dea0_5163,RIfcc6878_7281,RIee3ba10_5137,RIee3a930_5125,RIfe97290_8064,RIe172b00_2682,RIf16f958_5729,
        RIf16ee18_5721,RIf16da68_5707,RIf16d360_5702,RIfe96e58_8061,RIe222a50_4684,RIfe96cf0_8060,RIe21fd50_4652,RIf16a660_5670,RIe21d050_4620,RIe217650_4556,
        RIe214950_4524,RIf169f58_5665,RIe211c50_4492,RIf168770_5648,RIe20ef50_4460,RIf1677f8_5637,RIe20c250_4428,RIe209550_4396,RIe206850_4364,RIf166880_5626,
        RIf1657a0_5614,RIe201dc8_4311,RIe2005e0_4294,RIfe96b88_8059,RIf163b80_5594,RIf162c08_5583,RIf161420_5566,RIf15f530_5544,RIf15d7a8_5523,RIfe968b8_8057,
        RIfe96a20_8058,RIfcb3fc0_7070,RIfc7cf70_6444,RIfc579c8_6019,RIf159590_5476,RIf1584b0_5464,RIf157268_5451,RIf1569f8_5445,RIfe965e8_8055,RIf155d50_5436,
        RIf155210_5428,RIf153e60_5414,RIfe96750_8056,RIf1527e0_5398,RIf151430_5384,RIfcd2650_7416,RIe1f2648_4135,RIf14f108_5359,RIfc7f298_6469,RIf14d4e8_5339,
        RIe1ed350_4076,RIe1ea7b8_4045,RIe1e7ab8_4013,RIe1e4db8_3981,RIe1e20b8_3949,RIe1df3b8_3917,RIe1dc6b8_3885,RIe1d99b8_3853,RIe1d6cb8_3821,RIe1d12b8_3757,
        RIe1ce5b8_3725,RIe1cb8b8_3693,RIe1c8bb8_3661,RIe1c5eb8_3629,RIe1c31b8_3597,RIe1c04b8_3565,RIe1bd7b8_3533,RIf14c138_5325,RIf14ad88_5311,RIe1b8790_3476,
        RIfe96480_8054,RIf14a0e0_5302,RIf149870_5296,RIfe97128_8063,RIfe96318_8053,RIf148628_5283,RIfc58d78_6033,RIe1b20e8_3403,RIe1b04c8_3383,RIf146cd8_5265,
        RIfc591b0_6036,RIfe961b0_8052,RIfe96fc0_8062,RIe1a7af8_3285,RIe1a4df8_3253,RIe1a20f8_3221,RIe19f3f8_3189,RIe18b8f8_2965,RIe177df8_2741,RIe225750_4716,
        RIe21a350_4588,RIe203b50_4332,RIe1fdbb0_4264,RIe1f6f68_4187,RIe1efab0_4104,RIe1d3fb8_3789,RIe1baab8_3501,RIe1ad930_3352,RIe16ff68_2651,RIdec42f8_696,
        RIdec15f8_664,RIfcc6cb0_7284,RIdebe8f8_632,RIfe93780_8022,RIdebbbf8_600,RIdeb8ef8_568,RIdeb61f8_536,RIee1ea00_4807,RIdeb07f8_472,RIee1e2f8_4802,
        RIdeadaf8_440,RIfc5d3c8_6083,RIdea7cc0_408,RIdea13c0_376,RIde9aac0_344,RIfc58238_6025,RIfcc3b78_7249,RIfc7d0d8_6445,RIfc59750_6040,RIfe93a50_8024,
        RIfe938e8_8023,RIde88370_254,RIde83e88_233,RIfc5f420_6106,RIfc976b8_6745,RIfc90a70_6668,RIfc60500_6118,RIee38a40_5103,RIe16ab08_2591,RIe169488_2575,
        RIe166ff8_2549,RIe1642f8_2517,RIe1615f8_2485,RIee369e8_5080,RIe15e8f8_2453,RIee35bd8_5070,RIe15bbf8_2421,RIe1561f8_2357,RIe1534f8_2325,RIfc3ee28_5741,
        RIe1507f8_2293,RIfce6c90_7648,RIe14daf8_2261,RIfcca7c0_7326,RIe14adf8_2229,RIe1480f8_2197,RIe1453f8_2165,RIee33b80_5047,RIee32938_5034,RIee316f0_5021,
        RIee30bb0_5013,RIe1403d0_2108,RIfe93618_8021,RIdf3bfb0_2059,RIfe934b0_8020,RIfcd0d00_7398,RIee2ecc0_4991,RIee2e720_4987,RIee2cb00_4967,RIfe93bb8_8025,
        RIdf32938_1952,RIdf30340_1925,RIdf2e450_1903,RIee2b048_4948,RIee29b30_4933,RIfc67148_6195,RIfc6fb18_6293,RIdf29860_1849,RIfe931e0_8018,RIfe93348_8019,
        RIfe93078_8017,RIfc672b0_6196,RIfca8788_6939,RIdf22510_1767,RIfcea7a0_7690,RIdf20ff8_1752,RIdf1ecd0_1727,RIdf1aab8_1680,RIfea7c58_8225,RIdf15ec8_1626,
        RIdf131c8_1594,RIdf104c8_1562,RIdf0d7c8_1530,RIdf0aac8_1498,RIdf07dc8_1466,RIdf050c8_1434,RIdf023c8_1402,RIdefc9c8_1338,RIdef9cc8_1306,RIdef6fc8_1274,
        RIdef42c8_1242,RIdef15c8_1210,RIdeee8c8_1178,RIdeebbc8_1146,RIdee8ec8_1114,RIee24f40_4879,RIee24130_4869,RIee235f0_4861,RIee22c18_4854,RIfe93d20_8026,
        RIdee1fb0_1035,RIdee0228_1014,RIdeddc30_987,RIfc684f8_6209,RIee21ca0_4843,RIfc68390_6208,RIee20d28_4832,RIded8aa0_929,RIfe93ff0_8028,RIded45b8_880,
        RIfe93e88_8027,RIdecf6f8_824,RIdecc9f8_792,RIdec9cf8_760,RIdec6ff8_728,RIdeb34f8_504,RIde941c0_312,RIe16d100_2618,RIe158ef8_2389,RIe1426f8_2133,
        RIdf370f0_2003,RIdf2b750_1871,RIdf1bfd0_1695,RIdeff6c8_1370,RIdee61c8_1082,RIdedaf30_955,RIde7a108_185,RIe19c590_3156,RIe199890_3124,RIf144f50_5244,
        RIe196b90_3092,RIfc76058_6365,RIe193e90_3060,RIe191190_3028,RIe18e490_2996,RIe188a90_2932,RIe185d90_2900,RIfccd8f8_7361,RIe183090_2868,RIfc76e68_6375,
        RIe180390_2836,RIe17d690_2804,RIe17a990_2772,RIf1419e0_5206,RIf140630_5192,RIe176bb0_2728,RIe1750f8_2709,RIfcd1840_7406,RIfc5f6f0_6108,RIee3dd38_5162,
        RIee3cc58_5150,RIee3b8a8_5136,RIee3a7c8_5124,RIee39580_5111,RIfea9008_8239,RIf16f7f0_5728,RIf16ecb0_5720,RIf16d900_5706,RIfc78ec0_6398,RIfcc8060_7298,
        RIe2228e8_4683,RIfc5a3f8_6049,RIe21fbe8_4651,RIfc74000_6342,RIe21cee8_4619,RIe2174e8_4555,RIe2147e8_4523,RIfca2c20_6874,RIe211ae8_4491,RIfca2950_6872,
        RIe20ede8_4459,RIfcc24f8_7233,RIe20c0e8_4427,RIe2093e8_4395,RIe2066e8_4363,RIfc45110_5808,RIfcc6f80_7286,RIfe92f10_8016,RIfe92970_8012,RIf164af8_5605,
        RIf163a18_5593,RIf162aa0_5582,RIfe92ad8_8013,RIf15f3c8_5543,RIf15d640_5522,RIfe92808_8011,RIfe92c40_8014,RIfe926a0_8010,RIfe92da8_8015,RIfe92538_8009,
        RIfcb5a78_7089,RIf158348_5463,RIf157100_5450,RIfc53be8_5975,RIfec38b8_8345,RIfcc5ea0_7274,RIf1550a8_5427,RIf153cf8_5413,RIfec3a20_8346,RIf152678_5397,
        RIfec3750_8344,RIf14ff18_5369,RIfe923d0_8008,RIf14efa0_5358,RIf14e898_5353,RIf14d380_5338,RIfe92268_8007,RIe1ea650_4044,RIe1e7950_4012,RIe1e4c50_3980,
        RIe1e1f50_3948,RIe1df250_3916,RIe1dc550_3884,RIe1d9850_3852,RIe1d6b50_3820,RIe1d1150_3756,RIe1ce450_3724,RIe1cb750_3692,RIe1c8a50_3660,RIe1c5d50_3628,
        RIe1c3050_3596,RIe1c0350_3564,RIe1bd650_3532,RIfcda4e0_7506,RIfc9d220_6810,RIe1b8628_3475,RIe1b6738_3453,RIfc4f2c8_5923,RIfce16c8_7587,RIfe91cc8_8003,
        RIfe91e30_8004,RIf1484c0_5282,RIf147548_5271,RIfe91f98_8005,RIfe91b60_8002,RIf146b70_5264,RIfc9f548_6835,RIfe92100_8006,RIfe919f8_8001,RIe1a7990_3284,
        RIe1a4c90_3252,RIe1a1f90_3220,RIe19f290_3188,RIe18b790_2964,RIe177c90_2740,RIe2255e8_4715,RIe21a1e8_4587,RIe2039e8_4331,RIe1fda48_4263,RIe1f6e00_4186,
        RIe1ef948_4103,RIe1d3e50_3788,RIe1ba950_3500,RIe1ad7c8_3351,RIe16fe00_2650,RIdec4730_699,RIdec1a30_667,RIfce3f90_7616,RIdebed30_635,RIfcc3308_7243,
        RIdebc030_603,RIdeb9330_571,RIdeb6630_539,RIfc8c588_6619,RIdeb0c30_475,RIfc5a998_6053,RIdeadf30_443,RIfc99b48_6771,RIdea8698_411,RIdea1d98_379,
        RIde9b498_347,RIfc78bf0_6396,RIfcbc558_7165,RIfca12d0_6856,RIfca3fd0_6888,RIfec2670_8332,RIfec2508_8331,RIde88a00_256,RIde84518_235,RIfcc35d8_7245,
        RIfcb57a8_7087,RIfc5a290_6048,RIfca3058_6877,RIee38e78_5106,RIfec27d8_8333,RIfca3328_6879,RIe1672c8_2551,RIe164730_2520,RIe161a30_2488,RIee36cb8_5082,
        RIe15ed30_2456,RIfcc7250_7288,RIe15c030_2424,RIe156630_2360,RIe153930_2328,RIfcc7688_7291,RIe150c30_2296,RIfc8af08_6603,RIe14df30_2264,RIfc9a250_6776,
        RIe14b230_2232,RIe148530_2200,RIe145830_2168,RIfc9aac0_6782,RIfc56bb8_6009,RIfca1ca8_6863,RIfcec960_7714,RIe1406a0_2110,RIdf3e440_2085,RIdf3c280_2061,
        RIdf39f58_2036,RIfc9a958_6781,RIee2f0f8_4994,RIfcdb458_7517,RIee2cf38_4970,RIdf34c60_1977,RIfec2940_8334,RIdf30778_1928,RIdf2e888_1906,RIee2b480_4951,
        RIfec23a0_8330,RIee288e8_4920,RIfec2238_8329,RIdf29b30_1851,RIdf27808_1826,RIdf25a80_1805,RIdf23e60_1785,RIfc55100_5990,RIfcd9f40_7502,RIfc54f98_5989,
        RIfc54cc8_5987,RIfc4b218_5877,RIdf1efa0_1729,RIfcc69e0_7282,RIdf18bc8_1658,RIdf16300_1629,RIdf13600_1597,RIdf10900_1565,RIdf0dc00_1533,RIdf0af00_1501,
        RIdf08200_1469,RIdf05500_1437,RIdf02800_1405,RIdefce00_1341,RIdefa100_1309,RIdef7400_1277,RIdef4700_1245,RIdef1a00_1213,RIdeeed00_1181,RIdeec000_1149,
        RIdee9300_1117,RIfce4ad0_7624,RIfc9e8a0_6826,RIfcc46b8_7257,RIfcd4108_7435,RIdee4440_1061,RIdee2280_1037,RIdee0390_1015,RIdede068_990,RIfcda0a8_7503,
        RIfce54a8_7631,RIfca0790_6848,RIfc50ee8_5943,RIded8d70_931,RIded68e0_905,RIded4888_882,RIded2560_857,RIdecfb30_827,RIdecce30_795,RIdeca130_763,
        RIdec7430_731,RIdeb3930_507,RIde94b98_315,RIe16d538_2621,RIe159330_2392,RIe142b30_2136,RIdf37528_2006,RIdf2bb88_1874,RIdf1c408_1698,RIdeffb00_1373,
        RIdee6600_1085,RIdedb368_958,RIde7aae0_188,RIe19c9c8_3159,RIe199cc8_3127,RIfe8ea28_7967,RIe196fc8_3095,RIfec20d0_8328,RIe1942c8_3063,RIe1915c8_3031,
        RIe18e8c8_2999,RIe188ec8_2935,RIe1861c8_2903,RIfc68228_6207,RIe1834c8_2871,RIfccb5d0_7336,RIe1807c8_2839,RIe17dac8_2807,RIe17adc8_2775,RIf141e18_5209,
        RIf140900_5194,RIf140090_5188,RIe1753c8_2711,RIf13f988_5183,RIf13ece0_5174,RIee3e170_5165,RIee3cf28_5152,RIee3bce0_5139,RIee3ac00_5127,RIee39850_5113,
        RIe172dd0_2684,RIf16fc28_5731,RIf16f0e8_5723,RIf16dd38_5709,RIfce9120_7674,RIfc404a8_5757,RIe222d20_4686,RIf16b8a8_5683,RIe220020_4654,RIf16a930_5672,
        RIe21d320_4622,RIe217920_4558,RIe214c20_4526,RIfc5b910_6064,RIe211f20_4494,RIfe8e8c0_7966,RIe20f220_4462,RIfe8e758_7965,RIe20c520_4430,RIe209820_4398,
        RIe206b20_4366,RIf166b50_5628,RIf165a70_5616,RIfe8dd80_7958,RIfe8dab0_7956,RIf164c60_5606,RIf163e50_5596,RIf162ed8_5585,RIf1616f0_5568,RIf15f800_5546,
        RIf15da78_5525,RIfe8d948_7955,RIfe8dc18_7957,RIf15c560_5510,RIf15b048_5495,RIfc62828_6143,RIf159860_5478,RIf158780_5466,RIf157538_5453,RIfca6e38_6921,
        RIe1f9b00_4218,RIfc61e50_6136,RIfc61748_6131,RIf154130_5416,RIe1f4ad8_4161,RIf152ab0_5400,RIf151700_5386,RIf1501e8_5371,RIe1f27b0_4136,RIfc60ed8_6125,
        RIfc7b620_6426,RIf14d7b8_5341,RIe1ed4b8_4077,RIe1eaa88_4047,RIe1e7d88_4015,RIe1e5088_3983,RIe1e2388_3951,RIe1df688_3919,RIe1dc988_3887,RIe1d9c88_3855,
        RIe1d6f88_3823,RIe1d1588_3759,RIe1ce888_3727,RIe1cbb88_3695,RIe1c8e88_3663,RIe1c6188_3631,RIe1c3488_3599,RIe1c0788_3567,RIe1bda88_3535,RIfca4de0_6898,
        RIfc5ea48_6099,RIe1b8a60_3478,RIe1b6a08_3455,RIfcbd638_7177,RIfc44fa8_5807,RIfe8e5f0_7964,RIfe8e1b8_7961,RIf1488f8_5285,RIf147818_5273,RIfe8e050_7960,
        RIfe8e488_7963,RIf146e40_5266,RIf146030_5256,RIfe8dee8_7959,RIfe8e320_7962,RIe1a7dc8_3287,RIe1a50c8_3255,RIe1a23c8_3223,RIe19f6c8_3191,RIe18bbc8_2967,
        RIe1780c8_2743,RIe225a20_4718,RIe21a620_4590,RIe203e20_4334,RIe1fde80_4266,RIe1f7238_4189,RIe1efd80_4106,RIe1d4288_3791,RIe1bad88_3503,RIe1adc00_3354,
        RIe170238_2653,RIdec45c8_698,RIdec18c8_666,RIfce85e0_7666,RIdebebc8_634,RIfcb8bb0_7124,RIdebbec8_602,RIdeb91c8_570,RIdeb64c8_538,RIfc85d78_6545,
        RIdeb0ac8_474,RIfc85aa8_6543,RIdeaddc8_442,RIfc4d3d8_5901,RIdea8350_410,RIdea1a50_378,RIde9b150_346,RIfc85ee0_6546,RIfc9c9b0_6804,RIfce13f8_7585,
        RIfcb8778_7121,RIfe8d510_7952,RIfe8d3a8_7951,RIde886b8_255,RIde841d0_234,RIde806c0_216,RIfcb8070_7116,RIfce1128_7583,RIfc9c140_6798,RIee38d10_5105,
        RIe16ac70_2592,RIfc850d0_6536,RIe167160_2550,RIe1645c8_2519,RIe1618c8_2487,RIee36b50_5081,RIe15ebc8_2455,RIee35d40_5071,RIe15bec8_2423,RIe1564c8_2359,
        RIe1537c8_2327,RIfc3ef90_5742,RIe150ac8_2295,RIfe8d7e0_7954,RIe14ddc8_2263,RIfce0fc0_7582,RIe14b0c8_2231,RIe1483c8_2199,RIe1456c8_2167,RIee33e50_5049,
        RIee32c08_5036,RIee319c0_5023,RIee30d18_5014,RIfe8cf70_7948,RIfe8ce08_7947,RIfe8d240_7950,RIfe8d0d8_7949,RIfce9dc8_7683,RIee2ef90_4993,RIfce51d8_7629,
        RIee2cdd0_4969,RIdf34af8_1976,RIfe8d678_7953,RIdf30610_1927,RIdf2e720_1905,RIee2b318_4950,RIee29c98_4934,RIee28780_4919,RIee27538_4906,RIdf299c8_1850,
        RIdf276a0_1825,RIdf25918_1804,RIdf23cf8_1784,RIfc83ff0_6524,RIfcb73c8_7107,RIfc51320_5946,RIfcdaa80_7510,RIfc83d20_6522,RIdf1ee38_1728,RIfc51b90_5952,
        RIdf18a60_1657,RIdf16198_1628,RIdf13498_1596,RIdf10798_1564,RIdf0da98_1532,RIdf0ad98_1500,RIdf08098_1468,RIdf05398_1436,RIdf02698_1404,RIdefcc98_1340,
        RIdef9f98_1308,RIdef7298_1276,RIdef4598_1244,RIdef1898_1212,RIdeeeb98_1180,RIdeebe98_1148,RIdee9198_1116,RIee25210_4881,RIee24400_4871,RIee238c0_4863,
        RIee22ee8_4856,RIfe8cca0_7946,RIdee2118_1036,RIfe8cb38_7945,RIdeddf00_989,RIfcc5a68_7271,RIee21f70_4845,RIfcb6cc0_7102,RIee20e90_4833,RIded8c08_930,
        RIded6778_904,RIded4720_881,RIded23f8_856,RIdecf9c8_826,RIdecccc8_794,RIdec9fc8_762,RIdec72c8_730,RIdeb37c8_506,RIde94850_314,RIe16d3d0_2620,
        RIe1591c8_2391,RIe1429c8_2135,RIdf373c0_2005,RIdf2ba20_1873,RIdf1c2a0_1697,RIdeff998_1372,RIdee6498_1084,RIdedb200_957,RIde7a798_187,RIe19c860_3158,
        RIe199b60_3126,RIf145220_5246,RIe196e60_3094,RIf144140_5234,RIe194160_3062,RIe191460_3030,RIe18e760_2998,RIe188d60_2934,RIe186060_2902,RIf1431c8_5223,
        RIe183360_2870,RIf142ac0_5218,RIe180660_2838,RIe17d960_2806,RIe17ac60_2774,RIf141cb0_5208,RIf140798_5193,RIf13ff28_5187,RIfe8be90_7936,RIfceb880_7702,
        RIf13eb78_5173,RIee3e008_5164,RIee3cdc0_5151,RIee3bb78_5138,RIee3aa98_5126,RIee396e8_5112,RIe172c68_2683,RIf16fac0_5730,RIf16ef80_5722,RIf16dbd0_5708,
        RIfcc4af0_7260,RIf16c820_5694,RIe222bb8_4685,RIf16b740_5682,RIe21feb8_4653,RIf16a7c8_5671,RIe21d1b8_4621,RIe2177b8_4557,RIe214ab8_4525,RIfe8c430_7940,
        RIe211db8_4493,RIf1688d8_5649,RIe20f0b8_4461,RIf167960_5638,RIe20c3b8_4429,RIe2096b8_4397,RIe2069b8_4365,RIf1669e8_5627,RIf165908_5615,RIfe8c9d0_7944,
        RIfe8c700_7942,RIfc9c578_6801,RIf163ce8_5595,RIf162d70_5584,RIf161588_5567,RIf15f698_5545,RIf15d910_5524,RIfe8c598_7941,RIfe8c868_7943,RIf15c3f8_5509,
        RIf15aee0_5494,RIf15a0d0_5484,RIf1596f8_5477,RIf158618_5465,RIf1573d0_5452,RIf156b60_5446,RIfec1f68_8327,RIf155eb8_5437,RIf155378_5429,RIf153fc8_5415,
        RIfe8bff8_7937,RIf152948_5399,RIf151598_5385,RIf150080_5370,RIfe8c2c8_7939,RIf14f270_5360,RIfc503a8_5935,RIf14d650_5340,RIfe8c160_7938,RIe1ea920_4046,
        RIe1e7c20_4014,RIe1e4f20_3982,RIe1e2220_3950,RIe1df520_3918,RIe1dc820_3886,RIe1d9b20_3854,RIe1d6e20_3822,RIe1d1420_3758,RIe1ce720_3726,RIe1cba20_3694,
        RIe1c8d20_3662,RIe1c6020_3630,RIe1c3320_3598,RIe1c0620_3566,RIe1bd920_3534,RIf14c2a0_5326,RIf14aef0_5312,RIe1b88f8_3477,RIe1b68a0_3454,RIfcd4db0_7444,
        RIfc4ebc0_5918,RIfec1e00_8326,RIfe8bd28_7935,RIf148790_5284,RIf1476b0_5272,RIfe8ba58_7933,RIfec1b30_8324,RIfc4e788_5915,RIfcb8e80_7126,RIfe8bbc0_7934,
        RIfec1c98_8325,RIe1a7c60_3286,RIe1a4f60_3254,RIe1a2260_3222,RIe19f560_3190,RIe18ba60_2966,RIe177f60_2742,RIe2258b8_4717,RIe21a4b8_4589,RIe203cb8_4333,
        RIe1fdd18_4265,RIe1f70d0_4188,RIe1efc18_4105,RIe1d4120_3790,RIe1bac20_3502,RIe1ada98_3353,RIe1700d0_2652,RIdec4a00_701,RIdec1d00_669,RIfcad7b0_6996,
        RIdebf000_637,RIfc64cb8_6169,RIdebc300_605,RIdeb9600_573,RIdeb6900_541,RIfc6f9b0_6292,RIdeb0f00_477,RIfc657f8_6177,RIdeae200_445,RIfce69c0_7646,
        RIdea8d28_413,RIdea2428_381,RIde9bb28_349,RIfc6fc80_6294,RIee1b760_4771,RIfca8080_6934,RIfe8b8f0_7932,RIde90020_292,RIde8c510_274,RIde89090_258,
        RIde84ba8_237,RIfc65ac8_6179,RIfcad210_6992,RIfcce168_7367,RIfcce2d0_7368,RIfc51488_5947,RIe16af40_2594,RIfc65c30_6180,RIe167598_2553,RIe164a00_2522,
        RIe161d00_2490,RIfc66e78_6193,RIe15f000_2458,RIfc6e498_6277,RIe15c300_2426,RIe156900_2362,RIe153c00_2330,RIfc6e330_6276,RIe150f00_2298,RIfccda60_7362,
        RIe14e200_2266,RIfc6e1c8_6275,RIe14b500_2234,RIe148800_2202,RIe145b00_2170,RIee33fb8_5050,RIee32d70_5037,RIee31c90_5025,RIee30fe8_5016,RIfea8630_8232,
        RIdf3e5a8_2086,RIdf3c550_2063,RIfea8798_8233,RIfc6e060_6274,RIfcac6d0_6984,RIfc56078_6001,RIfc6e600_6278,RIdf34dc8_1978,RIdf32d70_1955,RIfea84c8_8231,
        RIdf2eb58_1908,RIee2b750_4953,RIfc6ee70_6284,RIfc6efd8_6285,RIee27808_4908,RIfe8b788_7931,RIdf27ad8_1828,RIdf25d50_1807,RIdf24130_1787,RIfc66608_6187,
        RIfccde98_7365,RIfc66a40_6190,RIfc668d8_6189,RIfcacf40_6990,RIfeaaef8_8261,RIfc6e8d0_6280,RIdf18d30_1659,RIdf165d0_1631,RIdf138d0_1599,RIdf10bd0_1567,
        RIdf0ded0_1535,RIdf0b1d0_1503,RIdf084d0_1471,RIdf057d0_1439,RIdf02ad0_1407,RIdefd0d0_1343,RIdefa3d0_1311,RIdef76d0_1279,RIdef49d0_1247,RIdef1cd0_1215,
        RIdeeefd0_1183,RIdeec2d0_1151,RIdee95d0_1119,RIfc6dc28_6271,RIfc67c88_6203,RIfccb300_7334,RIfccd4c0_7358,RIfea81f8_8229,RIfea8360_8230,RIdee04f8_1016,
        RIdede338_992,RIfc6def8_6273,RIfcac130_6980,RIfc67b20_6202,RIfc67df0_6204,RIded9040_933,RIded6a48_906,RIded4b58_884,RIded26c8_858,RIdecfe00_829,
        RIdecd100_797,RIdeca400_765,RIdec7700_733,RIdeb3c00_509,RIde95228_317,RIe16d808_2623,RIe159600_2394,RIe142e00_2138,RIdf377f8_2008,RIdf2be58_1876,
        RIdf1c6d8_1700,RIdeffdd0_1375,RIdee68d0_1087,RIdedb638_960,RIde7b170_190,RIe19cc98_3161,RIe199f98_3129,RIfc73088_6331,RIe197298_3097,RIf1442a8_5235,
        RIe194598_3065,RIe191898_3033,RIe18eb98_3001,RIe189198_2937,RIe186498_2905,RIfc72278_6321,RIe183798_2873,RIfc61ce8_6135,RIe180a98_2841,RIe17dd98_2809,
        RIe17b098_2777,RIfcaf268_7015,RIfca6a00_6918,RIfcc9b18_7317,RIe175530_2712,RIfc72818_6325,RIfc726b0_6324,RIfccf7e8_7383,RIfc72548_6323,RIee3be48_5140,
        RIee3ad68_5128,RIfc71fa8_6319,RIe1730a0_2686,RIfcaef98_7013,RIfccf518_7381,RIfc71e40_6318,RIfc62120_6138,RIfe8b350_7928,RIe222ff0_4688,RIfcc9f50_7320,
        RIe2202f0_4656,RIfc4a570_5868,RIe21d5f0_4624,RIe217bf0_4560,RIe214ef0_4528,RIfccf3b0_7380,RIe2121f0_4496,RIf168ba8_5651,RIe20f4f0_4464,RIfc71300_6310,
        RIe20c7f0_4432,RIe209af0_4400,RIe206df0_4368,RIfc718a0_6314,RIfc71a08_6315,RIe202098_4313,RIfe8b1e8_7927,RIfc715d0_6312,RIfce6588_7643,RIfc62c60_6146,
        RIf161858_5569,RIf15fad0_5548,RIf15dbe0_5526,RIe1fc698_4249,RIfe8b4b8_7929,RIfcae5c0_7006,RIfc63098_6149,RIfc63200_6150,RIfc71198_6309,RIf158a50_5468,
        RIf1576a0_5454,RIfcdc808_7531,RIfe8b620_7930,RIfc634d0_6152,RIfcceb40_7374,RIf154400_5418,RIe1f4da8_4163,RIf152c18_5401,RIf151868_5387,RIfc4d108_5899,
        RIe1f2a80_4138,RIfc70a90_6304,RIfc63bd8_6157,RIfca7810_6928,RIe1ed788_4079,RIe1ead58_4049,RIe1e8058_4017,RIe1e5358_3985,RIe1e2658_3953,RIe1df958_3921,
        RIe1dcc58_3889,RIe1d9f58_3857,RIe1d7258_3825,RIe1d1858_3761,RIe1ceb58_3729,RIe1cbe58_3697,RIe1c9158_3665,RIe1c6458_3633,RIe1c3758_3601,RIe1c0a58_3569,
        RIe1bdd58_3537,RIf14c408_5327,RIf14b1c0_5314,RIe1b8d30_3480,RIe1b6cd8_3457,RIfc707c0_6302,RIfca7c48_6931,RIe1b4de8_3435,RIe1b3a38_3421,RIfc70220_6298,
        RIfcce870_7372,RIe1b23b8_3405,RIe1b0630_3384,RIfc645b0_6164,RIfc700b8_6297,RIfeaac28_8259,RIe1aa690_3316,RIe1a8098_3289,RIe1a5398_3257,RIe1a2698_3225,
        RIe19f998_3193,RIe18be98_2969,RIe178398_2745,RIe225cf0_4720,RIe21a8f0_4592,RIe2040f0_4336,RIe1fe150_4268,RIe1f7508_4191,RIe1f0050_4108,RIe1d4558_3793,
        RIe1bb058_3505,RIe1aded0_3356,RIe170508_2655,RIdec4898_700,RIdec1b98_668,RIfc661d0_6184,RIdebee98_636,RIfce6b28_7647,RIdebc198_604,RIdeb9498_572,
        RIdeb6798_540,RIfc40d18_5763,RIdeb0d98_476,RIfcad648_6995,RIdeae098_444,RIfcaa510_6960,RIdea89e0_412,RIdea20e0_380,RIde9b7e0_348,RIfcab320_6970,
        RIfca8350_6936,RIfc6f6e0_6290,RIfcaa240_6958,RIde8fcd8_291,RIfe8aae0_7922,RIde88d48_257,RIde84860_236,RIde80a08_217,RIfc64718_6165,RIfcae020_7002,
        RIfcadeb8_7001,RIee38fe0_5107,RIe16add8_2593,RIe1695f0_2576,RIe167430_2552,RIe164898_2521,RIe161b98_2489,RIfe8a3d8_7917,RIe15ee98_2457,RIfe8a270_7916,
        RIe15c198_2425,RIe156798_2361,RIe153a98_2329,RIfc3f0f8_5743,RIe150d98_2297,RIfcab050_6968,RIe14e098_2265,RIfcca658_7325,RIe14b398_2233,RIe148698_2201,
        RIe145998_2169,RIfe8a810_7920,RIfe8a6a8_7919,RIee31b28_5024,RIee30e80_5015,RIe140808_2111,RIfe8a540_7918,RIdf3c3e8_2062,RIdf3a0c0_2037,RIfc6b1f8_6241,
        RIee2f260_4995,RIfc70d60_6306,RIee2d0a0_4971,RIfe8a978_7921,RIdf32c08_1954,RIdf308e0_1929,RIdf2e9f0_1907,RIee2b5e8_4952,RIee29e00_4935,RIee28a50_4921,
        RIee276a0_4907,RIdf29c98_1852,RIdf27970_1827,RIdf25be8_1806,RIdf23fc8_1786,RIfc6aaf0_6236,RIfc6ac58_6237,RIdf22678_1768,RIfcdd4b0_7540,RIdf21160_1753,
        RIdf1f108_1730,RIdf1ac20_1681,RIfeaa7f0_8256,RIdf16468_1630,RIdf13768_1598,RIdf10a68_1566,RIdf0dd68_1534,RIdf0b068_1502,RIdf08368_1470,RIdf05668_1438,
        RIdf02968_1406,RIdefcf68_1342,RIdefa268_1310,RIdef7568_1278,RIdef4868_1246,RIdef1b68_1214,RIdeeee68_1182,RIdeec168_1150,RIdee9468_1118,RIee25378_4882,
        RIee24568_4872,RIee23a28_4864,RIee23050_4857,RIfe8adb0_7924,RIdee23e8_1038,RIfe8ac48_7923,RIdede1d0_991,RIfca5650_6904,RIee220d8_4846,RIfceeb20_7738,
        RIee20ff8_4834,RIded8ed8_932,RIfe8af18_7925,RIded49f0_883,RIfe8b080_7926,RIdecfc98_828,RIdeccf98_796,RIdeca298_764,RIdec7598_732,RIdeb3a98_508,
        RIde94ee0_316,RIe16d6a0_2622,RIe159498_2393,RIe142c98_2137,RIdf37690_2007,RIdf2bcf0_1875,RIdf1c570_1699,RIdeffc68_1374,RIdee6768_1086,RIdedb4d0_959,
        RIde7ae28_189,RIe19cb30_3160,RIe199e30_3128,RIf145388_5247,RIe197130_3096,RIfe8a108_7915,RIe194430_3064,RIe191730_3032,RIe18ea30_3000,RIe189030_2936,
        RIe186330_2904,RIfc6c878_6257,RIe183630_2872,RIfcabcf8_6977,RIe180930_2840,RIe17dc30_2808,RIe17af30_2776,RIfcccc50_7352,RIfcccdb8_7353,RIe176d18_2729,
        RIfea7af0_8224,RIfe89fa0_7914,RIfe89e38_7913,RIfcdd078_7537,RIfccb738_7337,RIfca9868_6951,RIfcabb90_6976,RIfca99d0_6952,RIe172f38_2685,RIf16fd90_5732,
        RIf16f250_5724,RIfc6c440_6254,RIfcaba28_6975,RIfc40610_5758,RIe222e88_4687,RIfc5d260_6082,RIe220188_4655,RIfcab758_6973,RIe21d488_4623,RIe217a88_4559,
        RIe214d88_4527,RIfe892f8_7905,RIe212088_4495,RIf168a40_5650,RIe20f388_4463,RIf167ac8_5639,RIe20c688_4431,RIe209988_4399,RIe206c88_4367,RIfc6c2d8_6253,
        RIfceec88_7739,RIe201f30_4312,RIe200748_4295,RIf164dc8_5607,RIf163fb8_5597,RIf163040_5586,RIfe895c8_7907,RIf15f968_5547,RIfe89898_7909,RIfe89460_7906,
        RIe1fb5b8_4237,RIf15c6c8_5511,RIfe89730_7908,RIf15a238_5485,RIf1599c8_5479,RIf1588e8_5467,RIfe89cd0_7912,RIfc5ba78_6065,RIe1f9c68_4219,RIfc5bd48_6067,
        RIf1554e0_5430,RIf154298_5417,RIe1f4c40_4162,RIfe89b68_7911,RIfe89a00_7910,RIf150350_5372,RIe1f2918_4137,RIf14f3d8_5361,RIfccc818_7349,RIf14d920_5342,
        RIe1ed620_4078,RIe1eabf0_4048,RIe1e7ef0_4016,RIe1e51f0_3984,RIe1e24f0_3952,RIe1df7f0_3920,RIe1dcaf0_3888,RIe1d9df0_3856,RIe1d70f0_3824,RIe1d16f0_3760,
        RIe1ce9f0_3728,RIe1cbcf0_3696,RIe1c8ff0_3664,RIe1c62f0_3632,RIe1c35f0_3600,RIe1c08f0_3568,RIe1bdbf0_3536,RIfc680c0_6206,RIf14b058_5313,RIe1b8bc8_3479,
        RIe1b6b70_3456,RIfcac298_6981,RIf1499d8_5297,RIfe89190_7904,RIfec19c8_8323,RIf148a60_5286,RIfccdd30_7364,RIe1b2250_3404,RIfec1860_8322,RIfc6e768_6279,
        RIfc54728_5983,RIe1abfe0_3334,RIe1aa528_3315,RIe1a7f30_3288,RIe1a5230_3256,RIe1a2530_3224,RIe19f830_3192,RIe18bd30_2968,RIe178230_2744,RIe225b88_4719,
        RIe21a788_4591,RIe203f88_4335,RIe1fdfe8_4267,RIe1f73a0_4190,RIe1efee8_4107,RIe1d43f0_3792,RIe1baef0_3504,RIe1add68_3355,RIe1703a0_2654,RIdec4cd0_703,
        RIdec1fd0_671,RIfc7b4b8_6425,RIdebf2d0_639,RIfc7b1e8_6423,RIdebc5d0_607,RIdeb98d0_575,RIdeb6bd0_543,RIfe83358_7837,RIdeb11d0_479,RIee1e5c8_4804,
        RIdeae4d0_447,RIfc437c0_5790,RIdea93b8_415,RIdea2ab8_383,RIde9c1b8_351,RIfc90ea8_6671,RIfc7af18_6421,RIfe83088_7835,RIee1a950_4761,RIde906b0_294,
        RIde8cba0_276,RIfe82f20_7834,RIfe82db8_7833,RIee1a248_4756,RIfe831f0_7836,RIfcc2390_7232,RIee195a0_4747,RIfcbe718_7189,RIfea9e18_8249,RIfc43220_5786,
        RIe167868_2555,RIe164cd0_2524,RIe161fd0_2492,RIee36f88_5084,RIe15f2d0_2460,RIee35ea8_5072,RIe15c5d0_2428,RIe156bd0_2364,RIe153ed0_2332,RIfe83628_7839,
        RIe1511d0_2300,RIfebfda8_8303,RIe14e4d0_2268,RIfebfc40_8302,RIe14b7d0_2236,RIe148ad0_2204,RIe145dd0_2172,RIee34120_5051,RIee32ed8_5038,RIee31df8_5026,
        RIfcc1f58_7229,RIe140ad8_2113,RIdf3e878_2088,RIfe834c0_7838,RIdf3a390_2039,RIfc5a6c8_6051,RIfc91e20_6682,RIee2e888_4988,RIfc96a10_6736,RIdf35098_1980,
        RIfeab600_8266,RIdf30bb0_1931,RIfeab768_8267,RIfcbe9e8_7191,RIfc79fa0_6410,RIfc96740_6734,RIfc92258_6685,RIfea7118_8217,RIfea95a8_8243,RIdf26020_1809,
        RIdf24400_1789,RIfc79a00_6406,RIfc5add0_6056,RIfce5d18_7637,RIfc92690_6688,RIfce3018_7605,RIdf1f270_1731,RIfc79730_6404,RIdf19000_1661,RIdf168a0_1633,
        RIdf13ba0_1601,RIdf10ea0_1569,RIdf0e1a0_1537,RIdf0b4a0_1505,RIdf087a0_1473,RIdf05aa0_1441,RIdf02da0_1409,RIdefd3a0_1345,RIdefa6a0_1313,RIdef79a0_1281,
        RIdef4ca0_1249,RIdef1fa0_1217,RIdeef2a0_1185,RIdeec5a0_1153,RIdee98a0_1121,RIfc5b7a8_6063,RIfc5b640_6062,RIfc931d0_6696,RIfcecac8_7715,RIdee4710_1063,
        RIdee26b8_1040,RIdee07c8_1018,RIdede4a0_993,RIfcbf0f0_7196,RIfcbf528_7199,RIfc792f8_6401,RIfc93068_6695,RIded91a8_934,RIded6d18_908,RIded4e28_886,
        RIded2998_860,RIded00d0_831,RIdecd3d0_799,RIdeca6d0_767,RIdec79d0_735,RIdeb3ed0_511,RIde958b8_319,RIe16dad8_2625,RIe1598d0_2396,RIe1430d0_2140,
        RIdf37ac8_2010,RIdf2c128_1878,RIdf1c9a8_1702,RIdf000a0_1377,RIdee6ba0_1089,RIdedb908_962,RIde7b800_192,RIe19cf68_3163,RIe19a268_3131,RIfc8d7d0_6632,
        RIe197568_3099,RIfc561e0_6002,RIe194868_3067,RIe191b68_3035,RIe18ee68_3003,RIe189468_2939,RIe186768_2907,RIf143330_5224,RIe183a68_2875,RIfc7d948_6451,
        RIe180d68_2843,RIe17e068_2811,RIe17b368_2779,RIfc564b0_6004,RIfcd6700_7462,RIfc461f0_5820,RIe175698_2713,RIfc46088_5819,RIfc45f20_5818,RIfc7dc18_6453,
        RIfcd69d0_7464,RIfc98630_6756,RIfcc2a98_7237,RIfc7d510_6448,RIe173208_2687,RIfc8e478_6641,RIfc45ae8_5815,RIfc8e8b0_6644,RIfc45980_5814,RIfe82ae8_7831,
        RIe2232c0_4690,RIf16ba10_5684,RIe2205c0_4658,RIfcd24e8_7415,RIe21d8c0_4626,RIe217ec0_4562,RIe2151c0_4530,RIfebf268_8295,RIe2124c0_4498,RIf168d10_5652,
        RIe20f7c0_4466,RIfc7d240_6446,RIe20cac0_4434,RIe209dc0_4402,RIe2070c0_4370,RIf166e20_5630,RIfebf6a0_8298,RIfebf808_8299,RIfebf538_8297,RIfc8eb80_6646,
        RIf164120_5598,RIfc453e0_5810,RIf161b28_5571,RIf15fc38_5549,RIf15dd48_5527,RIe1fc968_4251,RIe1fb888_4239,RIfebf3d0_8296,RIf15b318_5497,RIfca2518_6869,
        RIfc8f120_6650,RIfebfad8_8301,RIfebf970_8300,RIfc7cca0_6442,RIe1f9dd0_4220,RIfe82c50_7832,RIf155648_5431,RIfc8f288_6651,RIe1f4f10_4164,RIf152d80_5402,
        RIfc8f828_6655,RIfcb3b88_7067,RIe1f2d50_4140,RIfc445d0_5800,RIfc8faf8_6657,RIf14da88_5343,RIe1eda58_4081,RIe1eb028_4051,RIe1e8328_4019,RIe1e5628_3987,
        RIe1e2928_3955,RIe1dfc28_3923,RIe1dcf28_3891,RIe1da228_3859,RIe1d7528_3827,RIe1d1b28_3763,RIe1cee28_3731,RIe1cc128_3699,RIe1c9428_3667,RIe1c6728_3635,
        RIe1c3a28_3603,RIe1c0d28_3571,RIe1be028_3539,RIfc7bff8_6433,RIfc44030_5796,RIe1b9000_3482,RIe1b6fa8_3459,RIfcbdd40_7182,RIfc8ff30_6660,RIe1b50b8_3437,
        RIe1b3d08_3423,RIfcbe178_7185,RIfc43d60_5794,RIe1b2520_3406,RIe1b0798_3385,RIfcdb5c0_7518,RIfc7ba58_6429,RIe1ac148_3335,RIe1aa960_3318,RIe1a8368_3291,
        RIe1a5668_3259,RIe1a2968_3227,RIe19fc68_3195,RIe18c168_2971,RIe178668_2747,RIe225fc0_4722,RIe21abc0_4594,RIe2043c0_4338,RIe1fe420_4270,RIe1f77d8_4193,
        RIe1f0320_4110,RIe1d4828_3795,RIe1bb328_3507,RIe1ae1a0_3358,RIe1707d8_2657,RIdec4b68_702,RIdec1e68_670,RIfc5df08_6091,RIdebf168_638,RIfce6df8_7649,
        RIdebc468_606,RIdeb9768_574,RIdeb6a68_542,RIfc75ef0_6364,RIdeb1068_478,RIfcc12b0_7220,RIdeae368_446,RIfc5e340_6094,RIdea9070_414,RIdea2770_382,
        RIde9be70_350,RIfced4a0_7722,RIfcc1418_7221,RIfc95930_6724,RIfcec0f0_7708,RIde90368_293,RIde8c858_275,RIde893d8_259,RIde84ef0_238,RIde80d50_218,
        RIfc95a98_6725,RIfced068_7719,RIfced1d0_7720,RIfcedfe0_7730,RIe16b0a8_2595,RIe169758_2577,RIe167700_2554,RIe164b68_2523,RIe161e68_2491,RIee36e20_5083,
        RIe15f168_2459,RIfc426e0_5778,RIe15c468_2427,RIe156a68_2363,RIe153d68_2331,RIfe82818_7829,RIe151068_2299,RIee34c60_5059,RIe14e368_2267,RIfc5f9c0_6110,
        RIe14b668_2235,RIe148968_2203,RIe145c68_2171,RIfccfef0_7388,RIfca57b8_6905,RIfc600c8_6115,RIfcafda8_7023,RIe140970_2112,RIdf3e710_2087,RIdf3c6b8_2064,
        RIdf3a228_2038,RIfc5fc90_6112,RIee2f3c8_4996,RIfc742d0_6344,RIee2d208_4972,RIdf34f30_1979,RIfebf100_8294,RIdf30a48_1930,RIdf2ecc0_1909,RIfcb08e8_7031,
        RIfcee418_7733,RIfc95ed0_6728,RIfcdef68_7559,RIdf29e00_1853,RIdf27c40_1829,RIdf25eb8_1808,RIdf24298_1788,RIfc5ed18_6101,RIfcee850_7736,RIdf227e0_1769,
        RIfc5efe8_6103,RIdf212c8_1754,RIfeaa520_8254,RIdf1ad88_1682,RIdf18e98_1660,RIdf16738_1632,RIdf13a38_1600,RIdf10d38_1568,RIdf0e038_1536,RIdf0b338_1504,
        RIdf08638_1472,RIdf05938_1440,RIdf02c38_1408,RIdefd238_1344,RIdefa538_1312,RIdef7838_1280,RIdef4b38_1248,RIdef1e38_1216,RIdeef138_1184,RIdeec438_1152,
        RIdee9738_1120,RIfcc96e0_7314,RIfccfd88_7387,RIfc60aa0_6122,RIfca5ec0_6910,RIdee45a8_1062,RIdee2550_1039,RIdee0660_1017,RIfe826b0_7828,RIfcdeb30_7556,
        RIfc73bc8_6339,RIfca5bf0_6908,RIfc73a60_6338,RIfe82980_7830,RIded6bb0_907,RIded4cc0_885,RIded2830_859,RIdecff68_830,RIdecd268_798,RIdeca568_766,
        RIdec7868_734,RIdeb3d68_510,RIde95570_318,RIe16d970_2624,RIe159768_2395,RIe142f68_2139,RIdf37960_2009,RIdf2bfc0_1877,RIdf1c840_1701,RIdefff38_1376,
        RIdee6a38_1088,RIdedb7a0_961,RIde7b4b8_191,RIe19ce00_3162,RIe19a100_3130,RIfce96c0_7678,RIe197400_3098,RIf144410_5236,RIe194700_3066,RIe191a00_3034,
        RIe18ed00_3002,RIe189300_2938,RIe186600_2906,RIfebee30_8292,RIe183900_2874,RIfcdbcc8_7523,RIe180c00_2842,RIe17df00_2810,RIe17b200_2778,RIf141f80_5210,
        RIfce7398_7653,RIfcb1e00_7046,RIfe82548_7827,RIfca42a0_6890,RIfcbff00_7206,RIfcaaee8_6967,RIee3d090_5153,RIfc5c180_6070,RIfce35b8_7609,RIee399b8_5114,
        RIfea8a68_8235,RIf16fef8_5733,RIfebecc8_8291,RIfc5c450_6072,RIfce9288_7675,RIfc40778_5759,RIe223158_4689,RIfce77d0_7656,RIe220458_4657,RIfce24d8_7597,
        RIe21d758_4625,RIe217d58_4561,RIe215058_4529,RIfce8a18_7669,RIe212358_4497,RIfce1998_7589,RIe20f658_4465,RIfc77840_6382,RIe20c958_4433,RIe209c58_4401,
        RIe206f58_4369,RIf166cb8_5629,RIf165bd8_5617,RIfe81fa8_7823,RIfe81e40_7822,RIfc5c888_6075,RIfceb178_7697,RIf1631a8_5587,RIf1619c0_5570,RIfccf248_7379,
        RIfc77570_6380,RIe1fc800_4250,RIe1fb720_4238,RIf15c830_5512,RIf15b1b0_5496,RIfcd0fd0_7400,RIfccc6b0_7348,RIf158bb8_5469,RIf157808_5455,RIfc5d0f8_6081,
        RIfebef98_8293,RIfcc8a38_7305,RIfcd7ab0_7476,RIfcb1428_7039,RIfeaa0e8_8251,RIfccc548_7347,RIfce3450_7608,RIf1504b8_5373,RIe1f2be8_4139,RIf14f540_5362,
        RIfc772a0_6378,RIfcec258_7709,RIe1ed8f0_4080,RIe1eaec0_4050,RIe1e81c0_4018,RIe1e54c0_3986,RIe1e27c0_3954,RIe1dfac0_3922,RIe1dcdc0_3890,RIe1da0c0_3858,
        RIe1d73c0_3826,RIe1d19c0_3762,RIe1cecc0_3730,RIe1cbfc0_3698,RIe1c92c0_3666,RIe1c65c0_3634,RIe1c38c0_3602,RIe1c0bc0_3570,RIe1bdec0_3538,RIf14c570_5328,
        RIf14b328_5315,RIe1b8e98_3481,RIe1b6e40_3458,RIfc76760_6370,RIfc94b20_6714,RIe1b4f50_3436,RIe1b3ba0_3422,RIfcec3c0_7710,RIfceb010_7696,RIfe823e0_7826,
        RIfe82110_7824,RIfcdd8e8_7543,RIfcc0ba8_7215,RIfe82278_7825,RIe1aa7f8_3317,RIe1a8200_3290,RIe1a5500_3258,RIe1a2800_3226,RIe19fb00_3194,RIe18c000_2970,
        RIe178500_2746,RIe225e58_4721,RIe21aa58_4593,RIe204258_4337,RIe1fe2b8_4269,RIe1f7670_4192,RIe1f01b8_4109,RIe1d46c0_3794,RIe1bb1c0_3506,RIe1ae038_3357,
        RIe170670_2656,RIdec4fa0_705,RIdec22a0_673,RIee1fdb0_4821,RIdebf5a0_641,RIee1f270_4813,RIdebc8a0_609,RIdeb9ba0_577,RIdeb6ea0_545,RIee1ecd0_4809,
        RIdeb14a0_481,RIee1e730_4805,RIdeae7a0_449,RIee1d920_4795,RIdea9a48_417,RIdea3148_385,RIde9c848_353,RIee1cb10_4785,RIee1ba30_4773,RIee1b1c0_4767,
        RIfec04b0_8308,RIfe850e0_7858,RIde8d230_278,RIfea9cb0_8248,RIfe84f78_7857,RIee1a3b0_4757,RIfe853b0_7860,RIee199d8_4750,RIfe85248_7859,RIee39148_5108,
        RIe16b378_2597,RIee38608_5100,RIe167b38_2557,RIe164fa0_2526,RIe1622a0_2494,RIfe85950_7864,RIe15f5a0_2462,RIee36010_5073,RIe15c8a0_2430,RIe156ea0_2366,
        RIe1541a0_2334,RIfe85c20_7866,RIe1514a0_2302,RIee34dc8_5060,RIe14e7a0_2270,RIfc861b0_6548,RIe14baa0_2238,RIe148da0_2206,RIe1460a0_2174,RIee343f0_5053,
        RIfe85518_7861,RIfe857e8_7863,RIfe85680_7862,RIe140c40_2114,RIdf3eb48_2090,RIdf3c820_2065,RIdf3a660_2041,RIfc9d4f0_6812,RIee2f698_4998,RIfc52298_5957,
        RIee2d4d8_4974,RIdf35368_1982,RIdf32ed8_1956,RIdf30e80_1933,RIfe85ab8_7865,RIee2b8b8_4954,RIee29f68_4936,RIee28bb8_4922,RIee27970_4909,RIdf2a0d0_1855,
        RIfe84e10_7856,RIdf262f0_1811,RIfe84ca8_7855,RIee27100_4903,RIee26b60_4899,RIfcd32f8_7425,RIee265c0_4895,RIfc9e300_6822,RIdf1f540_1733,RIee25eb8_4890,
        RIfe84b40_7854,RIdf16b70_1635,RIdf13e70_1603,RIdf11170_1571,RIdf0e470_1539,RIdf0b770_1507,RIdf08a70_1475,RIdf05d70_1443,RIdf03070_1411,RIdefd670_1347,
        RIdefa970_1315,RIdef7c70_1283,RIdef4f70_1251,RIdef2270_1219,RIdeef570_1187,RIdeec870_1155,RIdee9b70_1123,RIfec0348_8307,RIfcb54d8_7085,RIee23cf8_4866,
        RIfc54e30_5988,RIfec0078_8305,RIdee2988_1042,RIfec01e0_8306,RIdede770_995,RIfcd7ee8_7479,RIfcd43d8_7437,RIfc88eb0_6580,RIfc9e5d0_6824,RIded9478_936,
        RIded6fe8_910,RIded50f8_888,RIfeab330_8264,RIded03a0_833,RIdecd6a0_801,RIdeca9a0_769,RIdec7ca0_737,RIdeb41a0_513,RIde95f48_321,RIe16dda8_2627,
        RIe159ba0_2398,RIe1433a0_2142,RIdf37d98_2012,RIdf2c3f8_1880,RIdf1cc78_1704,RIdf00370_1379,RIdee6e70_1091,RIdedbbd8_964,RIde7be90_194,RIe19d238_3165,
        RIe19a538_3133,RIf145658_5249,RIe197838_3101,RIf1446e0_5238,RIe194b38_3069,RIe191e38_3037,RIe18f138_3005,RIe189738_2941,RIe186a38_2909,RIf143600_5226,
        RIe183d38_2877,RIf142c28_5219,RIe181038_2845,RIe17e338_2813,RIe17b638_2781,RIf1420e8_5211,RIf140a68_5195,RIf1401f8_5189,RIfebff10_8304,RIf13faf0_5184,
        RIf13ee48_5175,RIee3e2d8_5166,RIee3d1f8_5154,RIee3c118_5142,RIee3b038_5130,RIee39c88_5116,RIfe838f8_7841,RIf1701c8_5735,RIfc5ab00_6054,RIf16e008_5711,
        RIfcb0e88_7035,RIf16caf0_5696,RIe223590_4692,RIf16bce0_5686,RIe220890_4660,RIf16ac00_5674,RIe21db90_4628,RIe218190_4564,RIe215490_4532,RIf16a228_5667,
        RIe212790_4500,RIf168fe0_5654,RIe20fa90_4468,RIf167d98_5641,RIe20cd90_4436,RIe20a090_4404,RIe207390_4372,RIf1670f0_5632,RIf165ea8_5619,RIe202200_4314,
        RIfe83e98_7845,RIf164f30_5608,RIf1643f0_5600,RIfce8310_7664,RIf161df8_5573,RIf15ff08_5551,RIf15e018_5529,RIfe83d30_7844,RIfe84000_7846,RIf15cb00_5514,
        RIf15b5e8_5499,RIf15a508_5487,RIfc887a8_6575,RIf158d20_5470,RIf157970_5456,RIf156cc8_5447,RIfe84438_7849,RIf156020_5438,RIfc51fc8_5955,RIf154568_5419,
        RIe1f51e0_4166,RIf153050_5404,RIf1519d0_5388,RIf150788_5375,RIfe842d0_7848,RIf14f810_5364,RIf14eb68_5355,RIf14dd58_5345,RIfe84168_7847,RIe1eb2f8_4053,
        RIe1e85f8_4021,RIe1e58f8_3989,RIe1e2bf8_3957,RIe1dfef8_3925,RIe1dd1f8_3893,RIe1da4f8_3861,RIe1d77f8_3829,RIe1d1df8_3765,RIe1cf0f8_3733,RIe1cc3f8_3701,
        RIe1c96f8_3669,RIe1c69f8_3637,RIe1c3cf8_3605,RIe1c0ff8_3573,RIe1be2f8_3541,RIf14c840_5330,RIf14b5f8_5317,RIfe83a60_7842,RIfe849d8_7853,RIfc74168_6343,
        RIf149b40_5298,RIfe83bc8_7843,RIfe84708_7851,RIf148d30_5288,RIf147ae8_5275,RIfe84870_7852,RIe1b0900_3386,RIf146fa8_5267,RIf146300_5258,RIfe845a0_7850,
        RIfe83790_7840,RIe1a8638_3293,RIe1a5938_3261,RIe1a2c38_3229,RIe19ff38_3197,RIe18c438_2973,RIe178938_2749,RIe226290_4724,RIe21ae90_4596,RIe204690_4340,
        RIe1fe6f0_4272,RIe1f7aa8_4195,RIe1f05f0_4112,RIe1d4af8_3797,RIe1bb5f8_3509,RIe1ae470_3360,RIe170aa8_2659,RIdec4e38_704,RIdec2138_672,RIee1fc48_4820,
        RIdebf438_640,RIfc49490_5856,RIdebc738_608,RIdeb9a38_576,RIdeb6d38_544,RIfc48ef0_5852,RIdeb1338_480,RIfcd9b08_7499,RIdeae638_448,RIfc8b610_6608,
        RIdea9700_416,RIdea2e00_384,RIde9c500_352,RIee1c9a8_4784,RIee1b8c8_4772,RIfc80918_6485,RIfcdad50_7512,RIfe86e68_7879,RIde8cee8_277,RIfe86d00_7878,
        RIfec0d20_8314,RIde81098_219,RIfc8b8e0_6610,RIfcd2d58_7421,RIfce4530_7620,RIfc8ba48_6611,RIe16b210_2596,RIe1698c0_2578,RIe1679d0_2556,RIe164e38_2525,
        RIe162138_2493,RIee370f0_5085,RIe15f438_2461,RIfc999e0_6770,RIe15c738_2429,RIe156d38_2365,RIe154038_2333,RIfc3f260_5744,RIe151338_2301,RIfc48518_5845,
        RIe14e638_2269,RIfc99e18_6773,RIe14b938_2237,RIe148c38_2205,RIe145f38_2173,RIee34288_5052,RIee33040_5039,RIee31f60_5027,RIfcd99a0_7498,RIfe86b98_7877,
        RIdf3e9e0_2089,RIfe86a30_7876,RIdf3a4f8_2040,RIfcc3470_7244,RIee2f530_4997,RIfc7fdd8_6477,RIee2d370_4973,RIdf35200_1981,RIfec0ff0_8316,RIdf30d18_1932,
        RIfec0e88_8315,RIfcd2a88_7419,RIfc8c858_6621,RIfc47ca8_5839,RIfcd6430_7460,RIdf29f68_1854,RIdf27da8_1830,RIdf26188_1810,RIdf24568_1790,RIfc8cb28_6623,
        RIfcdb188_7515,RIdf22948_1770,RIfc475a0_5834,RIdf21430_1755,RIdf1f3d8_1732,RIfec0bb8_8313,RIfe868c8_7875,RIdf16a08_1634,RIdf13d08_1602,RIdf11008_1570,
        RIdf0e308_1538,RIdf0b608_1506,RIdf08908_1474,RIdf05c08_1442,RIdf02f08_1410,RIdefd508_1346,RIdefa808_1314,RIdef7b08_1282,RIdef4e08_1250,RIdef2108_1218,
        RIdeef408_1186,RIdeec708_1154,RIdee9a08_1122,RIee254e0_4883,RIee246d0_4873,RIee23b90_4865,RIee231b8_4858,RIfe86fd0_7880,RIdee2820_1041,RIdee0930_1019,
        RIdede608_994,RIfc55da8_5999,RIfc98a68_6759,RIfcc3038_7241,RIfc464c0_5822,RIded9310_935,RIded6e80_909,RIded4f90_887,RIded2b00_861,RIded0238_832,
        RIdecd538_800,RIdeca838_768,RIdec7b38_736,RIdeb4038_512,RIde95c00_320,RIe16dc40_2626,RIe159a38_2397,RIe143238_2141,RIdf37c30_2011,RIdf2c290_1879,
        RIdf1cb10_1703,RIdf00208_1378,RIdee6d08_1090,RIdedba70_963,RIde7bb48_193,RIe19d0d0_3164,RIe19a3d0_3132,RIf1454f0_5248,RIe1976d0_3100,RIf144578_5237,
        RIe1949d0_3068,RIe191cd0_3036,RIe18efd0_3004,RIe1895d0_2940,RIe1868d0_2908,RIf143498_5225,RIe183bd0_2876,RIfc51758_5949,RIe180ed0_2844,RIe17e1d0_2812,
        RIe17b4d0_2780,RIfc9b060_6786,RIfc9ee40_6830,RIe176e80_2730,RIe175800_2714,RIfcb70f8_7105,RIfce0cf0_7580,RIfcc4280_7254,RIfcba7d0_7144,RIee3bfb0_5141,
        RIee3aed0_5129,RIee39b20_5115,RIe173370_2688,RIf170060_5734,RIf16f3b8_5725,RIf16dea0_5710,RIf16d4c8_5703,RIf16c988_5695,RIe223428_4691,RIf16bb78_5685,
        RIe220728_4659,RIf16aa98_5673,RIe21da28_4627,RIe218028_4563,RIe215328_4531,RIf16a0c0_5666,RIe212628_4499,RIf168e78_5653,RIe20f928_4467,RIf167c30_5640,
        RIe20cc28_4435,RIe209f28_4403,RIe207228_4371,RIf166f88_5631,RIf165d40_5618,RIfec0618_8309,RIfe86760_7874,RIfc52b08_5963,RIf164288_5599,RIf163310_5588,
        RIf161c90_5572,RIf15fda0_5550,RIf15deb0_5528,RIfe865f8_7873,RIfe85d88_7867,RIf15c998_5513,RIf15b480_5498,RIf15a3a0_5486,RIf159b30_5480,RIfc83348_6515,
        RIfc4ade0_5874,RIfc89720_6586,RIe1f9f38_4221,RIfc4ac78_5873,RIfc9f110_6832,RIfc4ab10_5872,RIe1f5078_4165,RIf152ee8_5403,RIfc899f0_6588,RIf150620_5374,
        RIe1f2eb8_4141,RIf14f6a8_5363,RIf14ea00_5354,RIf14dbf0_5344,RIe1edbc0_4082,RIe1eb190_4052,RIe1e8490_4020,RIe1e5790_3988,RIe1e2a90_3956,RIe1dfd90_3924,
        RIe1dd090_3892,RIe1da390_3860,RIe1d7690_3828,RIe1d1c90_3764,RIe1cef90_3732,RIe1cc290_3700,RIe1c9590_3668,RIe1c6890_3636,RIe1c3b90_3604,RIe1c0e90_3572,
        RIe1be190_3540,RIf14c6d8_5329,RIf14b490_5316,RIfe85ef0_7868,RIfe86490_7872,RIf14a248_5303,RIfc819f8_6497,RIfec0a50_8312,RIfe861c0_7870,RIf148bc8_5287,
        RIf147980_5274,RIfe86328_7871,RIfec0780_8310,RIfcbb478_7153,RIf146198_5257,RIfe86058_7869,RIfec08e8_8311,RIe1a84d0_3292,RIe1a57d0_3260,RIe1a2ad0_3228,
        RIe19fdd0_3196,RIe18c2d0_2972,RIe1787d0_2748,RIe226128_4723,RIe21ad28_4595,RIe204528_4339,RIe1fe588_4271,RIe1f7940_4194,RIe1f0488_4111,RIe1d4990_3796,
        RIe1bb490_3508,RIe1ae308_3359,RIe170940_2658,RIdec53d8_708,RIdec26d8_676,RIee20080_4823,RIdebf9d8_644,RIee1f3d8_4814,RIdebccd8_612,RIdeb9fd8_580,
        RIdeb72d8_548,RIee1ee38_4810,RIdeb18d8_484,RIee1e898_4806,RIdeaebd8_452,RIee1da88_4796,RIdeaa420_420,RIdea3b20_388,RIde9d220_356,RIee1cde0_4787,
        RIee1bd00_4775,RIee1b490_4769,RIfcd8a28_7487,RIde91088_297,RIde8d8c0_280,RIfe7dac0_7774,RIfe7d958_7773,RIee1a518_4758,RIee19e10_4753,RIee19b40_4751,
        RIfc768c8_6371,RIfcd05f8_7393,RIfe7dd90_7776,RIee38770_5101,RIfe7dc28_7775,RIe1653d8_2529,RIe1626d8_2497,RIee373c0_5087,RIe15f9d8_2465,RIee362e0_5075,
        RIe15ccd8_2433,RIe1572d8_2369,RIe1545d8_2337,RIfe7def8_7777,RIe1518d8_2305,RIfebdeb8_8281,RIe14ebd8_2273,RIfc649e8_6167,RIe14bed8_2241,RIe1491d8_2209,
        RIe1464d8_2177,RIfe7d7f0_7772,RIfe7d688_7771,RIee32230_5029,RIfceb9e8_7703,RIfebdd50_8280,RIfe7d520_7770,RIfebdbe8_8279,RIfe7d3b8_7769,RIfc734c0_6334,
        RIee2f968_5000,RIfccfab8_7385,RIee2d7a8_4976,RIdf357a0_1985,RIdf33310_1959,RIdf312b8_1936,RIdf2f0f8_1912,RIee2bcf0_4957,RIee2a238_4938,RIee28e88_4924,
        RIee27c40_4911,RIfe7ce18_7765,RIfe7ccb0_7764,RIfe7cf80_7766,RIfe7cb48_7763,RIee27268_4904,RIee26e30_4901,RIee26890_4897,RIfcaa0d8_6957,RIee262f0_4893,
        RIfe7d250_7768,RIee26020_4891,RIfe7d0e8_7767,RIdf16fa8_1638,RIdf142a8_1606,RIdf115a8_1574,RIdf0e8a8_1542,RIdf0bba8_1510,RIdf08ea8_1478,RIdf061a8_1446,
        RIdf034a8_1414,RIdefdaa8_1350,RIdefada8_1318,RIdef80a8_1286,RIdef53a8_1254,RIdef26a8_1222,RIdeef9a8_1190,RIdeecca8_1158,RIdee9fa8_1126,RIee25648_4884,
        RIee249a0_4875,RIfebe020_8282,RIee23488_4860,RIfebe2f0_8284,RIfebe188_8283,RIfe7e1c8_7779,RIfe7e060_7778,RIfcbf7f8_7201,RIfc7aae0_6418,RIfc787b8_6393,
        RIfc618b0_6132,RIded98b0_939,RIded72b8_912,RIded5530_891,RIded2dd0_863,RIded07d8_836,RIdecdad8_804,RIdecadd8_772,RIdec80d8_740,RIdeb45d8_516,
        RIde96920_324,RIe16e1e0_2630,RIe159fd8_2401,RIe1437d8_2145,RIdf381d0_2015,RIdf2c830_1883,RIdf1d0b0_1707,RIdf007a8_1382,RIdee72a8_1094,RIdedc010_967,
        RIde7c868_197,RIe19d670_3168,RIe19a970_3136,RIfe7b630_7748,RIe197c70_3104,RIfe7b4c8_7747,RIe194f70_3072,RIe192270_3040,RIe18f570_3008,RIe189b70_2944,
        RIe186e70_2912,RIfe7b360_7746,RIe184170_2880,RIfe7b1f8_7745,RIe181470_2848,RIe17e770_2816,RIe17ba70_2784,RIf1423b8_5213,RIf140ea0_5198,RIf140360_5190,
        RIfe7b798_7749,RIf13fc58_5185,RIf13f280_5178,RIfc79460_6402,RIee3d4c8_5156,RIfe7b090_7744,RIfe7af28_7743,RIee39df0_5117,RIe1737a8_2691,RIfe7adc0_7742,
        RIfe7ac58_7741,RIf16e440_5714,RIfcb20d0_7048,RIfe7bd38_7753,RIe2239c8_4695,RIf16be48_5687,RIe220cc8_4663,RIf16aed0_5676,RIe21dfc8_4631,RIe2185c8_4567,
        RIe2158c8_4535,RIfebd7b0_8276,RIe212bc8_4503,RIfebd648_8275,RIe20fec8_4471,RIfe7b900_7750,RIe20d1c8_4439,RIe20a4c8_4407,RIe2077c8_4375,RIf167258_5633,
        RIf166178_5621,RIe2024d0_4316,RIfe7bbd0_7752,RIf165368_5611,RIf1646c0_5602,RIfcd0a30_7396,RIf1620c8_5575,RIf1601d8_5553,RIf15e2e8_5531,RIfe7ba68_7751,
        RIfe7bea0_7754,RIf15cdd0_5516,RIf15b8b8_5501,RIf15a7d8_5489,RIfca4840_6894,RIf158ff0_5472,RIf157c40_5458,RIf156f98_5449,RIfe7c170_7756,RIf156458_5441,
        RIf155918_5433,RIf1549a0_5422,RIe1f54b0_4168,RIfe7c008_7755,RIf151b38_5389,RIf150bc0_5378,RIe1f32f0_4144,RIf14fae0_5366,RIf14ee38_5357,RIf14e028_5347,
        RIe1edff8_4085,RIe1eb730_4056,RIe1e8a30_4024,RIe1e5d30_3992,RIe1e3030_3960,RIe1e0330_3928,RIe1dd630_3896,RIe1da930_3864,RIe1d7c30_3832,RIe1d2230_3768,
        RIe1cf530_3736,RIe1cc830_3704,RIe1c9b30_3672,RIe1c6e30_3640,RIe1c4130_3608,RIe1c1430_3576,RIe1be730_3544,RIf14cb10_5332,RIf14b8c8_5319,RIfebda80_8278,
        RIfe7c878_7761,RIf14a680_5306,RIfe7c2d8_7757,RIfe7c9e0_7762,RIfe7c440_7758,RIf149000_5290,RIf147db8_5277,RIe1b2688_3407,RIfebd918_8277,RIfe7c5a8_7759,
        RIf146738_5261,RIfe7c710_7760,RIe1aad98_3321,RIe1a8a70_3296,RIe1a5d70_3264,RIe1a3070_3232,RIe1a0370_3200,RIe18c870_2976,RIe178d70_2752,RIe2266c8_4727,
        RIe21b2c8_4599,RIe204ac8_4343,RIe1feb28_4275,RIe1f7ee0_4198,RIe1f0a28_4115,RIe1d4f30_3800,RIe1bba30_3512,RIe1ae8a8_3363,RIe170ee0_2662,RIdec5270_707,
        RIdec2570_675,RIee1ff18_4822,RIdebf870_643,RIfe7f848_7795,RIdebcb70_611,RIdeb9e70_579,RIdeb7170_547,RIfe7fc80_7798,RIdeb1770_483,RIfca5d58_6909,
        RIdeaea70_451,RIfcaf808_7019,RIdeaa0d8_419,RIdea37d8_387,RIde9ced8_355,RIfcdc3d0_7528,RIfcce438_7369,RIfcb0a50_7032,RIfc75680_6358,RIde90d40_296,
        RIfe7f9b0_7796,RIde89720_260,RIde85580_240,RIde81728_221,RIfc52f40_5966,RIfc82100_6502,RIfca7108_6923,RIfe7fb18_7797,RIe16b648_2599,RIe169a28_2579,
        RIe167ca0_2558,RIe165270_2528,RIe162570_2496,RIee37258_5086,RIe15f870_2464,RIee36178_5074,RIe15cb70_2432,RIe157170_2368,RIe154470_2336,RIfc86fc0_6558,
        RIe151770_2304,RIfc4eff8_5921,RIe14ea70_2272,RIfce1290_7584,RIe14bd70_2240,RIe149070_2208,RIe146370_2176,RIee34558_5054,RIee331a8_5040,RIee320c8_5028,
        RIee31150_5017,RIfe800b8_7801,RIfe7ff50_7800,RIdf3caf0_2067,RIfe7fde8_7799,RIfcc8330_7300,RIee2f800_4999,RIfca0d30_6852,RIee2d640_4975,RIdf35638_1984,
        RIdf331a8_1958,RIdf31150_1935,RIdf2ef90_1911,RIee2bb88_4956,RIee2a0d0_4937,RIee28d20_4923,RIfe7f578_7793,RIdf2a238_1856,RIdf27f10_1831,RIfe7f6e0_7794,
        RIdf246d0_1791,RIfcce9d8_7373,RIfc63638_6153,RIdf22c18_1772,RIfc62990_6144,RIdf21700_1757,RIdf1f810_1735,RIfeaa958_8257,RIdf19168_1662,RIdf16e40_1637,
        RIdf14140_1605,RIdf11440_1573,RIdf0e740_1541,RIdf0ba40_1509,RIdf08d40_1477,RIdf06040_1445,RIdf03340_1413,RIdefd940_1349,RIdefac40_1317,RIdef7f40_1285,
        RIdef5240_1253,RIdef2540_1221,RIdeef840_1189,RIdeecb40_1157,RIdee9e40_1125,RIfcb7800_7110,RIee24838_4874,RIfc4cb68_5895,RIee23320_4859,RIfe80388_7803,
        RIdee2c58_1044,RIfe80220_7802,RIdedea40_997,RIfc98900_6758,RIee223a8_4848,RIfcc8600_7302,RIee212c8_4836,RIded9748_938,RIfe804f0_7804,RIded53c8_890,
        RIded2c68_862,RIded0670_835,RIdecd970_803,RIdecac70_771,RIdec7f70_739,RIdeb4470_515,RIde965d8_323,RIe16e078_2629,RIe159e70_2400,RIe143670_2144,
        RIdf38068_2014,RIdf2c6c8_1882,RIdf1cf48_1706,RIdf00640_1381,RIdee7140_1093,RIdedbea8_966,RIde7c520_196,RIe19d508_3167,RIe19a808_3135,RIfe7ee70_7788,
        RIe197b08_3103,RIfe7efd8_7789,RIe194e08_3071,RIe192108_3039,RIe18f408_3007,RIe189a08_2943,RIe186d08_2911,RIf143768_5227,RIe184008_2879,RIfc4bbf0_5884,
        RIe181308_2847,RIe17e608_2815,RIe17b908_2783,RIfe7f410_7792,RIf140d38_5197,RIe176fe8_2731,RIe175ad0_2716,RIfe7f2a8_7791,RIf13f118_5177,RIee3e440_5167,
        RIee3d360_5155,RIee3c280_5143,RIee3b1a0_5131,RIfe7f140_7790,RIe173640_2690,RIf170330_5736,RIf16f520_5726,RIf16e2d8_5713,RIf16d630_5704,RIfe7ea38_7785,
        RIe223860_4694,RIfc9c410_6800,RIe220b60_4662,RIfcb8340_7118,RIe21de60_4630,RIe218460_4566,RIe215760_4534,RIfc9cc80_6806,RIe212a60_4502,RIfc4ddb0_5908,
        RIe20fd60_4470,RIfc873f8_6561,RIe20d060_4438,RIe20a360_4406,RIe207660_4374,RIfc86750_6552,RIfc4e4b8_5913,RIe202368_4315,RIe200a18_4297,RIf165200_5610,
        RIf164558_5601,RIf163478_5589,RIf161f60_5574,RIf160070_5552,RIf15e180_5530,RIe1fcc38_4253,RIe1fb9f0_4240,RIf15cc68_5515,RIf15b750_5500,RIf15a670_5488,
        RIf159c98_5481,RIf158e88_5471,RIf157ad8_5457,RIf156e30_5448,RIfe7e768_7783,RIf1562f0_5440,RIf1557b0_5432,RIf154838_5421,RIfe7e8d0_7784,RIf1531b8_5405,
        RIfc52400_5958,RIf150a58_5377,RIe1f3188_4143,RIf14f978_5365,RIf14ecd0_5356,RIf14dec0_5346,RIe1ede90_4084,RIe1eb5c8_4055,RIe1e88c8_4023,RIe1e5bc8_3991,
        RIe1e2ec8_3959,RIe1e01c8_3927,RIe1dd4c8_3895,RIe1da7c8_3863,RIe1d7ac8_3831,RIe1d20c8_3767,RIe1cf3c8_3735,RIe1cc6c8_3703,RIe1c99c8_3671,RIe1c6cc8_3639,
        RIe1c3fc8_3607,RIe1c12c8_3575,RIe1be5c8_3543,RIf14c9a8_5331,RIf14b760_5318,RIfe7ed08_7787,RIfe7e600_7782,RIf14a518_5305,RIfca1f78_6865,RIfe7eba0_7786,
        RIfe7e498_7781,RIf148e98_5289,RIf147c50_5276,RIfe7e330_7780,RIe1b0a68_3387,RIf147278_5269,RIf1465d0_5260,RIe1ac418_3337,RIe1aac30_3320,RIe1a8908_3295,
        RIe1a5c08_3263,RIe1a2f08_3231,RIe1a0208_3199,RIe18c708_2975,RIe178c08_2751,RIe226560_4726,RIe21b160_4598,RIe204960_4342,RIe1fe9c0_4274,RIe1f7d78_4197,
        RIe1f08c0_4114,RIe1d4dc8_3799,RIe1bb8c8_3511,RIe1ae740_3362,RIe170d78_2661,RIdec56a8_710,RIdec29a8_678,RIfc54020_5978,RIdebfca8_646,RIee1f540_4815,
        RIdebcfa8_614,RIdeba2a8_582,RIdeb75a8_550,RIfc4fe08_5931,RIdeb1ba8_486,RIfc6b630_6244,RIdeaeea8_454,RIfc6a118_6229,RIdeaaab0_422,RIdea41b0_390,
        RIde9d8b0_358,RIfc69ce0_6226,RIee1be68_4776,RIfc653c0_6174,RIee1ac20_4763,RIde91718_299,RIde8df50_282,RIde89db0_262,RIde85c10_242,RIde81db8_223,
        RIfca76a8_6927,RIfcca4f0_7324,RIfc4ce38_5897,RIfc6b360_6242,RIe16b918_2601,RIe169cf8_2581,RIe167f70_2560,RIe1656a8_2531,RIe1629a8_2499,RIee37690_5089,
        RIe15fca8_2467,RIfce93f0_7676,RIe15cfa8_2435,RIe1575a8_2371,RIe1548a8_2339,RIee35908_5068,RIe151ba8_2307,RIee34f30_5061,RIe14eea8_2275,RIfce32e8_7607,
        RIe14c1a8_2243,RIe1494a8_2211,RIe1467a8_2179,RIfcde2c0_7550,RIfc687c8_6211,RIfca9160_6946,RIfcb1590_7040,RIe141078_2117,RIdf3ef80_2093,RIdf3cdc0_2069,
        RIfebeb60_8290,RIfc64448_6163,RIee2fad0_5001,RIfca7978_6929,RIfc676e8_6199,RIdf35a70_1987,RIdf335e0_1961,RIdf31420_1937,RIdf2f3c8_1914,RIfccef78_7377,
        RIfca6fa0_6922,RIfc62558_6141,RIfc61fb8_6137,RIfe81b70_7820,RIdf281e0_1833,RIfe81cd8_7821,RIdf249a0_1793,RIfc44300_5798,RIfcafc40_7022,RIdf22ee8_1774,
        RIfcaac18_6965,RIdf219d0_1759,RIdf1fae0_1737,RIdf1b1c0_1685,RIdf19438_1664,RIdf17278_1640,RIdf14578_1608,RIdf11878_1576,RIdf0eb78_1544,RIdf0be78_1512,
        RIdf09178_1480,RIdf06478_1448,RIdf03778_1416,RIdefdd78_1352,RIdefb078_1320,RIdef8378_1288,RIdef5678_1256,RIdef2978_1224,RIdeefc78_1192,RIdeecf78_1160,
        RIdeea278_1128,RIfc611a8_6127,RIfc61a18_6133,RIfca65c8_6915,RIfca6b68_6919,RIdee4b48_1066,RIdee2dc0_1045,RIdee0c00_1021,RIdedeba8_998,RIfc626c0_6142,
        RIfc738f8_6337,RIfcb31b0_7060,RIee21430_4837,RIded9a18_940,RIded7588_914,RIded5698_892,RIded30a0_865,RIded0aa8_838,RIdecdda8_806,RIdecb0a8_774,
        RIdec83a8_742,RIdeb48a8_518,RIde96fb0_326,RIe16e4b0_2632,RIe15a2a8_2403,RIe143aa8_2147,RIdf384a0_2017,RIdf2cb00_1885,RIdf1d380_1709,RIdf00a78_1384,
        RIdee7578_1096,RIdedc2e0_969,RIde7cef8_199,RIe19d940_3170,RIe19ac40_3138,RIfc64880_6166,RIe197f40_3106,RIf144848_5239,RIe195240_3074,RIe192540_3042,
        RIe18f840_3010,RIe189e40_2946,RIe187140_2914,RIf143a38_5229,RIe184440_2882,RIfc6f140_6286,RIe181740_2850,RIe17ea40_2818,RIe17bd40_2786,RIfc64f88_6171,
        RIf141008_5199,RIe177150_2732,RIfe81738_7817,RIfccabf8_7329,RIf13f3e8_5179,RIfca81e8_6935,RIee3d630_5157,RIfc66068_6183,RIfc6ed08_6283,RIfcdde88_7547,
        RIe173a78_2693,RIfc66338_6185,RIfc6eba0_6282,RIfc664a0_6186,RIfcacdd8_6989,RIfe81468_7815,RIe223c98_4697,RIfc66d10_6192,RIe220f98_4665,RIf16b038_5677,
        RIe21e298_4633,RIe218898_4569,RIe215b98_4537,RIfc3fc38_5751,RIe212e98_4505,RIfc67850_6200,RIe210198_4473,RIf167f00_5642,RIe20d498_4441,RIe20a798_4409,
        RIe207a98_4377,RIfcacb08_6987,RIfcac9a0_6986,RIfea8900_8234,RIfe818a0_7818,RIfca8a58_6941,RIfccad60_7330,RIfcac838_6985,RIfc67418_6197,RIf160340_5554,
        RIf15e450_5532,RIfe81a08_7819,RIfe81300_7814,RIfc6dac0_6270,RIf15ba20_5502,RIfc6d958_6269,RIfc6d7f0_6268,RIfc587d8_6029,RIfc6cf80_6262,RIfc6d3b8_6265,
        RIfe815d0_7816,RIfc6d520_6266,RIfcabe60_6978,RIfc6d0e8_6263,RIe1f5780_4170,RIfc6c5a8_6255,RIfc68d68_6215,RIfc68c00_6214,RIe1f3458_4145,RIfc68a98_6213,
        RIfccb8a0_7338,RIfca9b38_6953,RIe1ee160_4086,RIe1eba00_4058,RIe1e8d00_4026,RIe1e6000_3994,RIe1e3300_3962,RIe1e0600_3930,RIe1dd900_3898,RIe1dac00_3866,
        RIe1d7f00_3834,RIe1d2500_3770,RIe1cf800_3738,RIe1ccb00_3706,RIe1c9e00_3674,RIe1c7100_3642,RIe1c4400_3610,RIe1c1700_3578,RIe1bea00_3546,RIfc6bbd0_6248,
        RIfcdd348_7539,RIe1b9438_3485,RIe1b73e0_3462,RIfcab5f0_6972,RIfccbb70_7340,RIe1b5220_3438,RIe1b3e70_3424,RIfc6c9e0_6258,RIfcab488_6971,RIfea7dc0_8226,
        RIe1b0bd0_3388,RIfc6ce18_6261,RIfcabfc8_6979,RIe1ac580_3338,RIe1aaf00_3322,RIe1a8d40_3298,RIe1a6040_3266,RIe1a3340_3234,RIe1a0640_3202,RIe18cb40_2978,
        RIe179040_2754,RIe226998_4729,RIe21b598_4601,RIe204d98_4345,RIe1fedf8_4277,RIe1f81b0_4200,RIe1f0cf8_4117,RIe1d5200_3802,RIe1bbd00_3514,RIe1aeb78_3365,
        RIe1711b0_2664,RIdec5540_709,RIdec2840_677,RIfcc4dc0_7262,RIdebfb40_645,RIfc9d7c0_6814,RIdebce40_613,RIdeba140_581,RIdeb7440_549,RIfc4d978_5905,
        RIdeb1a40_485,RIfc9dbf8_6817,RIdeaed40_453,RIfcb8610_7120,RIdeaa768_421,RIdea3e68_389,RIde9d568_357,RIfc50678_5937,RIfc507e0_5938,RIfc9dec8_6819,
        RIfc853a0_6538,RIde913d0_298,RIde8dc08_281,RIde89a68_261,RIde858c8_241,RIde81a70_222,RIfc84860_6530,RIfc50948_5939,RIfc84c98_6533,RIfcb7da0_7114,
        RIe16b7b0_2600,RIe169b90_2580,RIe167e08_2559,RIe165540_2530,RIe162840_2498,RIee37528_5088,RIe15fb40_2466,RIfcb5be0_7090,RIe15ce40_2434,RIe157440_2370,
        RIe154740_2338,RIfcd35c8_7427,RIe151a40_2306,RIfc53a80_5974,RIe14ed40_2274,RIfcc6170_7276,RIe14c040_2242,RIe149340_2210,RIe146640_2178,RIfc7f130_6468,
        RIee33310_5041,RIfcb4f38_7081,RIfc47f78_5841,RIe140f10_2116,RIdf3ee18_2092,RIdf3cc58_2068,RIdf3a7c8_2042,RIfc7fc70_6476,RIfcd27b8_7417,RIfca1000_6854,
        RIfcc6b48_7283,RIdf35908_1986,RIdf33478_1960,RIfebe9f8_8289,RIdf2f260_1913,RIfcb7968_7111,RIee2a3a0_4939,RIfc51050_5944,RIfcd3fa0_7434,RIdf2a3a0_1857,
        RIdf28078_1832,RIfe81198_7813,RIdf24838_1792,RIfc84428_6527,RIfce7ed8_7661,RIdf22d80_1773,RIfc515f0_5948,RIdf21868_1758,RIdf1f978_1736,RIdf1b058_1684,
        RIdf192d0_1663,RIdf17110_1639,RIdf14410_1607,RIdf11710_1575,RIdf0ea10_1543,RIdf0bd10_1511,RIdf09010_1479,RIdf06310_1447,RIdf03610_1415,RIdefdc10_1351,
        RIdefaf10_1319,RIdef8210_1287,RIdef5510_1255,RIdef2810_1223,RIdeefb10_1191,RIdeece10_1159,RIdeea110_1127,RIfc7e1b8_6457,RIfca19d8_6861,RIfc7dab0_6452,
        RIfc7e488_6459,RIdee49e0_1065,RIfe80d60_7810,RIfeabba0_8270,RIfe80bf8_7809,RIfcb3750_7064,RIfce9f30_7684,RIfc7e5f0_6460,RIfc56a50_6008,RIfe81030_7812,
        RIded7420_913,RIfe80ec8_7811,RIded2f38_864,RIded0940_837,RIdecdc40_805,RIdecaf40_773,RIdec8240_741,RIdeb4740_517,RIde96c68_325,RIe16e348_2631,
        RIe15a140_2402,RIe143940_2146,RIdf38338_2016,RIdf2c998_1884,RIdf1d218_1708,RIdf00910_1383,RIdee7410_1095,RIdedc178_968,RIde7cbb0_198,RIe19d7d8_3169,
        RIe19aad8_3137,RIfcc2d68_7239,RIe197dd8_3105,RIfc5c5b8_6073,RIe1950d8_3073,RIe1923d8_3041,RIe18f6d8_3009,RIe189cd8_2945,RIe186fd8_2913,RIf1438d0_5228,
        RIe1842d8_2881,RIfc5b370_6060,RIe1815d8_2849,RIe17e8d8_2817,RIe17bbd8_2785,RIfcbb748_7155,RIfc59480_6038,RIfcbbce8_7159,RIe175c38_2717,RIfcdb890_7520,
        RIfc59b88_6043,RIfc8ada0_6602,RIfcb5eb0_7092,RIfc57c98_6021,RIfc57158_6013,RIfc58aa8_6031,RIe173910_2692,RIfcc62d8_7277,RIfc8a968_6599,RIfc57428_6015,
        RIfc56d20_6010,RIfc408e0_5760,RIe223b30_4696,RIfc82970_6508,RIe220e30_4664,RIfcecc30_7716,RIe21e130_4632,RIe218730_4568,RIe215a30_4536,RIfc3fad0_5750,
        RIe212d30_4504,RIf169148_5655,RIe210030_4472,RIfc545c0_5982,RIe20d330_4440,RIe20a630_4408,RIe207930_4376,RIfc88d48_6579,RIfc4bec0_5886,RIe202638_4317,
        RIe200b80_4298,RIfc88910_6576,RIfc4c190_5888,RIfc4c2f8_5889,RIfcba398_7141,RIfcd4270_7436,RIfcba0c8_7139,RIe1fcda0_4254,RIe1fbb58_4241,RIfc53d50_5976,
        RIfc9b768_6791,RIfc537b0_5972,RIfc4c5c8_5891,RIfc9e468_6823,RIf157da8_5459,RIfcb9f60_7138,RIe1fa208_4223,RIfc849c8_6531,RIfc529a0_5962,RIfc9f6b0_6836,
        RIe1f5618_4169,RIf153320_5406,RIfcc4988_7259,RIf150d28_5379,RIfebe458_8285,RIfc87f38_6569,RIfcb7f08_7115,RIf14e190_5348,RIfe80658_7805,RIe1eb898_4057,
        RIe1e8b98_4025,RIe1e5e98_3993,RIe1e3198_3961,RIe1e0498_3929,RIe1dd798_3897,RIe1daa98_3865,RIe1d7d98_3833,RIe1d2398_3769,RIe1cf698_3737,RIe1cc998_3705,
        RIe1c9c98_3673,RIe1c6f98_3641,RIe1c4298_3609,RIe1c1598_3577,RIe1be898_3545,RIf14cc78_5333,RIf14ba30_5320,RIe1b92d0_3484,RIe1b7278_3461,RIf14a7e8_5307,
        RIf149ca8_5299,RIfebe5c0_8286,RIfe807c0_7806,RIfc50510_5936,RIfce4f08_7627,RIfe80a90_7808,RIfebe890_8288,RIfc9cde8_6807,RIfc87560_6562,RIfe80928_7807,
        RIfebe728_8287,RIe1a8bd8_3297,RIe1a5ed8_3265,RIe1a31d8_3233,RIe1a04d8_3201,RIe18c9d8_2977,RIe178ed8_2753,RIe226830_4728,RIe21b430_4600,RIe204c30_4344,
        RIe1fec90_4276,RIe1f8048_4199,RIe1f0b90_4116,RIe1d5098_3801,RIe1bbb98_3513,RIe1aea10_3364,RIe171048_2663,RIdec5978_712,RIdec2c78_680,RIfc8aad0_6600,
        RIdebff78_648,RIfc8ac38_6601,RIdebd278_616,RIdeba578_584,RIdeb7878_552,RIfc40e80_5764,RIdeb1e78_488,RIfcdaeb8_7513,RIdeaf178_456,RIee1dbf0_4797,
        RIdeab140_424,RIdea4840_392,RIde9df40_360,RIfc8b070_6604,RIfcc38a8_7247,RIfc807b0_6484,RIfcbb8b0_7156,RIde91a60_300,RIde8e298_283,RIde8a440_264,
        RIde862a0_244,RIde82100_224,RIfcbbb80_7158,RIfc8c150_6616,RIfcbbfb8_7161,RIfc54458_5981,RIe16bbe8_2603,RIfc8c2b8_6617,RIe168240_2562,RIe165978_2533,
        RIe162c78_2501,RIee37960_5091,RIe15ff78_2469,RIfcd6b38_7465,RIe15d278_2437,RIe157878_2373,RIe154b78_2341,RIfc8e5e0_6642,RIe151e78_2309,RIfcb4290_7072,
        RIe14f178_2277,RIfc56ff0_6012,RIe14c478_2245,RIe149778_2213,RIe146a78_2181,RIee346c0_5055,RIee335e0_5043,RIee32398_5030,RIee31420_5019,RIe141348_2119,
        RIe13f020_2094,RIfec16f8_8321,RIdf3a930_2043,RIfce3e28_7615,RIfc56780_6006,RIfcb4128_7071,RIfce2eb0_7604,RIdf35d40_1989,RIfe88218_7893,RIdf316f0_1939,
        RIdf2f698_1916,RIfc7f9a0_6474,RIfce4260_7618,RIfcd62c8_7459,RIfce9990_7680,RIdf2a670_1859,RIdf284b0_1835,RIdf26728_1814,RIdf24c70_1795,RIfc7ecf8_6465,
        RIfcc31a0_7242,RIfc99008_6763,RIfc46e98_5829,RIfce2a78_7601,RIdf1fdb0_1739,RIfcc6e18_7285,RIdf19708_1666,RIdf17548_1642,RIdf14848_1610,RIdf11b48_1578,
        RIdf0ee48_1546,RIdf0c148_1514,RIdf09448_1482,RIdf06748_1450,RIdf03a48_1418,RIdefe048_1354,RIdefb348_1322,RIdef8648_1290,RIdef5948_1258,RIdef2c48_1226,
        RIdeeff48_1194,RIdeed248_1162,RIdeea548_1130,RIfcd9130_7492,RIfc7cb38_6441,RIfc97af0_6748,RIfcb3e58_7069,RIdee4e18_1068,RIdee3090_1047,RIdee0ed0_1023,
        RIfe88380_7894,RIfc97dc0_6750,RIfcc2930_7236,RIfcd9298_7493,RIfc7c868_6439,RIded9ce8_942,RIded76f0_915,RIded5968_894,RIded3370_867,RIded0d78_840,
        RIdece078_808,RIdecb378_776,RIdec8678_744,RIdeb4b78_520,RIde97640_328,RIe16e780_2634,RIe15a578_2405,RIe143d78_2149,RIdf38770_2019,RIdf2cdd0_1887,
        RIdf1d650_1711,RIdf00d48_1386,RIdee7848_1098,RIdedc5b0_971,RIde7d588_201,RIe19dc10_3172,RIe19af10_3140,RIfec1590_8320,RIe198210_3108,RIfec1428_8319,
        RIe195510_3076,RIe192810_3044,RIe18fb10_3012,RIe18a110_2948,RIe187410_2916,RIfec12c0_8318,RIe184710_2884,RIfc88370_6572,RIe181a10_2852,RIe17ed10_2820,
        RIe17c010_2788,RIfc6ccb0_6260,RIfc5f858_6109,RIfca88f0_6940,RIe175f08_2719,RIfc81020_6490,RIfcc6008_7275,RIfc4ea58_5917,RIfc42140_5774,RIfca3b98_6885,
        RIfc5ac68_6055,RIfc984c8_6755,RIe173d48_2695,RIfc9b330_6788,RIf16f688_5727,RIfc42410_5776,RIfc5f588_6107,RIfe880b0_7892,RIe223f68_4699,RIf16bfb0_5688,
        RIe221268_4667,RIfc86cf0_6556,RIe21e568_4635,RIe218b68_4571,RIe215e68_4539,RIfe87de0_7890,RIe213168_4507,RIf1692b0_5656,RIe210468_4475,RIfcdf670_7564,
        RIe20d768_4443,RIe20aa68_4411,RIe207d68_4379,RIfca6460_6914,RIf1662e0_5622,RIe202908_4319,RIfe87b10_7888,RIfc58c10_6032,RIfc50ab0_5940,RIfccd790_7360,
        RIfccd1f0_7356,RIf160610_5556,RIf15e720_5534,RIfe87c78_7889,RIfe87f48_7891,RIfce7668_7655,RIfc86480_6550,RIfcd2218_7413,RIfcb01e0_7026,RIfc47b40_5838,
        RIfc84158_6525,RIfc4b920_5882,RIe1fa4d8_4225,RIfc4ba88_5883,RIfcb7530_7108,RIfcd58f0_7452,RIe1f5a50_4172,RIf153488_5407,RIf151ca0_5390,RIfc51e60_5954,
        RIe1f3728_4147,RIfc9aef8_6785,RIfcbaaa0_7146,RIfc52130_5956,RIe1ee430_4088,RIe1ebcd0_4060,RIe1e8fd0_4028,RIe1e62d0_3996,RIe1e35d0_3964,RIe1e08d0_3932,
        RIe1ddbd0_3900,RIe1daed0_3868,RIe1d81d0_3836,RIe1d27d0_3772,RIe1cfad0_3740,RIe1ccdd0_3708,RIe1ca0d0_3676,RIe1c73d0_3644,RIe1c46d0_3612,RIe1c19d0_3580,
        RIe1becd0_3548,RIfce0b88_7579,RIfc82808_6507,RIe1b9708_3487,RIe1b76b0_3464,RIfcd5bc0_7454,RIfcb69f0_7100,RIe1b54f0_3440,RIe1b4140_3426,RIfc89f90_6592,
        RIfce9af8_7681,RIe1b2958_3409,RIe1b0ea0_3390,RIfc4a138_5865,RIfc8a260_6594,RIe1ac850_3340,RIe1ab1d0_3324,RIe1a9010_3300,RIe1a6310_3268,RIe1a3610_3236,
        RIe1a0910_3204,RIe18ce10_2980,RIe179310_2756,RIe226c68_4731,RIe21b868_4603,RIe205068_4347,RIe1ff0c8_4279,RIe1f8480_4202,RIe1f0fc8_4119,RIe1d54d0_3804,
        RIe1bbfd0_3516,RIe1aee48_3367,RIe171480_2666,RIdec5810_711,RIdec2b10_679,RIfce6f60_7650,RIdebfe10_647,RIfc95228_6719,RIdebd110_615,RIdeba410_583,
        RIdeb7710_551,RIfe879a8_7887,RIdeb1d10_487,RIfcc16e8_7223,RIdeaf010_455,RIfca4f48_6899,RIdeaadf8_423,RIdea44f8_391,RIde9dbf8_359,RIee1cf48_4788,
        RIee1bfd0_4777,RIfc95660_6722,RIfcee148_7731,RIfe87840_7886,RIfe876d8_7885,RIde8a0f8_263,RIde85f58_243,RIfcb0780_7030,RIfcee9b8_7737,RIfc5f150_6104,
        RIfcdee00_7558,RIfcd8050_7480,RIe16ba80_2602,RIfca5380_6902,RIe1680d8_2561,RIe165810_2532,RIe162b10_2500,RIee377f8_5090,RIe15fe10_2468,RIee36448_5076,
        RIe15d110_2436,RIe157710_2372,RIe154a10_2340,RIfc3f3c8_5745,RIe151d10_2308,RIfcde9c8_7555,RIe14f010_2276,RIfc4a2a0_5866,RIe14c310_2244,RIe149610_2212,
        RIe146910_2180,RIfc62288_6139,RIee33478_5042,RIfc71b70_6316,RIee312b8_5018,RIe1411e0_2118,RIfe87570_7884,RIdf3cf28_2070,RIfe87408_7883,RIfcc99b0_7316,
        RIfccf0e0_7378,RIfcaeb60_7010,RIfcca220_7322,RIdf35bd8_1988,RIdf33748_1962,RIdf31588_1938,RIdf2f530_1915,RIee2be58_4958,RIee2a508_4940,RIee28ff0_4925,
        RIee27da8_4912,RIdf2a508_1858,RIdf28348_1834,RIdf265c0_1813,RIdf24b08_1794,RIfc74708_6347,RIfc42578_5777,RIfc43388_5787,RIfc745a0_6346,RIfcb0078_7025,
        RIdf1fc48_1738,RIfcaff10_7024,RIdf195a0_1665,RIdf173e0_1641,RIdf146e0_1609,RIdf119e0_1577,RIdf0ece0_1545,RIdf0bfe0_1513,RIdf092e0_1481,RIdf065e0_1449,
        RIdf038e0_1417,RIdefdee0_1353,RIdefb1e0_1321,RIdef84e0_1289,RIdef57e0_1257,RIdef2ae0_1225,RIdeefde0_1193,RIdeed0e0_1161,RIdeea3e0_1129,RIee257b0_4885,
        RIfca73d8_6925,RIee23e60_4867,RIfce66f0_7644,RIdee4cb0_1067,RIdee2f28_1046,RIdee0d68_1022,RIdeded10_999,RIfcca388_7323,RIfce6858_7645,RIfcceca8_7375,
        RIfcdc970_7532,RIded9b80_941,RIfeaaac0_8258,RIded5800_893,RIded3208_866,RIded0c10_839,RIdecdf10_807,RIdecb210_775,RIdec8510_743,RIdeb4a10_519,
        RIde972f8_327,RIe16e618_2633,RIe15a410_2404,RIe143c10_2148,RIdf38608_2018,RIdf2cc68_1886,RIdf1d4e8_1710,RIdf00be0_1385,RIdee76e0_1097,RIdedc448_970,
        RIde7d240_200,RIe19daa8_3171,RIe19ada8_3139,RIf1457c0_5250,RIe1980a8_3107,RIf1449b0_5240,RIe1953a8_3075,RIe1926a8_3043,RIe18f9a8_3011,RIe189fa8_2947,
        RIe1872a8_2915,RIf143ba0_5230,RIe1845a8_2883,RIfc912e0_6674,RIe1818a8_2851,RIe17eba8_2819,RIe17bea8_2787,RIfc915b0_6676,RIfcbe5b0_7188,RIfce3b58_7613,
        RIe175da0_2718,RIfceb448_7699,RIfcc7958_7293,RIfc42de8_5783,RIfc96e48_6739,RIfc7a810_6416,RIfc96ce0_6738,RIfcc7ac0_7294,RIe173be0_2694,RIfce39f0_7612,
        RIfc7a540_6414,RIfc91b50_6680,RIfc429b0_5780,RIfea9710_8244,RIe223e00_4698,RIfcd8488_7483,RIe221100_4666,RIfc920f0_6684,RIe21e400_4634,RIe218a00_4570,
        RIe215d00_4538,RIfc79e38_6409,RIe213000_4506,RIfcbee20_7194,RIe210300_4474,RIf168068_5643,RIe20d600_4442,RIe20a900_4410,RIe207c00_4378,RIfc5af38_6057,
        RIfcd73a8_7471,RIe2027a0_4318,RIe200ce8_4299,RIfcb2670_7052,RIfcdf940_7566,RIfc5b208_6059,RIfcbf3c0_7198,RIf1604a8_5555,RIf15e5b8_5533,RIfe872a0_7882,
        RIfe87138_7881,RIfc78920_6394,RIfec1158_8317,RIfc93338_6697,RIfcea368_7687,RIfcb23a0_7050,RIfc5bbe0_6066,RIfcede78_7729,RIe1fa370_4224,RIfcd4c48_7443,
        RIfce1dd0_7592,RIfcbf960_7202,RIe1f58e8_4171,RIfcbfc30_7204,RIfc78380_6390,RIfc93770_6700,RIe1f35c0_4146,RIfcb1f68_7047,RIfce1b00_7590,RIfc93a40_6702,
        RIe1ee2c8_4087,RIe1ebb68_4059,RIe1e8e68_4027,RIe1e6168_3995,RIe1e3468_3963,RIe1e0768_3931,RIe1dda68_3899,RIe1dad68_3867,RIe1d8068_3835,RIe1d2668_3771,
        RIe1cf968_3739,RIe1ccc68_3707,RIe1c9f68_3675,RIe1c7268_3643,RIe1c4568_3611,RIe1c1868_3579,RIe1beb68_3547,RIfcdec98_7557,RIfc94148_6707,RIe1b95a0_3486,
        RIe1b7548_3463,RIfcd12a0_7402,RIfceabd8_7693,RIe1b5388_3439,RIe1b3fd8_3425,RIfc94850_6712,RIfcd7c18_7477,RIe1b27f0_3408,RIe1b0d38_3389,RIfc76a30_6372,
        RIfce2640_7598,RIe1ac6e8_3339,RIe1ab068_3323,RIe1a8ea8_3299,RIe1a61a8_3267,RIe1a34a8_3235,RIe1a07a8_3203,RIe18cca8_2979,RIe1791a8_2755,RIe226b00_4730,
        RIe21b700_4602,RIe204f00_4346,RIe1fef60_4278,RIe1f8318_4201,RIe1f0e60_4118,RIe1d5368_3803,RIe1bbe68_3515,RIe1aece0_3366,RIe171318_2665,RIdec5c48_714,
        RIdec2f48_682,RIfc7c160_6434,RIdec0248_650,RIfcb38b8_7065,RIdebd548_618,RIdeba848_586,RIdeb7b48_554,RIfce7c08_7659,RIdeb2148_490,RIfce7aa0_7658,
        RIdeaf448_458,RIfca38c8_6883,RIdeab7d0_426,RIdea4ed0_394,RIde9e5d0_362,RIfc41e70_5772,RIfc5b0a0_6058,RIfcdbb60_7522,RIfc78650_6392,RIfea92d8_8241,
        RIde8e5e0_284,RIfea0d40_8174,RIfea0bd8_8173,RIfcdf508_7563,RIfcb1b30_7044,RIfc5ccc0_6078,RIfcb16f8_7041,RIfc77b10_6384,RIe16beb8_2605,RIe169e60_2582,
        RIe168510_2564,RIe165c48_2535,RIe162f48_2503,RIfc4f9d0_5928,RIe160248_2471,RIfc4e8f0_5916,RIe15d548_2439,RIe157b48_2375,RIe154e48_2343,RIfc4e1e8_5911,
        RIe152148_2311,RIfc868b8_6553,RIe14f448_2279,RIfc865e8_6551,RIe14c748_2247,RIe149a48_2215,RIe146d48_2183,RIfc9eb70_6828,RIfc9ecd8_6829,RIfcc5630_7268,
        RIfc83bb8_6521,RIe141618_2121,RIfea0ea8_8175,RIdf3d1f8_2072,RIdf3ac00_2045,RIee308e0_5011,RIfcd3cd0_7432,RIfc84e00_6534,RIfc834b0_6516,RIdf36010_1991,
        RIdf33a18_1964,RIdf31858_1940,RIdf2f968_1918,RIee2c128_4960,RIee2a7d8_4942,RIee292c0_4927,RIee28078_4914,RIdf2a940_1861,RIdf28780_1837,RIfea0a70_8172,
        RIfea0908_8171,RIfcd4f18_7445,RIfca0628_6847,RIdf23050_1775,RIfcd3190_7424,RIdf21b38_1760,RIdf20080_1741,RIdf1b328_1686,RIdf199d8_1668,RIdf17818_1644,
        RIdf14b18_1612,RIdf11e18_1580,RIdf0f118_1548,RIdf0c418_1516,RIdf09718_1484,RIdf06a18_1452,RIdf03d18_1420,RIdefe318_1356,RIdefb618_1324,RIdef8918_1292,
        RIdef5c18_1260,RIdef2f18_1228,RIdef0218_1196,RIdeed518_1164,RIdeea818_1132,RIfcdf3a0_7562,RIfca5218_6901,RIfcdc538_7529,RIfcdc6a0_7530,RIdee50e8_1070,
        RIdee3360_1049,RIfea07a0_8170,RIdedefe0_1001,RIfcb0d20_7034,RIfcd4978_7441,RIfca49a8_6895,RIfca1708_6859,RIded9fb8_944,RIded79c0_917,RIded5ad0_895,
        RIfeab498_8265,RIded1048_842,RIdece348_810,RIdecb648_778,RIdec8948_746,RIdeb4e48_522,RIde97cd0_330,RIe16ea50_2636,RIe15a848_2407,RIe144048_2151,
        RIdf38a40_2021,RIdf2d0a0_1889,RIdf1d920_1713,RIdf01018_1388,RIdee7b18_1100,RIdedc880_973,RIde7dc18_203,RIe19dee0_3174,RIe19b1e0_3142,RIfc67580_6198,
        RIe1984e0_3110,RIfccb030_7332,RIe1957e0_3078,RIe192ae0_3046,RIe18fde0_3014,RIe18a3e0_2950,RIe1876e0_2918,RIfc6a550_6232,RIe1849e0_2886,RIfcaa7e0_6962,
        RIe181ce0_2854,RIe17efe0_2822,RIe17c2e0_2790,RIfc65d98_6181,RIfc65690_6176,RIe1772b8_2733,RIfea0638_8169,RIfcca928_7327,RIfc607d0_6120,RIfc65258_6173,
        RIee3d798_5158,RIee3c3e8_5144,RIfca9430_6948,RIee39f58_5118,RIe174018_2697,RIfcecf00_7718,RIfc650f0_6172,RIf16e5a8_5715,RIfc43a90_5792,RIfc65528_6175,
        RIe224238_4701,RIfca9f70_6956,RIe221538_4669,RIfc6b4c8_6243,RIe21e838_4637,RIe218e38_4573,RIe216138_4541,RIfc3fda0_5752,RIe213438_4509,RIfc61310_6128,
        RIe210738_4477,RIfc60c08_6123,RIe20da38_4445,RIe20ad38_4413,RIe208038_4381,RIfc66ba8_6191,RIfccbcd8_7341,RIe202bd8_4321,RIe200fb8_4301,RIfcadbe8_6999,
        RIfccbe40_7342,RIfca7540_6926,RIfc6a3e8_6231,RIfca6898_6917,RIfc73358_6333,RIe1fd070_4256,RIe1fbe28_4243,RIfcc2660_7234,RIfc44468_5799,RIf15a940_5490,
        RIfca7270_6924,RIfc5e070_6092,RIfc5dda0_6090,RIfc7e050_6456,RIe1fa7a8_4227,RIfc5d968_6087,RIfcd9568_7495,RIfc8d668_6631,RIe1f5d20_4174,RIfca4138_6889,
        RIfc8cdf8_6625,RIfcc7c28_7295,RIe1f39f8_4149,RIfc99440_6766,RIfcbc3f0_7164,RIfc5a128_6047,RIe1ee700_4090,RIe1ebfa0_4062,RIe1e92a0_4030,RIe1e65a0_3998,
        RIe1e38a0_3966,RIe1e0ba0_3934,RIe1ddea0_3902,RIe1db1a0_3870,RIe1d84a0_3838,RIe1d2aa0_3774,RIe1cfda0_3742,RIe1cd0a0_3710,RIe1ca3a0_3678,RIe1c76a0_3646,
        RIe1c49a0_3614,RIe1c1ca0_3582,RIe1befa0_3550,RIf14cde0_5334,RIf14bb98_5321,RIe1b99d8_3489,RIe1b7980_3466,RIfc4c460_5890,RIfc9e738_6825,RIe1b5658_3441,
        RIfec54d8_8365,RIf149168_5291,RIf147f20_5278,RIe1b2ac0_3410,RIe1b1170_3392,RIf1473e0_5270,RIf1468a0_5262,RIe1acb20_3342,RIe1ab338_3325,RIe1a92e0_3302,
        RIe1a65e0_3270,RIe1a38e0_3238,RIe1a0be0_3206,RIe18d0e0_2982,RIe1795e0_2758,RIe226f38_4733,RIe21bb38_4605,RIe205338_4349,RIe1ff398_4281,RIe1f8750_4204,
        RIe1f1298_4121,RIe1d57a0_3806,RIe1bc2a0_3518,RIe1af118_3369,RIe171750_2668,RIdec5ae0_713,RIdec2de0_681,RIfc82268_6503,RIdec00e0_649,RIfcb8d18_7125,
        RIdebd3e0_617,RIdeba6e0_585,RIdeb79e0_553,RIfcb9858_7133,RIdeb1fe0_489,RIfc9efa8_6831,RIdeaf2e0_457,RIfce0750_7576,RIdeab488_425,RIdea4b88_393,
        RIde9e288_361,RIee1d0b0_4789,RIee1c138_4778,RIfcd0e68_7399,RIfc76d00_6374,RIfe89028_7903,RIfe88d58_7901,RIfe88ec0_7902,RIfe88bf0_7900,RIfcda7b0_7508,
        RIfc4d810_5904,RIfc52dd8_5965,RIfcde590_7552,RIfc4f868_5927,RIe16bd50_2604,RIfc68930_6212,RIe1683a8_2563,RIe165ae0_2534,RIe162de0_2502,RIfe88a88_7899,
        RIe1600e0_2470,RIfcc9140_7310,RIe15d3e0_2438,RIe1579e0_2374,RIe154ce0_2342,RIfc698a8_6223,RIe151fe0_2310,RIee35098_5062,RIe14f2e0_2278,RIfcc0338_7209,
        RIe14c5e0_2246,RIe1498e0_2214,RIe146be0_2182,RIfc88208_6571,RIfc85670_6540,RIfc81f98_6501,RIfcc4f28_7263,RIe1414b0_2120,RIe13f188_2095,RIdf3d090_2071,
        RIdf3aa98_2044,RIfcd2920_7418,RIfc7d7e0_6450,RIfc49760_5858,RIfce5a48_7635,RIdf35ea8_1990,RIdf338b0_1963,RIfe88920_7898,RIdf2f800_1917,RIee2bfc0_4959,
        RIee2a670_4941,RIee29158_4926,RIee27f10_4913,RIdf2a7d8_1860,RIdf28618_1836,RIdf26890_1815,RIdf24dd8_1796,RIfcad918_6997,RIfc69fb0_6228,RIfc63368_6151,
        RIfc623f0_6140,RIfc60938_6121,RIdf1ff18_1740,RIfcba500_7142,RIdf19870_1667,RIdf176b0_1643,RIdf149b0_1611,RIdf11cb0_1579,RIdf0efb0_1547,RIdf0c2b0_1515,
        RIdf095b0_1483,RIdf068b0_1451,RIdf03bb0_1419,RIdefe1b0_1355,RIdefb4b0_1323,RIdef87b0_1291,RIdef5ab0_1259,RIdef2db0_1227,RIdef00b0_1195,RIdeed3b0_1163,
        RIdeea6b0_1131,RIfcc9848_7315,RIfc69a10_6224,RIfcacc70_6988,RIfccbfa8_7343,RIdee4f80_1069,RIdee31f8_1048,RIdee1038_1024,RIdedee78_1000,RIfc84590_6528,
        RIfc9bba0_6794,RIee21b38_4842,RIfc47168_5831,RIded9e50_943,RIded7858_916,RIfe887b8_7897,RIded34d8_868,RIded0ee0_841,RIdece1e0_809,RIdecb4e0_777,
        RIdec87e0_745,RIdeb4ce0_521,RIde97988_329,RIe16e8e8_2635,RIe15a6e0_2406,RIe143ee0_2150,RIdf388d8_2020,RIdf2cf38_1888,RIdf1d7b8_1712,RIdf00eb0_1387,
        RIdee79b0_1099,RIdedc718_972,RIde7d8d0_202,RIe19dd78_3173,RIe19b078_3141,RIfca1438_6857,RIe198378_3109,RIfca35f8_6881,RIe195678_3077,RIe192978_3045,
        RIe18fc78_3013,RIe18a278_2949,RIe187578_2917,RIfcba230_7140,RIe184878_2885,RIf142d90_5220,RIe181b78_2853,RIe17ee78_2821,RIe17c178_2789,RIfc9be70_6796,
        RIfc9bd08_6795,RIfc4ccd0_5896,RIe176070_2720,RIfc87c68_6567,RIfc87b00_6566,RIfcc4c58_7261,RIfc4fca0_5930,RIfc4f598_5925,RIfc876c8_6563,RIfc4dae0_5906,
        RIe173eb0_2696,RIfcb9420_7130,RIfc4e080_5910,RIfc4e350_5912,RIfc9d388_6811,RIfc40a48_5761,RIe2240d0_4700,RIfc85508_6539,RIe2213d0_4668,RIfc9ba38_6793,
        RIe21e6d0_4636,RIe218cd0_4572,RIe215fd0_4540,RIfc52c70_5964,RIe2132d0_4508,RIfca3760_6882,RIe2105d0_4476,RIfc97988_6747,RIe20d8d0_4444,RIe20abd0_4412,
        RIe207ed0_4380,RIfceb5b0_7700,RIfcddbb8_7545,RIe202a70_4320,RIe200e50_4300,RIfc73d30_6340,RIfcaf100_7014,RIfc71468_6311,RIfcdcad8_7533,RIfcdda50_7544,
        RIfca8620_6938,RIe1fcf08_4255,RIe1fbcc0_4242,RIfc6c008_6251,RIfcdd1e0_7538,RIfca9700_6950,RIfca92c8_6947,RIfcce5a0_7370,RIfc6ba68_6247,RIfc6f410_6288,
        RIe1fa640_4226,RIfcce000_7366,RIfc53918_5973,RIfcce708_7371,RIe1f5bb8_4173,RIf1535f0_5408,RIf151e08_5391,RIfc72db8_6329,RIe1f3890_4148,RIf14fc48_5367,
        RIfc72c50_6328,RIfc73e98_6341,RIe1ee598_4089,RIe1ebe38_4061,RIe1e9138_4029,RIe1e6438_3997,RIe1e3738_3965,RIe1e0a38_3933,RIe1ddd38_3901,RIe1db038_3869,
        RIe1d8338_3837,RIe1d2938_3773,RIe1cfc38_3741,RIe1ccf38_3709,RIe1ca238_3677,RIe1c7538_3645,RIe1c4838_3613,RIe1c1b38_3581,RIe1bee38_3549,RIfcb8a48_7123,
        RIfcb84a8_7119,RIe1b9870_3488,RIe1b7818_3465,RIfc85940_6542,RIfc9e198_6821,RIfeac140_8274,RIe1b42a8_3427,RIfc518c0_5950,RIfc838e8_6519,RIfe884e8_7895,
        RIe1b1008_3391,RIfcc5900_7270,RIfc82ad8_6509,RIe1ac9b8_3341,RIfe88650_7896,RIe1a9178_3301,RIe1a6478_3269,RIe1a3778_3237,RIe1a0a78_3205,RIe18cf78_2981,
        RIe179478_2757,RIe226dd0_4732,RIe21b9d0_4604,RIe2051d0_4348,RIe1ff230_4280,RIe1f85e8_4203,RIe1f1130_4120,RIe1d5638_3805,RIe1bc138_3517,RIe1aefb0_3368,
        RIe1715e8_2667,RIdec5f18_716,RIdec3218_684,RIee20350_4825,RIdec0518_652,RIee1f6a8_4816,RIdebd818_620,RIdebab18_588,RIdeb7e18_556,RIfce4da0_7626,
        RIdeb2418_492,RIfcea908_7691,RIdeaf718_460,RIfce20a0_7594,RIdeabe60_428,RIdea5560_396,RIde9ec60_364,RIfce6420_7642,RIee1c2a0_4779,RIfc75950_6360,
        RIee1ad88_4764,RIde920f0_302,RIfea4148_8211,RIfeaa688_8255,RIfea3fe0_8210,RIde82790_226,RIfc6f848_6291,RIfc5dc38_6089,RIfc76b98_6373,RIfcae2f0_7004,
        RIe16c020_2606,RIe16a130_2584,RIe1687e0_2566,RIe165f18_2537,RIe163218_2505,RIfcadd50_7000,RIe160518_2473,RIfc55268_5991,RIe15d818_2441,RIe157e18_2377,
        RIe155118_2345,RIfc45548_5811,RIe152418_2313,RIfc498c8_5859,RIe14f718_2281,RIfcbda70_7180,RIe14ca18_2249,RIe149d18_2217,RIe147018_2185,RIee34828_5056,
        RIee33748_5044,RIee32668_5032,RIee31588_5020,RIe1418e8_2123,RIe13f458_2097,RIdf3d360_2073,RIdf3aed0_2047,RIfc526d0_5960,RIfc42848_5779,RIfcae9f8_7009,
        RIfcb7260_7106,RIfea42b0_8212,RIdf33ce8_1966,RIdf31b28_1942,RIdf2fc38_1920,RIee2c3f8_4962,RIfc4cfa0_5898,RIfc572c0_6014,RIfc4f430_5924,RIfea3e78_8209,
        RIdf28a50_1839,RIdf26b60_1817,RIdf250a8_1798,RIfc9b600_6790,RIfcb9df8_7137,RIdf23320_1777,RIfc86318_6549,RIfeabfd8_8273,RIdf201e8_1742,RIdf1b5f8_1688,
        RIdf19ca8_1670,RIdf17ae8_1646,RIdf14de8_1614,RIdf120e8_1582,RIdf0f3e8_1550,RIdf0c6e8_1518,RIdf099e8_1486,RIdf06ce8_1454,RIdf03fe8_1422,RIdefe5e8_1358,
        RIdefb8e8_1326,RIdef8be8_1294,RIdef5ee8_1262,RIdef31e8_1230,RIdef04e8_1198,RIdeed7e8_1166,RIdeeaae8_1134,RIfc89018_6581,RIfcc54c8_7267,RIfc89180_6582,
        RIfc4b380_5878,RIdee53b8_1072,RIdee34c8_1050,RIfea3d10_8208,RIdedf148_1002,RIfcae188_7003,RIfc4b0b0_5876,RIfc74870_6348,RIfce4968_7623,RIdeda288_946,
        RIded7c90_919,RIded5da0_897,RIded3640_869,RIded1318_844,RIdece618_812,RIdecb918_780,RIdec8c18_748,RIdeb5118_524,RIde98360_332,RIe16ed20_2638,
        RIe15ab18_2409,RIe144318_2153,RIdf38d10_2023,RIdf2d370_1891,RIdf1dbf0_1715,RIdf012e8_1390,RIdee7de8_1102,RIdedcb50_975,RIde7e2a8_205,RIe19e1b0_3176,
        RIe19b4b0_3144,RIfc9cf50_6808,RIe1987b0_3112,RIfc87290_6560,RIe195ab0_3080,RIe192db0_3048,RIe1900b0_3016,RIe18a6b0_2952,RIe1879b0_2920,RIfc842c0_6526,
        RIe184cb0_2888,RIfc83a50_6520,RIe181fb0_2856,RIe17f2b0_2824,RIe17c5b0_2792,RIfc9d0b8_6809,RIfc9e030_6820,RIe177420_2734,RIe176340_2722,RIfc4f700_5926,
        RIfcc4820_7258,RIfc4fb38_5929,RIfce8040_7662,RIee3c6b8_5146,RIee3b308_5132,RIfc812f0_6492,RIe174180_2698,RIfcd3028_7423,RIfc7f400_6470,RIfc46a60_5826,
        RIfc472d0_5832,RIf16cc58_5697,RIe224508_4703,RIfc7d3a8_6447,RIe221808_4671,RIfc97c58_6749,RIe21eb08_4639,RIe219108_4575,RIe216408_4543,RIfcdbe30_7524,
        RIe213708_4511,RIf169580_5658,RIe210a08_4479,RIfca4570_6892,RIe20dd08_4447,RIe20b008_4415,RIe208308_4383,RIfc7b080_6422,RIfc59cf0_6044,RIfea9b48_8247,
        RIfea4418_8213,RIfc79cd0_6408,RIfcd19a8_7407,RIfcc81c8_7299,RIf162230_5576,RIf160778_5557,RIf15e888_5535,RIfea4580_8214,RIfea46e8_8215,RIfc77f48_6387,
        RIfc41fd8_5773,RIf15aaa8_5491,RIfc7c430_6436,RIf159158_5473,RIf157f10_5460,RIfcae890_7008,RIe1faa78_4229,RIfc4a840_5870,RIfc4ed28_5919,RIfce0e58_7581,
        RIe1f5ff0_4176,RIf153758_5409,RIf151f70_5392,RIfccb468_7335,RIe1f3cc8_4151,RIfc68ed0_6216,RIfc6d250_6264,RIfca9ca0_6954,RIe1ee9d0_4092,RIe1ec270_4064,
        RIe1e9570_4032,RIe1e6870_4000,RIe1e3b70_3968,RIe1e0e70_3936,RIe1de170_3904,RIe1db470_3872,RIe1d8770_3840,RIe1d2d70_3776,RIe1d0070_3744,RIe1cd370_3712,
        RIe1ca670_3680,RIe1c7970_3648,RIe1c4c70_3616,RIe1c1f70_3584,RIe1bf270_3552,RIfc784e8_6391,RIfcbef88_7195,RIe1b9ca8_3491,RIe1b7ae8_3467,RIfcc20c0_7230,
        RIfca6190_6912,RIe1b5928_3443,RIe1b4410_3428,RIfcb81d8_7117,RIfcc5090_7264,RIe1b2d90_3412,RIe1b1440_3394,RIfcd5350_7448,RIfcb9588_7131,RIe1acc88_3343,
        RIe1ab4a0_3326,RIe1a95b0_3304,RIe1a68b0_3272,RIe1a3bb0_3240,RIe1a0eb0_3208,RIe18d3b0_2984,RIe1798b0_2760,RIe227208_4735,RIe21be08_4607,RIe205608_4351,
        RIe1ff668_4283,RIe1f8a20_4206,RIe1f1568_4123,RIe1d5a70_3808,RIe1bc570_3520,RIe1af3e8_3371,RIe171a20_2670,RIdec5db0_715,RIdec30b0_683,RIee201e8_4824,
        RIdec03b0_651,RIfcaf538_7017,RIdebd6b0_619,RIdeba9b0_587,RIdeb7cb0_555,RIfc40fe8_5765,RIdeb22b0_491,RIfcd08c8_7395,RIdeaf5b0_459,RIee1dd58_4798,
        RIdeabb18_427,RIdea5218_395,RIde9e918_363,RIee1d218_4790,RIfcedd10_7728,RIfce62b8_7641,RIfcc92a8_7311,RIde91da8_301,RIde8e928_285,RIde8a788_265,
        RIde865e8_245,RIde82448_225,RIfea1448_8179,RIfc750e0_6354,RIfcc19b8_7225,RIfced8d8_7725,RIfec5eb0_8372,RIe169fc8_2583,RIe168678_2565,RIe165db0_2536,
        RIe1630b0_2504,RIfccfc20_7386,RIe1603b0_2472,RIee365b0_5077,RIe15d6b0_2440,RIe157cb0_2376,RIe154fb0_2344,RIfea1718_8181,RIe1522b0_2312,RIee35200_5063,
        RIe14f5b0_2280,RIfcb0348_7027,RIe14c8b0_2248,RIe149bb0_2216,RIe146eb0_2184,RIfc73790_6336,RIfcdf238_7561,RIee32500_5031,RIfc94f58_6717,RIe141780_2122,
        RIe13f2f0_2096,RIfec5be0_8370,RIdf3ad68_2046,RIfea15b0_8180,RIfc5fb28_6111,RIfcae728_7007,RIfc74438_6345,RIdf36178_1992,RIdf33b80_1965,RIdf319c0_1941,
        RIdf2fad0_1919,RIee2c290_4961,RIee2a940_4943,RIfc70658_6301,RIfc704f0_6300,RIdf2aaa8_1862,RIdf288e8_1838,RIdf269f8_1816,RIdf24f40_1797,RIfc64b50_6168,
        RIfccaa90_7328,RIdf231b8_1776,RIfcad4e0_6994,RIdf21ca0_1761,RIfeaad90_8260,RIdf1b490_1687,RIdf19b40_1669,RIdf17980_1645,RIdf14c80_1613,RIdf11f80_1581,
        RIdf0f280_1549,RIdf0c580_1517,RIdf09880_1485,RIdf06b80_1453,RIdf03e80_1421,RIdefe480_1357,RIdefb780_1325,RIdef8a80_1293,RIdef5d80_1261,RIdef3080_1229,
        RIdef0380_1197,RIdeed680_1165,RIdeea980_1133,RIfc595e8_6039,RIfcac568_6983,RIfcccf20_7354,RIfccd358_7357,RIdee5250_1071,RIfea7f28_8227,RIdee11a0_1025,
        RIfea12e0_8178,RIfc679b8_6201,RIee22510_4849,RIfc6dd90_6272,RIfc6cb48_6259,RIdeda120_945,RIded7b28_918,RIded5c38_896,RIfec5d48_8371,RIded11b0_843,
        RIdece4b0_811,RIdecb7b0_779,RIdec8ab0_747,RIdeb4fb0_523,RIde98018_331,RIe16ebb8_2637,RIe15a9b0_2408,RIe1441b0_2152,RIdf38ba8_2022,RIdf2d208_1890,
        RIdf1da88_1714,RIdf01180_1389,RIdee7c80_1101,RIdedc9e8_974,RIde7df60_204,RIe19e048_3175,RIe19b348_3143,RIfcc3ce0_7250,RIe198648_3111,RIfc7efc8_6467,
        RIe195948_3079,RIe192c48_3047,RIe18ff48_3015,RIe18a548_2951,RIe187848_2919,RIfc46790_5824,RIe184b48_2887,RIfc98d38_6761,RIe181e48_2855,RIe17f148_2823,
        RIe17c448_2791,RIfcb5d48_7091,RIfc995a8_6767,RIfc9a3b8_6777,RIe1761d8_2721,RIfc54188_5979,RIfcd2bf0_7420,RIfc8b778_6609,RIfc7dee8_6455,RIee3c550_5145,
        RIfc8c420_6618,RIee3a0c0_5119,RIfeaba38_8269,RIfc46628_5823,RIfcbc288_7163,RIf16e710_5716,RIfc8fdc8_6659,RIfc48c20_5850,RIe2243a0_4702,RIfca0358_6845,
        RIe2216a0_4670,RIfc9a688_6779,RIe21e9a0_4638,RIe218fa0_4574,RIe2162a0_4542,RIfc456b0_5812,RIe2135a0_4510,RIf169418_5657,RIe2108a0_4478,RIfc8bfe8_6615,
        RIe20dba0_4446,RIe20aea0_4414,RIe2081a0_4382,RIfc8c9c0_6622,RIfc7f568_6471,RIe202d40_4322,RIe201120_4302,RIfce2910_7600,RIfc487e8_5847,RIfc46d30_5828,
        RIfc992d8_6765,RIfca2680_6870,RIfc44a08_5803,RIe1fd1d8_4257,RIe1fbf90_4244,RIfc580d0_6024,RIfcbdbd8_7181,RIfc8dd70_6636,RIfce01b0_7572,RIfc7bbc0_6430,
        RIfc90368_6663,RIfc7b8f0_6428,RIe1fa910_4228,RIfcd8b90_7488,RIfc43ec8_5795,RIfc7b788_6427,RIe1f5e88_4175,RIfc7b350_6424,RIfc90d40_6670,RIfca3490_6880,
        RIe1f3b60_4150,RIfc91010_6672,RIfcdb728_7519,RIfcd8758_7485,RIe1ee868_4091,RIe1ec108_4063,RIe1e9408_4031,RIe1e6708_3999,RIe1e3a08_3967,RIe1e0d08_3935,
        RIe1de008_3903,RIe1db308_3871,RIe1d8608_3839,RIe1d2c08_3775,RIe1cff08_3743,RIe1cd208_3711,RIe1ca508_3679,RIe1c7808_3647,RIe1c4b08_3615,RIe1c1e08_3583,
        RIe1bf108_3551,RIf14cf48_5335,RIfc78d58_6397,RIe1b9b40_3490,RIfec5910_8368,RIfc78a88_6395,RIfcd51e8_7447,RIe1b57c0_3442,RIfea1010_8176,RIf1492d0_5292,
        RIfec5a78_8369,RIe1b2c28_3411,RIe1b12d8_3393,RIfec5640_8366,RIf146a08_5263,RIfec57a8_8367,RIfea1178_8177,RIe1a9448_3303,RIe1a6748_3271,RIe1a3a48_3239,
        RIe1a0d48_3207,RIe18d248_2983,RIe179748_2759,RIe2270a0_4734,RIe21bca0_4606,RIe2054a0_4350,RIe1ff500_4282,RIe1f88b8_4205,RIe1f1400_4122,RIe1d5908_3807,
        RIe1bc408_3519,RIe1af280_3370,RIe1718b8_2669,RIdec6350_719,RIdec3650_687,RIfcaf3d0_7016,RIdec0950_655,RIfc6a280_6230,RIdebdc50_623,RIdebaf50_591,
        RIdeb8250_559,RIfc42f50_5784,RIdeb2850_495,RIfc981f8_6753,RIdeafb50_463,RIfc8c6f0_6620,RIdeac838_431,RIdea5f38_399,RIde9f638_367,RIee1d4e8_4792,
        RIfcda648_7507,RIfcc6440_7278,RIfcd5620_7450,RIde92ac8_305,RIfea34a0_8202,RIfea31d0_8200,RIfea3338_8201,RIfcb6b58_7101,RIfcb6888_7099,RIfc9dd60_6818,
        RIee19708_4748,RIfc50c18_5941,RIe16c458_2609,RIfc80a80_6486,RIfec62e8_8375,RIe166350_2540,RIe163650_2508,RIee37d98_5094,RIe160950_2476,RIfcaa678_6961,
        RIe15dc50_2444,RIe158250_2380,RIe155550_2348,RIfea3ba8_8207,RIe152850_2316,RIee35638_5066,RIe14fb50_2284,RIfc62f30_6148,RIe14ce50_2252,RIe14a150_2220,
        RIe147450_2188,RIfc97f28_6751,RIfc89888_6587,RIfc8f558_6653,RIfc52838_5961,RIe141bb8_2125,RIe13f890_2100,RIdf3d798_2076,RIdf3b308_2050,RIee30a48_5012,
        RIfc568e8_6007,RIee2e9f0_4989,RIee2dbe0_4979,RIdf365b0_1995,RIfea38d8_8205,RIfea3a40_8206,RIdf2ff08_1922,RIee2c6c8_4964,RIee2ac10_4945,RIee29590_4929,
        RIee28348_4916,RIdf2ad78_1864,RIdf28e88_1842,RIfea3608_8203,RIfea3770_8204,RIfcc0d10_7216,RIfc75c20_6362,RIfca50b0_6900,RIfc74e10_6352,RIfcc9410_7312,
        RIdf20620_1745,RIfc73628_6335,RIdf1a0e0_1673,RIdf17f20_1649,RIdf15220_1617,RIdf12520_1585,RIdf0f820_1553,RIdf0cb20_1521,RIdf09e20_1489,RIdf07120_1457,
        RIdf04420_1425,RIdefea20_1361,RIdefbd20_1329,RIdef9020_1297,RIdef6320_1265,RIdef3620_1233,RIdef0920_1201,RIdeedc20_1169,RIdeeaf20_1137,RIfcab8c0_6974,
        RIfc7c598_6437,RIfc5beb0_6068,RIfc58ee0_6034,RIdee5688_1074,RIdee3798_1052,RIdee15d8_1028,RIdedf580_1005,RIfcb3048_7059,RIfc72ae8_6327,RIfca3d00_6886,
        RIfcb6450_7096,RIdeda558_948,RIded7f60_921,RIfea3068_8199,RIded3a78_872,RIded1750_847,RIdecea50_815,RIdecbd50_783,RIdec9050_751,RIdeb5550_527,
        RIde98d38_335,RIe16f158_2641,RIe15af50_2412,RIe144750_2156,RIdf39148_2026,RIdf2d7a8_1894,RIdf1e028_1718,RIdf01720_1393,RIdee8220_1105,RIdedcf88_978,
        RIde7ec80_208,RIe19e5e8_3179,RIe19b8e8_3147,RIfca84b8_6937,RIe198be8_3115,RIfc846f8_6529,RIe195ee8_3083,RIe1931e8_3051,RIe1904e8_3019,RIe18aae8_2955,
        RIe187de8_2923,RIfce2be0_7602,RIe1850e8_2891,RIfc8e310_6640,RIe1823e8_2859,RIe17f6e8_2827,RIe17c9e8_2795,RIfcd1570_7404,RIfccc278_7345,RIf1404c8_5191,
        RIfea2d98_8197,RIfcc1b20_7226,RIfc60398_6117,RIee3e5a8_5168,RIee3da68_5160,RIfc642e0_6162,RIfca7f18_6933,RIee3a228_5120,RIfec6180_8374,RIfca9598_6949,
        RIfc5c720_6074,RIfc6bea0_6250,RIfccaec8_7331,RIfc44cd8_5805,RIe224940_4706,RIfcb6180_7094,RIe221c40_4674,RIfc55ad8_5997,RIe21ef40_4642,RIe219540_4578,
        RIe216840_4546,RIfc4dc48_5907,RIe213b40_4514,RIfcdcf10_7536,RIe210e40_4482,RIfcab1b8_6969,RIe20e140_4450,RIe20b440_4418,RIe208740_4386,RIfce3720_7610,
        RIfc64178_6161,RIe203178_4325,RIe201558_4305,RIfcd2ec0_7422,RIf164828_5603,RIfc7f838_6473,RIf162398_5577,RIfcc9c80_7318,RIfca8bc0_6942,RIfea2ac8_8195,
        RIfea2c30_8196,RIfc59318_6037,RIfc4f160_5922,RIf15ac10_5492,RIfcebf88_7707,RIfcbb040_7150,RIfca1870_6860,RIfc93d10_6704,RIe1faeb0_4232,RIf1565c0_5442,
        RIf155a80_5434,RIfc45c50_5816,RIe1f6428_4179,RIfccdbc8_7363,RIfcccae8_7351,RIfca6cd0_6920,RIfec6018_8373,RIfc64010_6160,RIfc434f0_5788,RIfc4c028_5887,
        RIe1eee08_4095,RIe1ec6a8_4067,RIe1e99a8_4035,RIe1e6ca8_4003,RIe1e3fa8_3971,RIe1e12a8_3939,RIe1de5a8_3907,RIe1db8a8_3875,RIe1d8ba8_3843,RIe1d31a8_3779,
        RIe1d04a8_3747,RIe1cd7a8_3715,RIe1caaa8_3683,RIe1c7da8_3651,RIe1c50a8_3619,RIe1c23a8_3587,RIe1bf6a8_3555,RIfc63908_6155,RIfc6bd38_6249,RIe1ba0e0_3494,
        RIe1b7f20_3470,RIfc66fe0_6194,RIfc92ac8_6691,RIe1b5d60_3446,RIfea2f00_8198,RIfc9bfd8_6797,RIfc50d80_5942,RIe1b31c8_3415,RIe1b1878_3397,RIfc4df18_5909,
        RIfc9d658_6813,RIe1ad0c0_3346,RIe1ab8d8_3329,RIe1a99e8_3307,RIe1a6ce8_3275,RIe1a3fe8_3243,RIe1a12e8_3211,RIe18d7e8_2987,RIe179ce8_2763,RIe227640_4738,
        RIe21c240_4610,RIe205a40_4354,RIe1ffaa0_4286,RIe1f8e58_4209,RIe1f19a0_4126,RIe1d5ea8_3811,RIe1bc9a8_3523,RIe1af820_3374,RIe171e58_2673,RIdec61e8_718,
        RIdec34e8_686,RIee20620_4827,RIdec07e8_654,RIfc4b7b8_5881,RIdebdae8_622,RIdebade8_590,RIdeb80e8_558,RIfc41150_5766,RIdeb26e8_494,RIfc87830_6564,
        RIdeaf9e8_462,RIee1dec0_4799,RIdeac4f0_430,RIdea5bf0_398,RIde9f2f0_366,RIee1d380_4791,RIfc77c78_6385,RIfc84f68_6535,RIfc6ff50_6296,RIde92780_304,
        RIde8efb8_287,RIde8ae18_267,RIde86c78_247,RIee1a680_4759,RIee19f78_4754,RIfcd7240_7470,RIfcbeb50_7192,RIfc76328_6367,RIe16c2f0_2608,RIee388d8_5102,
        RIfea20f0_8188,RIe1661e8_2539,RIe1634e8_2507,RIee37c30_5093,RIe1607e8_2475,RIfce7500_7654,RIe15dae8_2443,RIe1580e8_2379,RIe1553e8_2347,RIfc3f698_5747,
        RIe1526e8_2315,RIee354d0_5065,RIe14f9e8_2283,RIfc83e88_6523,RIe14cce8_2251,RIe149fe8_2219,RIe1472e8_2187,RIfcea4d0_7688,RIfcb7ad0_7112,RIfc695d8_6221,
        RIfc51a28_5951,RIe141a50_2124,RIe13f728_2099,RIdf3d630_2075,RIdf3b1a0_2049,RIfca9e08_6955,RIee2fda0_5003,RIfc88a78_6577,RIee2da78_4978,RIdf36448_1994,
        RIdf33fb8_1968,RIdf31df8_1944,RIfea2258_8189,RIee2c560_4963,RIee2aaa8_4944,RIee29428_4928,RIee281e0_4915,RIdf2ac10_1863,RIdf28d20_1841,RIfea27f8_8193,
        RIfea2960_8194,RIfcdabe8_7511,RIfca08f8_6849,RIfc8b1d8_6605,RIfc49058_5853,RIfca0a60_6850,RIdf204b8_1744,RIfc99cb0_6772,RIdf19f78_1672,RIdf17db8_1648,
        RIdf150b8_1616,RIdf123b8_1584,RIdf0f6b8_1552,RIdf0c9b8_1520,RIdf09cb8_1488,RIdf06fb8_1456,RIdf042b8_1424,RIdefe8b8_1360,RIdefbbb8_1328,RIdef8eb8_1296,
        RIdef61b8_1264,RIdef34b8_1232,RIdef07b8_1200,RIdeedab8_1168,RIdeeadb8_1136,RIfcd1f48_7411,RIfc57f68_6023,RIfcbe2e0_7186,RIfcd8fc8_7491,RIdee5520_1073,
        RIfea2690_8192,RIdee1470_1027,RIdedf418_1004,RIfc57b30_6020,RIfcb35e8_7063,RIfcbd7a0_7178,RIfc91178_6673,RIfea2528_8191,RIded7df8_920,RIfea23c0_8190,
        RIded3910_871,RIded15e8_846,RIdece8e8_814,RIdecbbe8_782,RIdec8ee8_750,RIdeb53e8_526,RIde989f0_334,RIe16eff0_2640,RIe15ade8_2411,RIe1445e8_2155,
        RIdf38fe0_2025,RIdf2d640_1893,RIdf1dec0_1717,RIdf015b8_1392,RIdee80b8_1104,RIdedce20_977,RIde7e938_207,RIe19e480_3178,RIe19b780_3146,RIfccc980_7350,
        RIe198a80_3114,RIfcc1148_7219,RIe195d80_3082,RIe193080_3050,RIe190380_3018,RIe18a980_2954,RIe187c80_2922,RIfcb2ee0_7058,RIe184f80_2890,RIfc615e0_6130,
        RIe182280_2858,RIe17f580_2826,RIe17c880_2794,RIfc69038_6217,RIfc4c898_5893,RIfc6f2a8_6287,RIe1764a8_2723,RIfcad0a8_6991,RIfc6adc0_6238,RIfc70388_6299,
        RIfea1b50_8184,RIfea1f88_8187,RIfc56e88_6011,RIfea1cb8_8185,RIe174450_2700,RIfc60d70_6124,RIfc6a820_6234,RIfea1e20_8186,RIf16d798_5705,RIfc40bb0_5762,
        RIe2247d8_4705,RIfc77138_6377,RIe221ad8_4673,RIfcd7d80_7478,RIe21edd8_4641,RIe2193d8_4577,RIe2166d8_4545,RIfc40070_5754,RIe2139d8_4513,RIf169850_5660,
        RIe210cd8_4481,RIfcc1580_7222,RIe20dfd8_4449,RIe20b2d8_4417,RIe2085d8_4385,RIfcd0058_7389,RIfc749d8_6349,RIe203010_4324,RIe2013f0_4304,RIfc60230_6116,
        RIfc60668_6119,RIfcaf970_7020,RIfc45818_5813,RIf160a48_5559,RIf15eb58_5537,RIfea1880_8182,RIfea19e8_8183,RIfc72110_6320,RIfc49b98_5861,RIfcca0b8_7321,
        RIfc71738_6313,RIfc4ca00_5894,RIfc71030_6308,RIfcde428_7551,RIe1fad48_4231,RIfc70bf8_6305,RIfc63a70_6156,RIfca7db0_6932,RIe1f62c0_4178,RIfcada80_6998,
        RIfc6fde8_6295,RIfc6f578_6289,RIe1f3f98_4153,RIfcde158_7549,RIfcad378_6993,RIfc65f00_6182,RIe1eeca0_4094,RIe1ec540_4066,RIe1e9840_4034,RIe1e6b40_4002,
        RIe1e3e40_3970,RIe1e1140_3938,RIe1de440_3906,RIe1db740_3874,RIe1d8a40_3842,RIe1d3040_3778,RIe1d0340_3746,RIe1cd640_3714,RIe1ca940_3682,RIe1c7c40_3650,
        RIe1c4f40_3618,RIe1c2240_3586,RIe1bf540_3554,RIfc69308_6219,RIfccba08_7339,RIe1b9f78_3493,RIe1b7db8_3469,RIfccd628_7359,RIfc69740_6222,RIe1b5bf8_3445,
        RIe1b4578_3429,RIfccf950_7384,RIf148088_5279,RIe1b3060_3414,RIe1b1710_3396,RIfc9f818_6837,RIfcb9c90_7136,RIe1acf58_3345,RIe1ab770_3328,RIe1a9880_3306,
        RIe1a6b80_3274,RIe1a3e80_3242,RIe1a1180_3210,RIe18d680_2986,RIe179b80_2762,RIe2274d8_4737,RIe21c0d8_4609,RIe2058d8_4353,RIe1ff938_4285,RIe1f8cf0_4208,
        RIe1f1838_4125,RIe1d5d40_3810,RIe1bc840_3522,RIe1af6b8_3373,RIe171cf0_2672;
output R_58_102f1b78,R_59_be1fc68,R_5a_10279198,R_5b_102299e8,R_5c_101d0448,R_5d_f7f82f0,R_5e_be21600,R_5f_f7fa5b8,R_60_1027d530,
        R_61_10205ae8,R_62_10283510,R_63_f82b578,R_64_ace4e68,R_65_f8204e0,R_66_1027a0b0,R_67_1022dc30,R_68_102478a8,R_69_10286f78,R_6a_f7edd80,
        R_6b_101c3628,R_6c_f7fbe00,R_6d_f7ce9f8,R_6e_f7c8830,R_6f_101ffc68,R_70_f7d4000,R_71_acee958,R_72_94046c0,R_73_101ee420,R_74_102eb268,
        R_75_b320c50,R_76_ad80a90,R_77_1027fd48,R_78_f7ce4b8,R_79_ad77048,R_7a_102a6ae0,R_7b_f7e4c78,R_7c_e2a6ce0,R_7d_101e86e0,R_7e_e2a9cc8,
        R_7f_10292be0,R_80_b33cde8,R_81_101e2908,R_82_102e9780,R_83_f8157a0,R_84_f819358,R_85_ace8b70,R_86_be142b0,R_87_f81b770,R_88_b330278,
        R_89_f7fe9f8,R_8a_101cf488,R_8b_f8225c0,R_8c_101d4738,R_8d_101c4000,R_8e_101fe960,R_8f_102a0330,R_90_f7f4bd0,R_91_1023e5a8,R_92_10248da8,
        R_93_be2c938,R_94_f7f5458,R_95_f7c6808,R_96_be316a8,R_97_e2a0328,R_98_be2d850,R_99_10217db0,R_9a_f7ec340,R_9b_be23ec0,R_9c_101d4540,
        R_9d_f800828,R_9e_102970c8,R_9f_10221de0,R_a0_ad8d568,R_a1_be4eb58,R_a2_f7c5500,R_a3_ad88f30,R_a4_f82f088,R_a5_f7dcbc8,R_a6_10292940,
        R_a7_be138d8,R_a8_acee418,R_a9_ad84450,R_aa_be10838,R_ab_be31fd8,R_ac_acdaef0,R_ad_acea908,R_ae_101f8830,R_af_f7dec98,R_b0_101e2c50,
        R_b1_f801b30,R_b2_be16e00,R_b3_102e3cf0,R_b4_10291788;

wire \8308 , \8309 , \8310 , \8311 , \8312 , \8313 , \8314 , \8315 , \8316 ,
         \8317 , \8318 , \8319 , \8320 , \8321 , \8322 , \8323 , \8324 , \8325 , \8326 ,
         \8327 , \8328 , \8329 , \8330 , \8331 , \8332 , \8333 , \8334 , \8335 , \8336 ,
         \8337 , \8338 , \8339 , \8340 , \8341 , \8342 , \8343 , \8344 , \8345 , \8346 ,
         \8347 , \8348 , \8349 , \8350 , \8351 , \8352 , \8353 , \8354 , \8355 , \8356 ,
         \8357 , \8358 , \8359 , \8360 , \8361 , \8362 , \8363 , \8364 , \8365 , \8366 ,
         \8367 , \8368 , \8369 , \8370 , \8371 , \8372 , \8373 , \8374 , \8375 , \8376 ,
         \8377 , \8378 , \8379 , \8380 , \8381 , \8382 , \8383 , \8384 , \8385 , \8386 ,
         \8387 , \8388 , \8389 , \8390 , \8391 , \8392 , \8393 , \8394 , \8395 , \8396 ,
         \8397 , \8398 , \8399 , \8400 , \8401 , \8402 , \8403 , \8404 , \8405 , \8406 ,
         \8407 , \8408 , \8409 , \8410 , \8411 , \8412 , \8413 , \8414 , \8415 , \8416 ,
         \8417 , \8418 , \8419 , \8420 , \8421 , \8422 , \8423 , \8424 , \8425 , \8426 ,
         \8427 , \8428 , \8429 , \8430 , \8431 , \8432 , \8433 , \8434 , \8435 , \8436 ,
         \8437 , \8438 , \8439 , \8440 , \8441 , \8442 , \8443 , \8444 , \8445 , \8446 ,
         \8447 , \8448 , \8449 , \8450 , \8451 , \8452 , \8453 , \8454 , \8455 , \8456 ,
         \8457 , \8458 , \8459 , \8460 , \8461 , \8462 , \8463 , \8464 , \8465 , \8466 ,
         \8467 , \8468 , \8469 , \8470 , \8471 , \8472 , \8473 , \8474 , \8475 , \8476 ,
         \8477 , \8478 , \8479 , \8480 , \8481 , \8482 , \8483 , \8484 , \8485 , \8486 ,
         \8487 , \8488 , \8489 , \8490 , \8491 , \8492 , \8493 , \8494 , \8495 , \8496 ,
         \8497 , \8498 , \8499 , \8500 , \8501 , \8502 , \8503 , \8504 , \8505 , \8506 ,
         \8507 , \8508 , \8509 , \8510 , \8511 , \8512 , \8513 , \8514 , \8515 , \8516 ,
         \8517 , \8518 , \8519 , \8520 , \8521 , \8522 , \8523 , \8524 , \8525 , \8526 ,
         \8527 , \8528 , \8529 , \8530 , \8531 , \8532 , \8533 , \8534 , \8535 , \8536 ,
         \8537 , \8538 , \8539 , \8540 , \8541 , \8542 , \8543 , \8544 , \8545 , \8546 ,
         \8547 , \8548 , \8549 , \8550 , \8551 , \8552 , \8553 , \8554 , \8555 , \8556 ,
         \8557 , \8558 , \8559 , \8560 , \8561 , \8562 , \8563 , \8564 , \8565 , \8566 ,
         \8567 , \8568 , \8569 , \8570 , \8571 , \8572 , \8573 , \8574 , \8575 , \8576 ,
         \8577 , \8578 , \8579 , \8580 , \8581 , \8582 , \8583 , \8584 , \8585 , \8586 ,
         \8587 , \8588 , \8589 , \8590 , \8591 , \8592 , \8593 , \8594 , \8595 , \8596 ,
         \8597 , \8598 , \8599 , \8600 , \8601 , \8602 , \8603 , \8604 , \8605 , \8606 ,
         \8607 , \8608 , \8609 , \8610 , \8611 , \8612 , \8613 , \8614 , \8615 , \8616 ,
         \8617 , \8618 , \8619 , \8620 , \8621 , \8622 , \8623 , \8624 , \8625 , \8626 ,
         \8627 , \8628 , \8629 , \8630 , \8631 , \8632 , \8633 , \8634 , \8635 , \8636 ,
         \8637 , \8638 , \8639 , \8640 , \8641 , \8642 , \8643 , \8644 , \8645 , \8646 ,
         \8647 , \8648 , \8649 , \8650 , \8651 , \8652 , \8653 , \8654 , \8655 , \8656 ,
         \8657 , \8658 , \8659 , \8660 , \8661 , \8662 , \8663 , \8664 , \8665 , \8666 ,
         \8667 , \8668 , \8669 , \8670 , \8671 , \8672 , \8673 , \8674 , \8675 , \8676 ,
         \8677 , \8678 , \8679 , \8680 , \8681 , \8682 , \8683 , \8684 , \8685 , \8686 ,
         \8687 , \8688 , \8689 , \8690 , \8691 , \8692 , \8693 , \8694 , \8695 , \8696 ,
         \8697 , \8698 , \8699 , \8700 , \8701 , \8702 , \8703 , \8704 , \8705 , \8706 ,
         \8707 , \8708 , \8709 , \8710 , \8711 , \8712 , \8713 , \8714 , \8715 , \8716 ,
         \8717 , \8718 , \8719 , \8720 , \8721 , \8722 , \8723 , \8724 , \8725 , \8726 ,
         \8727 , \8728 , \8729 , \8730 , \8731 , \8732 , \8733 , \8734 , \8735 , \8736 ,
         \8737 , \8738 , \8739 , \8740 , \8741 , \8742 , \8743 , \8744 , \8745 , \8746 ,
         \8747 , \8748 , \8749 , \8750 , \8751 , \8752 , \8753 , \8754 , \8755 , \8756 ,
         \8757 , \8758 , \8759 , \8760 , \8761 , \8762 , \8763 , \8764 , \8765 , \8766 ,
         \8767 , \8768 , \8769 , \8770 , \8771 , \8772 , \8773 , \8774 , \8775 , \8776 ,
         \8777 , \8778 , \8779 , \8780 , \8781 , \8782 , \8783 , \8784 , \8785 , \8786 ,
         \8787 , \8788 , \8789 , \8790 , \8791 , \8792 , \8793 , \8794 , \8795 , \8796 ,
         \8797 , \8798 , \8799 , \8800 , \8801 , \8802 , \8803 , \8804 , \8805 , \8806 ,
         \8807 , \8808 , \8809 , \8810 , \8811 , \8812 , \8813 , \8814 , \8815 , \8816 ,
         \8817 , \8818 , \8819 , \8820 , \8821 , \8822 , \8823 , \8824 , \8825 , \8826 ,
         \8827 , \8828 , \8829 , \8830 , \8831 , \8832 , \8833 , \8834 , \8835 , \8836 ,
         \8837 , \8838 , \8839 , \8840 , \8841 , \8842 , \8843 , \8844 , \8845 , \8846 ,
         \8847 , \8848 , \8849 , \8850 , \8851 , \8852 , \8853 , \8854 , \8855 , \8856 ,
         \8857 , \8858 , \8859 , \8860 , \8861 , \8862 , \8863 , \8864 , \8865 , \8866 ,
         \8867 , \8868 , \8869 , \8870 , \8871 , \8872 , \8873 , \8874 , \8875 , \8876 ,
         \8877 , \8878 , \8879 , \8880 , \8881 , \8882 , \8883 , \8884 , \8885 , \8886 ,
         \8887 , \8888 , \8889 , \8890 , \8891 , \8892 , \8893 , \8894 , \8895 , \8896 ,
         \8897 , \8898 , \8899 , \8900 , \8901 , \8902 , \8903 , \8904 , \8905 , \8906 ,
         \8907 , \8908 , \8909 , \8910 , \8911 , \8912 , \8913 , \8914 , \8915 , \8916 ,
         \8917 , \8918 , \8919 , \8920 , \8921 , \8922 , \8923 , \8924 , \8925 , \8926 ,
         \8927 , \8928 , \8929 , \8930 , \8931 , \8932 , \8933 , \8934 , \8935 , \8936 ,
         \8937 , \8938 , \8939 , \8940 , \8941 , \8942 , \8943 , \8944 , \8945 , \8946 ,
         \8947 , \8948 , \8949 , \8950 , \8951 , \8952 , \8953 , \8954 , \8955 , \8956 ,
         \8957 , \8958 , \8959 , \8960 , \8961 , \8962 , \8963 , \8964 , \8965 , \8966 ,
         \8967 , \8968 , \8969 , \8970 , \8971 , \8972 , \8973 , \8974 , \8975 , \8976 ,
         \8977 , \8978 , \8979 , \8980 , \8981 , \8982 , \8983 , \8984 , \8985 , \8986 ,
         \8987 , \8988 , \8989 , \8990 , \8991 , \8992 , \8993 , \8994 , \8995 , \8996 ,
         \8997 , \8998 , \8999 , \9000 , \9001 , \9002 , \9003 , \9004 , \9005 , \9006 ,
         \9007 , \9008 , \9009 , \9010 , \9011 , \9012 , \9013 , \9014 , \9015 , \9016 ,
         \9017 , \9018 , \9019 , \9020 , \9021 , \9022 , \9023 , \9024 , \9025 , \9026 ,
         \9027 , \9028 , \9029_N$6 , \9030_N$7 , \9031_N$8 , \9032 , \9033 , \9034 , \9035 , \9036_ZERO ,
         \9037 , \9038 , \9039 , \9040 , \9041 , \9042 , \9043 , \9044 , \9045 , \9046_N$1 ,
         \9047_N$2 , \9048_N$3 , \9049_N$4 , \9050_N$5 , \9051_ONE , \9052 , \9053 , \9054 , \9055 , \9056 ,
         \9057 , \9058 , \9059 , \9060 , \9061 , \9062 , \9063 , \9064 , \9065 , \9066 ,
         \9067 , \9068 , \9069 , \9070 , \9071 , \9072 , \9073 , \9074 , \9075 , \9076 ,
         \9077 , \9078 , \9079 , \9080 , \9081 , \9082 , \9083 , \9084 , \9085 , \9086 ,
         \9087 , \9088 , \9089 , \9090 , \9091 , \9092 , \9093 , \9094 , \9095 , \9096 ,
         \9097 , \9098 , \9099 , \9100 , \9101 , \9102 , \9103 , \9104 , \9105 , \9106 ,
         \9107 , \9108 , \9109 , \9110 , \9111 , \9112 , \9113 , \9114 , \9115 , \9116 ,
         \9117 , \9118 , \9119 , \9120 , \9121 , \9122 , \9123 , \9124 , \9125 , \9126 ,
         \9127 , \9128 , \9129 , \9130 , \9131 , \9132 , \9133 , \9134 , \9135 , \9136 ,
         \9137 , \9138 , \9139 , \9140 , \9141 , \9142 , \9143 , \9144 , \9145 , \9146 ,
         \9147 , \9148 , \9149 , \9150 , \9151 , \9152 , \9153 , \9154 , \9155 , \9156 ,
         \9157 , \9158 , \9159 , \9160 , \9161 , \9162 , \9163 , \9164 , \9165 , \9166 ,
         \9167 , \9168 , \9169 , \9170 , \9171 , \9172 , \9173 , \9174 , \9175 , \9176 ,
         \9177 , \9178 , \9179 , \9180 , \9181 , \9182 , \9183 , \9184 , \9185 , \9186 ,
         \9187 , \9188 , \9189 , \9190 , \9191 , \9192 , \9193 , \9194 , \9195 , \9196 ,
         \9197 , \9198 , \9199 , \9200 , \9201 , \9202 , \9203 , \9204 , \9205 , \9206 ,
         \9207 , \9208 , \9209 , \9210 , \9211 , \9212 , \9213 , \9214 , \9215 , \9216 ,
         \9217 , \9218 , \9219 , \9220 , \9221 , \9222 , \9223 , \9224 , \9225 , \9226 ,
         \9227 , \9228 , \9229 , \9230 , \9231 , \9232 , \9233 , \9234 , \9235 , \9236 ,
         \9237 , \9238 , \9239 , \9240 , \9241 , \9242 , \9243 , \9244 , \9245 , \9246 ,
         \9247 , \9248 , \9249 , \9250 , \9251 , \9252 , \9253 , \9254 , \9255 , \9256 ,
         \9257 , \9258 , \9259 , \9260 , \9261 , \9262 , \9263 , \9264 , \9265 , \9266 ,
         \9267 , \9268 , \9269 , \9270 , \9271 , \9272 , \9273 , \9274 , \9275 , \9276 ,
         \9277 , \9278 , \9279 , \9280 , \9281 , \9282 , \9283 , \9284 , \9285 , \9286 ,
         \9287 , \9288 , \9289 , \9290 , \9291 , \9292 , \9293 , \9294 , \9295 , \9296 ,
         \9297 , \9298 , \9299 , \9300 , \9301 , \9302 , \9303 , \9304 , \9305 , \9306 ,
         \9307 , \9308 , \9309 , \9310 , \9311 , \9312 , \9313 , \9314 , \9315 , \9316 ,
         \9317 , \9318 , \9319 , \9320 , \9321 , \9322 , \9323 , \9324_nG30c1 , \9325 , \9326 ,
         \9327 , \9328 , \9329 , \9330 , \9331 , \9332 , \9333 , \9334 , \9335 , \9336 ,
         \9337 , \9338 , \9339 , \9340 , \9341 , \9342 , \9343 , \9344 , \9345 , \9346 ,
         \9347 , \9348 , \9349 , \9350 , \9351 , \9352 , \9353 , \9354 , \9355 , \9356 ,
         \9357 , \9358 , \9359 , \9360 , \9361 , \9362 , \9363 , \9364 , \9365 , \9366 ,
         \9367 , \9368 , \9369 , \9370 , \9371 , \9372 , \9373 , \9374 , \9375 , \9376 ,
         \9377 , \9378 , \9379 , \9380 , \9381 , \9382 , \9383 , \9384 , \9385 , \9386 ,
         \9387 , \9388 , \9389 , \9390 , \9391 , \9392 , \9393 , \9394 , \9395 , \9396 ,
         \9397 , \9398 , \9399 , \9400 , \9401 , \9402 , \9403 , \9404 , \9405 , \9406 ,
         \9407 , \9408 , \9409 , \9410 , \9411 , \9412 , \9413 , \9414 , \9415 , \9416 ,
         \9417 , \9418 , \9419 , \9420 , \9421 , \9422 , \9423 , \9424 , \9425 , \9426 ,
         \9427 , \9428 , \9429 , \9430 , \9431 , \9432 , \9433 , \9434 , \9435 , \9436 ,
         \9437 , \9438 , \9439 , \9440 , \9441 , \9442 , \9443 , \9444 , \9445 , \9446 ,
         \9447 , \9448 , \9449 , \9450 , \9451 , \9452 , \9453 , \9454 , \9455 , \9456 ,
         \9457 , \9458 , \9459 , \9460 , \9461 , \9462 , \9463 , \9464 , \9465 , \9466 ,
         \9467 , \9468 , \9469 , \9470 , \9471 , \9472 , \9473 , \9474 , \9475 , \9476 ,
         \9477 , \9478 , \9479 , \9480 , \9481 , \9482 , \9483 , \9484 , \9485 , \9486 ,
         \9487 , \9488 , \9489 , \9490 , \9491 , \9492 , \9493 , \9494 , \9495 , \9496 ,
         \9497 , \9498 , \9499 , \9500 , \9501 , \9502 , \9503 , \9504 , \9505 , \9506 ,
         \9507 , \9508 , \9509 , \9510 , \9511 , \9512 , \9513 , \9514 , \9515 , \9516 ,
         \9517 , \9518 , \9519 , \9520 , \9521 , \9522 , \9523 , \9524 , \9525 , \9526 ,
         \9527 , \9528 , \9529 , \9530 , \9531 , \9532 , \9533 , \9534 , \9535 , \9536 ,
         \9537 , \9538 , \9539 , \9540 , \9541 , \9542 , \9543 , \9544 , \9545 , \9546 ,
         \9547 , \9548 , \9549 , \9550 , \9551 , \9552 , \9553 , \9554 , \9555 , \9556 ,
         \9557 , \9558 , \9559 , \9560 , \9561 , \9562 , \9563 , \9564 , \9565 , \9566 ,
         \9567 , \9568 , \9569 , \9570 , \9571 , \9572 , \9573 , \9574 , \9575 , \9576 ,
         \9577 , \9578 , \9579 , \9580 , \9581 , \9582 , \9583 , \9584 , \9585 , \9586 ,
         \9587 , \9588 , \9589 , \9590 , \9591 , \9592 , \9593 , \9594 , \9595 , \9596 ,
         \9597 , \9598_nG41ee , \9599 , \9600 , \9601 , \9602 , \9603 , \9604 , \9605 , \9606 ,
         \9607 , \9608 , \9609 , \9610 , \9611 , \9612 , \9613 , \9614 , \9615 , \9616 ,
         \9617 , \9618 , \9619 , \9620 , \9621 , \9622 , \9623 , \9624 , \9625 , \9626 ,
         \9627 , \9628 , \9629 , \9630 , \9631 , \9632 , \9633 , \9634 , \9635 , \9636 ,
         \9637 , \9638 , \9639 , \9640 , \9641 , \9642 , \9643 , \9644 , \9645 , \9646 ,
         \9647 , \9648 , \9649 , \9650 , \9651 , \9652 , \9653 , \9654 , \9655 , \9656 ,
         \9657 , \9658 , \9659 , \9660 , \9661 , \9662 , \9663 , \9664 , \9665 , \9666 ,
         \9667 , \9668 , \9669 , \9670 , \9671 , \9672 , \9673 , \9674 , \9675 , \9676 ,
         \9677 , \9678 , \9679 , \9680 , \9681 , \9682 , \9683 , \9684 , \9685 , \9686 ,
         \9687 , \9688 , \9689 , \9690 , \9691 , \9692 , \9693 , \9694 , \9695 , \9696 ,
         \9697 , \9698 , \9699 , \9700 , \9701 , \9702 , \9703 , \9704 , \9705 , \9706 ,
         \9707 , \9708 , \9709 , \9710 , \9711 , \9712 , \9713 , \9714 , \9715 , \9716 ,
         \9717 , \9718 , \9719 , \9720 , \9721 , \9722 , \9723 , \9724 , \9725 , \9726 ,
         \9727 , \9728 , \9729 , \9730 , \9731 , \9732_nG3146 , \9733 , \9734 , \9735 , \9736 ,
         \9737 , \9738 , \9739 , \9740 , \9741 , \9742 , \9743 , \9744 , \9745 , \9746 ,
         \9747 , \9748 , \9749 , \9750 , \9751 , \9752 , \9753 , \9754 , \9755 , \9756 ,
         \9757 , \9758 , \9759 , \9760 , \9761 , \9762 , \9763 , \9764 , \9765 , \9766 ,
         \9767 , \9768 , \9769 , \9770 , \9771 , \9772 , \9773 , \9774 , \9775 , \9776 ,
         \9777 , \9778 , \9779 , \9780 , \9781 , \9782 , \9783 , \9784 , \9785 , \9786 ,
         \9787 , \9788 , \9789 , \9790 , \9791 , \9792 , \9793 , \9794 , \9795 , \9796 ,
         \9797 , \9798 , \9799 , \9800 , \9801 , \9802 , \9803 , \9804 , \9805 , \9806 ,
         \9807 , \9808 , \9809 , \9810 , \9811 , \9812 , \9813 , \9814 , \9815 , \9816 ,
         \9817 , \9818 , \9819 , \9820 , \9821 , \9822 , \9823 , \9824 , \9825 , \9826 ,
         \9827 , \9828 , \9829 , \9830 , \9831 , \9832 , \9833 , \9834 , \9835 , \9836 ,
         \9837 , \9838 , \9839 , \9840 , \9841 , \9842 , \9843 , \9844 , \9845 , \9846 ,
         \9847 , \9848 , \9849 , \9850 , \9851 , \9852 , \9853 , \9854 , \9855 , \9856 ,
         \9857 , \9858 , \9859 , \9860 , \9861 , \9862 , \9863 , \9864 , \9865_nG4273 , \9866 ,
         \9867 , \9868 , \9869 , \9870 , \9871 , \9872 , \9873 , \9874 , \9875 , \9876 ,
         \9877 , \9878 , \9879 , \9880 , \9881 , \9882 , \9883 , \9884 , \9885 , \9886 ,
         \9887 , \9888 , \9889 , \9890 , \9891 , \9892 , \9893 , \9894 , \9895 , \9896 ,
         \9897 , \9898 , \9899 , \9900 , \9901 , \9902 , \9903 , \9904 , \9905 , \9906 ,
         \9907 , \9908 , \9909 , \9910 , \9911 , \9912 , \9913 , \9914 , \9915 , \9916 ,
         \9917 , \9918 , \9919 , \9920 , \9921 , \9922 , \9923 , \9924 , \9925 , \9926 ,
         \9927 , \9928 , \9929 , \9930 , \9931 , \9932 , \9933 , \9934 , \9935 , \9936 ,
         \9937 , \9938 , \9939 , \9940 , \9941 , \9942 , \9943 , \9944 , \9945 , \9946 ,
         \9947 , \9948 , \9949 , \9950 , \9951 , \9952 , \9953 , \9954 , \9955 , \9956 ,
         \9957 , \9958 , \9959 , \9960 , \9961 , \9962 , \9963 , \9964 , \9965 , \9966 ,
         \9967 , \9968 , \9969 , \9970 , \9971 , \9972 , \9973 , \9974 , \9975 , \9976 ,
         \9977 , \9978 , \9979 , \9980 , \9981 , \9982 , \9983 , \9984 , \9985 , \9986 ,
         \9987 , \9988 , \9989 , \9990 , \9991 , \9992 , \9993 , \9994 , \9995 , \9996 ,
         \9997 , \9998 , \9999_nG31cb , \10000 , \10001 , \10002 , \10003 , \10004 , \10005 , \10006 ,
         \10007 , \10008 , \10009 , \10010 , \10011 , \10012 , \10013 , \10014 , \10015 , \10016 ,
         \10017 , \10018 , \10019 , \10020 , \10021 , \10022 , \10023 , \10024 , \10025 , \10026 ,
         \10027 , \10028 , \10029 , \10030 , \10031 , \10032 , \10033 , \10034 , \10035 , \10036 ,
         \10037 , \10038 , \10039 , \10040 , \10041 , \10042 , \10043 , \10044 , \10045 , \10046 ,
         \10047 , \10048 , \10049 , \10050 , \10051 , \10052 , \10053 , \10054 , \10055 , \10056 ,
         \10057 , \10058 , \10059 , \10060 , \10061 , \10062 , \10063 , \10064 , \10065 , \10066 ,
         \10067 , \10068 , \10069 , \10070 , \10071 , \10072 , \10073 , \10074 , \10075 , \10076 ,
         \10077 , \10078 , \10079 , \10080 , \10081 , \10082 , \10083 , \10084 , \10085 , \10086 ,
         \10087 , \10088 , \10089 , \10090 , \10091 , \10092 , \10093 , \10094 , \10095 , \10096 ,
         \10097 , \10098 , \10099 , \10100 , \10101 , \10102 , \10103 , \10104 , \10105 , \10106 ,
         \10107 , \10108 , \10109 , \10110 , \10111 , \10112 , \10113 , \10114 , \10115 , \10116 ,
         \10117 , \10118 , \10119 , \10120 , \10121 , \10122 , \10123 , \10124 , \10125 , \10126 ,
         \10127 , \10128 , \10129 , \10130 , \10131 , \10132_nG42f8 , \10133 , \10134 , \10135 , \10136 ,
         \10137 , \10138 , \10139 , \10140 , \10141 , \10142 , \10143 , \10144 , \10145 , \10146 ,
         \10147 , \10148 , \10149 , \10150 , \10151 , \10152 , \10153 , \10154 , \10155 , \10156 ,
         \10157 , \10158 , \10159 , \10160 , \10161 , \10162 , \10163 , \10164 , \10165 , \10166 ,
         \10167 , \10168 , \10169 , \10170 , \10171 , \10172 , \10173 , \10174 , \10175 , \10176 ,
         \10177 , \10178 , \10179 , \10180 , \10181 , \10182 , \10183 , \10184 , \10185 , \10186 ,
         \10187 , \10188 , \10189 , \10190 , \10191 , \10192 , \10193 , \10194 , \10195 , \10196 ,
         \10197 , \10198 , \10199 , \10200 , \10201 , \10202 , \10203 , \10204 , \10205 , \10206 ,
         \10207 , \10208 , \10209 , \10210 , \10211 , \10212 , \10213 , \10214 , \10215 , \10216 ,
         \10217 , \10218 , \10219 , \10220 , \10221 , \10222 , \10223 , \10224 , \10225 , \10226 ,
         \10227 , \10228 , \10229 , \10230 , \10231 , \10232 , \10233 , \10234 , \10235 , \10236 ,
         \10237 , \10238 , \10239 , \10240 , \10241 , \10242 , \10243 , \10244 , \10245 , \10246 ,
         \10247 , \10248 , \10249 , \10250 , \10251 , \10252 , \10253 , \10254 , \10255 , \10256 ,
         \10257 , \10258 , \10259 , \10260 , \10261 , \10262 , \10263 , \10264 , \10265 , \10266_nG3250 ,
         \10267 , \10268 , \10269 , \10270 , \10271 , \10272 , \10273 , \10274 , \10275 , \10276 ,
         \10277 , \10278 , \10279 , \10280 , \10281 , \10282 , \10283 , \10284 , \10285 , \10286 ,
         \10287 , \10288 , \10289 , \10290 , \10291 , \10292 , \10293 , \10294 , \10295 , \10296 ,
         \10297 , \10298 , \10299 , \10300 , \10301 , \10302 , \10303 , \10304 , \10305 , \10306 ,
         \10307 , \10308 , \10309 , \10310 , \10311 , \10312 , \10313 , \10314 , \10315 , \10316 ,
         \10317 , \10318 , \10319 , \10320 , \10321 , \10322 , \10323 , \10324 , \10325 , \10326 ,
         \10327 , \10328 , \10329 , \10330 , \10331 , \10332 , \10333 , \10334 , \10335 , \10336 ,
         \10337 , \10338 , \10339 , \10340 , \10341 , \10342 , \10343 , \10344 , \10345 , \10346 ,
         \10347 , \10348 , \10349 , \10350 , \10351 , \10352 , \10353 , \10354 , \10355 , \10356 ,
         \10357 , \10358 , \10359 , \10360 , \10361 , \10362 , \10363 , \10364 , \10365 , \10366 ,
         \10367 , \10368 , \10369 , \10370 , \10371 , \10372 , \10373 , \10374 , \10375 , \10376 ,
         \10377 , \10378 , \10379 , \10380 , \10381 , \10382 , \10383 , \10384 , \10385 , \10386 ,
         \10387 , \10388 , \10389 , \10390 , \10391 , \10392 , \10393 , \10394 , \10395 , \10396 ,
         \10397 , \10398 , \10399_nG437d , \10400 , \10401 , \10402 , \10403 , \10404 , \10405 , \10406 ,
         \10407 , \10408 , \10409_nG444e , \10410 , \10411 , \10412_nG4451 , \10413 , \10414 , \10415_nG4454 , \10416 ,
         \10417 , \10418 , \10419 , \10420 , \10421 , \10422 , \10423 , \10424 , \10425 , \10426 ,
         \10427 , \10428 , \10429 , \10430 , \10431 , \10432 , \10433 , \10434 , \10435 , \10436 ,
         \10437 , \10438 , \10439 , \10440 , \10441 , \10442 , \10443 , \10444 , \10445 , \10446 ,
         \10447 , \10448 , \10449 , \10450 , \10451 , \10452 , \10453 , \10454 , \10455 , \10456 ,
         \10457 , \10458 , \10459 , \10460 , \10461 , \10462 , \10463 , \10464 , \10465 , \10466 ,
         \10467 , \10468 , \10469 , \10470 , \10471 , \10472 , \10473 , \10474 , \10475 , \10476 ,
         \10477 , \10478 , \10479 , \10480 , \10481 , \10482 , \10483 , \10484 , \10485 , \10486 ,
         \10487 , \10488 , \10489 , \10490 , \10491 , \10492 , \10493 , \10494 , \10495 , \10496 ,
         \10497 , \10498 , \10499 , \10500 , \10501 , \10502 , \10503 , \10504 , \10505 , \10506 ,
         \10507 , \10508 , \10509 , \10510 , \10511 , \10512 , \10513 , \10514 , \10515 , \10516 ,
         \10517 , \10518 , \10519 , \10520 , \10521 , \10522 , \10523 , \10524 , \10525 , \10526 ,
         \10527 , \10528 , \10529 , \10530 , \10531 , \10532 , \10533 , \10534 , \10535 , \10536 ,
         \10537 , \10538 , \10539 , \10540 , \10541 , \10542 , \10543 , \10544 , \10545 , \10546 ,
         \10547 , \10548 , \10549 , \10550 , \10551 , \10552 , \10553_nG6577 , \10554 , \10555 , \10556 ,
         \10557 , \10558 , \10559 , \10560 , \10561 , \10562 , \10563 , \10564 , \10565 , \10566 ,
         \10567 , \10568 , \10569 , \10570 , \10571 , \10572 , \10573 , \10574 , \10575 , \10576 ,
         \10577 , \10578 , \10579 , \10580 , \10581 , \10582 , \10583 , \10584 , \10585 , \10586 ,
         \10587 , \10588 , \10589 , \10590 , \10591 , \10592 , \10593 , \10594 , \10595 , \10596 ,
         \10597 , \10598 , \10599 , \10600 , \10601 , \10602 , \10603 , \10604 , \10605 , \10606 ,
         \10607 , \10608 , \10609 , \10610 , \10611 , \10612 , \10613 , \10614 , \10615 , \10616 ,
         \10617 , \10618 , \10619 , \10620 , \10621 , \10622 , \10623 , \10624 , \10625 , \10626 ,
         \10627 , \10628 , \10629 , \10630 , \10631 , \10632 , \10633 , \10634 , \10635 , \10636 ,
         \10637 , \10638 , \10639 , \10640 , \10641 , \10642 , \10643 , \10644 , \10645 , \10646 ,
         \10647 , \10648 , \10649 , \10650 , \10651 , \10652 , \10653 , \10654 , \10655 , \10656 ,
         \10657 , \10658 , \10659 , \10660 , \10661 , \10662 , \10663 , \10664 , \10665 , \10666 ,
         \10667 , \10668 , \10669 , \10670 , \10671 , \10672 , \10673 , \10674 , \10675 , \10676 ,
         \10677 , \10678 , \10679 , \10680 , \10681 , \10682 , \10683 , \10684 , \10685_nG6578 , \10686_nG6579 ,
         \10687 , \10688_nG44da , \10689_nG455e , \10690_nG455f , \10691 , \10692 , \10693 , \10694_nG9c0e , \10695 , \10696 ,
         \10697 , \10698 , \10699 , \10700 , \10701 , \10702_nG4456 , \10703 , \10704 , \10705 , \10706 ,
         \10707 , \10708 , \10709 , \10710 , \10711 , \10712 , \10713 , \10714 , \10715 , \10716 ,
         \10717 , \10718 , \10719 , \10720 , \10721 , \10722 , \10723 , \10724 , \10725 , \10726 ,
         \10727 , \10728 , \10729 , \10730 , \10731 , \10732 , \10733 , \10734 , \10735 , \10736 ,
         \10737 , \10738 , \10739 , \10740 , \10741 , \10742 , \10743 , \10744 , \10745 , \10746 ,
         \10747 , \10748 , \10749 , \10750 , \10751 , \10752 , \10753 , \10754 , \10755 , \10756 ,
         \10757 , \10758 , \10759 , \10760 , \10761 , \10762 , \10763 , \10764 , \10765 , \10766 ,
         \10767 , \10768 , \10769 , \10770 , \10771 , \10772 , \10773 , \10774 , \10775 , \10776 ,
         \10777 , \10778 , \10779 , \10780 , \10781 , \10782 , \10783 , \10784 , \10785 , \10786 ,
         \10787 , \10788 , \10789 , \10790 , \10791 , \10792 , \10793 , \10794 , \10795 , \10796 ,
         \10797 , \10798 , \10799 , \10800 , \10801 , \10802 , \10803 , \10804 , \10805 , \10806 ,
         \10807 , \10808 , \10809 , \10810 , \10811 , \10812 , \10813 , \10814 , \10815 , \10816 ,
         \10817 , \10818 , \10819 , \10820 , \10821 , \10822 , \10823 , \10824 , \10825 , \10826 ,
         \10827 , \10828 , \10829 , \10830 , \10831 , \10832 , \10833 , \10834 , \10835 , \10836 ,
         \10837 , \10838 , \10839 , \10840 , \10841 , \10842 , \10843 , \10844 , \10845 , \10846_nG45e3 ,
         \10847 , \10848 , \10849 , \10850 , \10851 , \10852 , \10853 , \10854 , \10855 , \10856 ,
         \10857 , \10858 , \10859 , \10860 , \10861 , \10862 , \10863 , \10864 , \10865 , \10866 ,
         \10867 , \10868 , \10869 , \10870 , \10871 , \10872 , \10873 , \10874 , \10875 , \10876 ,
         \10877 , \10878 , \10879 , \10880 , \10881 , \10882 , \10883 , \10884 , \10885 , \10886 ,
         \10887 , \10888 , \10889 , \10890 , \10891 , \10892 , \10893 , \10894 , \10895 , \10896 ,
         \10897 , \10898 , \10899 , \10900 , \10901 , \10902 , \10903 , \10904 , \10905 , \10906 ,
         \10907 , \10908 , \10909 , \10910 , \10911 , \10912 , \10913 , \10914 , \10915 , \10916 ,
         \10917 , \10918 , \10919 , \10920 , \10921 , \10922 , \10923 , \10924 , \10925 , \10926 ,
         \10927 , \10928 , \10929 , \10930 , \10931 , \10932 , \10933 , \10934 , \10935 , \10936 ,
         \10937 , \10938 , \10939 , \10940 , \10941 , \10942 , \10943 , \10944 , \10945 , \10946 ,
         \10947 , \10948 , \10949 , \10950 , \10951 , \10952 , \10953 , \10954 , \10955 , \10956 ,
         \10957 , \10958 , \10959 , \10960 , \10961 , \10962 , \10963 , \10964 , \10965 , \10966 ,
         \10967 , \10968 , \10969 , \10970 , \10971 , \10972 , \10973 , \10974 , \10975 , \10976 ,
         \10977 , \10978_nG4667 , \10979_nG4668 , \10980 , \10981 , \10982 , \10983 , \10984 , \10985_nG657a , \10986_nG657b ,
         \10987_nG657c , \10988 , \10989 , \10990 , \10991 , \10992 , \10993 , \10994 , \10995_nG9c0b , \10996 ,
         \10997 , \10998 , \10999 , \11000 , \11001 , \11002 , \11003 , \11004 , \11005 , \11006 ,
         \11007 , \11008 , \11009 , \11010 , \11011 , \11012 , \11013 , \11014 , \11015 , \11016 ,
         \11017 , \11018 , \11019 , \11020 , \11021 , \11022 , \11023 , \11024 , \11025 , \11026 ,
         \11027 , \11028 , \11029 , \11030 , \11031 , \11032 , \11033 , \11034 , \11035 , \11036 ,
         \11037 , \11038 , \11039 , \11040 , \11041 , \11042 , \11043 , \11044 , \11045 , \11046 ,
         \11047 , \11048 , \11049 , \11050 , \11051 , \11052 , \11053 , \11054 , \11055 , \11056 ,
         \11057 , \11058 , \11059 , \11060 , \11061 , \11062 , \11063 , \11064 , \11065 , \11066 ,
         \11067 , \11068 , \11069 , \11070 , \11071 , \11072 , \11073 , \11074 , \11075 , \11076 ,
         \11077 , \11078 , \11079 , \11080 , \11081 , \11082 , \11083 , \11084 , \11085 , \11086 ,
         \11087 , \11088 , \11089 , \11090 , \11091 , \11092 , \11093 , \11094 , \11095 , \11096 ,
         \11097 , \11098 , \11099 , \11100 , \11101 , \11102 , \11103 , \11104 , \11105 , \11106 ,
         \11107 , \11108 , \11109 , \11110 , \11111 , \11112 , \11113 , \11114 , \11115 , \11116 ,
         \11117 , \11118 , \11119 , \11120 , \11121 , \11122 , \11123 , \11124 , \11125 , \11126 ,
         \11127 , \11128 , \11129 , \11130 , \11131 , \11132 , \11133 , \11134 , \11135 , \11136_nG657d ,
         \11137 , \11138 , \11139 , \11140 , \11141 , \11142 , \11143 , \11144 , \11145 , \11146 ,
         \11147 , \11148 , \11149 , \11150 , \11151 , \11152 , \11153 , \11154 , \11155 , \11156 ,
         \11157 , \11158 , \11159 , \11160 , \11161 , \11162 , \11163 , \11164 , \11165 , \11166 ,
         \11167 , \11168 , \11169 , \11170 , \11171 , \11172 , \11173 , \11174 , \11175 , \11176 ,
         \11177 , \11178 , \11179 , \11180 , \11181 , \11182 , \11183 , \11184 , \11185 , \11186 ,
         \11187 , \11188 , \11189 , \11190 , \11191 , \11192 , \11193 , \11194 , \11195 , \11196 ,
         \11197 , \11198 , \11199 , \11200 , \11201 , \11202 , \11203 , \11204 , \11205 , \11206 ,
         \11207 , \11208 , \11209 , \11210 , \11211 , \11212 , \11213 , \11214 , \11215 , \11216 ,
         \11217 , \11218 , \11219 , \11220 , \11221 , \11222 , \11223 , \11224 , \11225 , \11226 ,
         \11227 , \11228 , \11229 , \11230 , \11231 , \11232 , \11233 , \11234 , \11235 , \11236 ,
         \11237 , \11238 , \11239 , \11240 , \11241 , \11242 , \11243 , \11244 , \11245 , \11246 ,
         \11247 , \11248 , \11249 , \11250 , \11251 , \11252 , \11253 , \11254 , \11255 , \11256 ,
         \11257 , \11258 , \11259 , \11260 , \11261 , \11262 , \11263 , \11264 , \11265 , \11266 ,
         \11267 , \11268_nG657e , \11269_nG657f , \11270 , \11271 , \11272 , \11273 , \11274_nG46ec , \11275_nG4770 , \11276_nG4771 ,
         \11277 , \11278 , \11279 , \11280 , \11281 , \11282 , \11283_nG9c08 , \11284 , \11285 , \11286 ,
         \11287 , \11288 , \11289 , \11290 , \11291 , \11292 , \11293 , \11294 , \11295 , \11296 ,
         \11297 , \11298 , \11299 , \11300 , \11301 , \11302 , \11303 , \11304 , \11305 , \11306 ,
         \11307 , \11308 , \11309 , \11310 , \11311 , \11312 , \11313 , \11314 , \11315 , \11316 ,
         \11317 , \11318 , \11319 , \11320 , \11321 , \11322 , \11323 , \11324 , \11325 , \11326 ,
         \11327 , \11328 , \11329 , \11330 , \11331 , \11332 , \11333 , \11334 , \11335 , \11336 ,
         \11337 , \11338 , \11339 , \11340 , \11341 , \11342 , \11343 , \11344 , \11345 , \11346 ,
         \11347 , \11348 , \11349 , \11350 , \11351 , \11352 , \11353 , \11354 , \11355 , \11356 ,
         \11357 , \11358 , \11359 , \11360 , \11361 , \11362 , \11363 , \11364 , \11365 , \11366 ,
         \11367 , \11368 , \11369 , \11370 , \11371 , \11372 , \11373 , \11374 , \11375 , \11376 ,
         \11377 , \11378 , \11379 , \11380 , \11381 , \11382 , \11383 , \11384 , \11385 , \11386 ,
         \11387 , \11388 , \11389 , \11390 , \11391 , \11392 , \11393 , \11394 , \11395 , \11396 ,
         \11397 , \11398 , \11399 , \11400 , \11401 , \11402 , \11403 , \11404 , \11405 , \11406 ,
         \11407 , \11408 , \11409 , \11410 , \11411 , \11412 , \11413 , \11414 , \11415 , \11416 ,
         \11417 , \11418 , \11419 , \11420 , \11421 , \11422 , \11423 , \11424 , \11425 , \11426 ,
         \11427 , \11428 , \11429 , \11430 , \11431 , \11432 , \11433 , \11434 , \11435 , \11436 ,
         \11437_nG47f5 , \11438 , \11439 , \11440 , \11441 , \11442 , \11443 , \11444 , \11445 , \11446 ,
         \11447 , \11448 , \11449 , \11450 , \11451 , \11452 , \11453 , \11454 , \11455 , \11456 ,
         \11457 , \11458 , \11459 , \11460 , \11461 , \11462 , \11463 , \11464 , \11465 , \11466 ,
         \11467 , \11468 , \11469 , \11470 , \11471 , \11472 , \11473 , \11474 , \11475 , \11476 ,
         \11477 , \11478 , \11479 , \11480 , \11481 , \11482 , \11483 , \11484 , \11485 , \11486 ,
         \11487 , \11488 , \11489 , \11490 , \11491 , \11492 , \11493 , \11494 , \11495 , \11496 ,
         \11497 , \11498 , \11499 , \11500 , \11501 , \11502 , \11503 , \11504 , \11505 , \11506 ,
         \11507 , \11508 , \11509 , \11510 , \11511 , \11512 , \11513 , \11514 , \11515 , \11516 ,
         \11517 , \11518 , \11519 , \11520 , \11521 , \11522 , \11523 , \11524 , \11525 , \11526 ,
         \11527 , \11528 , \11529 , \11530 , \11531 , \11532 , \11533 , \11534 , \11535 , \11536 ,
         \11537 , \11538 , \11539 , \11540 , \11541 , \11542 , \11543 , \11544 , \11545 , \11546 ,
         \11547 , \11548 , \11549 , \11550 , \11551 , \11552 , \11553 , \11554 , \11555 , \11556 ,
         \11557 , \11558 , \11559 , \11560 , \11561 , \11562 , \11563 , \11564 , \11565 , \11566 ,
         \11567 , \11568 , \11569_nG4879 , \11570_nG487a , \11571 , \11572 , \11573 , \11574 , \11575 , \11576 ,
         \11577 , \11578 , \11579 , \11580 , \11581 , \11582 , \11583_nG6580 , \11584_nG6581 , \11585_nG6582 , \11586 ,
         \11587 , \11588 , \11589 , \11590 , \11591 , \11592 , \11593 , \11594 , \11595 , \11596 ,
         \11597 , \11598_nG9c05 , \11599 , \11600 , \11601 , \11602 , \11603 , \11604 , \11605 , \11606 ,
         \11607 , \11608 , \11609 , \11610 , \11611 , \11612 , \11613 , \11614 , \11615 , \11616 ,
         \11617 , \11618 , \11619 , \11620 , \11621 , \11622 , \11623 , \11624 , \11625 , \11626 ,
         \11627 , \11628 , \11629 , \11630 , \11631 , \11632 , \11633 , \11634 , \11635 , \11636 ,
         \11637 , \11638 , \11639 , \11640 , \11641 , \11642 , \11643 , \11644 , \11645 , \11646 ,
         \11647 , \11648 , \11649 , \11650 , \11651 , \11652 , \11653 , \11654 , \11655 , \11656 ,
         \11657 , \11658 , \11659 , \11660 , \11661 , \11662 , \11663 , \11664 , \11665 , \11666 ,
         \11667 , \11668 , \11669 , \11670 , \11671 , \11672 , \11673 , \11674 , \11675 , \11676 ,
         \11677 , \11678 , \11679 , \11680 , \11681 , \11682 , \11683 , \11684 , \11685 , \11686 ,
         \11687 , \11688 , \11689 , \11690 , \11691 , \11692 , \11693 , \11694 , \11695 , \11696 ,
         \11697 , \11698 , \11699 , \11700 , \11701 , \11702 , \11703 , \11704 , \11705 , \11706 ,
         \11707 , \11708 , \11709 , \11710 , \11711 , \11712 , \11713 , \11714 , \11715 , \11716 ,
         \11717 , \11718 , \11719 , \11720 , \11721 , \11722 , \11723 , \11724 , \11725 , \11726 ,
         \11727 , \11728 , \11729 , \11730 , \11731 , \11732 , \11733 , \11734 , \11735 , \11736 ,
         \11737_nG2fb7 , \11738 , \11739 , \11740 , \11741 , \11742 , \11743 , \11744 , \11745 , \11746 ,
         \11747 , \11748 , \11749 , \11750 , \11751 , \11752 , \11753 , \11754 , \11755 , \11756 ,
         \11757 , \11758 , \11759 , \11760 , \11761 , \11762 , \11763 , \11764 , \11765 , \11766 ,
         \11767 , \11768 , \11769 , \11770 , \11771 , \11772 , \11773 , \11774 , \11775 , \11776 ,
         \11777 , \11778 , \11779 , \11780 , \11781 , \11782 , \11783 , \11784 , \11785 , \11786 ,
         \11787 , \11788 , \11789 , \11790 , \11791 , \11792 , \11793 , \11794 , \11795 , \11796 ,
         \11797 , \11798 , \11799 , \11800 , \11801 , \11802 , \11803 , \11804 , \11805 , \11806 ,
         \11807 , \11808 , \11809 , \11810 , \11811 , \11812 , \11813 , \11814 , \11815 , \11816 ,
         \11817 , \11818 , \11819 , \11820 , \11821 , \11822 , \11823 , \11824 , \11825 , \11826 ,
         \11827 , \11828 , \11829 , \11830 , \11831 , \11832 , \11833 , \11834 , \11835 , \11836 ,
         \11837 , \11838 , \11839 , \11840 , \11841 , \11842 , \11843 , \11844 , \11845 , \11846 ,
         \11847 , \11848 , \11849 , \11850 , \11851 , \11852 , \11853 , \11854 , \11855 , \11856 ,
         \11857 , \11858 , \11859 , \11860 , \11861 , \11862 , \11863 , \11864 , \11865 , \11866 ,
         \11867 , \11868 , \11869 , \11870_nG40e4 , \11871 , \11872 , \11873 , \11874 , \11875 , \11876 ,
         \11877 , \11878 , \11879 , \11880 , \11881 , \11882 , \11883 , \11884 , \11885 , \11886 ,
         \11887 , \11888 , \11889 , \11890 , \11891 , \11892 , \11893 , \11894 , \11895 , \11896 ,
         \11897 , \11898 , \11899 , \11900 , \11901 , \11902 , \11903 , \11904 , \11905 , \11906 ,
         \11907 , \11908 , \11909 , \11910 , \11911 , \11912 , \11913 , \11914 , \11915 , \11916 ,
         \11917 , \11918 , \11919 , \11920 , \11921 , \11922 , \11923 , \11924 , \11925 , \11926 ,
         \11927 , \11928 , \11929 , \11930 , \11931 , \11932 , \11933 , \11934 , \11935 , \11936 ,
         \11937 , \11938 , \11939 , \11940 , \11941 , \11942 , \11943 , \11944 , \11945 , \11946 ,
         \11947 , \11948 , \11949 , \11950 , \11951 , \11952 , \11953 , \11954 , \11955 , \11956 ,
         \11957 , \11958 , \11959 , \11960 , \11961 , \11962 , \11963 , \11964 , \11965 , \11966 ,
         \11967 , \11968 , \11969 , \11970 , \11971 , \11972 , \11973 , \11974 , \11975 , \11976 ,
         \11977 , \11978 , \11979 , \11980 , \11981 , \11982 , \11983 , \11984 , \11985 , \11986 ,
         \11987 , \11988 , \11989 , \11990 , \11991 , \11992 , \11993 , \11994 , \11995 , \11996 ,
         \11997 , \11998 , \11999 , \12000 , \12001 , \12002 , \12003 , \12004_nG303c , \12005 , \12006 ,
         \12007 , \12008 , \12009 , \12010 , \12011 , \12012 , \12013 , \12014 , \12015 , \12016 ,
         \12017 , \12018 , \12019 , \12020 , \12021 , \12022 , \12023 , \12024 , \12025 , \12026 ,
         \12027 , \12028 , \12029 , \12030 , \12031 , \12032 , \12033 , \12034 , \12035 , \12036 ,
         \12037 , \12038 , \12039 , \12040 , \12041 , \12042 , \12043 , \12044 , \12045 , \12046 ,
         \12047 , \12048 , \12049 , \12050 , \12051 , \12052 , \12053 , \12054 , \12055 , \12056 ,
         \12057 , \12058 , \12059 , \12060 , \12061 , \12062 , \12063 , \12064 , \12065 , \12066 ,
         \12067 , \12068 , \12069 , \12070 , \12071 , \12072 , \12073 , \12074 , \12075 , \12076 ,
         \12077 , \12078 , \12079 , \12080 , \12081 , \12082 , \12083 , \12084 , \12085 , \12086 ,
         \12087 , \12088 , \12089 , \12090 , \12091 , \12092 , \12093 , \12094 , \12095 , \12096 ,
         \12097 , \12098 , \12099 , \12100 , \12101 , \12102 , \12103 , \12104 , \12105 , \12106 ,
         \12107 , \12108 , \12109 , \12110 , \12111 , \12112 , \12113 , \12114 , \12115 , \12116 ,
         \12117 , \12118 , \12119 , \12120 , \12121 , \12122 , \12123 , \12124 , \12125 , \12126 ,
         \12127 , \12128 , \12129 , \12130 , \12131 , \12132 , \12133 , \12134 , \12135 , \12136 ,
         \12137_nG4169 , \12138 , \12139 , \12140 , \12141 , \12142 , \12143 , \12144 , \12145 , \12146 ,
         \12147 , \12148_nG4448 , \12149 , \12150 , \12151_nG444b , \12152 , \12153 , \12154 , \12155 , \12156 ,
         \12157 , \12158 , \12159 , \12160 , \12161 , \12162 , \12163 , \12164 , \12165 , \12166 ,
         \12167 , \12168 , \12169 , \12170 , \12171 , \12172 , \12173 , \12174 , \12175 , \12176 ,
         \12177 , \12178 , \12179 , \12180 , \12181 , \12182 , \12183 , \12184 , \12185 , \12186 ,
         \12187 , \12188 , \12189 , \12190 , \12191 , \12192 , \12193 , \12194 , \12195 , \12196 ,
         \12197 , \12198 , \12199 , \12200 , \12201 , \12202 , \12203 , \12204 , \12205 , \12206 ,
         \12207 , \12208 , \12209 , \12210 , \12211 , \12212 , \12213 , \12214 , \12215 , \12216 ,
         \12217 , \12218 , \12219 , \12220 , \12221 , \12222 , \12223 , \12224 , \12225 , \12226 ,
         \12227 , \12228 , \12229 , \12230 , \12231 , \12232 , \12233 , \12234 , \12235 , \12236 ,
         \12237 , \12238 , \12239 , \12240 , \12241 , \12242 , \12243 , \12244 , \12245 , \12246 ,
         \12247 , \12248 , \12249 , \12250 , \12251 , \12252 , \12253 , \12254 , \12255 , \12256 ,
         \12257 , \12258 , \12259 , \12260 , \12261 , \12262 , \12263 , \12264 , \12265 , \12266 ,
         \12267 , \12268 , \12269 , \12270 , \12271 , \12272 , \12273 , \12274 , \12275 , \12276 ,
         \12277 , \12278 , \12279 , \12280 , \12281 , \12282 , \12283 , \12284 , \12285 , \12286 ,
         \12287 , \12288 , \12289 , \12290 , \12291 , \12292 , \12293 , \12294 , \12295 , \12296 ,
         \12297 , \12298 , \12299 , \12300 , \12301 , \12302 , \12303 , \12304 , \12305 , \12306 ,
         \12307 , \12308 , \12309 , \12310 , \12311 , \12312 , \12313 , \12314_nG6583 , \12315 , \12316 ,
         \12317 , \12318 , \12319 , \12320 , \12321 , \12322 , \12323 , \12324 , \12325 , \12326 ,
         \12327 , \12328 , \12329 , \12330 , \12331 , \12332 , \12333 , \12334 , \12335 , \12336 ,
         \12337 , \12338 , \12339 , \12340 , \12341 , \12342 , \12343 , \12344 , \12345 , \12346 ,
         \12347 , \12348 , \12349 , \12350 , \12351 , \12352 , \12353 , \12354 , \12355 , \12356 ,
         \12357 , \12358 , \12359 , \12360 , \12361 , \12362 , \12363 , \12364 , \12365 , \12366 ,
         \12367 , \12368 , \12369 , \12370 , \12371 , \12372 , \12373 , \12374 , \12375 , \12376 ,
         \12377 , \12378 , \12379 , \12380 , \12381 , \12382 , \12383 , \12384 , \12385 , \12386 ,
         \12387 , \12388 , \12389 , \12390 , \12391 , \12392 , \12393 , \12394 , \12395 , \12396 ,
         \12397 , \12398 , \12399 , \12400 , \12401 , \12402 , \12403 , \12404 , \12405 , \12406 ,
         \12407 , \12408 , \12409 , \12410 , \12411 , \12412 , \12413 , \12414 , \12415 , \12416 ,
         \12417 , \12418 , \12419 , \12420 , \12421 , \12422 , \12423 , \12424 , \12425 , \12426 ,
         \12427 , \12428 , \12429 , \12430 , \12431 , \12432 , \12433 , \12434 , \12435 , \12436 ,
         \12437 , \12438 , \12439 , \12440 , \12441 , \12442 , \12443 , \12444 , \12445 , \12446_nG6584 ,
         \12447_nG6585 , \12448 , \12449 , \12450 , \12451 , \12452 , \12453 , \12454 , \12455 , \12456 ,
         \12457_nG48fe , \12458_nG4982 , \12459_nG4983 , \12460 , \12461 , \12462 , \12463 , \12464 , \12465 , \12466 ,
         \12467 , \12468 , \12469 , \12470_nG9c02 , \12471 , \12472 , \12473 , \12474 , \12475 , \12476 ,
         \12477 , \12478 , \12479 , \12480 , \12481 , \12482 , \12483 , \12484 , \12485 , \12486 ,
         \12487 , \12488 , \12489 , \12490 , \12491 , \12492 , \12493 , \12494 , \12495 , \12496 ,
         \12497 , \12498 , \12499 , \12500 , \12501 , \12502 , \12503 , \12504 , \12505 , \12506 ,
         \12507 , \12508 , \12509 , \12510 , \12511 , \12512 , \12513 , \12514 , \12515 , \12516 ,
         \12517 , \12518 , \12519 , \12520 , \12521 , \12522 , \12523 , \12524 , \12525 , \12526 ,
         \12527 , \12528 , \12529 , \12530 , \12531 , \12532 , \12533 , \12534 , \12535 , \12536 ,
         \12537 , \12538 , \12539 , \12540 , \12541 , \12542 , \12543 , \12544 , \12545 , \12546 ,
         \12547 , \12548 , \12549 , \12550 , \12551 , \12552 , \12553 , \12554 , \12555 , \12556 ,
         \12557 , \12558 , \12559 , \12560 , \12561 , \12562 , \12563 , \12564 , \12565 , \12566 ,
         \12567 , \12568 , \12569 , \12570 , \12571 , \12572 , \12573 , \12574 , \12575 , \12576 ,
         \12577 , \12578 , \12579 , \12580 , \12581 , \12582 , \12583 , \12584 , \12585 , \12586 ,
         \12587 , \12588 , \12589 , \12590 , \12591 , \12592 , \12593 , \12594 , \12595 , \12596 ,
         \12597 , \12598 , \12599 , \12600 , \12601 , \12602 , \12603 , \12604 , \12605 , \12606 ,
         \12607 , \12608 , \12609 , \12610 , \12611 , \12612 , \12613 , \12614 , \12615 , \12616 ,
         \12617 , \12618 , \12619 , \12620 , \12621 , \12622 , \12623 , \12624 , \12625 , \12626 ,
         \12627 , \12628 , \12629 , \12630 , \12631 , \12632 , \12633 , \12634 , \12635_nG6586 , \12636 ,
         \12637 , \12638 , \12639 , \12640 , \12641 , \12642 , \12643 , \12644 , \12645 , \12646 ,
         \12647 , \12648 , \12649 , \12650 , \12651 , \12652 , \12653 , \12654 , \12655 , \12656 ,
         \12657 , \12658 , \12659 , \12660 , \12661 , \12662 , \12663 , \12664 , \12665 , \12666 ,
         \12667 , \12668 , \12669 , \12670 , \12671 , \12672 , \12673 , \12674 , \12675 , \12676 ,
         \12677 , \12678 , \12679 , \12680 , \12681 , \12682 , \12683 , \12684 , \12685 , \12686 ,
         \12687 , \12688 , \12689 , \12690 , \12691 , \12692 , \12693 , \12694 , \12695 , \12696 ,
         \12697 , \12698 , \12699 , \12700 , \12701 , \12702 , \12703 , \12704 , \12705 , \12706 ,
         \12707 , \12708 , \12709 , \12710 , \12711 , \12712 , \12713 , \12714 , \12715 , \12716 ,
         \12717 , \12718 , \12719 , \12720 , \12721 , \12722 , \12723 , \12724 , \12725 , \12726 ,
         \12727 , \12728 , \12729 , \12730 , \12731 , \12732 , \12733 , \12734 , \12735 , \12736 ,
         \12737 , \12738 , \12739 , \12740 , \12741 , \12742 , \12743 , \12744 , \12745 , \12746 ,
         \12747 , \12748 , \12749 , \12750 , \12751 , \12752 , \12753 , \12754 , \12755 , \12756 ,
         \12757 , \12758 , \12759 , \12760 , \12761 , \12762 , \12763 , \12764 , \12765 , \12766 ,
         \12767_nG6587 , \12768_nG6588 , \12769 , \12770 , \12771 , \12772 , \12773 , \12774_nG4a07 , \12775_nG4a8b , \12776_nG4a8c ,
         \12777 , \12778 , \12779 , \12780 , \12781 , \12782 , \12783 , \12784 , \12785 , \12786 ,
         \12787 , \12788 , \12789 , \12790 , \12791 , \12792 , \12793 , \12794 , \12795 , \12796 ,
         \12797 , \12798 , \12799 , \12800 , \12801_nG9bff , \12802 , \12803 , \12804 , \12805 , \12806 ,
         \12807 , \12808 , \12809 , \12810 , \12811 , \12812 , \12813 , \12814 , \12815 , \12816 ,
         \12817 , \12818 , \12819 , \12820 , \12821 , \12822 , \12823 , \12824 , \12825 , \12826 ,
         \12827 , \12828 , \12829 , \12830 , \12831 , \12832 , \12833 , \12834 , \12835 , \12836 ,
         \12837 , \12838 , \12839 , \12840 , \12841 , \12842 , \12843 , \12844 , \12845 , \12846 ,
         \12847 , \12848 , \12849 , \12850 , \12851 , \12852 , \12853 , \12854 , \12855 , \12856 ,
         \12857 , \12858 , \12859 , \12860 , \12861 , \12862 , \12863 , \12864 , \12865 , \12866 ,
         \12867 , \12868 , \12869 , \12870 , \12871 , \12872 , \12873 , \12874 , \12875 , \12876 ,
         \12877 , \12878 , \12879 , \12880 , \12881 , \12882 , \12883 , \12884 , \12885 , \12886 ,
         \12887 , \12888 , \12889 , \12890 , \12891 , \12892 , \12893 , \12894 , \12895 , \12896 ,
         \12897 , \12898 , \12899 , \12900 , \12901 , \12902 , \12903 , \12904 , \12905 , \12906 ,
         \12907 , \12908 , \12909 , \12910 , \12911 , \12912 , \12913 , \12914 , \12915 , \12916 ,
         \12917 , \12918 , \12919 , \12920 , \12921 , \12922 , \12923 , \12924 , \12925 , \12926 ,
         \12927 , \12928 , \12929 , \12930 , \12931 , \12932 , \12933 , \12934 , \12935 , \12936 ,
         \12937 , \12938 , \12939 , \12940 , \12941 , \12942 , \12943 , \12944 , \12945 , \12946 ,
         \12947 , \12948 , \12949 , \12950_nG2ead , \12951 , \12952 , \12953 , \12954 , \12955 , \12956 ,
         \12957 , \12958 , \12959 , \12960 , \12961 , \12962 , \12963 , \12964 , \12965 , \12966 ,
         \12967 , \12968 , \12969 , \12970 , \12971 , \12972 , \12973 , \12974 , \12975 , \12976 ,
         \12977 , \12978 , \12979 , \12980 , \12981 , \12982 , \12983 , \12984 , \12985 , \12986 ,
         \12987 , \12988 , \12989 , \12990 , \12991 , \12992 , \12993 , \12994 , \12995 , \12996 ,
         \12997 , \12998 , \12999 , \13000 , \13001 , \13002 , \13003 , \13004 , \13005 , \13006 ,
         \13007 , \13008 , \13009 , \13010 , \13011 , \13012 , \13013 , \13014 , \13015 , \13016 ,
         \13017 , \13018 , \13019 , \13020 , \13021 , \13022 , \13023 , \13024 , \13025 , \13026 ,
         \13027 , \13028 , \13029 , \13030 , \13031 , \13032 , \13033 , \13034 , \13035 , \13036 ,
         \13037 , \13038 , \13039 , \13040 , \13041 , \13042 , \13043 , \13044 , \13045 , \13046 ,
         \13047 , \13048 , \13049 , \13050 , \13051 , \13052 , \13053 , \13054 , \13055 , \13056 ,
         \13057 , \13058 , \13059 , \13060 , \13061 , \13062 , \13063 , \13064 , \13065 , \13066 ,
         \13067 , \13068 , \13069 , \13070 , \13071 , \13072 , \13073 , \13074 , \13075 , \13076 ,
         \13077 , \13078 , \13079 , \13080 , \13081 , \13082 , \13083_nG3fda , \13084 , \13085 , \13086 ,
         \13087 , \13088 , \13089 , \13090 , \13091 , \13092 , \13093 , \13094 , \13095 , \13096 ,
         \13097 , \13098 , \13099 , \13100 , \13101 , \13102 , \13103 , \13104 , \13105 , \13106 ,
         \13107 , \13108 , \13109 , \13110 , \13111 , \13112 , \13113 , \13114 , \13115 , \13116 ,
         \13117 , \13118 , \13119 , \13120 , \13121 , \13122 , \13123 , \13124 , \13125 , \13126 ,
         \13127 , \13128 , \13129 , \13130 , \13131 , \13132 , \13133 , \13134 , \13135 , \13136 ,
         \13137 , \13138 , \13139 , \13140 , \13141 , \13142 , \13143 , \13144 , \13145 , \13146 ,
         \13147 , \13148 , \13149 , \13150 , \13151 , \13152 , \13153 , \13154 , \13155 , \13156 ,
         \13157 , \13158 , \13159 , \13160 , \13161 , \13162 , \13163 , \13164 , \13165 , \13166 ,
         \13167 , \13168 , \13169 , \13170 , \13171 , \13172 , \13173 , \13174 , \13175 , \13176 ,
         \13177 , \13178 , \13179 , \13180 , \13181 , \13182 , \13183 , \13184 , \13185 , \13186 ,
         \13187 , \13188 , \13189 , \13190 , \13191 , \13192 , \13193 , \13194 , \13195 , \13196 ,
         \13197 , \13198 , \13199 , \13200 , \13201 , \13202 , \13203 , \13204 , \13205 , \13206 ,
         \13207 , \13208 , \13209 , \13210 , \13211 , \13212 , \13213 , \13214 , \13215 , \13216 ,
         \13217_nG2f32 , \13218 , \13219 , \13220 , \13221 , \13222 , \13223 , \13224 , \13225 , \13226 ,
         \13227 , \13228 , \13229 , \13230 , \13231 , \13232 , \13233 , \13234 , \13235 , \13236 ,
         \13237 , \13238 , \13239 , \13240 , \13241 , \13242 , \13243 , \13244 , \13245 , \13246 ,
         \13247 , \13248 , \13249 , \13250 , \13251 , \13252 , \13253 , \13254 , \13255 , \13256 ,
         \13257 , \13258 , \13259 , \13260 , \13261 , \13262 , \13263 , \13264 , \13265 , \13266 ,
         \13267 , \13268 , \13269 , \13270 , \13271 , \13272 , \13273 , \13274 , \13275 , \13276 ,
         \13277 , \13278 , \13279 , \13280 , \13281 , \13282 , \13283 , \13284 , \13285 , \13286 ,
         \13287 , \13288 , \13289 , \13290 , \13291 , \13292 , \13293 , \13294 , \13295 , \13296 ,
         \13297 , \13298 , \13299 , \13300 , \13301 , \13302 , \13303 , \13304 , \13305 , \13306 ,
         \13307 , \13308 , \13309 , \13310 , \13311 , \13312 , \13313 , \13314 , \13315 , \13316 ,
         \13317 , \13318 , \13319 , \13320 , \13321 , \13322 , \13323 , \13324 , \13325 , \13326 ,
         \13327 , \13328 , \13329 , \13330 , \13331 , \13332 , \13333 , \13334 , \13335 , \13336 ,
         \13337 , \13338 , \13339 , \13340 , \13341 , \13342 , \13343 , \13344 , \13345 , \13346 ,
         \13347 , \13348 , \13349 , \13350_nG405f , \13351 , \13352 , \13353 , \13354 , \13355 , \13356 ,
         \13357 , \13358 , \13359 , \13360 , \13361_nG4442 , \13362 , \13363 , \13364_nG4445 , \13365 , \13366 ,
         \13367 , \13368 , \13369 , \13370 , \13371 , \13372 , \13373 , \13374 , \13375 , \13376 ,
         \13377 , \13378 , \13379 , \13380 , \13381 , \13382 , \13383 , \13384 , \13385 , \13386 ,
         \13387 , \13388 , \13389 , \13390 , \13391 , \13392 , \13393 , \13394 , \13395 , \13396 ,
         \13397 , \13398 , \13399 , \13400 , \13401 , \13402 , \13403 , \13404 , \13405 , \13406 ,
         \13407 , \13408 , \13409 , \13410 , \13411 , \13412 , \13413 , \13414 , \13415 , \13416 ,
         \13417 , \13418 , \13419 , \13420 , \13421 , \13422 , \13423 , \13424 , \13425 , \13426 ,
         \13427 , \13428 , \13429 , \13430 , \13431 , \13432 , \13433 , \13434 , \13435 , \13436 ,
         \13437 , \13438 , \13439 , \13440 , \13441 , \13442 , \13443 , \13444 , \13445 , \13446 ,
         \13447 , \13448 , \13449 , \13450 , \13451 , \13452 , \13453 , \13454 , \13455 , \13456 ,
         \13457 , \13458 , \13459 , \13460 , \13461 , \13462 , \13463 , \13464 , \13465 , \13466 ,
         \13467 , \13468 , \13469 , \13470 , \13471 , \13472 , \13473 , \13474 , \13475 , \13476 ,
         \13477 , \13478 , \13479 , \13480 , \13481 , \13482 , \13483 , \13484 , \13485 , \13486 ,
         \13487 , \13488 , \13489 , \13490 , \13491 , \13492 , \13493 , \13494 , \13495 , \13496 ,
         \13497 , \13498 , \13499 , \13500 , \13501 , \13502 , \13503 , \13504 , \13505 , \13506 ,
         \13507 , \13508 , \13509 , \13510 , \13511 , \13512 , \13513 , \13514 , \13515 , \13516 ,
         \13517 , \13518 , \13519 , \13520 , \13521 , \13522 , \13523 , \13524 , \13525 , \13526 ,
         \13527 , \13528 , \13529 , \13530 , \13531 , \13532 , \13533 , \13534 , \13535 , \13536 ,
         \13537 , \13538 , \13539 , \13540 , \13541 , \13542 , \13543 , \13544 , \13545_nG6589 , \13546 ,
         \13547 , \13548 , \13549 , \13550 , \13551 , \13552 , \13553 , \13554 , \13555 , \13556 ,
         \13557 , \13558 , \13559 , \13560 , \13561 , \13562 , \13563 , \13564 , \13565 , \13566 ,
         \13567 , \13568 , \13569 , \13570 , \13571 , \13572 , \13573 , \13574 , \13575 , \13576 ,
         \13577 , \13578 , \13579 , \13580 , \13581 , \13582 , \13583 , \13584 , \13585 , \13586 ,
         \13587 , \13588 , \13589 , \13590 , \13591 , \13592 , \13593 , \13594 , \13595 , \13596 ,
         \13597 , \13598 , \13599 , \13600 , \13601 , \13602 , \13603 , \13604 , \13605 , \13606 ,
         \13607 , \13608 , \13609 , \13610 , \13611 , \13612 , \13613 , \13614 , \13615 , \13616 ,
         \13617 , \13618 , \13619 , \13620 , \13621 , \13622 , \13623 , \13624 , \13625 , \13626 ,
         \13627 , \13628 , \13629 , \13630 , \13631 , \13632 , \13633 , \13634 , \13635 , \13636 ,
         \13637 , \13638 , \13639 , \13640 , \13641 , \13642 , \13643 , \13644 , \13645 , \13646 ,
         \13647 , \13648 , \13649 , \13650 , \13651 , \13652 , \13653 , \13654 , \13655 , \13656 ,
         \13657 , \13658 , \13659 , \13660 , \13661 , \13662 , \13663 , \13664 , \13665 , \13666 ,
         \13667 , \13668 , \13669 , \13670 , \13671 , \13672 , \13673 , \13674 , \13675 , \13676 ,
         \13677_nG658a , \13678_nG658b , \13679 , \13680 , \13681 , \13682 , \13683 , \13684 , \13685 , \13686 ,
         \13687 , \13688_nG4b10 , \13689_nG4b94 , \13690_nG4b95 , \13691 , \13692 , \13693 , \13694 , \13695 , \13696 ,
         \13697 , \13698 , \13699 , \13700 , \13701 , \13702 , \13703 , \13704 , \13705_nG9bfc , \13706 ,
         \13707 , \13708 , \13709 , \13710 , \13711 , \13712 , \13713 , \13714 , \13715 , \13716 ,
         \13717 , \13718 , \13719 , \13720 , \13721 , \13722 , \13723 , \13724 , \13725 , \13726 ,
         \13727 , \13728 , \13729 , \13730 , \13731 , \13732 , \13733 , \13734 , \13735 , \13736 ,
         \13737 , \13738 , \13739 , \13740 , \13741 , \13742 , \13743 , \13744 , \13745 , \13746 ,
         \13747 , \13748 , \13749 , \13750 , \13751 , \13752 , \13753 , \13754 , \13755 , \13756 ,
         \13757 , \13758 , \13759 , \13760 , \13761 , \13762 , \13763 , \13764 , \13765 , \13766 ,
         \13767 , \13768 , \13769 , \13770 , \13771 , \13772 , \13773 , \13774 , \13775 , \13776 ,
         \13777 , \13778 , \13779 , \13780 , \13781 , \13782 , \13783 , \13784 , \13785 , \13786 ,
         \13787 , \13788 , \13789 , \13790 , \13791 , \13792 , \13793 , \13794 , \13795 , \13796 ,
         \13797 , \13798 , \13799 , \13800 , \13801 , \13802 , \13803 , \13804 , \13805 , \13806 ,
         \13807 , \13808 , \13809 , \13810 , \13811 , \13812 , \13813 , \13814 , \13815 , \13816 ,
         \13817 , \13818 , \13819 , \13820 , \13821 , \13822 , \13823 , \13824 , \13825 , \13826 ,
         \13827 , \13828 , \13829 , \13830 , \13831 , \13832 , \13833 , \13834 , \13835 , \13836 ,
         \13837 , \13838 , \13839 , \13840 , \13841 , \13842 , \13843 , \13844 , \13845 , \13846 ,
         \13847 , \13848 , \13849 , \13850 , \13851 , \13852 , \13853 , \13854 , \13855 , \13856 ,
         \13857 , \13858 , \13859 , \13860 , \13861 , \13862 , \13863 , \13864 , \13865 , \13866 ,
         \13867 , \13868 , \13869 , \13870 , \13871 , \13872 , \13873 , \13874 , \13875 , \13876 ,
         \13877 , \13878 , \13879 , \13880 , \13881 , \13882 , \13883 , \13884 , \13885 , \13886 ,
         \13887 , \13888 , \13889 , \13890_nG658c , \13891 , \13892 , \13893 , \13894 , \13895 , \13896 ,
         \13897 , \13898 , \13899 , \13900 , \13901 , \13902 , \13903 , \13904 , \13905 , \13906 ,
         \13907 , \13908 , \13909 , \13910 , \13911 , \13912 , \13913 , \13914 , \13915 , \13916 ,
         \13917 , \13918 , \13919 , \13920 , \13921 , \13922 , \13923 , \13924 , \13925 , \13926 ,
         \13927 , \13928 , \13929 , \13930 , \13931 , \13932 , \13933 , \13934 , \13935 , \13936 ,
         \13937 , \13938 , \13939 , \13940 , \13941 , \13942 , \13943 , \13944 , \13945 , \13946 ,
         \13947 , \13948 , \13949 , \13950 , \13951 , \13952 , \13953 , \13954 , \13955 , \13956 ,
         \13957 , \13958 , \13959 , \13960 , \13961 , \13962 , \13963 , \13964 , \13965 , \13966 ,
         \13967 , \13968 , \13969 , \13970 , \13971 , \13972 , \13973 , \13974 , \13975 , \13976 ,
         \13977 , \13978 , \13979 , \13980 , \13981 , \13982 , \13983 , \13984 , \13985 , \13986 ,
         \13987 , \13988 , \13989 , \13990 , \13991 , \13992 , \13993 , \13994 , \13995 , \13996 ,
         \13997 , \13998 , \13999 , \14000 , \14001 , \14002 , \14003 , \14004 , \14005 , \14006 ,
         \14007 , \14008 , \14009 , \14010 , \14011 , \14012 , \14013 , \14014 , \14015 , \14016 ,
         \14017 , \14018 , \14019 , \14020 , \14021 , \14022_nG658d , \14023_nG658e , \14024 , \14025 , \14026 ,
         \14027 , \14028 , \14029_nG4c19 , \14030_nG4c9d , \14031_nG4c9e , \14032 , \14033 , \14034 , \14035 , \14036 ,
         \14037 , \14038 , \14039 , \14040 , \14041 , \14042 , \14043 , \14044 , \14045 , \14046 ,
         \14047 , \14048 , \14049 , \14050 , \14051 , \14052 , \14053 , \14054 , \14055 , \14056 ,
         \14057 , \14058 , \14059 , \14060 , \14061 , \14062 , \14063 , \14064 , \14065 , \14066 ,
         \14067 , \14068 , \14069 , \14070_nG9bf9 , \14071 , \14072 , \14073 , \14074 , \14075 , \14076 ,
         \14077 , \14078 , \14079 , \14080 , \14081 , \14082 , \14083 , \14084 , \14085 , \14086 ,
         \14087 , \14088 , \14089 , \14090 , \14091 , \14092 , \14093 , \14094 , \14095 , \14096 ,
         \14097 , \14098 , \14099 , \14100 , \14101 , \14102 , \14103 , \14104 , \14105 , \14106 ,
         \14107 , \14108 , \14109 , \14110 , \14111 , \14112 , \14113 , \14114 , \14115 , \14116 ,
         \14117 , \14118 , \14119 , \14120 , \14121 , \14122 , \14123 , \14124 , \14125 , \14126 ,
         \14127 , \14128 , \14129 , \14130 , \14131 , \14132 , \14133 , \14134 , \14135 , \14136 ,
         \14137 , \14138 , \14139 , \14140 , \14141 , \14142 , \14143 , \14144 , \14145 , \14146 ,
         \14147 , \14148 , \14149 , \14150 , \14151 , \14152 , \14153 , \14154 , \14155 , \14156 ,
         \14157 , \14158 , \14159 , \14160 , \14161 , \14162 , \14163 , \14164 , \14165 , \14166 ,
         \14167 , \14168 , \14169 , \14170 , \14171 , \14172 , \14173 , \14174 , \14175 , \14176 ,
         \14177 , \14178 , \14179 , \14180 , \14181 , \14182 , \14183 , \14184 , \14185 , \14186 ,
         \14187 , \14188 , \14189 , \14190 , \14191 , \14192 , \14193 , \14194 , \14195 , \14196 ,
         \14197 , \14198 , \14199 , \14200 , \14201 , \14202 , \14203 , \14204 , \14205 , \14206 ,
         \14207 , \14208 , \14209 , \14210 , \14211_nG2da3 , \14212 , \14213 , \14214 , \14215 , \14216 ,
         \14217 , \14218 , \14219 , \14220 , \14221 , \14222 , \14223 , \14224 , \14225 , \14226 ,
         \14227 , \14228 , \14229 , \14230 , \14231 , \14232 , \14233 , \14234 , \14235 , \14236 ,
         \14237 , \14238 , \14239 , \14240 , \14241 , \14242 , \14243 , \14244 , \14245 , \14246 ,
         \14247 , \14248 , \14249 , \14250 , \14251 , \14252 , \14253 , \14254 , \14255 , \14256 ,
         \14257 , \14258 , \14259 , \14260 , \14261 , \14262 , \14263 , \14264 , \14265 , \14266 ,
         \14267 , \14268 , \14269 , \14270 , \14271 , \14272 , \14273 , \14274 , \14275 , \14276 ,
         \14277 , \14278 , \14279 , \14280 , \14281 , \14282 , \14283 , \14284 , \14285 , \14286 ,
         \14287 , \14288 , \14289 , \14290 , \14291 , \14292 , \14293 , \14294 , \14295 , \14296 ,
         \14297 , \14298 , \14299 , \14300 , \14301 , \14302 , \14303 , \14304 , \14305 , \14306 ,
         \14307 , \14308 , \14309 , \14310 , \14311 , \14312 , \14313 , \14314 , \14315 , \14316 ,
         \14317 , \14318 , \14319 , \14320 , \14321 , \14322 , \14323 , \14324 , \14325 , \14326 ,
         \14327 , \14328 , \14329 , \14330 , \14331 , \14332 , \14333 , \14334 , \14335 , \14336 ,
         \14337 , \14338 , \14339 , \14340 , \14341 , \14342 , \14343 , \14344_nG3ed0 , \14345 , \14346 ,
         \14347 , \14348 , \14349 , \14350 , \14351 , \14352 , \14353 , \14354 , \14355 , \14356 ,
         \14357 , \14358 , \14359 , \14360 , \14361 , \14362 , \14363 , \14364 , \14365 , \14366 ,
         \14367 , \14368 , \14369 , \14370 , \14371 , \14372 , \14373 , \14374 , \14375 , \14376 ,
         \14377 , \14378 , \14379 , \14380 , \14381 , \14382 , \14383 , \14384 , \14385 , \14386 ,
         \14387 , \14388 , \14389 , \14390 , \14391 , \14392 , \14393 , \14394 , \14395 , \14396 ,
         \14397 , \14398 , \14399 , \14400 , \14401 , \14402 , \14403 , \14404 , \14405 , \14406 ,
         \14407 , \14408 , \14409 , \14410 , \14411 , \14412 , \14413 , \14414 , \14415 , \14416 ,
         \14417 , \14418 , \14419 , \14420 , \14421 , \14422 , \14423 , \14424 , \14425 , \14426 ,
         \14427 , \14428 , \14429 , \14430 , \14431 , \14432 , \14433 , \14434 , \14435 , \14436 ,
         \14437 , \14438 , \14439 , \14440 , \14441 , \14442 , \14443 , \14444 , \14445 , \14446 ,
         \14447 , \14448 , \14449 , \14450 , \14451 , \14452 , \14453 , \14454 , \14455 , \14456 ,
         \14457 , \14458 , \14459 , \14460 , \14461 , \14462 , \14463 , \14464 , \14465 , \14466 ,
         \14467 , \14468 , \14469 , \14470 , \14471 , \14472 , \14473 , \14474 , \14475 , \14476 ,
         \14477 , \14478_nG2e28 , \14479 , \14480 , \14481 , \14482 , \14483 , \14484 , \14485 , \14486 ,
         \14487 , \14488 , \14489 , \14490 , \14491 , \14492 , \14493 , \14494 , \14495 , \14496 ,
         \14497 , \14498 , \14499 , \14500 , \14501 , \14502 , \14503 , \14504 , \14505 , \14506 ,
         \14507 , \14508 , \14509 , \14510 , \14511 , \14512 , \14513 , \14514 , \14515 , \14516 ,
         \14517 , \14518 , \14519 , \14520 , \14521 , \14522 , \14523 , \14524 , \14525 , \14526 ,
         \14527 , \14528 , \14529 , \14530 , \14531 , \14532 , \14533 , \14534 , \14535 , \14536 ,
         \14537 , \14538 , \14539 , \14540 , \14541 , \14542 , \14543 , \14544 , \14545 , \14546 ,
         \14547 , \14548 , \14549 , \14550 , \14551 , \14552 , \14553 , \14554 , \14555 , \14556 ,
         \14557 , \14558 , \14559 , \14560 , \14561 , \14562 , \14563 , \14564 , \14565 , \14566 ,
         \14567 , \14568 , \14569 , \14570 , \14571 , \14572 , \14573 , \14574 , \14575 , \14576 ,
         \14577 , \14578 , \14579 , \14580 , \14581 , \14582 , \14583 , \14584 , \14585 , \14586 ,
         \14587 , \14588 , \14589 , \14590 , \14591 , \14592 , \14593 , \14594 , \14595 , \14596 ,
         \14597 , \14598 , \14599 , \14600 , \14601 , \14602 , \14603 , \14604 , \14605 , \14606 ,
         \14607 , \14608 , \14609 , \14610 , \14611_nG3f55 , \14612 , \14613 , \14614 , \14615 , \14616 ,
         \14617 , \14618 , \14619 , \14620 , \14621 , \14622_nG443c , \14623 , \14624 , \14625_nG443f , \14626 ,
         \14627 , \14628 , \14629 , \14630 , \14631 , \14632 , \14633 , \14634 , \14635 , \14636 ,
         \14637 , \14638 , \14639 , \14640 , \14641 , \14642 , \14643 , \14644 , \14645 , \14646 ,
         \14647 , \14648 , \14649 , \14650 , \14651 , \14652 , \14653 , \14654 , \14655 , \14656 ,
         \14657 , \14658 , \14659 , \14660 , \14661 , \14662 , \14663 , \14664 , \14665 , \14666 ,
         \14667 , \14668 , \14669 , \14670 , \14671 , \14672 , \14673 , \14674 , \14675 , \14676 ,
         \14677 , \14678 , \14679 , \14680 , \14681 , \14682 , \14683 , \14684 , \14685 , \14686 ,
         \14687 , \14688 , \14689 , \14690 , \14691 , \14692 , \14693 , \14694 , \14695 , \14696 ,
         \14697 , \14698 , \14699 , \14700 , \14701 , \14702 , \14703 , \14704 , \14705 , \14706 ,
         \14707 , \14708 , \14709 , \14710 , \14711 , \14712 , \14713 , \14714 , \14715 , \14716 ,
         \14717 , \14718 , \14719 , \14720 , \14721 , \14722 , \14723 , \14724 , \14725 , \14726 ,
         \14727 , \14728 , \14729 , \14730 , \14731 , \14732 , \14733 , \14734 , \14735 , \14736 ,
         \14737 , \14738 , \14739 , \14740 , \14741 , \14742 , \14743 , \14744 , \14745 , \14746 ,
         \14747 , \14748 , \14749 , \14750 , \14751 , \14752 , \14753 , \14754 , \14755 , \14756 ,
         \14757 , \14758 , \14759 , \14760 , \14761 , \14762 , \14763 , \14764 , \14765 , \14766 ,
         \14767 , \14768 , \14769 , \14770 , \14771 , \14772 , \14773 , \14774 , \14775 , \14776 ,
         \14777 , \14778 , \14779 , \14780 , \14781 , \14782 , \14783 , \14784 , \14785 , \14786 ,
         \14787 , \14788 , \14789 , \14790 , \14791 , \14792 , \14793 , \14794 , \14795 , \14796 ,
         \14797 , \14798 , \14799 , \14800 , \14801 , \14802 , \14803 , \14804 , \14805 , \14806 ,
         \14807 , \14808 , \14809 , \14810 , \14811 , \14812 , \14813 , \14814 , \14815 , \14816_nG658f ,
         \14817 , \14818 , \14819 , \14820 , \14821 , \14822 , \14823 , \14824 , \14825 , \14826 ,
         \14827 , \14828 , \14829 , \14830 , \14831 , \14832 , \14833 , \14834 , \14835 , \14836 ,
         \14837 , \14838 , \14839 , \14840 , \14841 , \14842 , \14843 , \14844 , \14845 , \14846 ,
         \14847 , \14848 , \14849 , \14850 , \14851 , \14852 , \14853 , \14854 , \14855 , \14856 ,
         \14857 , \14858 , \14859 , \14860 , \14861 , \14862 , \14863 , \14864 , \14865 , \14866 ,
         \14867 , \14868 , \14869 , \14870 , \14871 , \14872 , \14873 , \14874 , \14875 , \14876 ,
         \14877 , \14878 , \14879 , \14880 , \14881 , \14882 , \14883 , \14884 , \14885 , \14886 ,
         \14887 , \14888 , \14889 , \14890 , \14891 , \14892 , \14893 , \14894 , \14895 , \14896 ,
         \14897 , \14898 , \14899 , \14900 , \14901 , \14902 , \14903 , \14904 , \14905 , \14906 ,
         \14907 , \14908 , \14909 , \14910 , \14911 , \14912 , \14913 , \14914 , \14915 , \14916 ,
         \14917 , \14918 , \14919 , \14920 , \14921 , \14922 , \14923 , \14924 , \14925 , \14926 ,
         \14927 , \14928 , \14929 , \14930 , \14931 , \14932 , \14933 , \14934 , \14935 , \14936 ,
         \14937 , \14938 , \14939 , \14940 , \14941 , \14942 , \14943 , \14944 , \14945 , \14946 ,
         \14947 , \14948_nG6590 , \14949_nG6591 , \14950 , \14951 , \14952 , \14953 , \14954 , \14955 , \14956 ,
         \14957 , \14958 , \14959_nG4d22 , \14960_nG4da6 , \14961_nG4da7 , \14962 , \14963 , \14964 , \14965 , \14966 ,
         \14967 , \14968 , \14969 , \14970 , \14971 , \14972 , \14973 , \14974 , \14975 , \14976 ,
         \14977 , \14978 , \14979 , \14980 , \14981 , \14982 , \14983 , \14984_nG9bf6 , \14985 , \14986 ,
         \14987 , \14988 , \14989 , \14990 , \14991 , \14992 , \14993 , \14994 , \14995 , \14996 ,
         \14997 , \14998 , \14999 , \15000 , \15001 , \15002 , \15003 , \15004 , \15005 , \15006 ,
         \15007 , \15008 , \15009 , \15010 , \15011 , \15012 , \15013 , \15014 , \15015 , \15016 ,
         \15017 , \15018 , \15019 , \15020 , \15021 , \15022 , \15023 , \15024 , \15025 , \15026 ,
         \15027 , \15028 , \15029 , \15030 , \15031 , \15032 , \15033 , \15034 , \15035 , \15036 ,
         \15037 , \15038 , \15039 , \15040 , \15041 , \15042 , \15043 , \15044 , \15045 , \15046 ,
         \15047 , \15048 , \15049 , \15050 , \15051 , \15052 , \15053 , \15054 , \15055 , \15056 ,
         \15057 , \15058 , \15059 , \15060 , \15061 , \15062 , \15063 , \15064 , \15065 , \15066 ,
         \15067 , \15068 , \15069 , \15070 , \15071 , \15072 , \15073 , \15074 , \15075 , \15076 ,
         \15077 , \15078 , \15079 , \15080 , \15081 , \15082 , \15083 , \15084 , \15085 , \15086 ,
         \15087 , \15088 , \15089 , \15090 , \15091 , \15092 , \15093 , \15094 , \15095 , \15096 ,
         \15097 , \15098 , \15099 , \15100 , \15101 , \15102 , \15103 , \15104 , \15105 , \15106 ,
         \15107 , \15108 , \15109 , \15110 , \15111 , \15112 , \15113 , \15114 , \15115 , \15116 ,
         \15117 , \15118 , \15119 , \15120 , \15121 , \15122 , \15123 , \15124 , \15125 , \15126 ,
         \15127 , \15128 , \15129 , \15130 , \15131 , \15132 , \15133 , \15134 , \15135 , \15136 ,
         \15137 , \15138 , \15139 , \15140 , \15141 , \15142 , \15143 , \15144 , \15145 , \15146 ,
         \15147 , \15148 , \15149 , \15150 , \15151 , \15152 , \15153 , \15154 , \15155 , \15156 ,
         \15157 , \15158 , \15159 , \15160 , \15161 , \15162 , \15163 , \15164 , \15165 , \15166 ,
         \15167 , \15168 , \15169 , \15170 , \15171 , \15172 , \15173 , \15174 , \15175 , \15176 ,
         \15177 , \15178 , \15179 , \15180 , \15181 , \15182 , \15183 , \15184 , \15185 , \15186 ,
         \15187_nG6592 , \15188 , \15189 , \15190 , \15191 , \15192 , \15193 , \15194 , \15195 , \15196 ,
         \15197 , \15198 , \15199 , \15200 , \15201 , \15202 , \15203 , \15204 , \15205 , \15206 ,
         \15207 , \15208 , \15209 , \15210 , \15211 , \15212 , \15213 , \15214 , \15215 , \15216 ,
         \15217 , \15218 , \15219 , \15220 , \15221 , \15222 , \15223 , \15224 , \15225 , \15226 ,
         \15227 , \15228 , \15229 , \15230 , \15231 , \15232 , \15233 , \15234 , \15235 , \15236 ,
         \15237 , \15238 , \15239 , \15240 , \15241 , \15242 , \15243 , \15244 , \15245 , \15246 ,
         \15247 , \15248 , \15249 , \15250 , \15251 , \15252 , \15253 , \15254 , \15255 , \15256 ,
         \15257 , \15258 , \15259 , \15260 , \15261 , \15262 , \15263 , \15264 , \15265 , \15266 ,
         \15267 , \15268 , \15269 , \15270 , \15271 , \15272 , \15273 , \15274 , \15275 , \15276 ,
         \15277 , \15278 , \15279 , \15280 , \15281 , \15282 , \15283 , \15284 , \15285 , \15286 ,
         \15287 , \15288 , \15289 , \15290 , \15291 , \15292 , \15293 , \15294 , \15295 , \15296 ,
         \15297 , \15298 , \15299 , \15300 , \15301 , \15302 , \15303 , \15304 , \15305 , \15306 ,
         \15307 , \15308 , \15309 , \15310 , \15311 , \15312 , \15313 , \15314 , \15315 , \15316 ,
         \15317 , \15318 , \15319_nG6593 , \15320_nG6594 , \15321 , \15322 , \15323 , \15324 , \15325 , \15326 ,
         \15327 , \15328 , \15329 , \15330_nG4e2b , \15331_nG4eaf , \15332_nG4eb0 , \15333 , \15334 , \15335 , \15336 ,
         \15337 , \15338 , \15339 , \15340 , \15341 , \15342 , \15343 , \15344 , \15345 , \15346 ,
         \15347 , \15348 , \15349 , \15350 , \15351 , \15352 , \15353 , \15354 , \15355 , \15356 ,
         \15357 , \15358 , \15359 , \15360 , \15361 , \15362 , \15363 , \15364 , \15365 , \15366 ,
         \15367 , \15368 , \15369 , \15370 , \15371 , \15372 , \15373_nG9bf3 , \15374 , \15375 , \15376 ,
         \15377 , \15378 , \15379 , \15380 , \15381 , \15382 , \15383 , \15384 , \15385 , \15386 ,
         \15387 , \15388 , \15389 , \15390 , \15391 , \15392 , \15393 , \15394 , \15395 , \15396 ,
         \15397 , \15398 , \15399 , \15400 , \15401 , \15402 , \15403 , \15404 , \15405 , \15406 ,
         \15407 , \15408 , \15409 , \15410 , \15411 , \15412 , \15413 , \15414 , \15415 , \15416 ,
         \15417 , \15418 , \15419 , \15420 , \15421 , \15422 , \15423 , \15424 , \15425 , \15426 ,
         \15427 , \15428 , \15429 , \15430 , \15431 , \15432 , \15433 , \15434 , \15435 , \15436 ,
         \15437 , \15438 , \15439 , \15440 , \15441 , \15442 , \15443 , \15444 , \15445 , \15446 ,
         \15447 , \15448 , \15449 , \15450 , \15451 , \15452 , \15453 , \15454 , \15455 , \15456 ,
         \15457 , \15458 , \15459 , \15460 , \15461 , \15462 , \15463 , \15464 , \15465 , \15466 ,
         \15467 , \15468 , \15469 , \15470 , \15471 , \15472 , \15473 , \15474 , \15475 , \15476 ,
         \15477 , \15478 , \15479 , \15480 , \15481 , \15482 , \15483 , \15484 , \15485 , \15486 ,
         \15487 , \15488 , \15489 , \15490 , \15491 , \15492 , \15493 , \15494 , \15495 , \15496 ,
         \15497 , \15498 , \15499 , \15500 , \15501 , \15502 , \15503 , \15504 , \15505 , \15506 ,
         \15507 , \15508 , \15509 , \15510 , \15511 , \15512 , \15513 , \15514 , \15515 , \15516 ,
         \15517 , \15518 , \15519 , \15520_nG2c99 , \15521 , \15522 , \15523 , \15524 , \15525 , \15526 ,
         \15527 , \15528 , \15529 , \15530 , \15531 , \15532 , \15533 , \15534 , \15535 , \15536 ,
         \15537 , \15538 , \15539 , \15540 , \15541 , \15542 , \15543 , \15544 , \15545 , \15546 ,
         \15547 , \15548 , \15549 , \15550 , \15551 , \15552 , \15553 , \15554 , \15555 , \15556 ,
         \15557 , \15558 , \15559 , \15560 , \15561 , \15562 , \15563 , \15564 , \15565 , \15566 ,
         \15567 , \15568 , \15569 , \15570 , \15571 , \15572 , \15573 , \15574 , \15575 , \15576 ,
         \15577 , \15578 , \15579 , \15580 , \15581 , \15582 , \15583 , \15584 , \15585 , \15586 ,
         \15587 , \15588 , \15589 , \15590 , \15591 , \15592 , \15593 , \15594 , \15595 , \15596 ,
         \15597 , \15598 , \15599 , \15600 , \15601 , \15602 , \15603 , \15604 , \15605 , \15606 ,
         \15607 , \15608 , \15609 , \15610 , \15611 , \15612 , \15613 , \15614 , \15615 , \15616 ,
         \15617 , \15618 , \15619 , \15620 , \15621 , \15622 , \15623 , \15624 , \15625 , \15626 ,
         \15627 , \15628 , \15629 , \15630 , \15631 , \15632 , \15633 , \15634 , \15635 , \15636 ,
         \15637 , \15638 , \15639 , \15640 , \15641 , \15642 , \15643 , \15644 , \15645 , \15646 ,
         \15647 , \15648 , \15649 , \15650 , \15651 , \15652 , \15653_nG3dc6 , \15654 , \15655 , \15656 ,
         \15657 , \15658 , \15659 , \15660 , \15661 , \15662 , \15663 , \15664 , \15665 , \15666 ,
         \15667 , \15668 , \15669 , \15670 , \15671 , \15672 , \15673 , \15674 , \15675 , \15676 ,
         \15677 , \15678 , \15679 , \15680 , \15681 , \15682 , \15683 , \15684 , \15685 , \15686 ,
         \15687 , \15688 , \15689 , \15690 , \15691 , \15692 , \15693 , \15694 , \15695 , \15696 ,
         \15697 , \15698 , \15699 , \15700 , \15701 , \15702 , \15703 , \15704 , \15705 , \15706 ,
         \15707 , \15708 , \15709 , \15710 , \15711 , \15712 , \15713 , \15714 , \15715 , \15716 ,
         \15717 , \15718 , \15719 , \15720 , \15721 , \15722 , \15723 , \15724 , \15725 , \15726 ,
         \15727 , \15728 , \15729 , \15730 , \15731 , \15732 , \15733 , \15734 , \15735 , \15736 ,
         \15737 , \15738 , \15739 , \15740 , \15741 , \15742 , \15743 , \15744 , \15745 , \15746 ,
         \15747 , \15748 , \15749 , \15750 , \15751 , \15752 , \15753 , \15754 , \15755 , \15756 ,
         \15757 , \15758 , \15759 , \15760 , \15761 , \15762 , \15763 , \15764 , \15765 , \15766 ,
         \15767 , \15768 , \15769 , \15770 , \15771 , \15772 , \15773 , \15774 , \15775 , \15776 ,
         \15777 , \15778 , \15779 , \15780 , \15781 , \15782 , \15783 , \15784 , \15785 , \15786 ,
         \15787_nG2d1e , \15788 , \15789 , \15790 , \15791 , \15792 , \15793 , \15794 , \15795 , \15796 ,
         \15797 , \15798 , \15799 , \15800 , \15801 , \15802 , \15803 , \15804 , \15805 , \15806 ,
         \15807 , \15808 , \15809 , \15810 , \15811 , \15812 , \15813 , \15814 , \15815 , \15816 ,
         \15817 , \15818 , \15819 , \15820 , \15821 , \15822 , \15823 , \15824 , \15825 , \15826 ,
         \15827 , \15828 , \15829 , \15830 , \15831 , \15832 , \15833 , \15834 , \15835 , \15836 ,
         \15837 , \15838 , \15839 , \15840 , \15841 , \15842 , \15843 , \15844 , \15845 , \15846 ,
         \15847 , \15848 , \15849 , \15850 , \15851 , \15852 , \15853 , \15854 , \15855 , \15856 ,
         \15857 , \15858 , \15859 , \15860 , \15861 , \15862 , \15863 , \15864 , \15865 , \15866 ,
         \15867 , \15868 , \15869 , \15870 , \15871 , \15872 , \15873 , \15874 , \15875 , \15876 ,
         \15877 , \15878 , \15879 , \15880 , \15881 , \15882 , \15883 , \15884 , \15885 , \15886 ,
         \15887 , \15888 , \15889 , \15890 , \15891 , \15892 , \15893 , \15894 , \15895 , \15896 ,
         \15897 , \15898 , \15899 , \15900 , \15901 , \15902 , \15903 , \15904 , \15905 , \15906 ,
         \15907 , \15908 , \15909 , \15910 , \15911 , \15912 , \15913 , \15914 , \15915 , \15916 ,
         \15917 , \15918 , \15919 , \15920_nG3e4b , \15921 , \15922 , \15923 , \15924 , \15925 , \15926 ,
         \15927 , \15928 , \15929 , \15930 , \15931_nG4436 , \15932 , \15933 , \15934_nG4439 , \15935 , \15936 ,
         \15937 , \15938 , \15939 , \15940 , \15941 , \15942 , \15943 , \15944 , \15945 , \15946 ,
         \15947 , \15948 , \15949 , \15950 , \15951 , \15952 , \15953 , \15954 , \15955 , \15956 ,
         \15957 , \15958 , \15959 , \15960 , \15961 , \15962 , \15963 , \15964 , \15965 , \15966 ,
         \15967 , \15968 , \15969 , \15970 , \15971 , \15972 , \15973 , \15974 , \15975 , \15976 ,
         \15977 , \15978 , \15979 , \15980 , \15981 , \15982 , \15983 , \15984 , \15985 , \15986 ,
         \15987 , \15988 , \15989 , \15990 , \15991 , \15992 , \15993 , \15994 , \15995 , \15996 ,
         \15997 , \15998 , \15999 , \16000 , \16001 , \16002 , \16003 , \16004 , \16005 , \16006 ,
         \16007 , \16008 , \16009 , \16010 , \16011 , \16012 , \16013 , \16014 , \16015 , \16016 ,
         \16017 , \16018 , \16019 , \16020 , \16021 , \16022 , \16023 , \16024 , \16025 , \16026 ,
         \16027 , \16028 , \16029 , \16030 , \16031 , \16032 , \16033 , \16034 , \16035 , \16036 ,
         \16037 , \16038 , \16039 , \16040 , \16041 , \16042 , \16043 , \16044 , \16045 , \16046 ,
         \16047 , \16048 , \16049 , \16050 , \16051 , \16052 , \16053 , \16054 , \16055 , \16056 ,
         \16057 , \16058 , \16059 , \16060 , \16061 , \16062 , \16063 , \16064 , \16065 , \16066 ,
         \16067 , \16068 , \16069 , \16070 , \16071 , \16072 , \16073 , \16074 , \16075 , \16076 ,
         \16077 , \16078 , \16079 , \16080 , \16081 , \16082 , \16083 , \16084 , \16085 , \16086 ,
         \16087 , \16088 , \16089 , \16090 , \16091 , \16092 , \16093 , \16094 , \16095 , \16096 ,
         \16097 , \16098 , \16099 , \16100 , \16101 , \16102 , \16103 , \16104 , \16105 , \16106 ,
         \16107 , \16108 , \16109 , \16110 , \16111 , \16112 , \16113 , \16114 , \16115 , \16116 ,
         \16117 , \16118 , \16119 , \16120 , \16121 , \16122 , \16123 , \16124 , \16125 , \16126 ,
         \16127 , \16128 , \16129 , \16130 , \16131 , \16132 , \16133_nG6595 , \16134 , \16135 , \16136 ,
         \16137 , \16138 , \16139 , \16140 , \16141 , \16142 , \16143 , \16144 , \16145 , \16146 ,
         \16147 , \16148 , \16149 , \16150 , \16151 , \16152 , \16153 , \16154 , \16155 , \16156 ,
         \16157 , \16158 , \16159 , \16160 , \16161 , \16162 , \16163 , \16164 , \16165 , \16166 ,
         \16167 , \16168 , \16169 , \16170 , \16171 , \16172 , \16173 , \16174 , \16175 , \16176 ,
         \16177 , \16178 , \16179 , \16180 , \16181 , \16182 , \16183 , \16184 , \16185 , \16186 ,
         \16187 , \16188 , \16189 , \16190 , \16191 , \16192 , \16193 , \16194 , \16195 , \16196 ,
         \16197 , \16198 , \16199 , \16200 , \16201 , \16202 , \16203 , \16204 , \16205 , \16206 ,
         \16207 , \16208 , \16209 , \16210 , \16211 , \16212 , \16213 , \16214 , \16215 , \16216 ,
         \16217 , \16218 , \16219 , \16220 , \16221 , \16222 , \16223 , \16224 , \16225 , \16226 ,
         \16227 , \16228 , \16229 , \16230 , \16231 , \16232 , \16233 , \16234 , \16235 , \16236 ,
         \16237 , \16238 , \16239 , \16240 , \16241 , \16242 , \16243 , \16244 , \16245 , \16246 ,
         \16247 , \16248 , \16249 , \16250 , \16251 , \16252 , \16253 , \16254 , \16255 , \16256 ,
         \16257 , \16258 , \16259 , \16260 , \16261 , \16262 , \16263 , \16264 , \16265_nG6596 , \16266_nG6597 ,
         \16267 , \16268 , \16269 , \16270 , \16271 , \16272 , \16273 , \16274 , \16275 , \16276 ,
         \16277 , \16278 , \16279 , \16280 , \16281 , \16282 , \16283 , \16284 , \16285 , \16286 ,
         \16287 , \16288 , \16289 , \16290 , \16291 , \16292 , \16293 , \16294 , \16295 , \16296 ,
         \16297_nG4f34 , \16298_nG4fb8 , \16299_nG4fb9 , \16300 , \16301 , \16302 , \16303 , \16304 , \16305 , \16306 ,
         \16307 , \16308 , \16309 , \16310 , \16311 , \16312 , \16313 , \16314 , \16315_nG9bf0 , \16316 ,
         \16317 , \16318 , \16319 , \16320 , \16321 , \16322 , \16323 , \16324 , \16325 , \16326 ,
         \16327 , \16328 , \16329 , \16330 , \16331 , \16332 , \16333 , \16334 , \16335 , \16336 ,
         \16337 , \16338 , \16339 , \16340 , \16341 , \16342 , \16343 , \16344 , \16345 , \16346 ,
         \16347 , \16348 , \16349 , \16350 , \16351 , \16352 , \16353 , \16354 , \16355 , \16356 ,
         \16357 , \16358 , \16359 , \16360 , \16361 , \16362 , \16363 , \16364 , \16365 , \16366 ,
         \16367 , \16368 , \16369 , \16370 , \16371 , \16372 , \16373 , \16374 , \16375 , \16376 ,
         \16377 , \16378 , \16379 , \16380 , \16381 , \16382 , \16383 , \16384 , \16385 , \16386 ,
         \16387 , \16388 , \16389 , \16390 , \16391 , \16392 , \16393 , \16394 , \16395 , \16396 ,
         \16397 , \16398 , \16399 , \16400 , \16401 , \16402 , \16403 , \16404 , \16405 , \16406 ,
         \16407 , \16408 , \16409 , \16410 , \16411 , \16412 , \16413 , \16414 , \16415 , \16416 ,
         \16417 , \16418 , \16419 , \16420 , \16421 , \16422 , \16423 , \16424 , \16425 , \16426 ,
         \16427 , \16428 , \16429 , \16430 , \16431 , \16432 , \16433 , \16434 , \16435 , \16436 ,
         \16437 , \16438 , \16439 , \16440 , \16441 , \16442 , \16443 , \16444 , \16445 , \16446 ,
         \16447 , \16448 , \16449 , \16450 , \16451 , \16452 , \16453 , \16454 , \16455 , \16456 ,
         \16457 , \16458 , \16459 , \16460 , \16461 , \16462 , \16463 , \16464 , \16465 , \16466 ,
         \16467 , \16468 , \16469 , \16470 , \16471 , \16472 , \16473 , \16474 , \16475 , \16476 ,
         \16477 , \16478 , \16479 , \16480 , \16481 , \16482 , \16483 , \16484 , \16485 , \16486 ,
         \16487 , \16488_nG503d , \16489 , \16490 , \16491 , \16492 , \16493 , \16494 , \16495 , \16496 ,
         \16497 , \16498 , \16499 , \16500 , \16501 , \16502 , \16503 , \16504 , \16505 , \16506 ,
         \16507 , \16508 , \16509 , \16510 , \16511 , \16512 , \16513 , \16514 , \16515 , \16516 ,
         \16517 , \16518 , \16519 , \16520 , \16521 , \16522 , \16523 , \16524 , \16525 , \16526 ,
         \16527 , \16528 , \16529 , \16530 , \16531 , \16532 , \16533 , \16534 , \16535 , \16536 ,
         \16537 , \16538 , \16539 , \16540 , \16541 , \16542 , \16543 , \16544 , \16545 , \16546 ,
         \16547 , \16548 , \16549 , \16550 , \16551 , \16552 , \16553 , \16554 , \16555 , \16556 ,
         \16557 , \16558 , \16559 , \16560 , \16561 , \16562 , \16563 , \16564 , \16565 , \16566 ,
         \16567 , \16568 , \16569 , \16570 , \16571 , \16572 , \16573 , \16574 , \16575 , \16576 ,
         \16577 , \16578 , \16579 , \16580 , \16581 , \16582 , \16583 , \16584 , \16585 , \16586 ,
         \16587 , \16588 , \16589 , \16590 , \16591 , \16592 , \16593 , \16594 , \16595 , \16596 ,
         \16597 , \16598 , \16599 , \16600 , \16601 , \16602 , \16603 , \16604 , \16605 , \16606 ,
         \16607 , \16608 , \16609 , \16610 , \16611 , \16612 , \16613 , \16614 , \16615 , \16616 ,
         \16617 , \16618 , \16619 , \16620_nG50c1 , \16621_nG50c2 , \16622 , \16623 , \16624 , \16625 , \16626 ,
         \16627 , \16628 , \16629 , \16630 , \16631 , \16632 , \16633 , \16634 , \16635 , \16636 ,
         \16637 , \16638 , \16639 , \16640 , \16641 , \16642 , \16643 , \16644 , \16645 , \16646 ,
         \16647 , \16648 , \16649 , \16650 , \16651 , \16652_nG6598 , \16653_nG6599 , \16654_nG659a , \16655 , \16656 ,
         \16657 , \16658 , \16659 , \16660 , \16661 , \16662 , \16663 , \16664 , \16665 , \16666 ,
         \16667 , \16668 , \16669 , \16670 , \16671 , \16672 , \16673 , \16674 , \16675 , \16676 ,
         \16677 , \16678 , \16679 , \16680_nG9bed , \16681 , \16682 , \16683 , \16684 , \16685 , \16686 ,
         \16687 , \16688 , \16689 , \16690 , \16691 , \16692 , \16693 , \16694 , \16695 , \16696 ,
         \16697 , \16698 , \16699 , \16700 , \16701 , \16702 , \16703 , \16704 , \16705 , \16706 ,
         \16707 , \16708 , \16709 , \16710 , \16711 , \16712 , \16713 , \16714 , \16715 , \16716 ,
         \16717 , \16718 , \16719 , \16720 , \16721 , \16722 , \16723 , \16724 , \16725 , \16726 ,
         \16727 , \16728 , \16729 , \16730 , \16731 , \16732 , \16733 , \16734 , \16735 , \16736 ,
         \16737 , \16738 , \16739 , \16740 , \16741 , \16742 , \16743 , \16744 , \16745 , \16746 ,
         \16747 , \16748 , \16749 , \16750 , \16751 , \16752 , \16753 , \16754 , \16755 , \16756 ,
         \16757 , \16758 , \16759 , \16760 , \16761 , \16762 , \16763 , \16764 , \16765 , \16766 ,
         \16767 , \16768 , \16769 , \16770 , \16771 , \16772 , \16773 , \16774 , \16775 , \16776 ,
         \16777 , \16778 , \16779 , \16780 , \16781 , \16782 , \16783 , \16784 , \16785 , \16786 ,
         \16787 , \16788 , \16789 , \16790 , \16791 , \16792 , \16793 , \16794 , \16795 , \16796 ,
         \16797 , \16798 , \16799 , \16800 , \16801 , \16802 , \16803 , \16804 , \16805 , \16806 ,
         \16807 , \16808 , \16809 , \16810 , \16811 , \16812 , \16813 , \16814 , \16815 , \16816 ,
         \16817 , \16818 , \16819 , \16820 , \16821 , \16822 , \16823 , \16824 , \16825 , \16826 ,
         \16827 , \16828 , \16829 , \16830 , \16831 , \16832 , \16833 , \16834 , \16835 , \16836 ,
         \16837 , \16838 , \16839 , \16840 , \16841 , \16842 , \16843 , \16844 , \16845 , \16846 ,
         \16847 , \16848 , \16849 , \16850 , \16851 , \16852 , \16853 , \16854 , \16855 , \16856 ,
         \16857 , \16858 , \16859 , \16860 , \16861 , \16862 , \16863 , \16864 , \16865 , \16866 ,
         \16867 , \16868 , \16869 , \16870 , \16871 , \16872 , \16873 , \16874 , \16875 , \16876 ,
         \16877_nG2b8f , \16878 , \16879 , \16880 , \16881 , \16882 , \16883 , \16884 , \16885 , \16886 ,
         \16887 , \16888 , \16889 , \16890 , \16891 , \16892 , \16893 , \16894 , \16895 , \16896 ,
         \16897 , \16898 , \16899 , \16900 , \16901 , \16902 , \16903 , \16904 , \16905 , \16906 ,
         \16907 , \16908 , \16909 , \16910 , \16911 , \16912 , \16913 , \16914 , \16915 , \16916 ,
         \16917 , \16918 , \16919 , \16920 , \16921 , \16922 , \16923 , \16924 , \16925 , \16926 ,
         \16927 , \16928 , \16929 , \16930 , \16931 , \16932 , \16933 , \16934 , \16935 , \16936 ,
         \16937 , \16938 , \16939 , \16940 , \16941 , \16942 , \16943 , \16944 , \16945 , \16946 ,
         \16947 , \16948 , \16949 , \16950 , \16951 , \16952 , \16953 , \16954 , \16955 , \16956 ,
         \16957 , \16958 , \16959 , \16960 , \16961 , \16962 , \16963 , \16964 , \16965 , \16966 ,
         \16967 , \16968 , \16969 , \16970 , \16971 , \16972 , \16973 , \16974 , \16975 , \16976 ,
         \16977 , \16978 , \16979 , \16980 , \16981 , \16982 , \16983 , \16984 , \16985 , \16986 ,
         \16987 , \16988 , \16989 , \16990 , \16991 , \16992 , \16993 , \16994 , \16995 , \16996 ,
         \16997 , \16998 , \16999 , \17000 , \17001 , \17002 , \17003 , \17004 , \17005 , \17006 ,
         \17007 , \17008 , \17009 , \17010_nG3cbc , \17011 , \17012 , \17013 , \17014 , \17015 , \17016 ,
         \17017 , \17018 , \17019 , \17020 , \17021 , \17022 , \17023 , \17024 , \17025 , \17026 ,
         \17027 , \17028 , \17029 , \17030 , \17031 , \17032 , \17033 , \17034 , \17035 , \17036 ,
         \17037 , \17038 , \17039 , \17040 , \17041 , \17042 , \17043 , \17044 , \17045 , \17046 ,
         \17047 , \17048 , \17049 , \17050 , \17051 , \17052 , \17053 , \17054 , \17055 , \17056 ,
         \17057 , \17058 , \17059 , \17060 , \17061 , \17062 , \17063 , \17064 , \17065 , \17066 ,
         \17067 , \17068 , \17069 , \17070 , \17071 , \17072 , \17073 , \17074 , \17075 , \17076 ,
         \17077 , \17078 , \17079 , \17080 , \17081 , \17082 , \17083 , \17084 , \17085 , \17086 ,
         \17087 , \17088 , \17089 , \17090 , \17091 , \17092 , \17093 , \17094 , \17095 , \17096 ,
         \17097 , \17098 , \17099 , \17100 , \17101 , \17102 , \17103 , \17104 , \17105 , \17106 ,
         \17107 , \17108 , \17109 , \17110 , \17111 , \17112 , \17113 , \17114 , \17115 , \17116 ,
         \17117 , \17118 , \17119 , \17120 , \17121 , \17122 , \17123 , \17124 , \17125 , \17126 ,
         \17127 , \17128 , \17129 , \17130 , \17131 , \17132 , \17133 , \17134 , \17135 , \17136 ,
         \17137 , \17138 , \17139 , \17140 , \17141 , \17142 , \17143 , \17144_nG2c14 , \17145 , \17146 ,
         \17147 , \17148 , \17149 , \17150 , \17151 , \17152 , \17153 , \17154 , \17155 , \17156 ,
         \17157 , \17158 , \17159 , \17160 , \17161 , \17162 , \17163 , \17164 , \17165 , \17166 ,
         \17167 , \17168 , \17169 , \17170 , \17171 , \17172 , \17173 , \17174 , \17175 , \17176 ,
         \17177 , \17178 , \17179 , \17180 , \17181 , \17182 , \17183 , \17184 , \17185 , \17186 ,
         \17187 , \17188 , \17189 , \17190 , \17191 , \17192 , \17193 , \17194 , \17195 , \17196 ,
         \17197 , \17198 , \17199 , \17200 , \17201 , \17202 , \17203 , \17204 , \17205 , \17206 ,
         \17207 , \17208 , \17209 , \17210 , \17211 , \17212 , \17213 , \17214 , \17215 , \17216 ,
         \17217 , \17218 , \17219 , \17220 , \17221 , \17222 , \17223 , \17224 , \17225 , \17226 ,
         \17227 , \17228 , \17229 , \17230 , \17231 , \17232 , \17233 , \17234 , \17235 , \17236 ,
         \17237 , \17238 , \17239 , \17240 , \17241 , \17242 , \17243 , \17244 , \17245 , \17246 ,
         \17247 , \17248 , \17249 , \17250 , \17251 , \17252 , \17253 , \17254 , \17255 , \17256 ,
         \17257 , \17258 , \17259 , \17260 , \17261 , \17262 , \17263 , \17264 , \17265 , \17266 ,
         \17267 , \17268 , \17269 , \17270 , \17271 , \17272 , \17273 , \17274 , \17275 , \17276 ,
         \17277_nG3d41 , \17278 , \17279 , \17280 , \17281 , \17282 , \17283 , \17284 , \17285 , \17286 ,
         \17287 , \17288_nG4430 , \17289 , \17290 , \17291_nG4433 , \17292 , \17293 , \17294 , \17295 , \17296 ,
         \17297 , \17298 , \17299 , \17300 , \17301 , \17302 , \17303 , \17304 , \17305 , \17306 ,
         \17307 , \17308 , \17309 , \17310 , \17311 , \17312 , \17313 , \17314 , \17315 , \17316 ,
         \17317 , \17318 , \17319 , \17320 , \17321 , \17322 , \17323 , \17324 , \17325 , \17326 ,
         \17327 , \17328 , \17329 , \17330 , \17331 , \17332 , \17333 , \17334 , \17335 , \17336 ,
         \17337 , \17338 , \17339 , \17340 , \17341 , \17342 , \17343 , \17344 , \17345 , \17346 ,
         \17347 , \17348 , \17349 , \17350 , \17351 , \17352 , \17353 , \17354 , \17355 , \17356 ,
         \17357 , \17358 , \17359 , \17360 , \17361 , \17362 , \17363 , \17364 , \17365 , \17366 ,
         \17367 , \17368 , \17369 , \17370 , \17371 , \17372 , \17373 , \17374 , \17375 , \17376 ,
         \17377 , \17378 , \17379 , \17380 , \17381 , \17382 , \17383 , \17384 , \17385 , \17386 ,
         \17387 , \17388 , \17389 , \17390 , \17391 , \17392 , \17393 , \17394 , \17395 , \17396 ,
         \17397 , \17398 , \17399 , \17400 , \17401 , \17402 , \17403 , \17404 , \17405 , \17406 ,
         \17407 , \17408 , \17409 , \17410 , \17411 , \17412 , \17413 , \17414 , \17415 , \17416 ,
         \17417 , \17418 , \17419 , \17420 , \17421 , \17422 , \17423 , \17424 , \17425 , \17426 ,
         \17427 , \17428 , \17429 , \17430 , \17431 , \17432 , \17433 , \17434 , \17435 , \17436 ,
         \17437 , \17438 , \17439 , \17440 , \17441 , \17442 , \17443 , \17444 , \17445 , \17446 ,
         \17447 , \17448 , \17449 , \17450 , \17451 , \17452 , \17453 , \17454 , \17455 , \17456 ,
         \17457 , \17458 , \17459 , \17460 , \17461 , \17462 , \17463 , \17464 , \17465 , \17466 ,
         \17467 , \17468 , \17469 , \17470 , \17471 , \17472 , \17473 , \17474 , \17475 , \17476 ,
         \17477 , \17478 , \17479 , \17480 , \17481 , \17482 , \17483 , \17484 , \17485 , \17486 ,
         \17487 , \17488 , \17489 , \17490 , \17491 , \17492 , \17493_nG659b , \17494 , \17495 , \17496 ,
         \17497 , \17498 , \17499 , \17500 , \17501 , \17502 , \17503 , \17504 , \17505 , \17506 ,
         \17507 , \17508 , \17509 , \17510 , \17511 , \17512 , \17513 , \17514 , \17515 , \17516 ,
         \17517 , \17518 , \17519 , \17520 , \17521 , \17522 , \17523 , \17524 , \17525 , \17526 ,
         \17527 , \17528 , \17529 , \17530 , \17531 , \17532 , \17533 , \17534 , \17535 , \17536 ,
         \17537 , \17538 , \17539 , \17540 , \17541 , \17542 , \17543 , \17544 , \17545 , \17546 ,
         \17547 , \17548 , \17549 , \17550 , \17551 , \17552 , \17553 , \17554 , \17555 , \17556 ,
         \17557 , \17558 , \17559 , \17560 , \17561 , \17562 , \17563 , \17564 , \17565 , \17566 ,
         \17567 , \17568 , \17569 , \17570 , \17571 , \17572 , \17573 , \17574 , \17575 , \17576 ,
         \17577 , \17578 , \17579 , \17580 , \17581 , \17582 , \17583 , \17584 , \17585 , \17586 ,
         \17587 , \17588 , \17589 , \17590 , \17591 , \17592 , \17593 , \17594 , \17595 , \17596 ,
         \17597 , \17598 , \17599 , \17600 , \17601 , \17602 , \17603 , \17604 , \17605 , \17606 ,
         \17607 , \17608 , \17609 , \17610 , \17611 , \17612 , \17613 , \17614 , \17615 , \17616 ,
         \17617 , \17618 , \17619 , \17620 , \17621 , \17622 , \17623 , \17624 , \17625_nG659c , \17626_nG659d ,
         \17627 , \17628 , \17629 , \17630 , \17631 , \17632 , \17633 , \17634 , \17635 , \17636 ,
         \17637 , \17638 , \17639 , \17640 , \17641 , \17642 , \17643 , \17644 , \17645 , \17646 ,
         \17647 , \17648 , \17649 , \17650 , \17651_nG5146 , \17652_nG51ca , \17653_nG51cb , \17654 , \17655 , \17656 ,
         \17657 , \17658 , \17659 , \17660 , \17661 , \17662 , \17663 , \17664 , \17665_nG9bea , \17666 ,
         \17667 , \17668 , \17669 , \17670 , \17671 , \17672 , \17673 , \17674 , \17675 , \17676 ,
         \17677 , \17678 , \17679 , \17680 , \17681 , \17682 , \17683 , \17684 , \17685 , \17686 ,
         \17687 , \17688 , \17689 , \17690 , \17691 , \17692 , \17693 , \17694 , \17695 , \17696 ,
         \17697 , \17698 , \17699 , \17700 , \17701 , \17702 , \17703 , \17704 , \17705 , \17706 ,
         \17707 , \17708 , \17709 , \17710 , \17711 , \17712 , \17713 , \17714 , \17715 , \17716 ,
         \17717 , \17718 , \17719 , \17720 , \17721 , \17722 , \17723 , \17724 , \17725 , \17726 ,
         \17727 , \17728 , \17729 , \17730 , \17731 , \17732 , \17733 , \17734 , \17735 , \17736 ,
         \17737 , \17738 , \17739 , \17740 , \17741 , \17742 , \17743 , \17744 , \17745 , \17746 ,
         \17747 , \17748 , \17749 , \17750 , \17751 , \17752 , \17753 , \17754 , \17755 , \17756 ,
         \17757 , \17758 , \17759 , \17760 , \17761 , \17762 , \17763 , \17764 , \17765 , \17766 ,
         \17767 , \17768 , \17769 , \17770 , \17771 , \17772 , \17773 , \17774 , \17775 , \17776 ,
         \17777 , \17778 , \17779 , \17780 , \17781 , \17782 , \17783 , \17784 , \17785 , \17786 ,
         \17787 , \17788 , \17789 , \17790 , \17791 , \17792 , \17793 , \17794 , \17795 , \17796 ,
         \17797 , \17798 , \17799 , \17800 , \17801 , \17802 , \17803 , \17804 , \17805 , \17806 ,
         \17807 , \17808 , \17809 , \17810 , \17811 , \17812 , \17813 , \17814 , \17815 , \17816 ,
         \17817 , \17818 , \17819 , \17820 , \17821 , \17822 , \17823 , \17824 , \17825 , \17826 ,
         \17827 , \17828 , \17829 , \17830 , \17831 , \17832 , \17833 , \17834 , \17835 , \17836 ,
         \17837 , \17838 , \17839 , \17840 , \17841 , \17842 , \17843 , \17844 , \17845 , \17846 ,
         \17847 , \17848 , \17849 , \17850 , \17851 , \17852 , \17853 , \17854 , \17855 , \17856 ,
         \17857 , \17858 , \17859 , \17860 , \17861 , \17862 , \17863 , \17864 , \17865 , \17866 ,
         \17867 , \17868 , \17869 , \17870 , \17871 , \17872 , \17873 , \17874 , \17875 , \17876 ,
         \17877 , \17878 , \17879 , \17880 , \17881 , \17882 , \17883 , \17884 , \17885 , \17886 ,
         \17887 , \17888 , \17889 , \17890 , \17891 , \17892 , \17893 , \17894 , \17895 , \17896 ,
         \17897 , \17898 , \17899 , \17900 , \17901_nG659e , \17902 , \17903 , \17904 , \17905 , \17906 ,
         \17907 , \17908 , \17909 , \17910 , \17911 , \17912 , \17913 , \17914 , \17915 , \17916 ,
         \17917 , \17918 , \17919 , \17920 , \17921 , \17922 , \17923 , \17924 , \17925 , \17926 ,
         \17927 , \17928 , \17929 , \17930 , \17931 , \17932 , \17933 , \17934 , \17935 , \17936 ,
         \17937 , \17938 , \17939 , \17940 , \17941 , \17942 , \17943 , \17944 , \17945 , \17946 ,
         \17947 , \17948 , \17949 , \17950 , \17951 , \17952 , \17953 , \17954 , \17955 , \17956 ,
         \17957 , \17958 , \17959 , \17960 , \17961 , \17962 , \17963 , \17964 , \17965 , \17966 ,
         \17967 , \17968 , \17969 , \17970 , \17971 , \17972 , \17973 , \17974 , \17975 , \17976 ,
         \17977 , \17978 , \17979 , \17980 , \17981 , \17982 , \17983 , \17984 , \17985 , \17986 ,
         \17987 , \17988 , \17989 , \17990 , \17991 , \17992 , \17993 , \17994 , \17995 , \17996 ,
         \17997 , \17998 , \17999 , \18000 , \18001 , \18002 , \18003 , \18004 , \18005 , \18006 ,
         \18007 , \18008 , \18009 , \18010 , \18011 , \18012 , \18013 , \18014 , \18015 , \18016 ,
         \18017 , \18018 , \18019 , \18020 , \18021 , \18022 , \18023 , \18024 , \18025 , \18026 ,
         \18027 , \18028 , \18029 , \18030 , \18031 , \18032 , \18033_nG659f , \18034_nG65a0 , \18035 , \18036 ,
         \18037 , \18038 , \18039 , \18040_nG524f , \18041_nG52d3 , \18042_nG52d4 , \18043 , \18044 , \18045 , \18046 ,
         \18047 , \18048 , \18049 , \18050 , \18051 , \18052 , \18053 , \18054 , \18055 , \18056 ,
         \18057 , \18058 , \18059 , \18060 , \18061 , \18062 , \18063 , \18064 , \18065 , \18066 ,
         \18067 , \18068 , \18069 , \18070 , \18071 , \18072 , \18073 , \18074 , \18075 , \18076 ,
         \18077 , \18078 , \18079 , \18080 , \18081 , \18082 , \18083 , \18084 , \18085 , \18086 ,
         \18087 , \18088 , \18089 , \18090 , \18091 , \18092 , \18093 , \18094 , \18095 , \18096 ,
         \18097 , \18098 , \18099 , \18100 , \18101 , \18102 , \18103 , \18104 , \18105 , \18106 ,
         \18107_nG9be7 , \18108 , \18109 , \18110 , \18111 , \18112 , \18113 , \18114 , \18115 , \18116 ,
         \18117 , \18118 , \18119 , \18120 , \18121 , \18122 , \18123 , \18124 , \18125 , \18126 ,
         \18127 , \18128 , \18129 , \18130 , \18131 , \18132 , \18133 , \18134 , \18135 , \18136 ,
         \18137 , \18138 , \18139 , \18140 , \18141 , \18142 , \18143 , \18144 , \18145 , \18146 ,
         \18147 , \18148 , \18149 , \18150 , \18151 , \18152 , \18153 , \18154 , \18155 , \18156 ,
         \18157 , \18158 , \18159 , \18160 , \18161 , \18162 , \18163 , \18164 , \18165 , \18166 ,
         \18167 , \18168 , \18169 , \18170 , \18171 , \18172 , \18173 , \18174 , \18175 , \18176 ,
         \18177 , \18178 , \18179 , \18180 , \18181 , \18182 , \18183 , \18184 , \18185 , \18186 ,
         \18187 , \18188 , \18189 , \18190 , \18191 , \18192 , \18193 , \18194 , \18195 , \18196 ,
         \18197 , \18198 , \18199 , \18200 , \18201 , \18202 , \18203 , \18204 , \18205 , \18206 ,
         \18207 , \18208 , \18209 , \18210 , \18211 , \18212 , \18213 , \18214 , \18215 , \18216 ,
         \18217 , \18218 , \18219 , \18220 , \18221 , \18222 , \18223 , \18224 , \18225 , \18226 ,
         \18227 , \18228 , \18229 , \18230 , \18231 , \18232 , \18233 , \18234 , \18235 , \18236 ,
         \18237 , \18238 , \18239 , \18240 , \18241 , \18242 , \18243 , \18244 , \18245 , \18246 ,
         \18247 , \18248 , \18249 , \18250 , \18251 , \18252 , \18253 , \18254 , \18255 , \18256 ,
         \18257 , \18258 , \18259 , \18260 , \18261 , \18262 , \18263 , \18264 , \18265 , \18266 ,
         \18267 , \18268 , \18269 , \18270 , \18271 , \18272 , \18273 , \18274 , \18275 , \18276 ,
         \18277 , \18278 , \18279 , \18280 , \18281 , \18282_nG2a85 , \18283 , \18284 , \18285 , \18286 ,
         \18287 , \18288 , \18289 , \18290 , \18291 , \18292 , \18293 , \18294 , \18295 , \18296 ,
         \18297 , \18298 , \18299 , \18300 , \18301 , \18302 , \18303 , \18304 , \18305 , \18306 ,
         \18307 , \18308 , \18309 , \18310 , \18311 , \18312 , \18313 , \18314 , \18315 , \18316 ,
         \18317 , \18318 , \18319 , \18320 , \18321 , \18322 , \18323 , \18324 , \18325 , \18326 ,
         \18327 , \18328 , \18329 , \18330 , \18331 , \18332 , \18333 , \18334 , \18335 , \18336 ,
         \18337 , \18338 , \18339 , \18340 , \18341 , \18342 , \18343 , \18344 , \18345 , \18346 ,
         \18347 , \18348 , \18349 , \18350 , \18351 , \18352 , \18353 , \18354 , \18355 , \18356 ,
         \18357 , \18358 , \18359 , \18360 , \18361 , \18362 , \18363 , \18364 , \18365 , \18366 ,
         \18367 , \18368 , \18369 , \18370 , \18371 , \18372 , \18373 , \18374 , \18375 , \18376 ,
         \18377 , \18378 , \18379 , \18380 , \18381 , \18382 , \18383 , \18384 , \18385 , \18386 ,
         \18387 , \18388 , \18389 , \18390 , \18391 , \18392 , \18393 , \18394 , \18395 , \18396 ,
         \18397 , \18398 , \18399 , \18400 , \18401 , \18402 , \18403 , \18404 , \18405 , \18406 ,
         \18407 , \18408 , \18409 , \18410 , \18411 , \18412 , \18413 , \18414 , \18415_nG3bb2 , \18416 ,
         \18417 , \18418 , \18419 , \18420 , \18421 , \18422 , \18423 , \18424 , \18425 , \18426 ,
         \18427 , \18428 , \18429 , \18430 , \18431 , \18432 , \18433 , \18434 , \18435 , \18436 ,
         \18437 , \18438 , \18439 , \18440 , \18441 , \18442 , \18443 , \18444 , \18445 , \18446 ,
         \18447 , \18448 , \18449 , \18450 , \18451 , \18452 , \18453 , \18454 , \18455 , \18456 ,
         \18457 , \18458 , \18459 , \18460 , \18461 , \18462 , \18463 , \18464 , \18465 , \18466 ,
         \18467 , \18468 , \18469 , \18470 , \18471 , \18472 , \18473 , \18474 , \18475 , \18476 ,
         \18477 , \18478 , \18479 , \18480 , \18481 , \18482 , \18483 , \18484 , \18485 , \18486 ,
         \18487 , \18488 , \18489 , \18490 , \18491 , \18492 , \18493 , \18494 , \18495 , \18496 ,
         \18497 , \18498 , \18499 , \18500 , \18501 , \18502 , \18503 , \18504 , \18505 , \18506 ,
         \18507 , \18508 , \18509 , \18510 , \18511 , \18512 , \18513 , \18514 , \18515 , \18516 ,
         \18517 , \18518 , \18519 , \18520 , \18521 , \18522 , \18523 , \18524 , \18525 , \18526 ,
         \18527 , \18528 , \18529 , \18530 , \18531 , \18532 , \18533 , \18534 , \18535 , \18536 ,
         \18537 , \18538 , \18539 , \18540 , \18541 , \18542 , \18543 , \18544 , \18545 , \18546 ,
         \18547 , \18548 , \18549_nG2b0a , \18550 , \18551 , \18552 , \18553 , \18554 , \18555 , \18556 ,
         \18557 , \18558 , \18559 , \18560 , \18561 , \18562 , \18563 , \18564 , \18565 , \18566 ,
         \18567 , \18568 , \18569 , \18570 , \18571 , \18572 , \18573 , \18574 , \18575 , \18576 ,
         \18577 , \18578 , \18579 , \18580 , \18581 , \18582 , \18583 , \18584 , \18585 , \18586 ,
         \18587 , \18588 , \18589 , \18590 , \18591 , \18592 , \18593 , \18594 , \18595 , \18596 ,
         \18597 , \18598 , \18599 , \18600 , \18601 , \18602 , \18603 , \18604 , \18605 , \18606 ,
         \18607 , \18608 , \18609 , \18610 , \18611 , \18612 , \18613 , \18614 , \18615 , \18616 ,
         \18617 , \18618 , \18619 , \18620 , \18621 , \18622 , \18623 , \18624 , \18625 , \18626 ,
         \18627 , \18628 , \18629 , \18630 , \18631 , \18632 , \18633 , \18634 , \18635 , \18636 ,
         \18637 , \18638 , \18639 , \18640 , \18641 , \18642 , \18643 , \18644 , \18645 , \18646 ,
         \18647 , \18648 , \18649 , \18650 , \18651 , \18652 , \18653 , \18654 , \18655 , \18656 ,
         \18657 , \18658 , \18659 , \18660 , \18661 , \18662 , \18663 , \18664 , \18665 , \18666 ,
         \18667 , \18668 , \18669 , \18670 , \18671 , \18672 , \18673 , \18674 , \18675 , \18676 ,
         \18677 , \18678 , \18679 , \18680 , \18681 , \18682_nG3c37 , \18683 , \18684 , \18685 , \18686 ,
         \18687 , \18688 , \18689 , \18690 , \18691 , \18692 , \18693_nG442a , \18694 , \18695 , \18696_nG442d ,
         \18697 , \18698 , \18699 , \18700 , \18701 , \18702 , \18703 , \18704 , \18705 , \18706 ,
         \18707 , \18708 , \18709 , \18710 , \18711 , \18712 , \18713 , \18714 , \18715 , \18716 ,
         \18717 , \18718 , \18719 , \18720 , \18721 , \18722 , \18723 , \18724 , \18725 , \18726 ,
         \18727 , \18728 , \18729 , \18730 , \18731 , \18732 , \18733 , \18734 , \18735 , \18736 ,
         \18737 , \18738 , \18739 , \18740 , \18741 , \18742 , \18743 , \18744 , \18745 , \18746 ,
         \18747 , \18748 , \18749 , \18750 , \18751 , \18752 , \18753 , \18754 , \18755 , \18756 ,
         \18757 , \18758 , \18759 , \18760 , \18761 , \18762 , \18763 , \18764 , \18765 , \18766 ,
         \18767 , \18768 , \18769 , \18770 , \18771 , \18772 , \18773 , \18774 , \18775 , \18776 ,
         \18777 , \18778 , \18779 , \18780 , \18781 , \18782 , \18783 , \18784 , \18785 , \18786 ,
         \18787 , \18788 , \18789 , \18790 , \18791 , \18792 , \18793 , \18794 , \18795 , \18796 ,
         \18797 , \18798 , \18799 , \18800 , \18801 , \18802 , \18803 , \18804 , \18805 , \18806 ,
         \18807 , \18808 , \18809 , \18810 , \18811 , \18812 , \18813 , \18814 , \18815 , \18816 ,
         \18817 , \18818 , \18819 , \18820 , \18821 , \18822 , \18823 , \18824 , \18825 , \18826 ,
         \18827 , \18828 , \18829 , \18830 , \18831 , \18832 , \18833 , \18834 , \18835 , \18836 ,
         \18837 , \18838 , \18839 , \18840 , \18841 , \18842 , \18843 , \18844 , \18845 , \18846 ,
         \18847 , \18848 , \18849 , \18850 , \18851 , \18852 , \18853 , \18854 , \18855 , \18856 ,
         \18857 , \18858 , \18859 , \18860 , \18861 , \18862 , \18863 , \18864 , \18865 , \18866 ,
         \18867 , \18868 , \18869 , \18870 , \18871 , \18872 , \18873 , \18874 , \18875 , \18876 ,
         \18877 , \18878 , \18879 , \18880 , \18881 , \18882 , \18883 , \18884 , \18885 , \18886 ,
         \18887 , \18888 , \18889 , \18890 , \18891 , \18892 , \18893 , \18894 , \18895 , \18896 ,
         \18897 , \18898_nG65a1 , \18899 , \18900 , \18901 , \18902 , \18903 , \18904 , \18905 , \18906 ,
         \18907 , \18908 , \18909 , \18910 , \18911 , \18912 , \18913 , \18914 , \18915 , \18916 ,
         \18917 , \18918 , \18919 , \18920 , \18921 , \18922 , \18923 , \18924 , \18925 , \18926 ,
         \18927 , \18928 , \18929 , \18930 , \18931 , \18932 , \18933 , \18934 , \18935 , \18936 ,
         \18937 , \18938 , \18939 , \18940 , \18941 , \18942 , \18943 , \18944 , \18945 , \18946 ,
         \18947 , \18948 , \18949 , \18950 , \18951 , \18952 , \18953 , \18954 , \18955 , \18956 ,
         \18957 , \18958 , \18959 , \18960 , \18961 , \18962 , \18963 , \18964 , \18965 , \18966 ,
         \18967 , \18968 , \18969 , \18970 , \18971 , \18972 , \18973 , \18974 , \18975 , \18976 ,
         \18977 , \18978 , \18979 , \18980 , \18981 , \18982 , \18983 , \18984 , \18985 , \18986 ,
         \18987 , \18988 , \18989 , \18990 , \18991 , \18992 , \18993 , \18994 , \18995 , \18996 ,
         \18997 , \18998 , \18999 , \19000 , \19001 , \19002 , \19003 , \19004 , \19005 , \19006 ,
         \19007 , \19008 , \19009 , \19010 , \19011 , \19012 , \19013 , \19014 , \19015 , \19016 ,
         \19017 , \19018 , \19019 , \19020 , \19021 , \19022 , \19023 , \19024 , \19025 , \19026 ,
         \19027 , \19028 , \19029 , \19030_nG65a2 , \19031_nG65a3 , \19032 , \19033 , \19034 , \19035 , \19036 ,
         \19037 , \19038 , \19039 , \19040 , \19041_nG5358 , \19042_nG53dc , \19043_nG53dd , \19044 , \19045 , \19046 ,
         \19047 , \19048 , \19049 , \19050 , \19051 , \19052 , \19053 , \19054 , \19055 , \19056 ,
         \19057 , \19058 , \19059 , \19060 , \19061 , \19062 , \19063 , \19064 , \19065 , \19066 ,
         \19067 , \19068 , \19069 , \19070 , \19071 , \19072 , \19073 , \19074 , \19075 , \19076 ,
         \19077 , \19078 , \19079 , \19080 , \19081 , \19082 , \19083 , \19084 , \19085 , \19086 ,
         \19087 , \19088 , \19089 , \19090 , \19091_nG9be4 , \19092 , \19093 , \19094 , \19095 , \19096 ,
         \19097 , \19098 , \19099 , \19100 , \19101 , \19102 , \19103 , \19104 , \19105 , \19106 ,
         \19107 , \19108 , \19109 , \19110 , \19111 , \19112 , \19113 , \19114 , \19115 , \19116 ,
         \19117 , \19118 , \19119 , \19120 , \19121 , \19122 , \19123 , \19124 , \19125 , \19126 ,
         \19127 , \19128 , \19129 , \19130 , \19131 , \19132 , \19133 , \19134 , \19135 , \19136 ,
         \19137 , \19138 , \19139 , \19140 , \19141 , \19142 , \19143 , \19144 , \19145 , \19146 ,
         \19147 , \19148 , \19149 , \19150 , \19151 , \19152 , \19153 , \19154 , \19155 , \19156 ,
         \19157 , \19158 , \19159 , \19160 , \19161 , \19162 , \19163 , \19164 , \19165 , \19166 ,
         \19167 , \19168 , \19169 , \19170 , \19171 , \19172 , \19173 , \19174 , \19175 , \19176 ,
         \19177 , \19178 , \19179 , \19180 , \19181 , \19182 , \19183 , \19184 , \19185 , \19186 ,
         \19187 , \19188 , \19189 , \19190 , \19191 , \19192 , \19193 , \19194 , \19195 , \19196 ,
         \19197 , \19198 , \19199 , \19200 , \19201 , \19202 , \19203 , \19204 , \19205 , \19206 ,
         \19207 , \19208 , \19209 , \19210 , \19211 , \19212 , \19213 , \19214 , \19215 , \19216 ,
         \19217 , \19218 , \19219 , \19220 , \19221 , \19222 , \19223 , \19224 , \19225 , \19226 ,
         \19227 , \19228 , \19229 , \19230 , \19231 , \19232 , \19233 , \19234 , \19235 , \19236 ,
         \19237 , \19238 , \19239 , \19240 , \19241 , \19242 , \19243 , \19244 , \19245 , \19246 ,
         \19247 , \19248 , \19249 , \19250 , \19251 , \19252 , \19253 , \19254 , \19255 , \19256 ,
         \19257 , \19258 , \19259 , \19260 , \19261 , \19262 , \19263 , \19264 , \19265 , \19266 ,
         \19267 , \19268 , \19269 , \19270 , \19271 , \19272 , \19273 , \19274 , \19275 , \19276 ,
         \19277 , \19278 , \19279 , \19280 , \19281 , \19282 , \19283 , \19284 , \19285 , \19286 ,
         \19287 , \19288 , \19289 , \19290 , \19291 , \19292 , \19293 , \19294 , \19295 , \19296 ,
         \19297 , \19298 , \19299 , \19300 , \19301 , \19302 , \19303 , \19304 , \19305 , \19306 ,
         \19307 , \19308 , \19309 , \19310 , \19311 , \19312 , \19313 , \19314 , \19315 , \19316 ,
         \19317 , \19318 , \19319 , \19320 , \19321 , \19322 , \19323 , \19324 , \19325 , \19326 ,
         \19327 , \19328 , \19329 , \19330 , \19331 , \19332 , \19333 , \19334 , \19335 , \19336 ,
         \19337 , \19338 , \19339 , \19340 , \19341 , \19342 , \19343 , \19344 , \19345 , \19346 ,
         \19347 , \19348 , \19349 , \19350 , \19351 , \19352 , \19353 , \19354 , \19355 , \19356 ,
         \19357 , \19358 , \19359 , \19360 , \19361 , \19362 , \19363 , \19364 , \19365 , \19366 ,
         \19367 , \19368 , \19369 , \19370 , \19371 , \19372 , \19373 , \19374 , \19375 , \19376 ,
         \19377 , \19378 , \19379 , \19380 , \19381 , \19382 , \19383 , \19384 , \19385 , \19386 ,
         \19387 , \19388 , \19389 , \19390 , \19391 , \19392 , \19393 , \19394 , \19395 , \19396 ,
         \19397_nG5461 , \19398 , \19399 , \19400 , \19401 , \19402 , \19403 , \19404 , \19405 , \19406 ,
         \19407 , \19408 , \19409 , \19410 , \19411 , \19412 , \19413 , \19414 , \19415 , \19416 ,
         \19417 , \19418 , \19419 , \19420 , \19421 , \19422 , \19423 , \19424 , \19425 , \19426 ,
         \19427 , \19428 , \19429 , \19430 , \19431 , \19432 , \19433 , \19434 , \19435 , \19436 ,
         \19437 , \19438 , \19439 , \19440 , \19441 , \19442 , \19443 , \19444 , \19445 , \19446 ,
         \19447 , \19448 , \19449 , \19450 , \19451 , \19452 , \19453 , \19454 , \19455 , \19456 ,
         \19457 , \19458 , \19459 , \19460 , \19461 , \19462 , \19463 , \19464 , \19465 , \19466 ,
         \19467 , \19468 , \19469 , \19470 , \19471 , \19472 , \19473 , \19474 , \19475 , \19476 ,
         \19477 , \19478 , \19479 , \19480 , \19481 , \19482 , \19483 , \19484 , \19485 , \19486 ,
         \19487 , \19488 , \19489 , \19490 , \19491 , \19492 , \19493 , \19494 , \19495 , \19496 ,
         \19497 , \19498 , \19499 , \19500 , \19501 , \19502 , \19503 , \19504 , \19505 , \19506 ,
         \19507 , \19508 , \19509 , \19510 , \19511 , \19512 , \19513 , \19514 , \19515 , \19516 ,
         \19517 , \19518 , \19519 , \19520 , \19521 , \19522 , \19523 , \19524 , \19525 , \19526 ,
         \19527 , \19528 , \19529_nG54e5 , \19530_nG54e6 , \19531 , \19532 , \19533 , \19534 , \19535 , \19536 ,
         \19537 , \19538 , \19539 , \19540 , \19541 , \19542 , \19543 , \19544 , \19545 , \19546 ,
         \19547 , \19548 , \19549 , \19550 , \19551 , \19552 , \19553 , \19554 , \19555_nG65a4 , \19556_nG65a5 ,
         \19557_nG65a6 , \19558 , \19559 , \19560 , \19561 , \19562 , \19563 , \19564 , \19565 , \19566 ,
         \19567 , \19568 , \19569 , \19570 , \19571 , \19572 , \19573 , \19574 , \19575 , \19576 ,
         \19577 , \19578 , \19579 , \19580 , \19581 , \19582 , \19583 , \19584 , \19585 , \19586_nG9be1 ,
         \19587 , \19588 , \19589 , \19590 , \19591 , \19592 , \19593 , \19594 , \19595 , \19596 ,
         \19597 , \19598 , \19599 , \19600 , \19601 , \19602 , \19603 , \19604 , \19605 , \19606 ,
         \19607 , \19608 , \19609 , \19610 , \19611 , \19612 , \19613 , \19614 , \19615 , \19616 ,
         \19617 , \19618 , \19619 , \19620 , \19621 , \19622 , \19623 , \19624 , \19625 , \19626 ,
         \19627 , \19628 , \19629 , \19630 , \19631 , \19632 , \19633 , \19634 , \19635 , \19636 ,
         \19637 , \19638 , \19639 , \19640 , \19641 , \19642 , \19643 , \19644 , \19645 , \19646 ,
         \19647 , \19648 , \19649 , \19650 , \19651 , \19652 , \19653 , \19654 , \19655 , \19656 ,
         \19657 , \19658 , \19659 , \19660 , \19661 , \19662 , \19663 , \19664 , \19665 , \19666 ,
         \19667 , \19668 , \19669 , \19670 , \19671 , \19672 , \19673 , \19674 , \19675 , \19676 ,
         \19677 , \19678 , \19679 , \19680 , \19681 , \19682 , \19683 , \19684 , \19685 , \19686 ,
         \19687 , \19688 , \19689 , \19690 , \19691 , \19692 , \19693 , \19694 , \19695 , \19696 ,
         \19697 , \19698 , \19699 , \19700 , \19701 , \19702 , \19703 , \19704 , \19705 , \19706 ,
         \19707 , \19708 , \19709 , \19710 , \19711 , \19712 , \19713 , \19714 , \19715 , \19716 ,
         \19717 , \19718 , \19719 , \19720 , \19721 , \19722 , \19723 , \19724 , \19725 , \19726 ,
         \19727 , \19728 , \19729 , \19730 , \19731 , \19732 , \19733 , \19734 , \19735_nG297b , \19736 ,
         \19737 , \19738 , \19739 , \19740 , \19741 , \19742 , \19743 , \19744 , \19745 , \19746 ,
         \19747 , \19748 , \19749 , \19750 , \19751 , \19752 , \19753 , \19754 , \19755 , \19756 ,
         \19757 , \19758 , \19759 , \19760 , \19761 , \19762 , \19763 , \19764 , \19765 , \19766 ,
         \19767 , \19768 , \19769 , \19770 , \19771 , \19772 , \19773 , \19774 , \19775 , \19776 ,
         \19777 , \19778 , \19779 , \19780 , \19781 , \19782 , \19783 , \19784 , \19785 , \19786 ,
         \19787 , \19788 , \19789 , \19790 , \19791 , \19792 , \19793 , \19794 , \19795 , \19796 ,
         \19797 , \19798 , \19799 , \19800 , \19801 , \19802 , \19803 , \19804 , \19805 , \19806 ,
         \19807 , \19808 , \19809 , \19810 , \19811 , \19812 , \19813 , \19814 , \19815 , \19816 ,
         \19817 , \19818 , \19819 , \19820 , \19821 , \19822 , \19823 , \19824 , \19825 , \19826 ,
         \19827 , \19828 , \19829 , \19830 , \19831 , \19832 , \19833 , \19834 , \19835 , \19836 ,
         \19837 , \19838 , \19839 , \19840 , \19841 , \19842 , \19843 , \19844 , \19845 , \19846 ,
         \19847 , \19848 , \19849 , \19850 , \19851 , \19852 , \19853 , \19854 , \19855 , \19856 ,
         \19857 , \19858 , \19859 , \19860 , \19861 , \19862 , \19863 , \19864 , \19865 , \19866 ,
         \19867 , \19868_nG3aa8 , \19869 , \19870 , \19871 , \19872 , \19873 , \19874 , \19875 , \19876 ,
         \19877 , \19878 , \19879 , \19880 , \19881 , \19882 , \19883 , \19884 , \19885 , \19886 ,
         \19887 , \19888 , \19889 , \19890 , \19891 , \19892 , \19893 , \19894 , \19895 , \19896 ,
         \19897 , \19898 , \19899 , \19900 , \19901 , \19902 , \19903 , \19904 , \19905 , \19906 ,
         \19907 , \19908 , \19909 , \19910 , \19911 , \19912 , \19913 , \19914 , \19915 , \19916 ,
         \19917 , \19918 , \19919 , \19920 , \19921 , \19922 , \19923 , \19924 , \19925 , \19926 ,
         \19927 , \19928 , \19929 , \19930 , \19931 , \19932 , \19933 , \19934 , \19935 , \19936 ,
         \19937 , \19938 , \19939 , \19940 , \19941 , \19942 , \19943 , \19944 , \19945 , \19946 ,
         \19947 , \19948 , \19949 , \19950 , \19951 , \19952 , \19953 , \19954 , \19955 , \19956 ,
         \19957 , \19958 , \19959 , \19960 , \19961 , \19962 , \19963 , \19964 , \19965 , \19966 ,
         \19967 , \19968 , \19969 , \19970 , \19971 , \19972 , \19973 , \19974 , \19975 , \19976 ,
         \19977 , \19978 , \19979 , \19980 , \19981 , \19982 , \19983 , \19984 , \19985 , \19986 ,
         \19987 , \19988 , \19989 , \19990 , \19991 , \19992 , \19993 , \19994 , \19995 , \19996 ,
         \19997 , \19998 , \19999 , \20000 , \20001 , \20002_nG2a00 , \20003 , \20004 , \20005 , \20006 ,
         \20007 , \20008 , \20009 , \20010 , \20011 , \20012 , \20013 , \20014 , \20015 , \20016 ,
         \20017 , \20018 , \20019 , \20020 , \20021 , \20022 , \20023 , \20024 , \20025 , \20026 ,
         \20027 , \20028 , \20029 , \20030 , \20031 , \20032 , \20033 , \20034 , \20035 , \20036 ,
         \20037 , \20038 , \20039 , \20040 , \20041 , \20042 , \20043 , \20044 , \20045 , \20046 ,
         \20047 , \20048 , \20049 , \20050 , \20051 , \20052 , \20053 , \20054 , \20055 , \20056 ,
         \20057 , \20058 , \20059 , \20060 , \20061 , \20062 , \20063 , \20064 , \20065 , \20066 ,
         \20067 , \20068 , \20069 , \20070 , \20071 , \20072 , \20073 , \20074 , \20075 , \20076 ,
         \20077 , \20078 , \20079 , \20080 , \20081 , \20082 , \20083 , \20084 , \20085 , \20086 ,
         \20087 , \20088 , \20089 , \20090 , \20091 , \20092 , \20093 , \20094 , \20095 , \20096 ,
         \20097 , \20098 , \20099 , \20100 , \20101 , \20102 , \20103 , \20104 , \20105 , \20106 ,
         \20107 , \20108 , \20109 , \20110 , \20111 , \20112 , \20113 , \20114 , \20115 , \20116 ,
         \20117 , \20118 , \20119 , \20120 , \20121 , \20122 , \20123 , \20124 , \20125 , \20126 ,
         \20127 , \20128 , \20129 , \20130 , \20131 , \20132 , \20133 , \20134 , \20135_nG3b2d , \20136 ,
         \20137 , \20138 , \20139 , \20140 , \20141 , \20142 , \20143 , \20144 , \20145 , \20146_nG4424 ,
         \20147 , \20148 , \20149_nG4427 , \20150 , \20151 , \20152 , \20153 , \20154 , \20155 , \20156 ,
         \20157 , \20158 , \20159 , \20160 , \20161 , \20162 , \20163 , \20164 , \20165 , \20166 ,
         \20167 , \20168 , \20169 , \20170 , \20171 , \20172 , \20173 , \20174 , \20175 , \20176 ,
         \20177 , \20178 , \20179 , \20180 , \20181 , \20182 , \20183 , \20184 , \20185 , \20186 ,
         \20187 , \20188 , \20189 , \20190 , \20191 , \20192 , \20193 , \20194 , \20195 , \20196 ,
         \20197 , \20198 , \20199 , \20200 , \20201 , \20202 , \20203 , \20204 , \20205 , \20206 ,
         \20207 , \20208 , \20209 , \20210 , \20211 , \20212 , \20213 , \20214 , \20215 , \20216 ,
         \20217 , \20218 , \20219 , \20220 , \20221 , \20222 , \20223 , \20224 , \20225 , \20226 ,
         \20227 , \20228 , \20229 , \20230 , \20231 , \20232 , \20233 , \20234 , \20235 , \20236 ,
         \20237 , \20238 , \20239 , \20240 , \20241 , \20242 , \20243 , \20244 , \20245 , \20246 ,
         \20247 , \20248 , \20249 , \20250 , \20251 , \20252 , \20253 , \20254 , \20255 , \20256 ,
         \20257 , \20258 , \20259 , \20260 , \20261 , \20262 , \20263 , \20264 , \20265 , \20266 ,
         \20267 , \20268 , \20269 , \20270 , \20271 , \20272 , \20273 , \20274 , \20275 , \20276 ,
         \20277 , \20278 , \20279 , \20280 , \20281 , \20282 , \20283 , \20284 , \20285 , \20286 ,
         \20287 , \20288 , \20289 , \20290 , \20291 , \20292 , \20293 , \20294 , \20295 , \20296 ,
         \20297 , \20298 , \20299 , \20300 , \20301 , \20302 , \20303 , \20304 , \20305 , \20306 ,
         \20307 , \20308 , \20309 , \20310 , \20311 , \20312 , \20313 , \20314 , \20315 , \20316 ,
         \20317 , \20318 , \20319 , \20320 , \20321 , \20322 , \20323 , \20324 , \20325 , \20326 ,
         \20327 , \20328 , \20329 , \20330 , \20331 , \20332 , \20333 , \20334 , \20335 , \20336 ,
         \20337 , \20338 , \20339 , \20340 , \20341 , \20342 , \20343 , \20344 , \20345 , \20346 ,
         \20347 , \20348 , \20349 , \20350 , \20351 , \20352 , \20353 , \20354 , \20355 , \20356 ,
         \20357 , \20358 , \20359 , \20360 , \20361 , \20362 , \20363 , \20364 , \20365 , \20366 ,
         \20367 , \20368 , \20369 , \20370 , \20371 , \20372 , \20373 , \20374 , \20375 , \20376 ,
         \20377 , \20378 , \20379 , \20380 , \20381 , \20382 , \20383 , \20384 , \20385 , \20386 ,
         \20387 , \20388 , \20389 , \20390 , \20391 , \20392 , \20393 , \20394 , \20395 , \20396 ,
         \20397 , \20398 , \20399 , \20400 , \20401 , \20402 , \20403 , \20404 , \20405 , \20406 ,
         \20407 , \20408 , \20409 , \20410_nG65a7 , \20411 , \20412 , \20413 , \20414 , \20415 , \20416 ,
         \20417 , \20418 , \20419 , \20420 , \20421 , \20422 , \20423 , \20424 , \20425 , \20426 ,
         \20427 , \20428 , \20429 , \20430 , \20431 , \20432 , \20433 , \20434 , \20435 , \20436 ,
         \20437 , \20438 , \20439 , \20440 , \20441 , \20442 , \20443 , \20444 , \20445 , \20446 ,
         \20447 , \20448 , \20449 , \20450 , \20451 , \20452 , \20453 , \20454 , \20455 , \20456 ,
         \20457 , \20458 , \20459 , \20460 , \20461 , \20462 , \20463 , \20464 , \20465 , \20466 ,
         \20467 , \20468 , \20469 , \20470 , \20471 , \20472 , \20473 , \20474 , \20475 , \20476 ,
         \20477 , \20478 , \20479 , \20480 , \20481 , \20482 , \20483 , \20484 , \20485 , \20486 ,
         \20487 , \20488 , \20489 , \20490 , \20491 , \20492 , \20493 , \20494 , \20495 , \20496 ,
         \20497 , \20498 , \20499 , \20500 , \20501 , \20502 , \20503 , \20504 , \20505 , \20506 ,
         \20507 , \20508 , \20509 , \20510 , \20511 , \20512 , \20513 , \20514 , \20515 , \20516 ,
         \20517 , \20518 , \20519 , \20520 , \20521 , \20522 , \20523 , \20524 , \20525 , \20526 ,
         \20527 , \20528 , \20529 , \20530 , \20531 , \20532 , \20533 , \20534 , \20535 , \20536 ,
         \20537 , \20538 , \20539 , \20540 , \20541 , \20542_nG65a8 , \20543_nG65a9 , \20544 , \20545 , \20546 ,
         \20547 , \20548 , \20549 , \20550 , \20551 , \20552 , \20553_nG556a , \20554_nG55ee , \20555_nG55ef , \20556 ,
         \20557 , \20558 , \20559 , \20560 , \20561 , \20562 , \20563 , \20564 , \20565 , \20566 ,
         \20567 , \20568 , \20569 , \20570 , \20571 , \20572 , \20573 , \20574 , \20575 , \20576 ,
         \20577 , \20578 , \20579 , \20580 , \20581 , \20582 , \20583 , \20584 , \20585 , \20586 ,
         \20587 , \20588 , \20589 , \20590 , \20591 , \20592 , \20593 , \20594 , \20595 , \20596 ,
         \20597 , \20598 , \20599 , \20600 , \20601 , \20602 , \20603 , \20604 , \20605 , \20606 ,
         \20607 , \20608_nG9bde , \20609 , \20610 , \20611 , \20612 , \20613 , \20614 , \20615 , \20616 ,
         \20617 , \20618 , \20619 , \20620 , \20621 , \20622 , \20623 , \20624 , \20625 , \20626 ,
         \20627 , \20628 , \20629 , \20630 , \20631 , \20632 , \20633 , \20634 , \20635 , \20636 ,
         \20637 , \20638 , \20639 , \20640 , \20641 , \20642 , \20643 , \20644 , \20645 , \20646 ,
         \20647 , \20648 , \20649 , \20650 , \20651 , \20652 , \20653 , \20654 , \20655 , \20656 ,
         \20657 , \20658 , \20659 , \20660 , \20661 , \20662 , \20663 , \20664 , \20665 , \20666 ,
         \20667 , \20668 , \20669 , \20670 , \20671 , \20672 , \20673 , \20674 , \20675 , \20676 ,
         \20677 , \20678 , \20679 , \20680 , \20681 , \20682 , \20683 , \20684 , \20685 , \20686 ,
         \20687 , \20688 , \20689 , \20690 , \20691 , \20692 , \20693 , \20694 , \20695 , \20696 ,
         \20697 , \20698 , \20699 , \20700 , \20701 , \20702 , \20703 , \20704 , \20705 , \20706 ,
         \20707 , \20708 , \20709 , \20710 , \20711 , \20712 , \20713 , \20714 , \20715 , \20716 ,
         \20717 , \20718 , \20719 , \20720 , \20721 , \20722 , \20723 , \20724 , \20725 , \20726 ,
         \20727 , \20728 , \20729 , \20730 , \20731 , \20732 , \20733 , \20734 , \20735 , \20736 ,
         \20737 , \20738 , \20739 , \20740 , \20741 , \20742 , \20743 , \20744 , \20745 , \20746 ,
         \20747 , \20748 , \20749 , \20750 , \20751 , \20752 , \20753 , \20754 , \20755 , \20756 ,
         \20757 , \20758 , \20759 , \20760 , \20761 , \20762 , \20763 , \20764 , \20765 , \20766 ,
         \20767 , \20768 , \20769 , \20770 , \20771 , \20772 , \20773 , \20774 , \20775 , \20776 ,
         \20777 , \20778 , \20779 , \20780 , \20781 , \20782 , \20783 , \20784 , \20785 , \20786 ,
         \20787 , \20788 , \20789 , \20790 , \20791 , \20792 , \20793 , \20794 , \20795 , \20796 ,
         \20797 , \20798 , \20799 , \20800 , \20801 , \20802 , \20803 , \20804 , \20805 , \20806 ,
         \20807 , \20808 , \20809 , \20810 , \20811 , \20812 , \20813 , \20814 , \20815 , \20816 ,
         \20817 , \20818 , \20819 , \20820 , \20821 , \20822 , \20823 , \20824 , \20825 , \20826 ,
         \20827 , \20828 , \20829 , \20830 , \20831 , \20832 , \20833 , \20834 , \20835 , \20836 ,
         \20837 , \20838 , \20839 , \20840 , \20841 , \20842 , \20843 , \20844 , \20845 , \20846 ,
         \20847 , \20848 , \20849 , \20850 , \20851 , \20852 , \20853 , \20854 , \20855 , \20856 ,
         \20857 , \20858 , \20859 , \20860 , \20861 , \20862 , \20863 , \20864 , \20865 , \20866 ,
         \20867 , \20868_nG5673 , \20869 , \20870 , \20871 , \20872 , \20873 , \20874 , \20875 , \20876 ,
         \20877 , \20878 , \20879 , \20880 , \20881 , \20882 , \20883 , \20884 , \20885 , \20886 ,
         \20887 , \20888 , \20889 , \20890 , \20891 , \20892 , \20893 , \20894 , \20895 , \20896 ,
         \20897 , \20898 , \20899 , \20900 , \20901 , \20902 , \20903 , \20904 , \20905 , \20906 ,
         \20907 , \20908 , \20909 , \20910 , \20911 , \20912 , \20913 , \20914 , \20915 , \20916 ,
         \20917 , \20918 , \20919 , \20920 , \20921 , \20922 , \20923 , \20924 , \20925 , \20926 ,
         \20927 , \20928 , \20929 , \20930 , \20931 , \20932 , \20933 , \20934 , \20935 , \20936 ,
         \20937 , \20938 , \20939 , \20940 , \20941 , \20942 , \20943 , \20944 , \20945 , \20946 ,
         \20947 , \20948 , \20949 , \20950 , \20951 , \20952 , \20953 , \20954 , \20955 , \20956 ,
         \20957 , \20958 , \20959 , \20960 , \20961 , \20962 , \20963 , \20964 , \20965 , \20966 ,
         \20967 , \20968 , \20969 , \20970 , \20971 , \20972 , \20973 , \20974 , \20975 , \20976 ,
         \20977 , \20978 , \20979 , \20980 , \20981 , \20982 , \20983 , \20984 , \20985 , \20986 ,
         \20987 , \20988 , \20989 , \20990 , \20991 , \20992 , \20993 , \20994 , \20995 , \20996 ,
         \20997 , \20998 , \20999 , \21000_nG56f7 , \21001_nG56f8 , \21002 , \21003 , \21004 , \21005 , \21006 ,
         \21007 , \21008 , \21009 , \21010 , \21011 , \21012 , \21013 , \21014 , \21015 , \21016 ,
         \21017 , \21018 , \21019 , \21020 , \21021 , \21022 , \21023 , \21024 , \21025 , \21026 ,
         \21027 , \21028 , \21029 , \21030_nG65aa , \21031_nG65ab , \21032_nG65ac , \21033 , \21034 , \21035 , \21036 ,
         \21037 , \21038 , \21039 , \21040 , \21041 , \21042 , \21043 , \21044 , \21045 , \21046 ,
         \21047 , \21048 , \21049 , \21050 , \21051 , \21052 , \21053 , \21054 , \21055 , \21056 ,
         \21057 , \21058 , \21059 , \21060 , \21061 , \21062 , \21063 , \21064 , \21065 , \21066 ,
         \21067 , \21068 , \21069 , \21070 , \21071 , \21072 , \21073 , \21074 , \21075 , \21076 ,
         \21077 , \21078 , \21079 , \21080 , \21081 , \21082 , \21083 , \21084 , \21085 , \21086_nG9bdb ,
         \21087 , \21088 , \21089 , \21090 , \21091 , \21092 , \21093 , \21094 , \21095 , \21096 ,
         \21097 , \21098 , \21099 , \21100 , \21101 , \21102 , \21103 , \21104 , \21105 , \21106 ,
         \21107 , \21108 , \21109 , \21110 , \21111 , \21112 , \21113 , \21114 , \21115 , \21116 ,
         \21117 , \21118 , \21119 , \21120 , \21121 , \21122 , \21123 , \21124 , \21125 , \21126 ,
         \21127 , \21128 , \21129 , \21130 , \21131 , \21132 , \21133 , \21134 , \21135 , \21136 ,
         \21137 , \21138 , \21139 , \21140 , \21141 , \21142 , \21143 , \21144 , \21145 , \21146 ,
         \21147 , \21148 , \21149 , \21150 , \21151 , \21152 , \21153 , \21154 , \21155 , \21156 ,
         \21157 , \21158 , \21159 , \21160 , \21161 , \21162 , \21163 , \21164 , \21165 , \21166 ,
         \21167 , \21168 , \21169 , \21170 , \21171 , \21172 , \21173 , \21174 , \21175 , \21176 ,
         \21177 , \21178 , \21179 , \21180 , \21181 , \21182 , \21183 , \21184 , \21185 , \21186 ,
         \21187 , \21188 , \21189 , \21190 , \21191 , \21192 , \21193 , \21194 , \21195 , \21196 ,
         \21197 , \21198 , \21199 , \21200 , \21201 , \21202 , \21203 , \21204 , \21205 , \21206 ,
         \21207 , \21208 , \21209 , \21210 , \21211 , \21212 , \21213 , \21214 , \21215 , \21216 ,
         \21217 , \21218 , \21219 , \21220 , \21221 , \21222 , \21223 , \21224 , \21225 , \21226 ,
         \21227 , \21228 , \21229 , \21230 , \21231 , \21232 , \21233 , \21234 , \21235 , \21236 ,
         \21237 , \21238_nG2871 , \21239 , \21240 , \21241 , \21242 , \21243 , \21244 , \21245 , \21246 ,
         \21247 , \21248 , \21249 , \21250 , \21251 , \21252 , \21253 , \21254 , \21255 , \21256 ,
         \21257 , \21258 , \21259 , \21260 , \21261 , \21262 , \21263 , \21264 , \21265 , \21266 ,
         \21267 , \21268 , \21269 , \21270 , \21271 , \21272 , \21273 , \21274 , \21275 , \21276 ,
         \21277 , \21278 , \21279 , \21280 , \21281 , \21282 , \21283 , \21284 , \21285 , \21286 ,
         \21287 , \21288 , \21289 , \21290 , \21291 , \21292 , \21293 , \21294 , \21295 , \21296 ,
         \21297 , \21298 , \21299 , \21300 , \21301 , \21302 , \21303 , \21304 , \21305 , \21306 ,
         \21307 , \21308 , \21309 , \21310 , \21311 , \21312 , \21313 , \21314 , \21315 , \21316 ,
         \21317 , \21318 , \21319 , \21320 , \21321 , \21322 , \21323 , \21324 , \21325 , \21326 ,
         \21327 , \21328 , \21329 , \21330 , \21331 , \21332 , \21333 , \21334 , \21335 , \21336 ,
         \21337 , \21338 , \21339 , \21340 , \21341 , \21342 , \21343 , \21344 , \21345 , \21346 ,
         \21347 , \21348 , \21349 , \21350 , \21351 , \21352 , \21353 , \21354 , \21355 , \21356 ,
         \21357 , \21358 , \21359 , \21360 , \21361 , \21362 , \21363 , \21364 , \21365 , \21366 ,
         \21367 , \21368 , \21369 , \21370 , \21371_nG399e , \21372 , \21373 , \21374 , \21375 , \21376 ,
         \21377 , \21378 , \21379 , \21380 , \21381 , \21382 , \21383 , \21384 , \21385 , \21386 ,
         \21387 , \21388 , \21389 , \21390 , \21391 , \21392 , \21393 , \21394 , \21395 , \21396 ,
         \21397 , \21398 , \21399 , \21400 , \21401 , \21402 , \21403 , \21404 , \21405 , \21406 ,
         \21407 , \21408 , \21409 , \21410 , \21411 , \21412 , \21413 , \21414 , \21415 , \21416 ,
         \21417 , \21418 , \21419 , \21420 , \21421 , \21422 , \21423 , \21424 , \21425 , \21426 ,
         \21427 , \21428 , \21429 , \21430 , \21431 , \21432 , \21433 , \21434 , \21435 , \21436 ,
         \21437 , \21438 , \21439 , \21440 , \21441 , \21442 , \21443 , \21444 , \21445 , \21446 ,
         \21447 , \21448 , \21449 , \21450 , \21451 , \21452 , \21453 , \21454 , \21455 , \21456 ,
         \21457 , \21458 , \21459 , \21460 , \21461 , \21462 , \21463 , \21464 , \21465 , \21466 ,
         \21467 , \21468 , \21469 , \21470 , \21471 , \21472 , \21473 , \21474 , \21475 , \21476 ,
         \21477 , \21478 , \21479 , \21480 , \21481 , \21482 , \21483 , \21484 , \21485 , \21486 ,
         \21487 , \21488 , \21489 , \21490 , \21491 , \21492 , \21493 , \21494 , \21495 , \21496 ,
         \21497 , \21498 , \21499 , \21500 , \21501 , \21502 , \21503 , \21504 , \21505_nG28f6 , \21506 ,
         \21507 , \21508 , \21509 , \21510 , \21511 , \21512 , \21513 , \21514 , \21515 , \21516 ,
         \21517 , \21518 , \21519 , \21520 , \21521 , \21522 , \21523 , \21524 , \21525 , \21526 ,
         \21527 , \21528 , \21529 , \21530 , \21531 , \21532 , \21533 , \21534 , \21535 , \21536 ,
         \21537 , \21538 , \21539 , \21540 , \21541 , \21542 , \21543 , \21544 , \21545 , \21546 ,
         \21547 , \21548 , \21549 , \21550 , \21551 , \21552 , \21553 , \21554 , \21555 , \21556 ,
         \21557 , \21558 , \21559 , \21560 , \21561 , \21562 , \21563 , \21564 , \21565 , \21566 ,
         \21567 , \21568 , \21569 , \21570 , \21571 , \21572 , \21573 , \21574 , \21575 , \21576 ,
         \21577 , \21578 , \21579 , \21580 , \21581 , \21582 , \21583 , \21584 , \21585 , \21586 ,
         \21587 , \21588 , \21589 , \21590 , \21591 , \21592 , \21593 , \21594 , \21595 , \21596 ,
         \21597 , \21598 , \21599 , \21600 , \21601 , \21602 , \21603 , \21604 , \21605 , \21606 ,
         \21607 , \21608 , \21609 , \21610 , \21611 , \21612 , \21613 , \21614 , \21615 , \21616 ,
         \21617 , \21618 , \21619 , \21620 , \21621 , \21622 , \21623 , \21624 , \21625 , \21626 ,
         \21627 , \21628 , \21629 , \21630 , \21631 , \21632 , \21633 , \21634 , \21635 , \21636 ,
         \21637 , \21638_nG3a23 , \21639 , \21640 , \21641 , \21642 , \21643 , \21644 , \21645 , \21646 ,
         \21647 , \21648 , \21649_nG441e , \21650 , \21651 , \21652_nG4421 , \21653 , \21654 , \21655 , \21656 ,
         \21657 , \21658 , \21659 , \21660 , \21661 , \21662 , \21663 , \21664 , \21665 , \21666 ,
         \21667 , \21668 , \21669 , \21670 , \21671 , \21672 , \21673 , \21674 , \21675 , \21676 ,
         \21677 , \21678 , \21679 , \21680 , \21681 , \21682 , \21683 , \21684 , \21685 , \21686 ,
         \21687 , \21688 , \21689 , \21690 , \21691 , \21692 , \21693 , \21694 , \21695 , \21696 ,
         \21697 , \21698 , \21699 , \21700 , \21701 , \21702 , \21703 , \21704 , \21705 , \21706 ,
         \21707 , \21708 , \21709 , \21710 , \21711 , \21712 , \21713 , \21714 , \21715 , \21716 ,
         \21717 , \21718 , \21719 , \21720 , \21721 , \21722 , \21723 , \21724 , \21725 , \21726 ,
         \21727 , \21728 , \21729 , \21730 , \21731 , \21732 , \21733 , \21734 , \21735 , \21736 ,
         \21737 , \21738 , \21739 , \21740 , \21741 , \21742 , \21743 , \21744 , \21745 , \21746 ,
         \21747 , \21748 , \21749 , \21750 , \21751 , \21752 , \21753 , \21754 , \21755 , \21756 ,
         \21757 , \21758 , \21759 , \21760 , \21761 , \21762 , \21763 , \21764 , \21765 , \21766 ,
         \21767 , \21768 , \21769 , \21770 , \21771 , \21772 , \21773 , \21774 , \21775 , \21776 ,
         \21777 , \21778 , \21779 , \21780 , \21781 , \21782 , \21783 , \21784 , \21785 , \21786 ,
         \21787 , \21788 , \21789 , \21790 , \21791 , \21792 , \21793 , \21794 , \21795 , \21796 ,
         \21797 , \21798 , \21799 , \21800 , \21801 , \21802 , \21803 , \21804 , \21805 , \21806 ,
         \21807 , \21808 , \21809 , \21810 , \21811 , \21812 , \21813 , \21814 , \21815 , \21816 ,
         \21817 , \21818 , \21819 , \21820 , \21821 , \21822 , \21823 , \21824 , \21825 , \21826 ,
         \21827 , \21828 , \21829 , \21830 , \21831 , \21832 , \21833 , \21834 , \21835 , \21836 ,
         \21837 , \21838 , \21839 , \21840 , \21841 , \21842 , \21843 , \21844 , \21845 , \21846 ,
         \21847 , \21848 , \21849 , \21850 , \21851 , \21852 , \21853 , \21854 , \21855 , \21856 ,
         \21857 , \21858 , \21859 , \21860 , \21861 , \21862 , \21863 , \21864 , \21865 , \21866 ,
         \21867 , \21868 , \21869 , \21870 , \21871 , \21872 , \21873 , \21874 , \21875 , \21876 ,
         \21877 , \21878 , \21879 , \21880 , \21881 , \21882 , \21883 , \21884 , \21885 , \21886 ,
         \21887 , \21888 , \21889 , \21890 , \21891 , \21892 , \21893 , \21894 , \21895 , \21896 ,
         \21897 , \21898 , \21899 , \21900 , \21901 , \21902 , \21903 , \21904 , \21905 , \21906 ,
         \21907 , \21908 , \21909 , \21910 , \21911 , \21912 , \21913 , \21914 , \21915 , \21916 ,
         \21917 , \21918 , \21919 , \21920 , \21921 , \21922 , \21923 , \21924 , \21925 , \21926 ,
         \21927 , \21928 , \21929 , \21930 , \21931 , \21932 , \21933 , \21934 , \21935 , \21936 ,
         \21937 , \21938 , \21939 , \21940 , \21941 , \21942 , \21943 , \21944 , \21945 , \21946 ,
         \21947 , \21948 , \21949 , \21950 , \21951 , \21952 , \21953 , \21954 , \21955 , \21956_nG65ad ,
         \21957 , \21958 , \21959 , \21960 , \21961 , \21962 , \21963 , \21964 , \21965 , \21966 ,
         \21967 , \21968 , \21969 , \21970 , \21971 , \21972 , \21973 , \21974 , \21975 , \21976 ,
         \21977 , \21978 , \21979 , \21980 , \21981 , \21982 , \21983 , \21984 , \21985 , \21986 ,
         \21987 , \21988 , \21989 , \21990 , \21991 , \21992 , \21993 , \21994 , \21995 , \21996 ,
         \21997 , \21998 , \21999 , \22000 , \22001 , \22002 , \22003 , \22004 , \22005 , \22006 ,
         \22007 , \22008 , \22009 , \22010 , \22011 , \22012 , \22013 , \22014 , \22015 , \22016 ,
         \22017 , \22018 , \22019 , \22020 , \22021 , \22022 , \22023 , \22024 , \22025 , \22026 ,
         \22027 , \22028 , \22029 , \22030 , \22031 , \22032 , \22033 , \22034 , \22035 , \22036 ,
         \22037 , \22038 , \22039 , \22040 , \22041 , \22042 , \22043 , \22044 , \22045 , \22046 ,
         \22047 , \22048 , \22049 , \22050 , \22051 , \22052 , \22053 , \22054 , \22055 , \22056 ,
         \22057 , \22058 , \22059 , \22060 , \22061 , \22062 , \22063 , \22064 , \22065 , \22066 ,
         \22067 , \22068 , \22069 , \22070 , \22071 , \22072 , \22073 , \22074 , \22075 , \22076 ,
         \22077 , \22078 , \22079 , \22080 , \22081 , \22082 , \22083 , \22084 , \22085 , \22086 ,
         \22087 , \22088_nG65ae , \22089_nG65af , \22090 , \22091 , \22092 , \22093 , \22094 , \22095 , \22096 ,
         \22097 , \22098 , \22099_nG577c , \22100_nG5800 , \22101_nG5801 , \22102 , \22103 , \22104 , \22105 , \22106 ,
         \22107 , \22108 , \22109 , \22110 , \22111 , \22112 , \22113 , \22114 , \22115 , \22116 ,
         \22117 , \22118 , \22119 , \22120 , \22121 , \22122 , \22123 , \22124 , \22125 , \22126 ,
         \22127 , \22128 , \22129_nG9bd8 , \22130 , \22131 , \22132 , \22133 , \22134 , \22135 , \22136 ,
         \22137 , \22138 , \22139 , \22140 , \22141 , \22142 , \22143 , \22144 , \22145 , \22146 ,
         \22147 , \22148 , \22149 , \22150 , \22151 , \22152 , \22153 , \22154 , \22155 , \22156 ,
         \22157 , \22158 , \22159 , \22160 , \22161 , \22162 , \22163 , \22164 , \22165 , \22166 ,
         \22167 , \22168 , \22169 , \22170 , \22171 , \22172 , \22173 , \22174 , \22175 , \22176 ,
         \22177 , \22178 , \22179 , \22180 , \22181 , \22182 , \22183 , \22184 , \22185 , \22186 ,
         \22187 , \22188 , \22189 , \22190 , \22191 , \22192 , \22193 , \22194 , \22195 , \22196 ,
         \22197 , \22198 , \22199 , \22200 , \22201 , \22202 , \22203 , \22204 , \22205 , \22206 ,
         \22207 , \22208 , \22209 , \22210 , \22211 , \22212 , \22213 , \22214 , \22215 , \22216 ,
         \22217 , \22218 , \22219 , \22220 , \22221 , \22222 , \22223 , \22224 , \22225 , \22226 ,
         \22227 , \22228 , \22229 , \22230 , \22231 , \22232 , \22233 , \22234 , \22235 , \22236 ,
         \22237 , \22238 , \22239 , \22240 , \22241 , \22242 , \22243 , \22244 , \22245 , \22246 ,
         \22247 , \22248 , \22249 , \22250 , \22251 , \22252 , \22253 , \22254 , \22255 , \22256 ,
         \22257 , \22258 , \22259 , \22260 , \22261 , \22262 , \22263 , \22264 , \22265 , \22266 ,
         \22267 , \22268 , \22269 , \22270 , \22271 , \22272 , \22273 , \22274 , \22275 , \22276 ,
         \22277 , \22278 , \22279 , \22280 , \22281 , \22282 , \22283 , \22284 , \22285 , \22286 ,
         \22287 , \22288 , \22289 , \22290 , \22291 , \22292 , \22293 , \22294 , \22295 , \22296 ,
         \22297 , \22298 , \22299 , \22300 , \22301 , \22302 , \22303 , \22304 , \22305 , \22306 ,
         \22307 , \22308 , \22309 , \22310 , \22311 , \22312 , \22313 , \22314 , \22315 , \22316 ,
         \22317 , \22318 , \22319 , \22320 , \22321 , \22322 , \22323 , \22324 , \22325 , \22326 ,
         \22327 , \22328 , \22329 , \22330 , \22331 , \22332 , \22333 , \22334 , \22335 , \22336 ,
         \22337 , \22338 , \22339 , \22340 , \22341 , \22342 , \22343 , \22344 , \22345 , \22346 ,
         \22347 , \22348 , \22349 , \22350 , \22351 , \22352 , \22353 , \22354 , \22355 , \22356 ,
         \22357 , \22358 , \22359 , \22360 , \22361 , \22362 , \22363 , \22364 , \22365 , \22366 ,
         \22367 , \22368 , \22369 , \22370 , \22371 , \22372 , \22373 , \22374 , \22375 , \22376 ,
         \22377 , \22378 , \22379 , \22380 , \22381 , \22382 , \22383 , \22384 , \22385 , \22386 ,
         \22387 , \22388 , \22389 , \22390 , \22391 , \22392 , \22393 , \22394 , \22395 , \22396 ,
         \22397 , \22398 , \22399 , \22400 , \22401 , \22402 , \22403 , \22404 , \22405_nG5885 , \22406 ,
         \22407 , \22408 , \22409 , \22410 , \22411 , \22412 , \22413 , \22414 , \22415 , \22416 ,
         \22417 , \22418 , \22419 , \22420 , \22421 , \22422 , \22423 , \22424 , \22425 , \22426 ,
         \22427 , \22428 , \22429 , \22430 , \22431 , \22432 , \22433 , \22434 , \22435 , \22436 ,
         \22437 , \22438 , \22439 , \22440 , \22441 , \22442 , \22443 , \22444 , \22445 , \22446 ,
         \22447 , \22448 , \22449 , \22450 , \22451 , \22452 , \22453 , \22454 , \22455 , \22456 ,
         \22457 , \22458 , \22459 , \22460 , \22461 , \22462 , \22463 , \22464 , \22465 , \22466 ,
         \22467 , \22468 , \22469 , \22470 , \22471 , \22472 , \22473 , \22474 , \22475 , \22476 ,
         \22477 , \22478 , \22479 , \22480 , \22481 , \22482 , \22483 , \22484 , \22485 , \22486 ,
         \22487 , \22488 , \22489 , \22490 , \22491 , \22492 , \22493 , \22494 , \22495 , \22496 ,
         \22497 , \22498 , \22499 , \22500 , \22501 , \22502 , \22503 , \22504 , \22505 , \22506 ,
         \22507 , \22508 , \22509 , \22510 , \22511 , \22512 , \22513 , \22514 , \22515 , \22516 ,
         \22517 , \22518 , \22519 , \22520 , \22521 , \22522 , \22523 , \22524 , \22525 , \22526 ,
         \22527 , \22528 , \22529 , \22530 , \22531 , \22532 , \22533 , \22534 , \22535 , \22536 ,
         \22537_nG5909 , \22538_nG590a , \22539 , \22540 , \22541 , \22542 , \22543 , \22544 , \22545 , \22546 ,
         \22547 , \22548 , \22549 , \22550 , \22551 , \22552 , \22553_nG65b0 , \22554_nG65b1 , \22555_nG65b2 , \22556 ,
         \22557 , \22558 , \22559 , \22560 , \22561 , \22562 , \22563 , \22564 , \22565 , \22566 ,
         \22567 , \22568 , \22569 , \22570 , \22571 , \22572 , \22573 , \22574 , \22575 , \22576 ,
         \22577 , \22578 , \22579 , \22580 , \22581 , \22582 , \22583 , \22584 , \22585 , \22586 ,
         \22587 , \22588 , \22589 , \22590 , \22591 , \22592 , \22593 , \22594 , \22595 , \22596 ,
         \22597 , \22598 , \22599 , \22600 , \22601 , \22602 , \22603 , \22604 , \22605 , \22606 ,
         \22607 , \22608 , \22609 , \22610 , \22611 , \22612 , \22613 , \22614 , \22615 , \22616 ,
         \22617 , \22618 , \22619 , \22620 , \22621 , \22622 , \22623 , \22624 , \22625 , \22626 ,
         \22627 , \22628 , \22629_nG9bd5 , \22630 , \22631 , \22632 , \22633 , \22634 , \22635 , \22636 ,
         \22637 , \22638 , \22639 , \22640 , \22641 , \22642 , \22643 , \22644 , \22645 , \22646 ,
         \22647 , \22648 , \22649 , \22650 , \22651 , \22652 , \22653 , \22654 , \22655 , \22656 ,
         \22657 , \22658 , \22659 , \22660 , \22661 , \22662 , \22663 , \22664 , \22665 , \22666 ,
         \22667 , \22668 , \22669 , \22670 , \22671 , \22672 , \22673 , \22674 , \22675 , \22676 ,
         \22677 , \22678 , \22679 , \22680 , \22681 , \22682 , \22683 , \22684 , \22685 , \22686 ,
         \22687 , \22688 , \22689 , \22690 , \22691 , \22692 , \22693 , \22694 , \22695 , \22696 ,
         \22697 , \22698 , \22699 , \22700 , \22701 , \22702 , \22703 , \22704 , \22705 , \22706 ,
         \22707 , \22708 , \22709 , \22710 , \22711 , \22712 , \22713 , \22714 , \22715 , \22716 ,
         \22717 , \22718 , \22719 , \22720 , \22721 , \22722 , \22723 , \22724 , \22725 , \22726 ,
         \22727 , \22728 , \22729 , \22730 , \22731 , \22732 , \22733 , \22734 , \22735 , \22736 ,
         \22737 , \22738 , \22739 , \22740 , \22741 , \22742 , \22743 , \22744 , \22745 , \22746 ,
         \22747 , \22748 , \22749 , \22750 , \22751 , \22752 , \22753 , \22754 , \22755 , \22756 ,
         \22757 , \22758 , \22759 , \22760 , \22761 , \22762 , \22763 , \22764 , \22765 , \22766 ,
         \22767 , \22768 , \22769 , \22770 , \22771 , \22772 , \22773 , \22774 , \22775 , \22776 ,
         \22777 , \22778 , \22779 , \22780 , \22781_nG2767 , \22782 , \22783 , \22784 , \22785 , \22786 ,
         \22787 , \22788 , \22789 , \22790 , \22791 , \22792 , \22793 , \22794 , \22795 , \22796 ,
         \22797 , \22798 , \22799 , \22800 , \22801 , \22802 , \22803 , \22804 , \22805 , \22806 ,
         \22807 , \22808 , \22809 , \22810 , \22811 , \22812 , \22813 , \22814 , \22815 , \22816 ,
         \22817 , \22818 , \22819 , \22820 , \22821 , \22822 , \22823 , \22824 , \22825 , \22826 ,
         \22827 , \22828 , \22829 , \22830 , \22831 , \22832 , \22833 , \22834 , \22835 , \22836 ,
         \22837 , \22838 , \22839 , \22840 , \22841 , \22842 , \22843 , \22844 , \22845 , \22846 ,
         \22847 , \22848 , \22849 , \22850 , \22851 , \22852 , \22853 , \22854 , \22855 , \22856 ,
         \22857 , \22858 , \22859 , \22860 , \22861 , \22862 , \22863 , \22864 , \22865 , \22866 ,
         \22867 , \22868 , \22869 , \22870 , \22871 , \22872 , \22873 , \22874 , \22875 , \22876 ,
         \22877 , \22878 , \22879 , \22880 , \22881 , \22882 , \22883 , \22884 , \22885 , \22886 ,
         \22887 , \22888 , \22889 , \22890 , \22891 , \22892 , \22893 , \22894 , \22895 , \22896 ,
         \22897 , \22898 , \22899 , \22900 , \22901 , \22902 , \22903 , \22904 , \22905 , \22906 ,
         \22907 , \22908 , \22909 , \22910 , \22911 , \22912 , \22913 , \22914_nG3894 , \22915 , \22916 ,
         \22917 , \22918 , \22919 , \22920 , \22921 , \22922 , \22923 , \22924 , \22925 , \22926 ,
         \22927 , \22928 , \22929 , \22930 , \22931 , \22932 , \22933 , \22934 , \22935 , \22936 ,
         \22937 , \22938 , \22939 , \22940 , \22941 , \22942 , \22943 , \22944 , \22945 , \22946 ,
         \22947 , \22948 , \22949 , \22950 , \22951 , \22952 , \22953 , \22954 , \22955 , \22956 ,
         \22957 , \22958 , \22959 , \22960 , \22961 , \22962 , \22963 , \22964 , \22965 , \22966 ,
         \22967 , \22968 , \22969 , \22970 , \22971 , \22972 , \22973 , \22974 , \22975 , \22976 ,
         \22977 , \22978 , \22979 , \22980 , \22981 , \22982 , \22983 , \22984 , \22985 , \22986 ,
         \22987 , \22988 , \22989 , \22990 , \22991 , \22992 , \22993 , \22994 , \22995 , \22996 ,
         \22997 , \22998 , \22999 , \23000 , \23001 , \23002 , \23003 , \23004 , \23005 , \23006 ,
         \23007 , \23008 , \23009 , \23010 , \23011 , \23012 , \23013 , \23014 , \23015 , \23016 ,
         \23017 , \23018 , \23019 , \23020 , \23021 , \23022 , \23023 , \23024 , \23025 , \23026 ,
         \23027 , \23028 , \23029 , \23030 , \23031 , \23032 , \23033 , \23034 , \23035 , \23036 ,
         \23037 , \23038 , \23039 , \23040 , \23041 , \23042 , \23043 , \23044 , \23045 , \23046 ,
         \23047 , \23048_nG27ec , \23049 , \23050 , \23051 , \23052 , \23053 , \23054 , \23055 , \23056 ,
         \23057 , \23058 , \23059 , \23060 , \23061 , \23062 , \23063 , \23064 , \23065 , \23066 ,
         \23067 , \23068 , \23069 , \23070 , \23071 , \23072 , \23073 , \23074 , \23075 , \23076 ,
         \23077 , \23078 , \23079 , \23080 , \23081 , \23082 , \23083 , \23084 , \23085 , \23086 ,
         \23087 , \23088 , \23089 , \23090 , \23091 , \23092 , \23093 , \23094 , \23095 , \23096 ,
         \23097 , \23098 , \23099 , \23100 , \23101 , \23102 , \23103 , \23104 , \23105 , \23106 ,
         \23107 , \23108 , \23109 , \23110 , \23111 , \23112 , \23113 , \23114 , \23115 , \23116 ,
         \23117 , \23118 , \23119 , \23120 , \23121 , \23122 , \23123 , \23124 , \23125 , \23126 ,
         \23127 , \23128 , \23129 , \23130 , \23131 , \23132 , \23133 , \23134 , \23135 , \23136 ,
         \23137 , \23138 , \23139 , \23140 , \23141 , \23142 , \23143 , \23144 , \23145 , \23146 ,
         \23147 , \23148 , \23149 , \23150 , \23151 , \23152 , \23153 , \23154 , \23155 , \23156 ,
         \23157 , \23158 , \23159 , \23160 , \23161 , \23162 , \23163 , \23164 , \23165 , \23166 ,
         \23167 , \23168 , \23169 , \23170 , \23171 , \23172 , \23173 , \23174 , \23175 , \23176 ,
         \23177 , \23178 , \23179 , \23180 , \23181_nG3919 , \23182 , \23183 , \23184 , \23185 , \23186 ,
         \23187 , \23188 , \23189 , \23190 , \23191 , \23192_nG4418 , \23193 , \23194 , \23195_nG441b , \23196 ,
         \23197 , \23198 , \23199 , \23200 , \23201 , \23202 , \23203 , \23204 , \23205 , \23206 ,
         \23207 , \23208 , \23209 , \23210 , \23211 , \23212 , \23213 , \23214 , \23215 , \23216 ,
         \23217 , \23218 , \23219 , \23220 , \23221 , \23222 , \23223 , \23224 , \23225 , \23226 ,
         \23227 , \23228 , \23229 , \23230 , \23231 , \23232 , \23233 , \23234 , \23235 , \23236 ,
         \23237 , \23238 , \23239 , \23240 , \23241 , \23242 , \23243 , \23244 , \23245 , \23246 ,
         \23247 , \23248 , \23249 , \23250 , \23251 , \23252 , \23253 , \23254 , \23255 , \23256 ,
         \23257 , \23258 , \23259 , \23260 , \23261 , \23262 , \23263 , \23264 , \23265 , \23266 ,
         \23267 , \23268 , \23269 , \23270 , \23271 , \23272 , \23273 , \23274 , \23275 , \23276 ,
         \23277 , \23278 , \23279 , \23280 , \23281 , \23282 , \23283 , \23284 , \23285 , \23286 ,
         \23287 , \23288 , \23289 , \23290 , \23291 , \23292 , \23293 , \23294 , \23295 , \23296 ,
         \23297 , \23298 , \23299 , \23300 , \23301 , \23302 , \23303 , \23304 , \23305 , \23306 ,
         \23307 , \23308 , \23309 , \23310 , \23311 , \23312 , \23313 , \23314 , \23315 , \23316 ,
         \23317 , \23318 , \23319 , \23320 , \23321 , \23322 , \23323 , \23324 , \23325 , \23326 ,
         \23327 , \23328 , \23329 , \23330 , \23331 , \23332 , \23333 , \23334 , \23335 , \23336 ,
         \23337 , \23338 , \23339 , \23340 , \23341 , \23342 , \23343 , \23344 , \23345 , \23346 ,
         \23347 , \23348 , \23349 , \23350 , \23351 , \23352 , \23353 , \23354 , \23355 , \23356 ,
         \23357 , \23358 , \23359 , \23360 , \23361 , \23362 , \23363 , \23364 , \23365 , \23366 ,
         \23367 , \23368 , \23369 , \23370 , \23371 , \23372 , \23373 , \23374 , \23375 , \23376 ,
         \23377 , \23378 , \23379 , \23380 , \23381 , \23382 , \23383 , \23384 , \23385 , \23386 ,
         \23387 , \23388 , \23389 , \23390 , \23391 , \23392 , \23393 , \23394 , \23395 , \23396 ,
         \23397 , \23398 , \23399 , \23400 , \23401 , \23402 , \23403 , \23404 , \23405 , \23406 ,
         \23407 , \23408 , \23409 , \23410 , \23411 , \23412 , \23413 , \23414 , \23415 , \23416 ,
         \23417 , \23418 , \23419 , \23420 , \23421 , \23422 , \23423 , \23424 , \23425 , \23426 ,
         \23427 , \23428 , \23429 , \23430 , \23431 , \23432 , \23433 , \23434 , \23435 , \23436 ,
         \23437 , \23438 , \23439 , \23440 , \23441 , \23442 , \23443 , \23444 , \23445 , \23446 ,
         \23447 , \23448 , \23449 , \23450 , \23451 , \23452 , \23453 , \23454 , \23455 , \23456 ,
         \23457 , \23458 , \23459 , \23460 , \23461 , \23462 , \23463 , \23464 , \23465 , \23466 ,
         \23467 , \23468 , \23469 , \23470 , \23471 , \23472 , \23473 , \23474 , \23475 , \23476 ,
         \23477 , \23478 , \23479 , \23480 , \23481 , \23482 , \23483_nG65b3 , \23484 , \23485 , \23486 ,
         \23487 , \23488 , \23489 , \23490 , \23491 , \23492 , \23493 , \23494 , \23495 , \23496 ,
         \23497 , \23498 , \23499 , \23500 , \23501 , \23502 , \23503 , \23504 , \23505 , \23506 ,
         \23507 , \23508 , \23509 , \23510 , \23511 , \23512 , \23513 , \23514 , \23515 , \23516 ,
         \23517 , \23518 , \23519 , \23520 , \23521 , \23522 , \23523 , \23524 , \23525 , \23526 ,
         \23527 , \23528 , \23529 , \23530 , \23531 , \23532 , \23533 , \23534 , \23535 , \23536 ,
         \23537 , \23538 , \23539 , \23540 , \23541 , \23542 , \23543 , \23544 , \23545 , \23546 ,
         \23547 , \23548 , \23549 , \23550 , \23551 , \23552 , \23553 , \23554 , \23555 , \23556 ,
         \23557 , \23558 , \23559 , \23560 , \23561 , \23562 , \23563 , \23564 , \23565 , \23566 ,
         \23567 , \23568 , \23569 , \23570 , \23571 , \23572 , \23573 , \23574 , \23575 , \23576 ,
         \23577 , \23578 , \23579 , \23580 , \23581 , \23582 , \23583 , \23584 , \23585 , \23586 ,
         \23587 , \23588 , \23589 , \23590 , \23591 , \23592 , \23593 , \23594 , \23595 , \23596 ,
         \23597 , \23598 , \23599 , \23600 , \23601 , \23602 , \23603 , \23604 , \23605 , \23606 ,
         \23607 , \23608 , \23609 , \23610 , \23611 , \23612 , \23613 , \23614 , \23615_nG65b4 , \23616_nG65b5 ,
         \23617 , \23618 , \23619 , \23620 , \23621 , \23622 , \23623 , \23624 , \23625 , \23626_nG598e ,
         \23627_nG5a12 , \23628_nG5a13 , \23629 , \23630 , \23631 , \23632 , \23633 , \23634 , \23635 , \23636 ,
         \23637 , \23638 , \23639 , \23640 , \23641 , \23642 , \23643 , \23644 , \23645 , \23646 ,
         \23647 , \23648 , \23649 , \23650 , \23651 , \23652 , \23653 , \23654 , \23655 , \23656 ,
         \23657 , \23658 , \23659 , \23660 , \23661 , \23662 , \23663 , \23664 , \23665 , \23666 ,
         \23667 , \23668 , \23669 , \23670 , \23671 , \23672 , \23673 , \23674 , \23675 , \23676 ,
         \23677 , \23678 , \23679 , \23680 , \23681 , \23682 , \23683 , \23684 , \23685 , \23686 ,
         \23687 , \23688 , \23689 , \23690 , \23691 , \23692 , \23693 , \23694 , \23695 , \23696_nG9bd2 ,
         \23697 , \23698 , \23699 , \23700 , \23701 , \23702 , \23703 , \23704 , \23705 , \23706 ,
         \23707 , \23708 , \23709 , \23710 , \23711 , \23712 , \23713 , \23714 , \23715 , \23716 ,
         \23717 , \23718 , \23719 , \23720 , \23721 , \23722 , \23723 , \23724 , \23725 , \23726 ,
         \23727 , \23728 , \23729 , \23730 , \23731 , \23732 , \23733 , \23734 , \23735 , \23736 ,
         \23737 , \23738 , \23739 , \23740 , \23741 , \23742 , \23743 , \23744 , \23745 , \23746 ,
         \23747 , \23748 , \23749 , \23750 , \23751 , \23752 , \23753 , \23754 , \23755 , \23756 ,
         \23757 , \23758 , \23759 , \23760 , \23761 , \23762 , \23763 , \23764 , \23765 , \23766 ,
         \23767 , \23768 , \23769 , \23770 , \23771 , \23772 , \23773 , \23774 , \23775 , \23776 ,
         \23777 , \23778 , \23779 , \23780 , \23781 , \23782 , \23783 , \23784 , \23785 , \23786 ,
         \23787 , \23788 , \23789 , \23790 , \23791 , \23792 , \23793 , \23794 , \23795 , \23796 ,
         \23797 , \23798 , \23799 , \23800 , \23801 , \23802 , \23803 , \23804 , \23805 , \23806 ,
         \23807 , \23808 , \23809 , \23810 , \23811 , \23812 , \23813 , \23814 , \23815 , \23816 ,
         \23817 , \23818 , \23819 , \23820 , \23821 , \23822 , \23823 , \23824 , \23825 , \23826 ,
         \23827 , \23828 , \23829 , \23830 , \23831 , \23832 , \23833 , \23834 , \23835 , \23836 ,
         \23837 , \23838 , \23839 , \23840 , \23841 , \23842 , \23843 , \23844 , \23845 , \23846 ,
         \23847 , \23848 , \23849 , \23850 , \23851 , \23852 , \23853 , \23854 , \23855 , \23856 ,
         \23857 , \23858 , \23859 , \23860 , \23861 , \23862 , \23863 , \23864 , \23865 , \23866 ,
         \23867 , \23868 , \23869 , \23870 , \23871 , \23872 , \23873 , \23874 , \23875 , \23876 ,
         \23877 , \23878 , \23879 , \23880 , \23881 , \23882 , \23883 , \23884 , \23885 , \23886 ,
         \23887 , \23888 , \23889 , \23890 , \23891 , \23892 , \23893 , \23894 , \23895 , \23896 ,
         \23897 , \23898 , \23899 , \23900 , \23901 , \23902 , \23903 , \23904 , \23905 , \23906 ,
         \23907 , \23908 , \23909 , \23910 , \23911 , \23912 , \23913 , \23914 , \23915 , \23916 ,
         \23917 , \23918 , \23919 , \23920 , \23921 , \23922 , \23923 , \23924 , \23925 , \23926 ,
         \23927 , \23928 , \23929 , \23930 , \23931 , \23932 , \23933 , \23934 , \23935 , \23936 ,
         \23937 , \23938 , \23939 , \23940 , \23941 , \23942 , \23943 , \23944 , \23945 , \23946 ,
         \23947 , \23948 , \23949 , \23950 , \23951 , \23952 , \23953 , \23954 , \23955 , \23956 ,
         \23957 , \23958 , \23959 , \23960 , \23961 , \23962 , \23963 , \23964 , \23965 , \23966 ,
         \23967 , \23968 , \23969 , \23970 , \23971 , \23972 , \23973 , \23974 , \23975 , \23976 ,
         \23977 , \23978 , \23979 , \23980 , \23981 , \23982 , \23983 , \23984 , \23985 , \23986 ,
         \23987 , \23988 , \23989 , \23990 , \23991 , \23992 , \23993 , \23994 , \23995 , \23996 ,
         \23997 , \23998 , \23999 , \24000 , \24001_nG5a97 , \24002 , \24003 , \24004 , \24005 , \24006 ,
         \24007 , \24008 , \24009 , \24010 , \24011 , \24012 , \24013 , \24014 , \24015 , \24016 ,
         \24017 , \24018 , \24019 , \24020 , \24021 , \24022 , \24023 , \24024 , \24025 , \24026 ,
         \24027 , \24028 , \24029 , \24030 , \24031 , \24032 , \24033 , \24034 , \24035 , \24036 ,
         \24037 , \24038 , \24039 , \24040 , \24041 , \24042 , \24043 , \24044 , \24045 , \24046 ,
         \24047 , \24048 , \24049 , \24050 , \24051 , \24052 , \24053 , \24054 , \24055 , \24056 ,
         \24057 , \24058 , \24059 , \24060 , \24061 , \24062 , \24063 , \24064 , \24065 , \24066 ,
         \24067 , \24068 , \24069 , \24070 , \24071 , \24072 , \24073 , \24074 , \24075 , \24076 ,
         \24077 , \24078 , \24079 , \24080 , \24081 , \24082 , \24083 , \24084 , \24085 , \24086 ,
         \24087 , \24088 , \24089 , \24090 , \24091 , \24092 , \24093 , \24094 , \24095 , \24096 ,
         \24097 , \24098 , \24099 , \24100 , \24101 , \24102 , \24103 , \24104 , \24105 , \24106 ,
         \24107 , \24108 , \24109 , \24110 , \24111 , \24112 , \24113 , \24114 , \24115 , \24116 ,
         \24117 , \24118 , \24119 , \24120 , \24121 , \24122 , \24123 , \24124 , \24125 , \24126 ,
         \24127 , \24128 , \24129 , \24130 , \24131 , \24132 , \24133_nG5b1b , \24134_nG5b1c , \24135 , \24136 ,
         \24137 , \24138 , \24139 , \24140 , \24141 , \24142 , \24143 , \24144 , \24145 , \24146 ,
         \24147 , \24148 , \24149 , \24150 , \24151 , \24152 , \24153 , \24154 , \24155 , \24156 ,
         \24157 , \24158 , \24159 , \24160 , \24161 , \24162 , \24163 , \24164 , \24165 , \24166 ,
         \24167 , \24168 , \24169 , \24170 , \24171 , \24172 , \24173 , \24174 , \24175 , \24176 ,
         \24177 , \24178 , \24179 , \24180 , \24181 , \24182 , \24183 , \24184 , \24185 , \24186 ,
         \24187 , \24188 , \24189 , \24190 , \24191 , \24192 , \24193 , \24194 , \24195 , \24196_nG65b6 ,
         \24197_nG65b7 , \24198_nG65b8 , \24199 , \24200 , \24201 , \24202 , \24203 , \24204 , \24205 , \24206 ,
         \24207 , \24208 , \24209 , \24210 , \24211 , \24212 , \24213 , \24214 , \24215 , \24216 ,
         \24217 , \24218 , \24219 , \24220 , \24221 , \24222 , \24223 , \24224 , \24225 , \24226_nG9bcf ,
         \24227 , \24228 , \24229 , \24230 , \24231 , \24232 , \24233 , \24234 , \24235 , \24236 ,
         \24237 , \24238 , \24239 , \24240 , \24241 , \24242 , \24243 , \24244 , \24245 , \24246 ,
         \24247 , \24248 , \24249 , \24250 , \24251 , \24252 , \24253 , \24254 , \24255 , \24256 ,
         \24257 , \24258 , \24259 , \24260 , \24261 , \24262 , \24263 , \24264 , \24265 , \24266 ,
         \24267 , \24268 , \24269 , \24270 , \24271 , \24272 , \24273 , \24274 , \24275 , \24276 ,
         \24277 , \24278 , \24279 , \24280 , \24281 , \24282 , \24283 , \24284 , \24285 , \24286 ,
         \24287 , \24288 , \24289 , \24290 , \24291 , \24292 , \24293 , \24294 , \24295 , \24296 ,
         \24297 , \24298 , \24299 , \24300 , \24301 , \24302 , \24303 , \24304 , \24305 , \24306 ,
         \24307 , \24308 , \24309 , \24310 , \24311 , \24312 , \24313 , \24314 , \24315 , \24316 ,
         \24317 , \24318 , \24319 , \24320 , \24321 , \24322 , \24323 , \24324 , \24325 , \24326 ,
         \24327 , \24328 , \24329 , \24330 , \24331 , \24332 , \24333 , \24334 , \24335 , \24336 ,
         \24337 , \24338 , \24339 , \24340 , \24341 , \24342 , \24343 , \24344 , \24345 , \24346 ,
         \24347 , \24348 , \24349 , \24350 , \24351 , \24352 , \24353 , \24354 , \24355 , \24356 ,
         \24357 , \24358 , \24359 , \24360 , \24361 , \24362 , \24363 , \24364 , \24365 , \24366 ,
         \24367 , \24368 , \24369 , \24370 , \24371 , \24372_nG265d , \24373 , \24374 , \24375 , \24376 ,
         \24377 , \24378 , \24379 , \24380 , \24381 , \24382 , \24383 , \24384 , \24385 , \24386 ,
         \24387 , \24388 , \24389 , \24390 , \24391 , \24392 , \24393 , \24394 , \24395 , \24396 ,
         \24397 , \24398 , \24399 , \24400 , \24401 , \24402 , \24403 , \24404 , \24405 , \24406 ,
         \24407 , \24408 , \24409 , \24410 , \24411 , \24412 , \24413 , \24414 , \24415 , \24416 ,
         \24417 , \24418 , \24419 , \24420 , \24421 , \24422 , \24423 , \24424 , \24425 , \24426 ,
         \24427 , \24428 , \24429 , \24430 , \24431 , \24432 , \24433 , \24434 , \24435 , \24436 ,
         \24437 , \24438 , \24439 , \24440 , \24441 , \24442 , \24443 , \24444 , \24445 , \24446 ,
         \24447 , \24448 , \24449 , \24450 , \24451 , \24452 , \24453 , \24454 , \24455 , \24456 ,
         \24457 , \24458 , \24459 , \24460 , \24461 , \24462 , \24463 , \24464 , \24465 , \24466 ,
         \24467 , \24468 , \24469 , \24470 , \24471 , \24472 , \24473 , \24474 , \24475 , \24476 ,
         \24477 , \24478 , \24479 , \24480 , \24481 , \24482 , \24483 , \24484 , \24485 , \24486 ,
         \24487 , \24488 , \24489 , \24490 , \24491 , \24492 , \24493 , \24494 , \24495 , \24496 ,
         \24497 , \24498 , \24499 , \24500 , \24501 , \24502 , \24503 , \24504 , \24505_nG378a , \24506 ,
         \24507 , \24508 , \24509 , \24510 , \24511 , \24512 , \24513 , \24514 , \24515 , \24516 ,
         \24517 , \24518 , \24519 , \24520 , \24521 , \24522 , \24523 , \24524 , \24525 , \24526 ,
         \24527 , \24528 , \24529 , \24530 , \24531 , \24532 , \24533 , \24534 , \24535 , \24536 ,
         \24537 , \24538 , \24539 , \24540 , \24541 , \24542 , \24543 , \24544 , \24545 , \24546 ,
         \24547 , \24548 , \24549 , \24550 , \24551 , \24552 , \24553 , \24554 , \24555 , \24556 ,
         \24557 , \24558 , \24559 , \24560 , \24561 , \24562 , \24563 , \24564 , \24565 , \24566 ,
         \24567 , \24568 , \24569 , \24570 , \24571 , \24572 , \24573 , \24574 , \24575 , \24576 ,
         \24577 , \24578 , \24579 , \24580 , \24581 , \24582 , \24583 , \24584 , \24585 , \24586 ,
         \24587 , \24588 , \24589 , \24590 , \24591 , \24592 , \24593 , \24594 , \24595 , \24596 ,
         \24597 , \24598 , \24599 , \24600 , \24601 , \24602 , \24603 , \24604 , \24605 , \24606 ,
         \24607 , \24608 , \24609 , \24610 , \24611 , \24612 , \24613 , \24614 , \24615 , \24616 ,
         \24617 , \24618 , \24619 , \24620 , \24621 , \24622 , \24623 , \24624 , \24625 , \24626 ,
         \24627 , \24628 , \24629 , \24630 , \24631 , \24632 , \24633 , \24634 , \24635 , \24636 ,
         \24637 , \24638 , \24639_nG26e2 , \24640 , \24641 , \24642 , \24643 , \24644 , \24645 , \24646 ,
         \24647 , \24648 , \24649 , \24650 , \24651 , \24652 , \24653 , \24654 , \24655 , \24656 ,
         \24657 , \24658 , \24659 , \24660 , \24661 , \24662 , \24663 , \24664 , \24665 , \24666 ,
         \24667 , \24668 , \24669 , \24670 , \24671 , \24672 , \24673 , \24674 , \24675 , \24676 ,
         \24677 , \24678 , \24679 , \24680 , \24681 , \24682 , \24683 , \24684 , \24685 , \24686 ,
         \24687 , \24688 , \24689 , \24690 , \24691 , \24692 , \24693 , \24694 , \24695 , \24696 ,
         \24697 , \24698 , \24699 , \24700 , \24701 , \24702 , \24703 , \24704 , \24705 , \24706 ,
         \24707 , \24708 , \24709 , \24710 , \24711 , \24712 , \24713 , \24714 , \24715 , \24716 ,
         \24717 , \24718 , \24719 , \24720 , \24721 , \24722 , \24723 , \24724 , \24725 , \24726 ,
         \24727 , \24728 , \24729 , \24730 , \24731 , \24732 , \24733 , \24734 , \24735 , \24736 ,
         \24737 , \24738 , \24739 , \24740 , \24741 , \24742 , \24743 , \24744 , \24745 , \24746 ,
         \24747 , \24748 , \24749 , \24750 , \24751 , \24752 , \24753 , \24754 , \24755 , \24756 ,
         \24757 , \24758 , \24759 , \24760 , \24761 , \24762 , \24763 , \24764 , \24765 , \24766 ,
         \24767 , \24768 , \24769 , \24770 , \24771 , \24772_nG380f , \24773 , \24774 , \24775 , \24776 ,
         \24777 , \24778 , \24779 , \24780 , \24781 , \24782 , \24783_nG4412 , \24784 , \24785 , \24786_nG4415 ,
         \24787 , \24788 , \24789 , \24790 , \24791 , \24792 , \24793 , \24794 , \24795 , \24796 ,
         \24797 , \24798 , \24799 , \24800 , \24801 , \24802 , \24803 , \24804 , \24805 , \24806 ,
         \24807 , \24808 , \24809 , \24810 , \24811 , \24812 , \24813 , \24814 , \24815 , \24816 ,
         \24817 , \24818 , \24819 , \24820 , \24821 , \24822 , \24823 , \24824 , \24825 , \24826 ,
         \24827 , \24828 , \24829 , \24830 , \24831 , \24832 , \24833 , \24834 , \24835 , \24836 ,
         \24837 , \24838 , \24839 , \24840 , \24841 , \24842 , \24843 , \24844 , \24845 , \24846 ,
         \24847 , \24848 , \24849 , \24850 , \24851 , \24852 , \24853 , \24854 , \24855 , \24856 ,
         \24857 , \24858 , \24859 , \24860 , \24861 , \24862 , \24863 , \24864 , \24865 , \24866 ,
         \24867 , \24868 , \24869 , \24870 , \24871 , \24872 , \24873 , \24874 , \24875 , \24876 ,
         \24877 , \24878 , \24879 , \24880 , \24881 , \24882 , \24883 , \24884 , \24885 , \24886 ,
         \24887 , \24888 , \24889 , \24890 , \24891 , \24892 , \24893 , \24894 , \24895 , \24896 ,
         \24897 , \24898 , \24899 , \24900 , \24901 , \24902 , \24903 , \24904 , \24905 , \24906 ,
         \24907 , \24908 , \24909 , \24910 , \24911 , \24912 , \24913 , \24914 , \24915 , \24916 ,
         \24917 , \24918 , \24919 , \24920 , \24921 , \24922 , \24923 , \24924 , \24925 , \24926 ,
         \24927 , \24928 , \24929 , \24930 , \24931 , \24932 , \24933 , \24934 , \24935 , \24936 ,
         \24937 , \24938 , \24939 , \24940 , \24941 , \24942 , \24943 , \24944 , \24945 , \24946 ,
         \24947 , \24948 , \24949 , \24950 , \24951 , \24952 , \24953 , \24954 , \24955 , \24956 ,
         \24957 , \24958 , \24959 , \24960 , \24961 , \24962 , \24963 , \24964 , \24965 , \24966 ,
         \24967 , \24968 , \24969 , \24970 , \24971 , \24972 , \24973 , \24974 , \24975 , \24976 ,
         \24977 , \24978 , \24979 , \24980 , \24981 , \24982 , \24983 , \24984 , \24985 , \24986 ,
         \24987 , \24988 , \24989 , \24990 , \24991 , \24992 , \24993 , \24994 , \24995 , \24996 ,
         \24997 , \24998 , \24999 , \25000 , \25001 , \25002 , \25003 , \25004 , \25005 , \25006 ,
         \25007 , \25008 , \25009 , \25010 , \25011 , \25012 , \25013 , \25014 , \25015 , \25016 ,
         \25017 , \25018 , \25019 , \25020 , \25021 , \25022 , \25023 , \25024 , \25025 , \25026 ,
         \25027 , \25028 , \25029 , \25030 , \25031 , \25032 , \25033 , \25034 , \25035 , \25036 ,
         \25037 , \25038 , \25039 , \25040 , \25041 , \25042 , \25043 , \25044 , \25045 , \25046 ,
         \25047 , \25048 , \25049 , \25050 , \25051 , \25052 , \25053 , \25054 , \25055 , \25056 ,
         \25057 , \25058 , \25059 , \25060 , \25061 , \25062 , \25063 , \25064 , \25065 , \25066 ,
         \25067 , \25068 , \25069 , \25070 , \25071 , \25072 , \25073 , \25074 , \25075 , \25076 ,
         \25077 , \25078 , \25079 , \25080 , \25081 , \25082 , \25083 , \25084 , \25085 , \25086 ,
         \25087 , \25088 , \25089 , \25090 , \25091 , \25092 , \25093 , \25094 , \25095 , \25096 ,
         \25097 , \25098 , \25099 , \25100 , \25101 , \25102 , \25103 , \25104 , \25105 , \25106 ,
         \25107 , \25108 , \25109 , \25110 , \25111 , \25112 , \25113 , \25114 , \25115 , \25116 ,
         \25117 , \25118 , \25119 , \25120 , \25121 , \25122 , \25123 , \25124 , \25125 , \25126 ,
         \25127 , \25128 , \25129_nG5ba0 , \25130 , \25131 , \25132 , \25133 , \25134 , \25135 , \25136 ,
         \25137 , \25138 , \25139 , \25140 , \25141 , \25142 , \25143 , \25144 , \25145 , \25146 ,
         \25147 , \25148 , \25149 , \25150 , \25151 , \25152 , \25153 , \25154 , \25155 , \25156 ,
         \25157 , \25158 , \25159 , \25160 , \25161 , \25162 , \25163 , \25164 , \25165 , \25166 ,
         \25167 , \25168 , \25169 , \25170 , \25171 , \25172 , \25173 , \25174 , \25175 , \25176 ,
         \25177 , \25178 , \25179 , \25180 , \25181 , \25182 , \25183 , \25184 , \25185 , \25186 ,
         \25187 , \25188 , \25189 , \25190 , \25191 , \25192 , \25193 , \25194 , \25195 , \25196 ,
         \25197 , \25198 , \25199 , \25200 , \25201 , \25202 , \25203 , \25204 , \25205 , \25206 ,
         \25207 , \25208 , \25209 , \25210 , \25211 , \25212 , \25213 , \25214 , \25215 , \25216 ,
         \25217 , \25218 , \25219 , \25220 , \25221 , \25222 , \25223 , \25224 , \25225 , \25226 ,
         \25227 , \25228 , \25229 , \25230 , \25231 , \25232 , \25233 , \25234 , \25235 , \25236 ,
         \25237 , \25238 , \25239 , \25240 , \25241 , \25242 , \25243 , \25244 , \25245 , \25246 ,
         \25247 , \25248 , \25249 , \25250 , \25251 , \25252 , \25253 , \25254 , \25255 , \25256 ,
         \25257 , \25258 , \25259 , \25260 , \25261_nG5c24 , \25262_nG5c25 , \25263 , \25264 , \25265 , \25266 ,
         \25267 , \25268 , \25269_nG65b9 , \25270_nG65ba , \25271_nG65bb , \25272 , \25273 , \25274 , \25275 , \25276 ,
         \25277 , \25278 , \25279 , \25280 , \25281 , \25282 , \25283 , \25284 , \25285 , \25286 ,
         \25287 , \25288 , \25289 , \25290 , \25291 , \25292 , \25293 , \25294 , \25295 , \25296 ,
         \25297 , \25298_nG9bcc , \25299 , \25300 , \25301 , \25302 , \25303 , \25304 , \25305 , \25306 ,
         \25307 , \25308 , \25309 , \25310 , \25311 , \25312 , \25313 , \25314 , \25315 , \25316 ,
         \25317 , \25318 , \25319 , \25320 , \25321 , \25322 , \25323 , \25324 , \25325 , \25326 ,
         \25327 , \25328 , \25329 , \25330 , \25331 , \25332 , \25333 , \25334 , \25335 , \25336 ,
         \25337 , \25338 , \25339 , \25340 , \25341 , \25342 , \25343 , \25344 , \25345 , \25346 ,
         \25347 , \25348 , \25349 , \25350 , \25351 , \25352 , \25353 , \25354 , \25355 , \25356 ,
         \25357 , \25358 , \25359 , \25360 , \25361 , \25362 , \25363 , \25364 , \25365 , \25366 ,
         \25367 , \25368 , \25369 , \25370 , \25371 , \25372 , \25373 , \25374 , \25375 , \25376 ,
         \25377 , \25378 , \25379 , \25380 , \25381 , \25382 , \25383 , \25384 , \25385 , \25386 ,
         \25387 , \25388 , \25389 , \25390 , \25391 , \25392 , \25393 , \25394 , \25395 , \25396 ,
         \25397 , \25398 , \25399 , \25400 , \25401 , \25402 , \25403 , \25404 , \25405 , \25406 ,
         \25407 , \25408 , \25409 , \25410 , \25411 , \25412 , \25413 , \25414 , \25415 , \25416 ,
         \25417 , \25418 , \25419 , \25420 , \25421 , \25422 , \25423 , \25424 , \25425 , \25426 ,
         \25427 , \25428 , \25429 , \25430 , \25431 , \25432 , \25433 , \25434 , \25435 , \25436 ,
         \25437 , \25438 , \25439 , \25440 , \25441 , \25442 , \25443 , \25444 , \25445 , \25446 ,
         \25447 , \25448 , \25449 , \25450 , \25451 , \25452 , \25453 , \25454 , \25455 , \25456 ,
         \25457 , \25458 , \25459 , \25460 , \25461 , \25462 , \25463 , \25464 , \25465 , \25466 ,
         \25467 , \25468 , \25469 , \25470 , \25471 , \25472 , \25473 , \25474 , \25475 , \25476 ,
         \25477 , \25478 , \25479 , \25480 , \25481 , \25482 , \25483 , \25484 , \25485 , \25486 ,
         \25487 , \25488 , \25489 , \25490 , \25491 , \25492 , \25493 , \25494 , \25495 , \25496 ,
         \25497 , \25498 , \25499 , \25500 , \25501 , \25502 , \25503 , \25504 , \25505 , \25506 ,
         \25507 , \25508 , \25509 , \25510 , \25511 , \25512 , \25513 , \25514 , \25515 , \25516 ,
         \25517 , \25518 , \25519 , \25520 , \25521 , \25522 , \25523 , \25524 , \25525 , \25526 ,
         \25527 , \25528 , \25529 , \25530 , \25531 , \25532 , \25533 , \25534 , \25535 , \25536 ,
         \25537 , \25538 , \25539 , \25540 , \25541 , \25542 , \25543 , \25544 , \25545 , \25546 ,
         \25547 , \25548 , \25549 , \25550 , \25551 , \25552 , \25553 , \25554 , \25555 , \25556 ,
         \25557 , \25558 , \25559 , \25560 , \25561 , \25562 , \25563 , \25564 , \25565 , \25566 ,
         \25567 , \25568 , \25569 , \25570 , \25571 , \25572 , \25573 , \25574 , \25575 , \25576 ,
         \25577 , \25578 , \25579 , \25580 , \25581 , \25582 , \25583 , \25584 , \25585 , \25586 ,
         \25587 , \25588 , \25589 , \25590 , \25591 , \25592 , \25593 , \25594 , \25595 , \25596 ,
         \25597 , \25598 , \25599 , \25600 , \25601 , \25602 , \25603 , \25604 , \25605 , \25606 ,
         \25607 , \25608 , \25609 , \25610 , \25611 , \25612 , \25613 , \25614 , \25615 , \25616 ,
         \25617 , \25618 , \25619 , \25620 , \25621 , \25622 , \25623 , \25624 , \25625 , \25626 ,
         \25627 , \25628 , \25629 , \25630 , \25631 , \25632 , \25633 , \25634 , \25635 , \25636_nG5ca9 ,
         \25637 , \25638 , \25639 , \25640 , \25641 , \25642 , \25643 , \25644 , \25645 , \25646 ,
         \25647 , \25648 , \25649 , \25650 , \25651 , \25652 , \25653 , \25654 , \25655 , \25656 ,
         \25657 , \25658 , \25659 , \25660 , \25661 , \25662 , \25663 , \25664 , \25665 , \25666 ,
         \25667 , \25668 , \25669 , \25670 , \25671 , \25672 , \25673 , \25674 , \25675 , \25676 ,
         \25677 , \25678 , \25679 , \25680 , \25681 , \25682 , \25683 , \25684 , \25685 , \25686 ,
         \25687 , \25688 , \25689 , \25690 , \25691 , \25692 , \25693 , \25694 , \25695 , \25696 ,
         \25697 , \25698 , \25699 , \25700 , \25701 , \25702 , \25703 , \25704 , \25705 , \25706 ,
         \25707 , \25708 , \25709 , \25710 , \25711 , \25712 , \25713 , \25714 , \25715 , \25716 ,
         \25717 , \25718 , \25719 , \25720 , \25721 , \25722 , \25723 , \25724 , \25725 , \25726 ,
         \25727 , \25728 , \25729 , \25730 , \25731 , \25732 , \25733 , \25734 , \25735 , \25736 ,
         \25737 , \25738 , \25739 , \25740 , \25741 , \25742 , \25743 , \25744 , \25745 , \25746 ,
         \25747 , \25748 , \25749 , \25750 , \25751 , \25752 , \25753 , \25754 , \25755 , \25756 ,
         \25757 , \25758 , \25759 , \25760 , \25761 , \25762 , \25763 , \25764 , \25765 , \25766 ,
         \25767 , \25768_nG5d2d , \25769_nG5d2e , \25770 , \25771 , \25772 , \25773 , \25774 , \25775 , \25776 ,
         \25777 , \25778 , \25779 , \25780 , \25781 , \25782 , \25783 , \25784 , \25785 , \25786 ,
         \25787 , \25788 , \25789 , \25790 , \25791 , \25792 , \25793 , \25794 , \25795 , \25796 ,
         \25797 , \25798 , \25799 , \25800 , \25801 , \25802 , \25803 , \25804 , \25805 , \25806 ,
         \25807 , \25808 , \25809 , \25810 , \25811 , \25812_nG65bc , \25813_nG65bd , \25814_nG65be , \25815 , \25816 ,
         \25817 , \25818 , \25819 , \25820 , \25821 , \25822 , \25823 , \25824 , \25825 , \25826 ,
         \25827 , \25828 , \25829 , \25830 , \25831 , \25832 , \25833 , \25834 , \25835 , \25836 ,
         \25837 , \25838 , \25839 , \25840 , \25841 , \25842 , \25843 , \25844 , \25845 , \25846 ,
         \25847 , \25848 , \25849 , \25850 , \25851 , \25852 , \25853 , \25854 , \25855 , \25856 ,
         \25857 , \25858 , \25859 , \25860_nG9bc9 , \25861 , \25862 , \25863 , \25864 , \25865 , \25866 ,
         \25867 , \25868 , \25869 , \25870 , \25871 , \25872 , \25873 , \25874 , \25875 , \25876 ,
         \25877 , \25878 , \25879 , \25880 , \25881 , \25882 , \25883 , \25884 , \25885 , \25886 ,
         \25887 , \25888 , \25889 , \25890 , \25891 , \25892 , \25893 , \25894 , \25895 , \25896 ,
         \25897 , \25898 , \25899 , \25900 , \25901 , \25902 , \25903 , \25904 , \25905 , \25906 ,
         \25907 , \25908 , \25909 , \25910 , \25911 , \25912 , \25913 , \25914 , \25915 , \25916 ,
         \25917 , \25918 , \25919 , \25920 , \25921 , \25922 , \25923 , \25924 , \25925 , \25926 ,
         \25927 , \25928 , \25929 , \25930 , \25931 , \25932 , \25933 , \25934 , \25935 , \25936 ,
         \25937 , \25938 , \25939 , \25940 , \25941 , \25942 , \25943 , \25944 , \25945 , \25946 ,
         \25947 , \25948 , \25949 , \25950 , \25951 , \25952 , \25953 , \25954 , \25955 , \25956 ,
         \25957 , \25958 , \25959 , \25960 , \25961 , \25962 , \25963 , \25964 , \25965 , \25966 ,
         \25967 , \25968 , \25969 , \25970 , \25971 , \25972 , \25973 , \25974 , \25975 , \25976 ,
         \25977 , \25978 , \25979 , \25980 , \25981 , \25982 , \25983 , \25984 , \25985 , \25986 ,
         \25987 , \25988 , \25989 , \25990 , \25991 , \25992 , \25993 , \25994 , \25995 , \25996 ,
         \25997 , \25998 , \25999 , \26000 , \26001 , \26002 , \26003 , \26004 , \26005 , \26006 ,
         \26007 , \26008 , \26009 , \26010 , \26011_nG2553 , \26012 , \26013 , \26014 , \26015 , \26016 ,
         \26017 , \26018 , \26019 , \26020 , \26021 , \26022 , \26023 , \26024 , \26025 , \26026 ,
         \26027 , \26028 , \26029 , \26030 , \26031 , \26032 , \26033 , \26034 , \26035 , \26036 ,
         \26037 , \26038 , \26039 , \26040 , \26041 , \26042 , \26043 , \26044 , \26045 , \26046 ,
         \26047 , \26048 , \26049 , \26050 , \26051 , \26052 , \26053 , \26054 , \26055 , \26056 ,
         \26057 , \26058 , \26059 , \26060 , \26061 , \26062 , \26063 , \26064 , \26065 , \26066 ,
         \26067 , \26068 , \26069 , \26070 , \26071 , \26072 , \26073 , \26074 , \26075 , \26076 ,
         \26077 , \26078 , \26079 , \26080 , \26081 , \26082 , \26083 , \26084 , \26085 , \26086 ,
         \26087 , \26088 , \26089 , \26090 , \26091 , \26092 , \26093 , \26094 , \26095 , \26096 ,
         \26097 , \26098 , \26099 , \26100 , \26101 , \26102 , \26103 , \26104 , \26105 , \26106 ,
         \26107 , \26108 , \26109 , \26110 , \26111 , \26112 , \26113 , \26114 , \26115 , \26116 ,
         \26117 , \26118 , \26119 , \26120 , \26121 , \26122 , \26123 , \26124 , \26125 , \26126 ,
         \26127 , \26128 , \26129 , \26130 , \26131 , \26132 , \26133 , \26134 , \26135 , \26136 ,
         \26137 , \26138 , \26139 , \26140 , \26141 , \26142 , \26143 , \26144_nG3680 , \26145 , \26146 ,
         \26147 , \26148 , \26149 , \26150 , \26151 , \26152 , \26153 , \26154 , \26155 , \26156 ,
         \26157 , \26158 , \26159 , \26160 , \26161 , \26162 , \26163 , \26164 , \26165 , \26166 ,
         \26167 , \26168 , \26169 , \26170 , \26171 , \26172 , \26173 , \26174 , \26175 , \26176 ,
         \26177 , \26178 , \26179 , \26180 , \26181 , \26182 , \26183 , \26184 , \26185 , \26186 ,
         \26187 , \26188 , \26189 , \26190 , \26191 , \26192 , \26193 , \26194 , \26195 , \26196 ,
         \26197 , \26198 , \26199 , \26200 , \26201 , \26202 , \26203 , \26204 , \26205 , \26206 ,
         \26207 , \26208 , \26209 , \26210 , \26211 , \26212 , \26213 , \26214 , \26215 , \26216 ,
         \26217 , \26218 , \26219 , \26220 , \26221 , \26222 , \26223 , \26224 , \26225 , \26226 ,
         \26227 , \26228 , \26229 , \26230 , \26231 , \26232 , \26233 , \26234 , \26235 , \26236 ,
         \26237 , \26238 , \26239 , \26240 , \26241 , \26242 , \26243 , \26244 , \26245 , \26246 ,
         \26247 , \26248 , \26249 , \26250 , \26251 , \26252 , \26253 , \26254 , \26255 , \26256 ,
         \26257 , \26258 , \26259 , \26260 , \26261 , \26262 , \26263 , \26264 , \26265 , \26266 ,
         \26267 , \26268 , \26269 , \26270 , \26271 , \26272 , \26273 , \26274 , \26275 , \26276 ,
         \26277 , \26278_nG25d8 , \26279 , \26280 , \26281 , \26282 , \26283 , \26284 , \26285 , \26286 ,
         \26287 , \26288 , \26289 , \26290 , \26291 , \26292 , \26293 , \26294 , \26295 , \26296 ,
         \26297 , \26298 , \26299 , \26300 , \26301 , \26302 , \26303 , \26304 , \26305 , \26306 ,
         \26307 , \26308 , \26309 , \26310 , \26311 , \26312 , \26313 , \26314 , \26315 , \26316 ,
         \26317 , \26318 , \26319 , \26320 , \26321 , \26322 , \26323 , \26324 , \26325 , \26326 ,
         \26327 , \26328 , \26329 , \26330 , \26331 , \26332 , \26333 , \26334 , \26335 , \26336 ,
         \26337 , \26338 , \26339 , \26340 , \26341 , \26342 , \26343 , \26344 , \26345 , \26346 ,
         \26347 , \26348 , \26349 , \26350 , \26351 , \26352 , \26353 , \26354 , \26355 , \26356 ,
         \26357 , \26358 , \26359 , \26360 , \26361 , \26362 , \26363 , \26364 , \26365 , \26366 ,
         \26367 , \26368 , \26369 , \26370 , \26371 , \26372 , \26373 , \26374 , \26375 , \26376 ,
         \26377 , \26378 , \26379 , \26380 , \26381 , \26382 , \26383 , \26384 , \26385 , \26386 ,
         \26387 , \26388 , \26389 , \26390 , \26391 , \26392 , \26393 , \26394 , \26395 , \26396 ,
         \26397 , \26398 , \26399 , \26400 , \26401 , \26402 , \26403 , \26404 , \26405 , \26406 ,
         \26407 , \26408 , \26409 , \26410 , \26411_nG3705 , \26412 , \26413 , \26414 , \26415 , \26416 ,
         \26417 , \26418 , \26419 , \26420 , \26421 , \26422_nG440c , \26423 , \26424 , \26425_nG440f , \26426 ,
         \26427 , \26428 , \26429 , \26430 , \26431 , \26432 , \26433 , \26434 , \26435 , \26436 ,
         \26437 , \26438 , \26439 , \26440 , \26441 , \26442 , \26443 , \26444 , \26445 , \26446 ,
         \26447 , \26448 , \26449 , \26450 , \26451 , \26452 , \26453 , \26454 , \26455 , \26456 ,
         \26457 , \26458 , \26459 , \26460 , \26461 , \26462 , \26463 , \26464 , \26465 , \26466 ,
         \26467 , \26468 , \26469 , \26470 , \26471 , \26472 , \26473 , \26474 , \26475 , \26476 ,
         \26477 , \26478 , \26479 , \26480 , \26481 , \26482 , \26483 , \26484 , \26485 , \26486 ,
         \26487 , \26488 , \26489 , \26490 , \26491 , \26492 , \26493 , \26494 , \26495 , \26496 ,
         \26497 , \26498 , \26499 , \26500 , \26501 , \26502 , \26503 , \26504 , \26505 , \26506 ,
         \26507 , \26508 , \26509 , \26510 , \26511 , \26512 , \26513 , \26514 , \26515 , \26516 ,
         \26517 , \26518 , \26519 , \26520 , \26521 , \26522 , \26523 , \26524 , \26525 , \26526 ,
         \26527 , \26528 , \26529 , \26530 , \26531 , \26532 , \26533 , \26534 , \26535 , \26536 ,
         \26537 , \26538 , \26539 , \26540 , \26541 , \26542 , \26543 , \26544 , \26545 , \26546 ,
         \26547 , \26548 , \26549 , \26550 , \26551 , \26552 , \26553 , \26554 , \26555 , \26556 ,
         \26557 , \26558 , \26559 , \26560 , \26561 , \26562 , \26563 , \26564 , \26565 , \26566 ,
         \26567 , \26568 , \26569 , \26570 , \26571 , \26572 , \26573 , \26574 , \26575 , \26576 ,
         \26577 , \26578 , \26579 , \26580 , \26581 , \26582 , \26583 , \26584 , \26585 , \26586 ,
         \26587 , \26588 , \26589 , \26590 , \26591 , \26592 , \26593 , \26594 , \26595 , \26596 ,
         \26597 , \26598 , \26599 , \26600 , \26601 , \26602 , \26603 , \26604 , \26605 , \26606 ,
         \26607 , \26608 , \26609 , \26610 , \26611 , \26612 , \26613 , \26614 , \26615 , \26616 ,
         \26617 , \26618 , \26619 , \26620 , \26621 , \26622 , \26623 , \26624 , \26625 , \26626 ,
         \26627 , \26628 , \26629 , \26630 , \26631 , \26632 , \26633 , \26634 , \26635 , \26636 ,
         \26637 , \26638 , \26639 , \26640 , \26641 , \26642 , \26643 , \26644 , \26645 , \26646 ,
         \26647 , \26648 , \26649 , \26650 , \26651 , \26652 , \26653 , \26654 , \26655 , \26656 ,
         \26657 , \26658 , \26659 , \26660 , \26661 , \26662 , \26663 , \26664 , \26665 , \26666 ,
         \26667 , \26668 , \26669 , \26670 , \26671 , \26672_nG5db2 , \26673 , \26674 , \26675 , \26676 ,
         \26677 , \26678 , \26679 , \26680 , \26681 , \26682 , \26683 , \26684 , \26685 , \26686 ,
         \26687 , \26688 , \26689 , \26690 , \26691 , \26692 , \26693 , \26694 , \26695 , \26696 ,
         \26697 , \26698 , \26699 , \26700 , \26701 , \26702 , \26703 , \26704 , \26705 , \26706 ,
         \26707 , \26708 , \26709 , \26710 , \26711 , \26712 , \26713 , \26714 , \26715 , \26716 ,
         \26717 , \26718 , \26719 , \26720 , \26721 , \26722 , \26723 , \26724 , \26725 , \26726 ,
         \26727 , \26728 , \26729 , \26730 , \26731 , \26732 , \26733 , \26734 , \26735 , \26736 ,
         \26737 , \26738 , \26739 , \26740 , \26741 , \26742 , \26743 , \26744 , \26745 , \26746 ,
         \26747 , \26748 , \26749 , \26750 , \26751 , \26752 , \26753 , \26754 , \26755 , \26756 ,
         \26757 , \26758 , \26759 , \26760 , \26761 , \26762 , \26763 , \26764 , \26765 , \26766 ,
         \26767 , \26768 , \26769 , \26770 , \26771 , \26772 , \26773 , \26774 , \26775 , \26776 ,
         \26777 , \26778 , \26779 , \26780 , \26781 , \26782 , \26783 , \26784 , \26785 , \26786 ,
         \26787 , \26788 , \26789 , \26790 , \26791 , \26792 , \26793 , \26794 , \26795 , \26796 ,
         \26797 , \26798 , \26799 , \26800 , \26801 , \26802 , \26803 , \26804_nG5e36 , \26805_nG5e37 , \26806 ,
         \26807 , \26808 , \26809 , \26810 , \26811 , \26812 , \26813 , \26814 , \26815 , \26816 ,
         \26817 , \26818 , \26819 , \26820 , \26821 , \26822 , \26823 , \26824 , \26825 , \26826_nG65bf ,
         \26827_nG65c0 , \26828_nG65c1 , \26829 , \26830 , \26831 , \26832 , \26833 , \26834 , \26835 , \26836 ,
         \26837 , \26838 , \26839 , \26840 , \26841 , \26842 , \26843 , \26844 , \26845 , \26846 ,
         \26847 , \26848 , \26849 , \26850 , \26851 , \26852 , \26853 , \26854 , \26855 , \26856 ,
         \26857 , \26858 , \26859 , \26860 , \26861 , \26862 , \26863 , \26864 , \26865 , \26866 ,
         \26867 , \26868 , \26869 , \26870 , \26871 , \26872 , \26873 , \26874 , \26875 , \26876 ,
         \26877 , \26878 , \26879 , \26880 , \26881 , \26882 , \26883 , \26884 , \26885 , \26886 ,
         \26887_nG9bc6 , \26888 , \26889 , \26890 , \26891 , \26892 , \26893 , \26894 , \26895 , \26896 ,
         \26897 , \26898 , \26899 , \26900 , \26901 , \26902 , \26903 , \26904 , \26905 , \26906 ,
         \26907 , \26908 , \26909 , \26910 , \26911 , \26912 , \26913 , \26914 , \26915 , \26916 ,
         \26917 , \26918 , \26919 , \26920 , \26921 , \26922 , \26923 , \26924 , \26925 , \26926 ,
         \26927 , \26928 , \26929 , \26930 , \26931 , \26932 , \26933 , \26934 , \26935 , \26936 ,
         \26937 , \26938 , \26939 , \26940 , \26941 , \26942 , \26943 , \26944 , \26945 , \26946 ,
         \26947 , \26948 , \26949 , \26950 , \26951 , \26952 , \26953 , \26954 , \26955 , \26956 ,
         \26957 , \26958 , \26959 , \26960 , \26961 , \26962 , \26963 , \26964 , \26965 , \26966 ,
         \26967 , \26968 , \26969 , \26970 , \26971 , \26972 , \26973 , \26974 , \26975 , \26976 ,
         \26977 , \26978 , \26979 , \26980 , \26981 , \26982 , \26983 , \26984 , \26985 , \26986 ,
         \26987 , \26988 , \26989 , \26990 , \26991 , \26992 , \26993 , \26994 , \26995 , \26996 ,
         \26997 , \26998 , \26999 , \27000 , \27001 , \27002 , \27003 , \27004 , \27005 , \27006 ,
         \27007 , \27008 , \27009 , \27010 , \27011 , \27012 , \27013 , \27014 , \27015 , \27016 ,
         \27017 , \27018 , \27019 , \27020 , \27021 , \27022 , \27023 , \27024 , \27025 , \27026 ,
         \27027 , \27028 , \27029 , \27030 , \27031 , \27032 , \27033 , \27034 , \27035 , \27036 ,
         \27037 , \27038 , \27039 , \27040 , \27041 , \27042 , \27043 , \27044 , \27045 , \27046 ,
         \27047 , \27048 , \27049 , \27050 , \27051 , \27052 , \27053 , \27054 , \27055 , \27056 ,
         \27057 , \27058 , \27059 , \27060 , \27061 , \27062 , \27063 , \27064 , \27065 , \27066 ,
         \27067 , \27068 , \27069 , \27070 , \27071 , \27072 , \27073 , \27074 , \27075 , \27076 ,
         \27077 , \27078 , \27079 , \27080 , \27081 , \27082 , \27083 , \27084 , \27085 , \27086 ,
         \27087 , \27088 , \27089 , \27090 , \27091 , \27092 , \27093 , \27094 , \27095 , \27096 ,
         \27097 , \27098 , \27099 , \27100 , \27101 , \27102 , \27103 , \27104 , \27105 , \27106 ,
         \27107 , \27108 , \27109 , \27110 , \27111 , \27112 , \27113 , \27114 , \27115 , \27116 ,
         \27117 , \27118 , \27119 , \27120 , \27121 , \27122 , \27123 , \27124 , \27125 , \27126 ,
         \27127 , \27128 , \27129 , \27130 , \27131 , \27132 , \27133 , \27134 , \27135 , \27136 ,
         \27137 , \27138 , \27139 , \27140 , \27141 , \27142 , \27143 , \27144 , \27145 , \27146 ,
         \27147 , \27148 , \27149 , \27150 , \27151 , \27152 , \27153 , \27154 , \27155 , \27156 ,
         \27157 , \27158_nG5ebb , \27159 , \27160 , \27161 , \27162 , \27163 , \27164 , \27165 , \27166 ,
         \27167 , \27168 , \27169 , \27170 , \27171 , \27172 , \27173 , \27174 , \27175 , \27176 ,
         \27177 , \27178 , \27179 , \27180 , \27181 , \27182 , \27183 , \27184 , \27185 , \27186 ,
         \27187 , \27188 , \27189 , \27190 , \27191 , \27192 , \27193 , \27194 , \27195 , \27196 ,
         \27197 , \27198 , \27199 , \27200 , \27201 , \27202 , \27203 , \27204 , \27205 , \27206 ,
         \27207 , \27208 , \27209 , \27210 , \27211 , \27212 , \27213 , \27214 , \27215 , \27216 ,
         \27217 , \27218 , \27219 , \27220 , \27221 , \27222 , \27223 , \27224 , \27225 , \27226 ,
         \27227 , \27228 , \27229 , \27230 , \27231 , \27232 , \27233 , \27234 , \27235 , \27236 ,
         \27237 , \27238 , \27239 , \27240 , \27241 , \27242 , \27243 , \27244 , \27245 , \27246 ,
         \27247 , \27248 , \27249 , \27250 , \27251 , \27252 , \27253 , \27254 , \27255 , \27256 ,
         \27257 , \27258 , \27259 , \27260 , \27261 , \27262 , \27263 , \27264 , \27265 , \27266 ,
         \27267 , \27268 , \27269 , \27270 , \27271 , \27272 , \27273 , \27274 , \27275 , \27276 ,
         \27277 , \27278 , \27279 , \27280 , \27281 , \27282 , \27283 , \27284 , \27285 , \27286 ,
         \27287 , \27288 , \27289 , \27290_nG5f3f , \27291_nG5f40 , \27292 , \27293 , \27294 , \27295 , \27296 ,
         \27297 , \27298 , \27299 , \27300 , \27301 , \27302 , \27303 , \27304 , \27305 , \27306 ,
         \27307 , \27308 , \27309 , \27310_nG65c2 , \27311_nG65c3 , \27312_nG65c4 , \27313 , \27314 , \27315 , \27316 ,
         \27317 , \27318 , \27319 , \27320 , \27321 , \27322 , \27323 , \27324 , \27325 , \27326 ,
         \27327 , \27328 , \27329 , \27330 , \27331 , \27332 , \27333 , \27334 , \27335 , \27336 ,
         \27337 , \27338 , \27339 , \27340 , \27341 , \27342 , \27343 , \27344 , \27345 , \27346 ,
         \27347 , \27348 , \27349 , \27350 , \27351 , \27352 , \27353 , \27354 , \27355 , \27356 ,
         \27357 , \27358 , \27359 , \27360 , \27361 , \27362 , \27363 , \27364 , \27365 , \27366 ,
         \27367 , \27368 , \27369 , \27370 , \27371 , \27372 , \27373 , \27374 , \27375 , \27376 ,
         \27377 , \27378 , \27379 , \27380 , \27381 , \27382 , \27383 , \27384 , \27385 , \27386 ,
         \27387 , \27388 , \27389 , \27390 , \27391 , \27392 , \27393 , \27394 , \27395 , \27396 ,
         \27397 , \27398 , \27399 , \27400 , \27401 , \27402 , \27403 , \27404 , \27405 , \27406 ,
         \27407 , \27408 , \27409 , \27410 , \27411 , \27412 , \27413 , \27414 , \27415 , \27416_nG9bc3 ,
         \27417 , \27418 , \27419 , \27420 , \27421 , \27422 , \27423 , \27424 , \27425 , \27426 ,
         \27427 , \27428 , \27429 , \27430 , \27431 , \27432 , \27433 , \27434 , \27435 , \27436 ,
         \27437 , \27438 , \27439 , \27440 , \27441 , \27442 , \27443 , \27444 , \27445 , \27446 ,
         \27447 , \27448 , \27449 , \27450 , \27451 , \27452 , \27453 , \27454 , \27455 , \27456 ,
         \27457 , \27458 , \27459 , \27460 , \27461 , \27462 , \27463 , \27464 , \27465 , \27466 ,
         \27467 , \27468 , \27469 , \27470 , \27471 , \27472 , \27473 , \27474 , \27475 , \27476 ,
         \27477 , \27478 , \27479 , \27480 , \27481 , \27482 , \27483 , \27484 , \27485 , \27486 ,
         \27487 , \27488 , \27489 , \27490 , \27491 , \27492 , \27493 , \27494 , \27495 , \27496 ,
         \27497 , \27498 , \27499 , \27500 , \27501 , \27502 , \27503 , \27504 , \27505 , \27506 ,
         \27507 , \27508 , \27509 , \27510 , \27511 , \27512 , \27513 , \27514 , \27515 , \27516 ,
         \27517 , \27518 , \27519 , \27520 , \27521 , \27522 , \27523 , \27524 , \27525 , \27526 ,
         \27527 , \27528 , \27529 , \27530 , \27531 , \27532 , \27533 , \27534 , \27535 , \27536 ,
         \27537 , \27538 , \27539 , \27540 , \27541 , \27542 , \27543 , \27544 , \27545 , \27546 ,
         \27547 , \27548 , \27549 , \27550 , \27551 , \27552 , \27553 , \27554 , \27555 , \27556 ,
         \27557 , \27558 , \27559 , \27560 , \27561 , \27562 , \27563 , \27564 , \27565 , \27566 ,
         \27567 , \27568 , \27569 , \27570 , \27571 , \27572 , \27573 , \27574 , \27575 , \27576 ,
         \27577 , \27578 , \27579 , \27580 , \27581 , \27582 , \27583 , \27584 , \27585 , \27586 ,
         \27587 , \27588 , \27589 , \27590 , \27591 , \27592 , \27593 , \27594 , \27595 , \27596 ,
         \27597 , \27598 , \27599 , \27600 , \27601 , \27602 , \27603 , \27604 , \27605 , \27606 ,
         \27607 , \27608 , \27609 , \27610 , \27611 , \27612 , \27613 , \27614 , \27615 , \27616 ,
         \27617 , \27618 , \27619 , \27620 , \27621 , \27622 , \27623 , \27624 , \27625 , \27626 ,
         \27627 , \27628 , \27629 , \27630 , \27631 , \27632 , \27633 , \27634 , \27635 , \27636 ,
         \27637 , \27638 , \27639 , \27640 , \27641 , \27642 , \27643 , \27644 , \27645 , \27646 ,
         \27647 , \27648 , \27649 , \27650 , \27651 , \27652 , \27653 , \27654 , \27655 , \27656 ,
         \27657 , \27658 , \27659 , \27660 , \27661 , \27662 , \27663 , \27664 , \27665 , \27666 ,
         \27667 , \27668 , \27669 , \27670 , \27671 , \27672 , \27673 , \27674 , \27675 , \27676 ,
         \27677 , \27678 , \27679 , \27680 , \27681 , \27682 , \27683 , \27684 , \27685 , \27686 ,
         \27687 , \27688 , \27689 , \27690 , \27691 , \27692 , \27693 , \27694 , \27695 , \27696 ,
         \27697 , \27698_nG2449 , \27699 , \27700 , \27701 , \27702 , \27703 , \27704 , \27705 , \27706 ,
         \27707 , \27708 , \27709 , \27710 , \27711 , \27712 , \27713 , \27714 , \27715 , \27716 ,
         \27717 , \27718 , \27719 , \27720 , \27721 , \27722 , \27723 , \27724 , \27725 , \27726 ,
         \27727 , \27728 , \27729 , \27730 , \27731 , \27732 , \27733 , \27734 , \27735 , \27736 ,
         \27737 , \27738 , \27739 , \27740 , \27741 , \27742 , \27743 , \27744 , \27745 , \27746 ,
         \27747 , \27748 , \27749 , \27750 , \27751 , \27752 , \27753 , \27754 , \27755 , \27756 ,
         \27757 , \27758 , \27759 , \27760 , \27761 , \27762 , \27763 , \27764 , \27765 , \27766 ,
         \27767 , \27768 , \27769 , \27770 , \27771 , \27772 , \27773 , \27774 , \27775 , \27776 ,
         \27777 , \27778 , \27779 , \27780 , \27781 , \27782 , \27783 , \27784 , \27785 , \27786 ,
         \27787 , \27788 , \27789 , \27790 , \27791 , \27792 , \27793 , \27794 , \27795 , \27796 ,
         \27797 , \27798 , \27799 , \27800 , \27801 , \27802 , \27803 , \27804 , \27805 , \27806 ,
         \27807 , \27808 , \27809 , \27810 , \27811 , \27812 , \27813 , \27814 , \27815 , \27816 ,
         \27817 , \27818 , \27819 , \27820 , \27821 , \27822 , \27823 , \27824 , \27825 , \27826 ,
         \27827 , \27828 , \27829 , \27830 , \27831_nG3576 , \27832 , \27833 , \27834 , \27835 , \27836 ,
         \27837 , \27838 , \27839 , \27840 , \27841 , \27842 , \27843 , \27844 , \27845 , \27846 ,
         \27847 , \27848 , \27849 , \27850 , \27851 , \27852 , \27853 , \27854 , \27855 , \27856 ,
         \27857 , \27858 , \27859 , \27860 , \27861 , \27862 , \27863 , \27864 , \27865 , \27866 ,
         \27867 , \27868 , \27869 , \27870 , \27871 , \27872 , \27873 , \27874 , \27875 , \27876 ,
         \27877 , \27878 , \27879 , \27880 , \27881 , \27882 , \27883 , \27884 , \27885 , \27886 ,
         \27887 , \27888 , \27889 , \27890 , \27891 , \27892 , \27893 , \27894 , \27895 , \27896 ,
         \27897 , \27898 , \27899 , \27900 , \27901 , \27902 , \27903 , \27904 , \27905 , \27906 ,
         \27907 , \27908 , \27909 , \27910 , \27911 , \27912 , \27913 , \27914 , \27915 , \27916 ,
         \27917 , \27918 , \27919 , \27920 , \27921 , \27922 , \27923 , \27924 , \27925 , \27926 ,
         \27927 , \27928 , \27929 , \27930 , \27931 , \27932 , \27933 , \27934 , \27935 , \27936 ,
         \27937 , \27938 , \27939 , \27940 , \27941 , \27942 , \27943 , \27944 , \27945 , \27946 ,
         \27947 , \27948 , \27949 , \27950 , \27951 , \27952 , \27953 , \27954 , \27955 , \27956 ,
         \27957 , \27958 , \27959 , \27960 , \27961 , \27962 , \27963 , \27964 , \27965_nG24ce , \27966 ,
         \27967 , \27968 , \27969 , \27970 , \27971 , \27972 , \27973 , \27974 , \27975 , \27976 ,
         \27977 , \27978 , \27979 , \27980 , \27981 , \27982 , \27983 , \27984 , \27985 , \27986 ,
         \27987 , \27988 , \27989 , \27990 , \27991 , \27992 , \27993 , \27994 , \27995 , \27996 ,
         \27997 , \27998 , \27999 , \28000 , \28001 , \28002 , \28003 , \28004 , \28005 , \28006 ,
         \28007 , \28008 , \28009 , \28010 , \28011 , \28012 , \28013 , \28014 , \28015 , \28016 ,
         \28017 , \28018 , \28019 , \28020 , \28021 , \28022 , \28023 , \28024 , \28025 , \28026 ,
         \28027 , \28028 , \28029 , \28030 , \28031 , \28032 , \28033 , \28034 , \28035 , \28036 ,
         \28037 , \28038 , \28039 , \28040 , \28041 , \28042 , \28043 , \28044 , \28045 , \28046 ,
         \28047 , \28048 , \28049 , \28050 , \28051 , \28052 , \28053 , \28054 , \28055 , \28056 ,
         \28057 , \28058 , \28059 , \28060 , \28061 , \28062 , \28063 , \28064 , \28065 , \28066 ,
         \28067 , \28068 , \28069 , \28070 , \28071 , \28072 , \28073 , \28074 , \28075 , \28076 ,
         \28077 , \28078 , \28079 , \28080 , \28081 , \28082 , \28083 , \28084 , \28085 , \28086 ,
         \28087 , \28088 , \28089 , \28090 , \28091 , \28092 , \28093 , \28094 , \28095 , \28096 ,
         \28097 , \28098_nG35fb , \28099 , \28100 , \28101 , \28102 , \28103 , \28104 , \28105 , \28106 ,
         \28107 , \28108 , \28109_nG4406 , \28110 , \28111 , \28112_nG4409 , \28113 , \28114 , \28115 , \28116 ,
         \28117 , \28118 , \28119 , \28120 , \28121 , \28122 , \28123 , \28124 , \28125 , \28126 ,
         \28127 , \28128 , \28129 , \28130 , \28131 , \28132 , \28133 , \28134 , \28135 , \28136 ,
         \28137 , \28138 , \28139 , \28140 , \28141 , \28142 , \28143 , \28144 , \28145 , \28146 ,
         \28147 , \28148 , \28149 , \28150 , \28151 , \28152 , \28153 , \28154 , \28155 , \28156 ,
         \28157 , \28158 , \28159 , \28160 , \28161 , \28162 , \28163 , \28164 , \28165 , \28166 ,
         \28167 , \28168 , \28169 , \28170 , \28171 , \28172 , \28173 , \28174 , \28175 , \28176 ,
         \28177 , \28178 , \28179 , \28180 , \28181 , \28182 , \28183 , \28184 , \28185 , \28186 ,
         \28187 , \28188 , \28189 , \28190 , \28191 , \28192 , \28193 , \28194 , \28195 , \28196 ,
         \28197 , \28198 , \28199 , \28200 , \28201 , \28202 , \28203 , \28204 , \28205 , \28206 ,
         \28207 , \28208 , \28209 , \28210 , \28211 , \28212 , \28213 , \28214 , \28215 , \28216 ,
         \28217 , \28218 , \28219 , \28220 , \28221 , \28222 , \28223 , \28224 , \28225 , \28226 ,
         \28227 , \28228 , \28229 , \28230 , \28231 , \28232 , \28233 , \28234 , \28235 , \28236 ,
         \28237 , \28238 , \28239 , \28240 , \28241 , \28242 , \28243 , \28244 , \28245 , \28246 ,
         \28247 , \28248 , \28249 , \28250 , \28251 , \28252 , \28253 , \28254 , \28255 , \28256 ,
         \28257 , \28258 , \28259 , \28260 , \28261 , \28262 , \28263 , \28264 , \28265 , \28266 ,
         \28267 , \28268 , \28269 , \28270 , \28271 , \28272 , \28273 , \28274 , \28275 , \28276 ,
         \28277 , \28278 , \28279 , \28280 , \28281 , \28282 , \28283 , \28284 , \28285 , \28286 ,
         \28287 , \28288 , \28289 , \28290 , \28291 , \28292 , \28293 , \28294 , \28295 , \28296 ,
         \28297 , \28298 , \28299 , \28300 , \28301 , \28302 , \28303 , \28304 , \28305 , \28306 ,
         \28307 , \28308 , \28309 , \28310 , \28311 , \28312 , \28313 , \28314 , \28315 , \28316 ,
         \28317 , \28318 , \28319 , \28320 , \28321 , \28322 , \28323 , \28324 , \28325 , \28326 ,
         \28327 , \28328 , \28329 , \28330 , \28331 , \28332 , \28333 , \28334 , \28335 , \28336 ,
         \28337 , \28338 , \28339 , \28340 , \28341 , \28342 , \28343 , \28344 , \28345 , \28346 ,
         \28347 , \28348 , \28349 , \28350 , \28351 , \28352 , \28353 , \28354 , \28355 , \28356 ,
         \28357 , \28358 , \28359 , \28360 , \28361 , \28362 , \28363 , \28364 , \28365 , \28366 ,
         \28367 , \28368 , \28369 , \28370 , \28371 , \28372 , \28373 , \28374 , \28375 , \28376 ,
         \28377 , \28378 , \28379 , \28380 , \28381 , \28382 , \28383 , \28384 , \28385 , \28386 ,
         \28387 , \28388 , \28389 , \28390 , \28391_nG5fc4 , \28392 , \28393 , \28394 , \28395 , \28396 ,
         \28397 , \28398 , \28399 , \28400 , \28401 , \28402 , \28403 , \28404 , \28405 , \28406 ,
         \28407 , \28408 , \28409 , \28410 , \28411 , \28412 , \28413 , \28414 , \28415 , \28416 ,
         \28417 , \28418 , \28419 , \28420 , \28421 , \28422 , \28423 , \28424 , \28425 , \28426 ,
         \28427 , \28428 , \28429 , \28430 , \28431 , \28432 , \28433 , \28434 , \28435 , \28436 ,
         \28437 , \28438 , \28439 , \28440 , \28441 , \28442 , \28443 , \28444 , \28445 , \28446 ,
         \28447 , \28448 , \28449 , \28450 , \28451 , \28452 , \28453 , \28454 , \28455 , \28456 ,
         \28457 , \28458 , \28459 , \28460 , \28461 , \28462 , \28463 , \28464 , \28465 , \28466 ,
         \28467 , \28468 , \28469 , \28470 , \28471 , \28472 , \28473 , \28474 , \28475 , \28476 ,
         \28477 , \28478 , \28479 , \28480 , \28481 , \28482 , \28483 , \28484 , \28485 , \28486 ,
         \28487 , \28488 , \28489 , \28490 , \28491 , \28492 , \28493 , \28494 , \28495 , \28496 ,
         \28497 , \28498 , \28499 , \28500 , \28501 , \28502 , \28503 , \28504 , \28505 , \28506 ,
         \28507 , \28508 , \28509 , \28510 , \28511 , \28512 , \28513 , \28514 , \28515 , \28516 ,
         \28517 , \28518 , \28519 , \28520 , \28521 , \28522 , \28523_nG6048 , \28524_nG6049 , \28525 , \28526 ,
         \28527 , \28528 , \28529 , \28530 , \28531_nG65c5 , \28532_nG65c6 , \28533_nG65c7 , \28534 , \28535 , \28536 ,
         \28537 , \28538 , \28539 , \28540 , \28541 , \28542 , \28543 , \28544 , \28545 , \28546 ,
         \28547 , \28548 , \28549 , \28550 , \28551 , \28552 , \28553 , \28554 , \28555 , \28556 ,
         \28557 , \28558 , \28559 , \28560 , \28561 , \28562 , \28563 , \28564 , \28565 , \28566 ,
         \28567 , \28568 , \28569 , \28570 , \28571 , \28572 , \28573 , \28574 , \28575 , \28576 ,
         \28577 , \28578 , \28579 , \28580 , \28581 , \28582 , \28583 , \28584 , \28585 , \28586 ,
         \28587 , \28588 , \28589 , \28590 , \28591 , \28592 , \28593 , \28594 , \28595 , \28596 ,
         \28597 , \28598 , \28599 , \28600 , \28601 , \28602_nG9bc0 , \28603 , \28604 , \28605 , \28606 ,
         \28607 , \28608 , \28609 , \28610 , \28611 , \28612 , \28613 , \28614 , \28615 , \28616 ,
         \28617 , \28618 , \28619 , \28620 , \28621 , \28622 , \28623 , \28624 , \28625 , \28626 ,
         \28627 , \28628 , \28629 , \28630 , \28631 , \28632 , \28633 , \28634 , \28635 , \28636 ,
         \28637 , \28638 , \28639 , \28640 , \28641 , \28642 , \28643 , \28644 , \28645 , \28646 ,
         \28647 , \28648 , \28649 , \28650 , \28651 , \28652 , \28653 , \28654 , \28655 , \28656 ,
         \28657 , \28658 , \28659 , \28660 , \28661 , \28662 , \28663 , \28664 , \28665 , \28666 ,
         \28667 , \28668 , \28669 , \28670 , \28671 , \28672 , \28673 , \28674 , \28675 , \28676 ,
         \28677 , \28678 , \28679 , \28680 , \28681 , \28682 , \28683 , \28684 , \28685 , \28686 ,
         \28687 , \28688 , \28689 , \28690 , \28691 , \28692 , \28693 , \28694 , \28695 , \28696 ,
         \28697 , \28698 , \28699 , \28700 , \28701 , \28702 , \28703 , \28704 , \28705 , \28706 ,
         \28707 , \28708 , \28709 , \28710 , \28711 , \28712 , \28713 , \28714 , \28715 , \28716 ,
         \28717 , \28718 , \28719 , \28720 , \28721 , \28722 , \28723 , \28724 , \28725 , \28726 ,
         \28727 , \28728 , \28729 , \28730 , \28731 , \28732 , \28733 , \28734 , \28735 , \28736 ,
         \28737 , \28738 , \28739 , \28740 , \28741 , \28742 , \28743 , \28744 , \28745 , \28746 ,
         \28747 , \28748 , \28749 , \28750 , \28751 , \28752 , \28753 , \28754 , \28755 , \28756 ,
         \28757 , \28758 , \28759 , \28760 , \28761 , \28762 , \28763 , \28764 , \28765 , \28766 ,
         \28767 , \28768 , \28769 , \28770 , \28771 , \28772 , \28773 , \28774 , \28775 , \28776 ,
         \28777 , \28778 , \28779 , \28780 , \28781 , \28782 , \28783 , \28784 , \28785 , \28786 ,
         \28787 , \28788 , \28789 , \28790 , \28791 , \28792 , \28793 , \28794 , \28795 , \28796 ,
         \28797 , \28798 , \28799 , \28800 , \28801 , \28802 , \28803 , \28804 , \28805 , \28806 ,
         \28807 , \28808 , \28809 , \28810 , \28811 , \28812 , \28813 , \28814 , \28815 , \28816 ,
         \28817 , \28818 , \28819 , \28820 , \28821 , \28822 , \28823 , \28824 , \28825 , \28826 ,
         \28827 , \28828 , \28829 , \28830 , \28831 , \28832 , \28833 , \28834 , \28835 , \28836 ,
         \28837 , \28838 , \28839 , \28840 , \28841 , \28842 , \28843 , \28844 , \28845 , \28846 ,
         \28847 , \28848 , \28849 , \28850 , \28851 , \28852 , \28853 , \28854 , \28855 , \28856 ,
         \28857 , \28858 , \28859 , \28860 , \28861 , \28862 , \28863 , \28864 , \28865 , \28866 ,
         \28867 , \28868 , \28869 , \28870 , \28871 , \28872 , \28873 , \28874 , \28875 , \28876 ,
         \28877 , \28878 , \28879 , \28880 , \28881 , \28882 , \28883 , \28884 , \28885 , \28886 ,
         \28887 , \28888 , \28889 , \28890 , \28891 , \28892 , \28893 , \28894 , \28895 , \28896 ,
         \28897 , \28898 , \28899 , \28900 , \28901 , \28902 , \28903 , \28904 , \28905 , \28906 ,
         \28907 , \28908 , \28909 , \28910 , \28911 , \28912 , \28913 , \28914 , \28915 , \28916 ,
         \28917 , \28918 , \28919 , \28920 , \28921 , \28922 , \28923 , \28924 , \28925 , \28926 ,
         \28927 , \28928 , \28929 , \28930 , \28931 , \28932 , \28933_nG60cd , \28934 , \28935 , \28936 ,
         \28937 , \28938 , \28939 , \28940 , \28941 , \28942 , \28943 , \28944 , \28945 , \28946 ,
         \28947 , \28948 , \28949 , \28950 , \28951 , \28952 , \28953 , \28954 , \28955 , \28956 ,
         \28957 , \28958 , \28959 , \28960 , \28961 , \28962 , \28963 , \28964 , \28965 , \28966 ,
         \28967 , \28968 , \28969 , \28970 , \28971 , \28972 , \28973 , \28974 , \28975 , \28976 ,
         \28977 , \28978 , \28979 , \28980 , \28981 , \28982 , \28983 , \28984 , \28985 , \28986 ,
         \28987 , \28988 , \28989 , \28990 , \28991 , \28992 , \28993 , \28994 , \28995 , \28996 ,
         \28997 , \28998 , \28999 , \29000 , \29001 , \29002 , \29003 , \29004 , \29005 , \29006 ,
         \29007 , \29008 , \29009 , \29010 , \29011 , \29012 , \29013 , \29014 , \29015 , \29016 ,
         \29017 , \29018 , \29019 , \29020 , \29021 , \29022 , \29023 , \29024 , \29025 , \29026 ,
         \29027 , \29028 , \29029 , \29030 , \29031 , \29032 , \29033 , \29034 , \29035 , \29036 ,
         \29037 , \29038 , \29039 , \29040 , \29041 , \29042 , \29043 , \29044 , \29045 , \29046 ,
         \29047 , \29048 , \29049 , \29050 , \29051 , \29052 , \29053 , \29054 , \29055 , \29056 ,
         \29057 , \29058 , \29059 , \29060 , \29061 , \29062 , \29063 , \29064 , \29065_nG6151 , \29066_nG6152 ,
         \29067 , \29068 , \29069 , \29070 , \29071 , \29072 , \29073 , \29074 , \29075 , \29076 ,
         \29077 , \29078 , \29079 , \29080 , \29081_nG65c8 , \29082_nG65c9 , \29083_nG65ca , \29084 , \29085 , \29086 ,
         \29087 , \29088 , \29089 , \29090 , \29091 , \29092 , \29093 , \29094 , \29095 , \29096 ,
         \29097 , \29098 , \29099 , \29100 , \29101 , \29102 , \29103 , \29104 , \29105 , \29106 ,
         \29107 , \29108 , \29109 , \29110 , \29111 , \29112 , \29113 , \29114 , \29115 , \29116 ,
         \29117 , \29118 , \29119 , \29120 , \29121 , \29122 , \29123 , \29124 , \29125 , \29126 ,
         \29127 , \29128 , \29129 , \29130 , \29131 , \29132 , \29133 , \29134 , \29135 , \29136 ,
         \29137 , \29138 , \29139 , \29140 , \29141 , \29142 , \29143 , \29144 , \29145 , \29146 ,
         \29147 , \29148 , \29149 , \29150 , \29151 , \29152 , \29153 , \29154 , \29155 , \29156 ,
         \29157 , \29158 , \29159 , \29160 , \29161 , \29162 , \29163 , \29164 , \29165 , \29166 ,
         \29167 , \29168 , \29169 , \29170 , \29171 , \29172 , \29173 , \29174 , \29175 , \29176 ,
         \29177 , \29178 , \29179_nG9bbd , \29180 , \29181 , \29182 , \29183 , \29184 , \29185 , \29186 ,
         \29187 , \29188 , \29189 , \29190 , \29191 , \29192 , \29193 , \29194 , \29195 , \29196 ,
         \29197 , \29198 , \29199 , \29200 , \29201 , \29202 , \29203 , \29204 , \29205 , \29206 ,
         \29207 , \29208 , \29209 , \29210 , \29211 , \29212 , \29213 , \29214 , \29215 , \29216 ,
         \29217 , \29218 , \29219 , \29220 , \29221 , \29222 , \29223 , \29224 , \29225 , \29226 ,
         \29227 , \29228 , \29229 , \29230 , \29231 , \29232 , \29233 , \29234 , \29235 , \29236 ,
         \29237 , \29238 , \29239 , \29240 , \29241 , \29242 , \29243 , \29244 , \29245 , \29246 ,
         \29247 , \29248 , \29249 , \29250 , \29251 , \29252 , \29253 , \29254 , \29255 , \29256 ,
         \29257 , \29258 , \29259 , \29260 , \29261 , \29262 , \29263 , \29264 , \29265 , \29266 ,
         \29267 , \29268 , \29269 , \29270 , \29271 , \29272 , \29273 , \29274 , \29275 , \29276 ,
         \29277 , \29278 , \29279 , \29280 , \29281 , \29282 , \29283 , \29284 , \29285 , \29286 ,
         \29287 , \29288 , \29289 , \29290 , \29291 , \29292 , \29293 , \29294 , \29295 , \29296 ,
         \29297 , \29298 , \29299 , \29300 , \29301 , \29302 , \29303 , \29304 , \29305 , \29306 ,
         \29307 , \29308 , \29309 , \29310 , \29311 , \29312 , \29313 , \29314 , \29315 , \29316 ,
         \29317 , \29318 , \29319 , \29320 , \29321 , \29322 , \29323 , \29324 , \29325 , \29326 ,
         \29327 , \29328 , \29329 , \29330 , \29331 , \29332 , \29333 , \29334 , \29335 , \29336 ,
         \29337 , \29338 , \29339 , \29340 , \29341 , \29342 , \29343 , \29344 , \29345 , \29346 ,
         \29347 , \29348 , \29349 , \29350 , \29351 , \29352 , \29353 , \29354 , \29355 , \29356 ,
         \29357 , \29358 , \29359 , \29360 , \29361 , \29362 , \29363 , \29364 , \29365 , \29366 ,
         \29367 , \29368 , \29369 , \29370 , \29371 , \29372 , \29373 , \29374 , \29375 , \29376 ,
         \29377 , \29378 , \29379 , \29380 , \29381 , \29382 , \29383 , \29384 , \29385 , \29386 ,
         \29387 , \29388 , \29389 , \29390 , \29391 , \29392 , \29393 , \29394 , \29395 , \29396 ,
         \29397 , \29398 , \29399 , \29400 , \29401 , \29402 , \29403 , \29404 , \29405 , \29406 ,
         \29407 , \29408 , \29409 , \29410 , \29411 , \29412 , \29413 , \29414 , \29415 , \29416 ,
         \29417 , \29418 , \29419 , \29420 , \29421 , \29422 , \29423 , \29424 , \29425 , \29426 ,
         \29427 , \29428 , \29429 , \29430 , \29431 , \29432 , \29433_nG233f , \29434 , \29435 , \29436 ,
         \29437 , \29438 , \29439 , \29440 , \29441 , \29442 , \29443 , \29444 , \29445 , \29446 ,
         \29447 , \29448 , \29449 , \29450 , \29451 , \29452 , \29453 , \29454 , \29455 , \29456 ,
         \29457 , \29458 , \29459 , \29460 , \29461 , \29462 , \29463 , \29464 , \29465 , \29466 ,
         \29467 , \29468 , \29469 , \29470 , \29471 , \29472 , \29473 , \29474 , \29475 , \29476 ,
         \29477 , \29478 , \29479 , \29480 , \29481 , \29482 , \29483 , \29484 , \29485 , \29486 ,
         \29487 , \29488 , \29489 , \29490 , \29491 , \29492 , \29493 , \29494 , \29495 , \29496 ,
         \29497 , \29498 , \29499 , \29500 , \29501 , \29502 , \29503 , \29504 , \29505 , \29506 ,
         \29507 , \29508 , \29509 , \29510 , \29511 , \29512 , \29513 , \29514 , \29515 , \29516 ,
         \29517 , \29518 , \29519 , \29520 , \29521 , \29522 , \29523 , \29524 , \29525 , \29526 ,
         \29527 , \29528 , \29529 , \29530 , \29531 , \29532 , \29533 , \29534 , \29535 , \29536 ,
         \29537 , \29538 , \29539 , \29540 , \29541 , \29542 , \29543 , \29544 , \29545 , \29546 ,
         \29547 , \29548 , \29549 , \29550 , \29551 , \29552 , \29553 , \29554 , \29555 , \29556 ,
         \29557 , \29558 , \29559 , \29560 , \29561 , \29562 , \29563 , \29564 , \29565 , \29566_nG346c ,
         \29567 , \29568 , \29569 , \29570 , \29571 , \29572 , \29573 , \29574 , \29575 , \29576 ,
         \29577 , \29578 , \29579 , \29580 , \29581 , \29582 , \29583 , \29584 , \29585 , \29586 ,
         \29587 , \29588 , \29589 , \29590 , \29591 , \29592 , \29593 , \29594 , \29595 , \29596 ,
         \29597 , \29598 , \29599 , \29600 , \29601 , \29602 , \29603 , \29604 , \29605 , \29606 ,
         \29607 , \29608 , \29609 , \29610 , \29611 , \29612 , \29613 , \29614 , \29615 , \29616 ,
         \29617 , \29618 , \29619 , \29620 , \29621 , \29622 , \29623 , \29624 , \29625 , \29626 ,
         \29627 , \29628 , \29629 , \29630 , \29631 , \29632 , \29633 , \29634 , \29635 , \29636 ,
         \29637 , \29638 , \29639 , \29640 , \29641 , \29642 , \29643 , \29644 , \29645 , \29646 ,
         \29647 , \29648 , \29649 , \29650 , \29651 , \29652 , \29653 , \29654 , \29655 , \29656 ,
         \29657 , \29658 , \29659 , \29660 , \29661 , \29662 , \29663 , \29664 , \29665 , \29666 ,
         \29667 , \29668 , \29669 , \29670 , \29671 , \29672 , \29673 , \29674 , \29675 , \29676 ,
         \29677 , \29678 , \29679 , \29680 , \29681 , \29682 , \29683 , \29684 , \29685 , \29686 ,
         \29687 , \29688 , \29689 , \29690 , \29691 , \29692 , \29693 , \29694 , \29695 , \29696 ,
         \29697 , \29698 , \29699 , \29700_nG23c4 , \29701 , \29702 , \29703 , \29704 , \29705 , \29706 ,
         \29707 , \29708 , \29709 , \29710 , \29711 , \29712 , \29713 , \29714 , \29715 , \29716 ,
         \29717 , \29718 , \29719 , \29720 , \29721 , \29722 , \29723 , \29724 , \29725 , \29726 ,
         \29727 , \29728 , \29729 , \29730 , \29731 , \29732 , \29733 , \29734 , \29735 , \29736 ,
         \29737 , \29738 , \29739 , \29740 , \29741 , \29742 , \29743 , \29744 , \29745 , \29746 ,
         \29747 , \29748 , \29749 , \29750 , \29751 , \29752 , \29753 , \29754 , \29755 , \29756 ,
         \29757 , \29758 , \29759 , \29760 , \29761 , \29762 , \29763 , \29764 , \29765 , \29766 ,
         \29767 , \29768 , \29769 , \29770 , \29771 , \29772 , \29773 , \29774 , \29775 , \29776 ,
         \29777 , \29778 , \29779 , \29780 , \29781 , \29782 , \29783 , \29784 , \29785 , \29786 ,
         \29787 , \29788 , \29789 , \29790 , \29791 , \29792 , \29793 , \29794 , \29795 , \29796 ,
         \29797 , \29798 , \29799 , \29800 , \29801 , \29802 , \29803 , \29804 , \29805 , \29806 ,
         \29807 , \29808 , \29809 , \29810 , \29811 , \29812 , \29813 , \29814 , \29815 , \29816 ,
         \29817 , \29818 , \29819 , \29820 , \29821 , \29822 , \29823 , \29824 , \29825 , \29826 ,
         \29827 , \29828 , \29829 , \29830 , \29831 , \29832 , \29833_nG34f1 , \29834 , \29835 , \29836 ,
         \29837 , \29838 , \29839 , \29840 , \29841 , \29842 , \29843 , \29844_nG4400 , \29845 , \29846 ,
         \29847_nG4403 , \29848 , \29849 , \29850 , \29851 , \29852 , \29853 , \29854 , \29855 , \29856 ,
         \29857 , \29858 , \29859 , \29860 , \29861 , \29862 , \29863 , \29864 , \29865 , \29866 ,
         \29867 , \29868 , \29869 , \29870 , \29871 , \29872 , \29873 , \29874 , \29875 , \29876 ,
         \29877 , \29878 , \29879 , \29880 , \29881 , \29882 , \29883 , \29884 , \29885 , \29886 ,
         \29887 , \29888 , \29889 , \29890 , \29891 , \29892 , \29893 , \29894 , \29895 , \29896 ,
         \29897 , \29898 , \29899 , \29900 , \29901 , \29902 , \29903 , \29904 , \29905 , \29906 ,
         \29907 , \29908 , \29909 , \29910 , \29911 , \29912 , \29913 , \29914 , \29915 , \29916 ,
         \29917 , \29918 , \29919 , \29920 , \29921 , \29922 , \29923 , \29924 , \29925 , \29926 ,
         \29927 , \29928 , \29929 , \29930 , \29931 , \29932 , \29933 , \29934 , \29935 , \29936 ,
         \29937 , \29938 , \29939 , \29940 , \29941 , \29942 , \29943 , \29944 , \29945 , \29946 ,
         \29947 , \29948 , \29949 , \29950 , \29951 , \29952 , \29953 , \29954 , \29955 , \29956 ,
         \29957 , \29958 , \29959 , \29960 , \29961 , \29962 , \29963 , \29964 , \29965 , \29966 ,
         \29967 , \29968 , \29969 , \29970 , \29971 , \29972 , \29973 , \29974 , \29975 , \29976 ,
         \29977 , \29978 , \29979 , \29980 , \29981 , \29982 , \29983 , \29984 , \29985 , \29986 ,
         \29987 , \29988 , \29989 , \29990 , \29991 , \29992 , \29993 , \29994 , \29995 , \29996 ,
         \29997 , \29998 , \29999 , \30000 , \30001 , \30002 , \30003 , \30004 , \30005 , \30006 ,
         \30007 , \30008 , \30009 , \30010 , \30011 , \30012 , \30013 , \30014 , \30015 , \30016 ,
         \30017 , \30018 , \30019 , \30020 , \30021 , \30022 , \30023 , \30024 , \30025 , \30026 ,
         \30027 , \30028 , \30029 , \30030 , \30031 , \30032 , \30033 , \30034 , \30035 , \30036 ,
         \30037 , \30038 , \30039 , \30040 , \30041 , \30042 , \30043 , \30044 , \30045 , \30046 ,
         \30047 , \30048 , \30049 , \30050 , \30051 , \30052 , \30053 , \30054 , \30055 , \30056 ,
         \30057 , \30058 , \30059 , \30060 , \30061 , \30062 , \30063 , \30064 , \30065 , \30066 ,
         \30067 , \30068 , \30069 , \30070 , \30071 , \30072 , \30073 , \30074 , \30075 , \30076 ,
         \30077 , \30078 , \30079 , \30080 , \30081 , \30082 , \30083 , \30084 , \30085 , \30086 ,
         \30087 , \30088 , \30089 , \30090 , \30091 , \30092 , \30093 , \30094 , \30095 , \30096 ,
         \30097 , \30098 , \30099 , \30100 , \30101 , \30102 , \30103 , \30104 , \30105 , \30106 ,
         \30107 , \30108 , \30109 , \30110 , \30111_nG61d6 , \30112 , \30113 , \30114 , \30115 , \30116 ,
         \30117 , \30118 , \30119 , \30120 , \30121 , \30122 , \30123 , \30124 , \30125 , \30126 ,
         \30127 , \30128 , \30129 , \30130 , \30131 , \30132 , \30133 , \30134 , \30135 , \30136 ,
         \30137 , \30138 , \30139 , \30140 , \30141 , \30142 , \30143 , \30144 , \30145 , \30146 ,
         \30147 , \30148 , \30149 , \30150 , \30151 , \30152 , \30153 , \30154 , \30155 , \30156 ,
         \30157 , \30158 , \30159 , \30160 , \30161 , \30162 , \30163 , \30164 , \30165 , \30166 ,
         \30167 , \30168 , \30169 , \30170 , \30171 , \30172 , \30173 , \30174 , \30175 , \30176 ,
         \30177 , \30178 , \30179 , \30180 , \30181 , \30182 , \30183 , \30184 , \30185 , \30186 ,
         \30187 , \30188 , \30189 , \30190 , \30191 , \30192 , \30193 , \30194 , \30195 , \30196 ,
         \30197 , \30198 , \30199 , \30200 , \30201 , \30202 , \30203 , \30204 , \30205 , \30206 ,
         \30207 , \30208 , \30209 , \30210 , \30211 , \30212 , \30213 , \30214 , \30215 , \30216 ,
         \30217 , \30218 , \30219 , \30220 , \30221 , \30222 , \30223 , \30224 , \30225 , \30226 ,
         \30227 , \30228 , \30229 , \30230 , \30231 , \30232 , \30233 , \30234 , \30235 , \30236 ,
         \30237 , \30238 , \30239 , \30240 , \30241 , \30242 , \30243_nG625a , \30244_nG625b , \30245 , \30246 ,
         \30247 , \30248 , \30249 , \30250 , \30251 , \30252 , \30253 , \30254 , \30255 , \30256 ,
         \30257 , \30258 , \30259 , \30260 , \30261 , \30262 , \30263 , \30264 , \30265_nG65cb , \30266_nG65cc ,
         \30267_nG65cd , \30268 , \30269 , \30270 , \30271 , \30272 , \30273 , \30274 , \30275 , \30276 ,
         \30277 , \30278 , \30279 , \30280 , \30281 , \30282 , \30283 , \30284 , \30285 , \30286 ,
         \30287 , \30288 , \30289 , \30290 , \30291 , \30292 , \30293 , \30294 , \30295 , \30296 ,
         \30297 , \30298 , \30299 , \30300 , \30301 , \30302 , \30303 , \30304 , \30305 , \30306 ,
         \30307 , \30308 , \30309 , \30310 , \30311 , \30312 , \30313 , \30314 , \30315 , \30316 ,
         \30317 , \30318 , \30319 , \30320 , \30321 , \30322 , \30323 , \30324 , \30325 , \30326 ,
         \30327 , \30328 , \30329 , \30330 , \30331 , \30332 , \30333 , \30334 , \30335 , \30336 ,
         \30337 , \30338 , \30339 , \30340 , \30341 , \30342 , \30343 , \30344 , \30345 , \30346 ,
         \30347 , \30348 , \30349 , \30350 , \30351 , \30352 , \30353 , \30354 , \30355 , \30356 ,
         \30357 , \30358 , \30359 , \30360 , \30361 , \30362 , \30363 , \30364 , \30365 , \30366_nG9bba ,
         \30367 , \30368 , \30369 , \30370 , \30371 , \30372 , \30373 , \30374 , \30375 , \30376 ,
         \30377 , \30378 , \30379 , \30380 , \30381 , \30382 , \30383 , \30384 , \30385 , \30386 ,
         \30387 , \30388 , \30389 , \30390 , \30391 , \30392 , \30393 , \30394 , \30395 , \30396 ,
         \30397 , \30398 , \30399 , \30400 , \30401 , \30402 , \30403 , \30404 , \30405 , \30406 ,
         \30407 , \30408 , \30409 , \30410 , \30411 , \30412 , \30413 , \30414 , \30415 , \30416 ,
         \30417 , \30418 , \30419 , \30420 , \30421 , \30422 , \30423 , \30424 , \30425 , \30426 ,
         \30427 , \30428 , \30429 , \30430 , \30431 , \30432 , \30433 , \30434 , \30435 , \30436 ,
         \30437 , \30438 , \30439 , \30440 , \30441 , \30442 , \30443 , \30444 , \30445 , \30446 ,
         \30447 , \30448 , \30449 , \30450 , \30451 , \30452 , \30453 , \30454 , \30455 , \30456 ,
         \30457 , \30458 , \30459 , \30460 , \30461 , \30462 , \30463 , \30464 , \30465 , \30466 ,
         \30467 , \30468 , \30469 , \30470 , \30471 , \30472 , \30473 , \30474 , \30475 , \30476 ,
         \30477 , \30478 , \30479 , \30480 , \30481 , \30482 , \30483 , \30484 , \30485 , \30486 ,
         \30487 , \30488 , \30489 , \30490 , \30491 , \30492 , \30493 , \30494 , \30495 , \30496 ,
         \30497 , \30498 , \30499 , \30500 , \30501 , \30502 , \30503 , \30504 , \30505 , \30506 ,
         \30507 , \30508 , \30509 , \30510 , \30511 , \30512 , \30513 , \30514 , \30515 , \30516 ,
         \30517 , \30518 , \30519 , \30520 , \30521 , \30522 , \30523 , \30524 , \30525 , \30526 ,
         \30527 , \30528 , \30529 , \30530 , \30531 , \30532 , \30533 , \30534 , \30535 , \30536 ,
         \30537 , \30538 , \30539 , \30540 , \30541 , \30542 , \30543 , \30544 , \30545 , \30546 ,
         \30547 , \30548 , \30549 , \30550 , \30551 , \30552 , \30553 , \30554 , \30555 , \30556 ,
         \30557 , \30558 , \30559 , \30560 , \30561 , \30562 , \30563 , \30564 , \30565 , \30566 ,
         \30567 , \30568 , \30569 , \30570 , \30571 , \30572 , \30573 , \30574 , \30575 , \30576 ,
         \30577 , \30578 , \30579 , \30580 , \30581 , \30582 , \30583 , \30584 , \30585 , \30586 ,
         \30587 , \30588 , \30589 , \30590 , \30591 , \30592 , \30593 , \30594 , \30595 , \30596 ,
         \30597 , \30598 , \30599 , \30600 , \30601 , \30602 , \30603 , \30604 , \30605 , \30606 ,
         \30607 , \30608 , \30609 , \30610 , \30611 , \30612 , \30613 , \30614 , \30615 , \30616 ,
         \30617 , \30618 , \30619 , \30620 , \30621 , \30622 , \30623 , \30624 , \30625 , \30626 ,
         \30627 , \30628 , \30629 , \30630 , \30631 , \30632 , \30633 , \30634 , \30635 , \30636 ,
         \30637 , \30638 , \30639 , \30640 , \30641 , \30642 , \30643 , \30644 , \30645 , \30646 ,
         \30647 , \30648 , \30649 , \30650 , \30651 , \30652 , \30653 , \30654 , \30655 , \30656 ,
         \30657 , \30658 , \30659 , \30660 , \30661 , \30662 , \30663 , \30664 , \30665 , \30666 ,
         \30667 , \30668_nG65ce , \30669 , \30670 , \30671 , \30672 , \30673 , \30674 , \30675 , \30676 ,
         \30677 , \30678 , \30679 , \30680 , \30681 , \30682 , \30683 , \30684 , \30685 , \30686 ,
         \30687 , \30688 , \30689 , \30690 , \30691 , \30692 , \30693 , \30694 , \30695 , \30696 ,
         \30697 , \30698 , \30699 , \30700 , \30701 , \30702 , \30703 , \30704 , \30705 , \30706 ,
         \30707 , \30708 , \30709 , \30710 , \30711 , \30712 , \30713 , \30714 , \30715 , \30716 ,
         \30717 , \30718 , \30719 , \30720 , \30721 , \30722 , \30723 , \30724 , \30725 , \30726 ,
         \30727 , \30728 , \30729 , \30730 , \30731 , \30732 , \30733 , \30734 , \30735 , \30736 ,
         \30737 , \30738 , \30739 , \30740 , \30741 , \30742 , \30743 , \30744 , \30745 , \30746 ,
         \30747 , \30748 , \30749 , \30750 , \30751 , \30752 , \30753 , \30754 , \30755 , \30756 ,
         \30757 , \30758 , \30759 , \30760 , \30761 , \30762 , \30763 , \30764 , \30765 , \30766 ,
         \30767 , \30768 , \30769 , \30770 , \30771 , \30772 , \30773 , \30774 , \30775 , \30776 ,
         \30777 , \30778 , \30779 , \30780 , \30781 , \30782 , \30783 , \30784 , \30785 , \30786 ,
         \30787 , \30788 , \30789 , \30790 , \30791 , \30792 , \30793 , \30794 , \30795 , \30796 ,
         \30797 , \30798 , \30799 , \30800_nG65cf , \30801_nG65d0 , \30802 , \30803 , \30804 , \30805 , \30806 ,
         \30807_nG62df , \30808_nG6363 , \30809_nG6364 , \30810 , \30811 , \30812 , \30813 , \30814 , \30815 , \30816 ,
         \30817 , \30818 , \30819 , \30820 , \30821 , \30822 , \30823 , \30824 , \30825 , \30826 ,
         \30827 , \30828 , \30829 , \30830 , \30831 , \30832 , \30833 , \30834 , \30835 , \30836 ,
         \30837 , \30838 , \30839 , \30840 , \30841 , \30842 , \30843 , \30844 , \30845 , \30846 ,
         \30847 , \30848 , \30849 , \30850 , \30851 , \30852 , \30853 , \30854 , \30855 , \30856 ,
         \30857 , \30858 , \30859 , \30860 , \30861 , \30862 , \30863 , \30864 , \30865 , \30866 ,
         \30867 , \30868 , \30869 , \30870 , \30871 , \30872 , \30873 , \30874 , \30875 , \30876 ,
         \30877 , \30878 , \30879 , \30880 , \30881 , \30882 , \30883 , \30884 , \30885 , \30886 ,
         \30887 , \30888 , \30889 , \30890 , \30891 , \30892 , \30893 , \30894 , \30895 , \30896 ,
         \30897 , \30898 , \30899 , \30900 , \30901 , \30902 , \30903 , \30904 , \30905 , \30906 ,
         \30907 , \30908 , \30909 , \30910 , \30911 , \30912 , \30913 , \30914 , \30915 , \30916 ,
         \30917 , \30918 , \30919 , \30920 , \30921 , \30922 , \30923 , \30924 , \30925 , \30926 ,
         \30927 , \30928 , \30929 , \30930 , \30931 , \30932 , \30933 , \30934 , \30935 , \30936 ,
         \30937 , \30938 , \30939 , \30940_nG9bb7 , \30941 , \30942 , \30943 , \30944 , \30945 , \30946 ,
         \30947 , \30948 , \30949 , \30950 , \30951 , \30952 , \30953 , \30954 , \30955 , \30956 ,
         \30957 , \30958 , \30959 , \30960 , \30961 , \30962 , \30963 , \30964 , \30965 , \30966 ,
         \30967 , \30968 , \30969 , \30970 , \30971 , \30972 , \30973 , \30974 , \30975 , \30976 ,
         \30977 , \30978 , \30979 , \30980 , \30981 , \30982 , \30983 , \30984 , \30985 , \30986 ,
         \30987 , \30988 , \30989 , \30990 , \30991 , \30992 , \30993 , \30994 , \30995 , \30996 ,
         \30997 , \30998 , \30999 , \31000 , \31001 , \31002 , \31003 , \31004 , \31005 , \31006 ,
         \31007 , \31008 , \31009 , \31010 , \31011 , \31012 , \31013 , \31014 , \31015 , \31016 ,
         \31017 , \31018 , \31019 , \31020 , \31021 , \31022 , \31023 , \31024 , \31025 , \31026 ,
         \31027 , \31028 , \31029 , \31030 , \31031 , \31032 , \31033 , \31034 , \31035 , \31036 ,
         \31037 , \31038 , \31039 , \31040 , \31041 , \31042 , \31043 , \31044 , \31045 , \31046 ,
         \31047 , \31048 , \31049 , \31050 , \31051 , \31052 , \31053 , \31054 , \31055 , \31056 ,
         \31057 , \31058 , \31059 , \31060 , \31061 , \31062 , \31063 , \31064 , \31065 , \31066 ,
         \31067 , \31068 , \31069 , \31070 , \31071 , \31072 , \31073 , \31074 , \31075 , \31076 ,
         \31077 , \31078 , \31079 , \31080 , \31081 , \31082 , \31083 , \31084 , \31085 , \31086 ,
         \31087 , \31088 , \31089 , \31090 , \31091 , \31092 , \31093 , \31094 , \31095 , \31096 ,
         \31097 , \31098 , \31099 , \31100 , \31101 , \31102 , \31103 , \31104 , \31105 , \31106 ,
         \31107 , \31108 , \31109 , \31110 , \31111 , \31112 , \31113 , \31114 , \31115 , \31116 ,
         \31117 , \31118 , \31119 , \31120 , \31121 , \31122 , \31123 , \31124 , \31125 , \31126 ,
         \31127 , \31128 , \31129 , \31130 , \31131 , \31132 , \31133 , \31134 , \31135 , \31136 ,
         \31137 , \31138 , \31139 , \31140 , \31141 , \31142 , \31143 , \31144 , \31145 , \31146 ,
         \31147 , \31148 , \31149 , \31150 , \31151 , \31152 , \31153 , \31154 , \31155 , \31156 ,
         \31157 , \31158 , \31159 , \31160 , \31161 , \31162 , \31163 , \31164 , \31165 , \31166 ,
         \31167 , \31168 , \31169 , \31170 , \31171 , \31172 , \31173 , \31174 , \31175 , \31176 ,
         \31177 , \31178 , \31179 , \31180 , \31181 , \31182 , \31183 , \31184 , \31185 , \31186 ,
         \31187 , \31188 , \31189 , \31190 , \31191 , \31192 , \31193 , \31194 , \31195 , \31196 ,
         \31197 , \31198 , \31199 , \31200 , \31201 , \31202 , \31203 , \31204 , \31205 , \31206 ,
         \31207 , \31208 , \31209 , \31210 , \31211 , \31212 , \31213 , \31214 , \31215 , \31216_nG2235 ,
         \31217 , \31218 , \31219 , \31220 , \31221 , \31222 , \31223 , \31224 , \31225 , \31226 ,
         \31227 , \31228 , \31229 , \31230 , \31231 , \31232 , \31233 , \31234 , \31235 , \31236 ,
         \31237 , \31238 , \31239 , \31240 , \31241 , \31242 , \31243 , \31244 , \31245 , \31246 ,
         \31247 , \31248 , \31249 , \31250 , \31251 , \31252 , \31253 , \31254 , \31255 , \31256 ,
         \31257 , \31258 , \31259 , \31260 , \31261 , \31262 , \31263 , \31264 , \31265 , \31266 ,
         \31267 , \31268 , \31269 , \31270 , \31271 , \31272 , \31273 , \31274 , \31275 , \31276 ,
         \31277 , \31278 , \31279 , \31280 , \31281 , \31282 , \31283 , \31284 , \31285 , \31286 ,
         \31287 , \31288 , \31289 , \31290 , \31291 , \31292 , \31293 , \31294 , \31295 , \31296 ,
         \31297 , \31298 , \31299 , \31300 , \31301 , \31302 , \31303 , \31304 , \31305 , \31306 ,
         \31307 , \31308 , \31309 , \31310 , \31311 , \31312 , \31313 , \31314 , \31315 , \31316 ,
         \31317 , \31318 , \31319 , \31320 , \31321 , \31322 , \31323 , \31324 , \31325 , \31326 ,
         \31327 , \31328 , \31329 , \31330 , \31331 , \31332 , \31333 , \31334 , \31335 , \31336 ,
         \31337 , \31338 , \31339 , \31340 , \31341 , \31342 , \31343 , \31344 , \31345 , \31346 ,
         \31347 , \31348 , \31349_nG3362 , \31350 , \31351 , \31352 , \31353 , \31354 , \31355 , \31356 ,
         \31357 , \31358 , \31359 , \31360 , \31361 , \31362 , \31363 , \31364 , \31365 , \31366 ,
         \31367 , \31368 , \31369 , \31370 , \31371 , \31372 , \31373 , \31374 , \31375 , \31376 ,
         \31377 , \31378 , \31379 , \31380 , \31381 , \31382 , \31383 , \31384 , \31385 , \31386 ,
         \31387 , \31388 , \31389 , \31390 , \31391 , \31392 , \31393 , \31394 , \31395 , \31396 ,
         \31397 , \31398 , \31399 , \31400 , \31401 , \31402 , \31403 , \31404 , \31405 , \31406 ,
         \31407 , \31408 , \31409 , \31410 , \31411 , \31412 , \31413 , \31414 , \31415 , \31416 ,
         \31417 , \31418 , \31419 , \31420 , \31421 , \31422 , \31423 , \31424 , \31425 , \31426 ,
         \31427 , \31428 , \31429 , \31430 , \31431 , \31432 , \31433 , \31434 , \31435 , \31436 ,
         \31437 , \31438 , \31439 , \31440 , \31441 , \31442 , \31443 , \31444 , \31445 , \31446 ,
         \31447 , \31448 , \31449 , \31450 , \31451 , \31452 , \31453 , \31454 , \31455 , \31456 ,
         \31457 , \31458 , \31459 , \31460 , \31461 , \31462 , \31463 , \31464 , \31465 , \31466 ,
         \31467 , \31468 , \31469 , \31470 , \31471 , \31472 , \31473 , \31474 , \31475 , \31476 ,
         \31477 , \31478 , \31479 , \31480 , \31481 , \31482 , \31483_nG22ba , \31484 , \31485 , \31486 ,
         \31487 , \31488 , \31489 , \31490 , \31491 , \31492 , \31493 , \31494 , \31495 , \31496 ,
         \31497 , \31498 , \31499 , \31500 , \31501 , \31502 , \31503 , \31504 , \31505 , \31506 ,
         \31507 , \31508 , \31509 , \31510 , \31511 , \31512 , \31513 , \31514 , \31515 , \31516 ,
         \31517 , \31518 , \31519 , \31520 , \31521 , \31522 , \31523 , \31524 , \31525 , \31526 ,
         \31527 , \31528 , \31529 , \31530 , \31531 , \31532 , \31533 , \31534 , \31535 , \31536 ,
         \31537 , \31538 , \31539 , \31540 , \31541 , \31542 , \31543 , \31544 , \31545 , \31546 ,
         \31547 , \31548 , \31549 , \31550 , \31551 , \31552 , \31553 , \31554 , \31555 , \31556 ,
         \31557 , \31558 , \31559 , \31560 , \31561 , \31562 , \31563 , \31564 , \31565 , \31566 ,
         \31567 , \31568 , \31569 , \31570 , \31571 , \31572 , \31573 , \31574 , \31575 , \31576 ,
         \31577 , \31578 , \31579 , \31580 , \31581 , \31582 , \31583 , \31584 , \31585 , \31586 ,
         \31587 , \31588 , \31589 , \31590 , \31591 , \31592 , \31593 , \31594 , \31595 , \31596 ,
         \31597 , \31598 , \31599 , \31600 , \31601 , \31602 , \31603 , \31604 , \31605 , \31606 ,
         \31607 , \31608 , \31609 , \31610 , \31611 , \31612 , \31613 , \31614 , \31615 , \31616_nG33e7 ,
         \31617 , \31618 , \31619 , \31620 , \31621 , \31622 , \31623 , \31624 , \31625 , \31626 ,
         \31627_nG43fa , \31628 , \31629 , \31630_nG43fd , \31631 , \31632 , \31633 , \31634 , \31635 , \31636 ,
         \31637 , \31638 , \31639 , \31640 , \31641 , \31642 , \31643 , \31644 , \31645 , \31646 ,
         \31647 , \31648 , \31649 , \31650 , \31651 , \31652 , \31653 , \31654 , \31655 , \31656 ,
         \31657 , \31658 , \31659 , \31660 , \31661 , \31662 , \31663 , \31664 , \31665 , \31666 ,
         \31667 , \31668 , \31669 , \31670 , \31671 , \31672 , \31673 , \31674 , \31675 , \31676 ,
         \31677 , \31678 , \31679 , \31680 , \31681 , \31682 , \31683 , \31684 , \31685 , \31686 ,
         \31687 , \31688 , \31689 , \31690 , \31691 , \31692 , \31693 , \31694 , \31695 , \31696 ,
         \31697 , \31698 , \31699 , \31700 , \31701 , \31702 , \31703 , \31704 , \31705 , \31706 ,
         \31707 , \31708 , \31709 , \31710 , \31711 , \31712 , \31713 , \31714 , \31715 , \31716 ,
         \31717 , \31718 , \31719 , \31720 , \31721 , \31722 , \31723 , \31724 , \31725 , \31726 ,
         \31727 , \31728 , \31729 , \31730 , \31731 , \31732 , \31733 , \31734 , \31735 , \31736 ,
         \31737 , \31738 , \31739 , \31740 , \31741 , \31742 , \31743 , \31744 , \31745 , \31746 ,
         \31747 , \31748 , \31749 , \31750 , \31751 , \31752 , \31753 , \31754 , \31755 , \31756 ,
         \31757 , \31758 , \31759 , \31760 , \31761 , \31762 , \31763 , \31764 , \31765 , \31766 ,
         \31767 , \31768 , \31769 , \31770 , \31771 , \31772 , \31773 , \31774 , \31775 , \31776 ,
         \31777 , \31778 , \31779 , \31780 , \31781 , \31782 , \31783 , \31784 , \31785 , \31786 ,
         \31787 , \31788 , \31789 , \31790 , \31791 , \31792 , \31793 , \31794 , \31795 , \31796 ,
         \31797 , \31798 , \31799 , \31800 , \31801 , \31802 , \31803 , \31804 , \31805 , \31806 ,
         \31807 , \31808 , \31809 , \31810 , \31811 , \31812 , \31813 , \31814 , \31815 , \31816 ,
         \31817 , \31818 , \31819 , \31820 , \31821 , \31822 , \31823 , \31824 , \31825 , \31826 ,
         \31827 , \31828 , \31829 , \31830 , \31831 , \31832 , \31833 , \31834 , \31835 , \31836 ,
         \31837 , \31838 , \31839 , \31840 , \31841 , \31842 , \31843 , \31844 , \31845 , \31846 ,
         \31847 , \31848 , \31849 , \31850 , \31851 , \31852 , \31853 , \31854 , \31855 , \31856 ,
         \31857 , \31858 , \31859 , \31860 , \31861 , \31862 , \31863 , \31864 , \31865 , \31866 ,
         \31867 , \31868 , \31869 , \31870 , \31871 , \31872 , \31873 , \31874 , \31875 , \31876 ,
         \31877 , \31878 , \31879 , \31880 , \31881 , \31882 , \31883 , \31884 , \31885 , \31886 ,
         \31887 , \31888 , \31889 , \31890 , \31891 , \31892 , \31893 , \31894 , \31895 , \31896 ,
         \31897 , \31898 , \31899 , \31900 , \31901 , \31902 , \31903 , \31904 , \31905 , \31906 ,
         \31907 , \31908 , \31909 , \31910 , \31911 , \31912 , \31913 , \31914 , \31915 , \31916 ,
         \31917 , \31918 , \31919 , \31920_nG65d1 , \31921 , \31922 , \31923 , \31924 , \31925 , \31926 ,
         \31927 , \31928 , \31929 , \31930 , \31931 , \31932 , \31933 , \31934 , \31935 , \31936 ,
         \31937 , \31938 , \31939 , \31940 , \31941 , \31942 , \31943 , \31944 , \31945 , \31946 ,
         \31947 , \31948 , \31949 , \31950 , \31951 , \31952 , \31953 , \31954 , \31955 , \31956 ,
         \31957 , \31958 , \31959 , \31960 , \31961 , \31962 , \31963 , \31964 , \31965 , \31966 ,
         \31967 , \31968 , \31969 , \31970 , \31971 , \31972 , \31973 , \31974 , \31975 , \31976 ,
         \31977 , \31978 , \31979 , \31980 , \31981 , \31982 , \31983 , \31984 , \31985 , \31986 ,
         \31987 , \31988 , \31989 , \31990 , \31991 , \31992 , \31993 , \31994 , \31995 , \31996 ,
         \31997 , \31998 , \31999 , \32000 , \32001 , \32002 , \32003 , \32004 , \32005 , \32006 ,
         \32007 , \32008 , \32009 , \32010 , \32011 , \32012 , \32013 , \32014 , \32015 , \32016 ,
         \32017 , \32018 , \32019 , \32020 , \32021 , \32022 , \32023 , \32024 , \32025 , \32026 ,
         \32027 , \32028 , \32029 , \32030 , \32031 , \32032 , \32033 , \32034 , \32035 , \32036 ,
         \32037 , \32038 , \32039 , \32040 , \32041 , \32042 , \32043 , \32044 , \32045 , \32046 ,
         \32047 , \32048 , \32049 , \32050 , \32051 , \32052_nG65d2 , \32053_nG65d3 , \32054 , \32055 , \32056 ,
         \32057 , \32058 , \32059 , \32060 , \32061 , \32062 , \32063_nG63e8 , \32064_nG646c , \32065_nG646d , \32066 ,
         \32067 , \32068 , \32069 , \32070 , \32071 , \32072 , \32073 , \32074 , \32075 , \32076 ,
         \32077 , \32078 , \32079 , \32080 , \32081 , \32082 , \32083 , \32084 , \32085 , \32086 ,
         \32087 , \32088 , \32089 , \32090 , \32091 , \32092 , \32093 , \32094 , \32095 , \32096 ,
         \32097 , \32098 , \32099 , \32100 , \32101 , \32102 , \32103 , \32104 , \32105 , \32106 ,
         \32107 , \32108 , \32109 , \32110 , \32111 , \32112 , \32113 , \32114 , \32115 , \32116 ,
         \32117 , \32118 , \32119 , \32120 , \32121 , \32122 , \32123 , \32124 , \32125 , \32126 ,
         \32127 , \32128 , \32129 , \32130 , \32131 , \32132 , \32133 , \32134 , \32135 , \32136 ,
         \32137 , \32138 , \32139 , \32140 , \32141 , \32142 , \32143 , \32144 , \32145 , \32146 ,
         \32147 , \32148 , \32149 , \32150 , \32151 , \32152 , \32153 , \32154 , \32155 , \32156 ,
         \32157 , \32158 , \32159 , \32160 , \32161 , \32162 , \32163 , \32164 , \32165 , \32166 ,
         \32167 , \32168 , \32169 , \32170 , \32171 , \32172 , \32173 , \32174 , \32175 , \32176 ,
         \32177 , \32178 , \32179_nG9bb4 , \32180 , \32181 , \32182 , \32183 , \32184 , \32185 , \32186 ,
         \32187 , \32188 , \32189 , \32190 , \32191 , \32192 , \32193 , \32194 , \32195 , \32196 ,
         \32197 , \32198 , \32199 , \32200 , \32201 , \32202 , \32203 , \32204 , \32205 , \32206 ,
         \32207 , \32208 , \32209 , \32210 , \32211 , \32212 , \32213 , \32214 , \32215 , \32216 ,
         \32217 , \32218 , \32219 , \32220 , \32221 , \32222 , \32223 , \32224 , \32225 , \32226 ,
         \32227 , \32228 , \32229 , \32230 , \32231 , \32232 , \32233 , \32234 , \32235 , \32236 ,
         \32237 , \32238 , \32239 , \32240 , \32241 , \32242 , \32243 , \32244 , \32245 , \32246 ,
         \32247 , \32248 , \32249 , \32250 , \32251 , \32252 , \32253 , \32254 , \32255 , \32256 ,
         \32257 , \32258 , \32259 , \32260 , \32261 , \32262 , \32263 , \32264 , \32265 , \32266 ,
         \32267 , \32268 , \32269 , \32270 , \32271 , \32272 , \32273 , \32274 , \32275 , \32276 ,
         \32277 , \32278 , \32279 , \32280 , \32281 , \32282 , \32283 , \32284 , \32285 , \32286 ,
         \32287 , \32288 , \32289 , \32290 , \32291 , \32292 , \32293 , \32294 , \32295 , \32296 ,
         \32297 , \32298 , \32299 , \32300 , \32301 , \32302 , \32303 , \32304 , \32305 , \32306 ,
         \32307 , \32308 , \32309 , \32310 , \32311 , \32312 , \32313 , \32314 , \32315 , \32316 ,
         \32317 , \32318 , \32319 , \32320 , \32321 , \32322 , \32323 , \32324 , \32325 , \32326 ,
         \32327 , \32328 , \32329 , \32330 , \32331 , \32332 , \32333 , \32334 , \32335 , \32336 ,
         \32337 , \32338 , \32339 , \32340 , \32341 , \32342 , \32343 , \32344 , \32345 , \32346 ,
         \32347 , \32348 , \32349 , \32350 , \32351 , \32352 , \32353 , \32354 , \32355 , \32356 ,
         \32357 , \32358 , \32359 , \32360 , \32361 , \32362 , \32363 , \32364 , \32365 , \32366 ,
         \32367 , \32368 , \32369 , \32370 , \32371 , \32372 , \32373 , \32374 , \32375 , \32376 ,
         \32377 , \32378 , \32379 , \32380 , \32381 , \32382 , \32383 , \32384 , \32385 , \32386 ,
         \32387 , \32388 , \32389 , \32390 , \32391 , \32392 , \32393 , \32394 , \32395 , \32396 ,
         \32397 , \32398 , \32399 , \32400 , \32401 , \32402 , \32403 , \32404 , \32405 , \32406 ,
         \32407 , \32408 , \32409 , \32410 , \32411 , \32412 , \32413 , \32414 , \32415 , \32416 ,
         \32417 , \32418 , \32419 , \32420 , \32421 , \32422 , \32423 , \32424 , \32425 , \32426 ,
         \32427 , \32428 , \32429 , \32430 , \32431 , \32432 , \32433 , \32434 , \32435 , \32436 ,
         \32437 , \32438 , \32439 , \32440 , \32441 , \32442 , \32443 , \32444 , \32445 , \32446 ,
         \32447 , \32448 , \32449 , \32450 , \32451 , \32452 , \32453 , \32454 , \32455 , \32456 ,
         \32457 , \32458 , \32459 , \32460 , \32461 , \32462 , \32463 , \32464 , \32465 , \32466 ,
         \32467 , \32468 , \32469 , \32470 , \32471 , \32472 , \32473 , \32474 , \32475 , \32476 ,
         \32477 , \32478 , \32479 , \32480 , \32481 , \32482 , \32483 , \32484 , \32485 , \32486 ,
         \32487 , \32488 , \32489 , \32490 , \32491 , \32492 , \32493 , \32494 , \32495 , \32496 ,
         \32497 , \32498 , \32499 , \32500 , \32501 , \32502 , \32503 , \32504 , \32505 , \32506 ,
         \32507 , \32508 , \32509 , \32510 , \32511 , \32512 , \32513 , \32514 , \32515 , \32516 ,
         \32517 , \32518 , \32519 , \32520 , \32521 , \32522 , \32523 , \32524 , \32525 , \32526 ,
         \32527 , \32528 , \32529 , \32530 , \32531 , \32532 , \32533 , \32534 , \32535 , \32536 ,
         \32537 , \32538 , \32539 , \32540 , \32541 , \32542 , \32543 , \32544 , \32545 , \32546 ,
         \32547 , \32548 , \32549 , \32550 , \32551 , \32552 , \32553 , \32554 , \32555 , \32556 ,
         \32557 , \32558 , \32559 , \32560 , \32561 , \32562 , \32563 , \32564 , \32565 , \32566 ,
         \32567 , \32568 , \32569 , \32570 , \32571 , \32572 , \32573 , \32574 , \32575 , \32576 ,
         \32577 , \32578 , \32579 , \32580 , \32581 , \32582 , \32583 , \32584 , \32585 , \32586 ,
         \32587 , \32588 , \32589 , \32590 , \32591 , \32592 , \32593 , \32594 , \32595 , \32596 ,
         \32597 , \32598 , \32599 , \32600 , \32601 , \32602 , \32603 , \32604 , \32605 , \32606 ,
         \32607 , \32608 , \32609 , \32610 , \32611 , \32612 , \32613 , \32614 , \32615 , \32616 ,
         \32617 , \32618 , \32619 , \32620 , \32621 , \32622 , \32623 , \32624 , \32625 , \32626 ,
         \32627 , \32628 , \32629 , \32630 , \32631 , \32632 , \32633 , \32634 , \32635 , \32636 ,
         \32637 , \32638 , \32639 , \32640 , \32641 , \32642 , \32643 , \32644 , \32645 , \32646 ,
         \32647 , \32648 , \32649 , \32650 , \32651 , \32652 , \32653 , \32654 , \32655 , \32656 ,
         \32657 , \32658 , \32659 , \32660_nG65d4 , \32661 , \32662 , \32663 , \32664 , \32665 , \32666 ,
         \32667 , \32668 , \32669 , \32670 , \32671 , \32672 , \32673 , \32674 , \32675 , \32676 ,
         \32677 , \32678 , \32679 , \32680 , \32681 , \32682 , \32683 , \32684 , \32685 , \32686 ,
         \32687 , \32688 , \32689 , \32690 , \32691 , \32692 , \32693 , \32694 , \32695 , \32696 ,
         \32697 , \32698 , \32699 , \32700 , \32701 , \32702 , \32703 , \32704 , \32705 , \32706 ,
         \32707 , \32708 , \32709 , \32710 , \32711 , \32712 , \32713 , \32714 , \32715 , \32716 ,
         \32717 , \32718 , \32719 , \32720 , \32721 , \32722 , \32723 , \32724 , \32725 , \32726 ,
         \32727 , \32728 , \32729 , \32730 , \32731 , \32732 , \32733 , \32734 , \32735 , \32736 ,
         \32737 , \32738 , \32739 , \32740 , \32741 , \32742 , \32743 , \32744 , \32745 , \32746 ,
         \32747 , \32748 , \32749 , \32750 , \32751 , \32752 , \32753 , \32754 , \32755 , \32756 ,
         \32757 , \32758 , \32759 , \32760 , \32761 , \32762 , \32763 , \32764 , \32765 , \32766 ,
         \32767 , \32768 , \32769 , \32770 , \32771 , \32772 , \32773 , \32774 , \32775 , \32776 ,
         \32777 , \32778 , \32779 , \32780 , \32781 , \32782 , \32783 , \32784 , \32785 , \32786 ,
         \32787 , \32788 , \32789 , \32790 , \32791 , \32792_nG65d5 , \32793_nG65d6 , \32794 , \32795 , \32796 ,
         \32797 , \32798 , \32799_nG64f1 , \32800_nG6575 , \32801_nG6576 , \32802 , \32803 , \32804 , \32805 , \32806 ,
         \32807 , \32808 , \32809 , \32810 , \32811 , \32812 , \32813 , \32814 , \32815 , \32816 ,
         \32817 , \32818 , \32819 , \32820 , \32821 , \32822 , \32823 , \32824 , \32825 , \32826 ,
         \32827 , \32828 , \32829 , \32830 , \32831 , \32832 , \32833 , \32834 , \32835 , \32836 ,
         \32837 , \32838 , \32839 , \32840 , \32841 , \32842 , \32843 , \32844 , \32845 , \32846 ,
         \32847 , \32848 , \32849 , \32850 , \32851 , \32852 , \32853 , \32854 , \32855 , \32856 ,
         \32857 , \32858 , \32859 , \32860 , \32861 , \32862 , \32863 , \32864 , \32865 , \32866 ,
         \32867 , \32868 , \32869 , \32870 , \32871 , \32872 , \32873 , \32874 , \32875 , \32876 ,
         \32877 , \32878 , \32879 , \32880 , \32881 , \32882 , \32883 , \32884 , \32885 , \32886 ,
         \32887 , \32888_nG9bb1 , \32889 , \32890 , \32891 , \32892 , \32893 , \32894 , \32895 , \32896 ,
         \32897 , \32898 , \32899 , \32900 , \32901 , \32902 , \32903 , \32904 , \32905 , \32906 ,
         \32907 , \32908 , \32909 , \32910 , \32911 , \32912 , \32913 , \32914 , \32915 , \32916 ,
         \32917 , \32918 , \32919 , \32920 , \32921 , \32922 , \32923 , \32924 , \32925 , \32926 ,
         \32927 , \32928 , \32929 , \32930 , \32931 , \32932 , \32933 , \32934 , \32935 , \32936 ,
         \32937 , \32938 , \32939 , \32940 , \32941 , \32942 , \32943 , \32944 , \32945 , \32946 ,
         \32947 , \32948 , \32949 , \32950 , \32951 , \32952 , \32953 , \32954 , \32955 , \32956 ,
         \32957 , \32958 , \32959 , \32960 , \32961 , \32962 , \32963 , \32964 , \32965 , \32966 ,
         \32967 , \32968 , \32969 , \32970 , \32971 , \32972 , \32973 , \32974 , \32975 , \32976 ,
         \32977 , \32978 , \32979 , \32980 , \32981 , \32982 , \32983 , \32984 , \32985 , \32986 ,
         \32987 , \32988 , \32989 , \32990 , \32991 , \32992 , \32993 , \32994 , \32995 , \32996 ,
         \32997 , \32998 , \32999 , \33000 , \33001 , \33002 , \33003 , \33004 , \33005 , \33006 ,
         \33007 , \33008 , \33009 , \33010 , \33011 , \33012 , \33013 , \33014 , \33015 , \33016 ,
         \33017 , \33018 , \33019 , \33020 , \33021 , \33022 , \33023 , \33024 , \33025 , \33026 ,
         \33027 , \33028 , \33029 , \33030 , \33031 , \33032 , \33033 , \33034 , \33035 , \33036 ,
         \33037 , \33038 , \33039 , \33040 , \33041 , \33042 , \33043 , \33044 , \33045 , \33046 ,
         \33047 , \33048 , \33049 , \33050 , \33051 , \33052 , \33053 , \33054 , \33055 , \33056 ,
         \33057 , \33058 , \33059 , \33060 , \33061 , \33062 , \33063 , \33064 , \33065 , \33066 ,
         \33067 , \33068 , \33069 , \33070 , \33071 , \33072 , \33073 , \33074 , \33075 , \33076 ,
         \33077 , \33078 , \33079 , \33080 , \33081 , \33082 , \33083 , \33084 , \33085 , \33086 ,
         \33087 , \33088 , \33089 , \33090 , \33091 , \33092 , \33093 , \33094 , \33095 , \33096 ,
         \33097 , \33098 , \33099 , \33100 , \33101 , \33102 , \33103 , \33104 , \33105 , \33106 ,
         \33107 , \33108 , \33109 , \33110 , \33111 , \33112 , \33113 , \33114 , \33115 , \33116 ,
         \33117 , \33118 , \33119 , \33120 , \33121 , \33122 , \33123 , \33124 , \33125 , \33126 ,
         \33127 , \33128 , \33129 , \33130 , \33131 , \33132 , \33133 , \33134 , \33135 , \33136 ,
         \33137 , \33138 , \33139 , \33140 , \33141 , \33142 , \33143 , \33144 , \33145 , \33146 ,
         \33147 , \33148 , \33149 , \33150 , \33151 , \33152 , \33153 , \33154 , \33155 , \33156 ,
         \33157 , \33158 , \33159 , \33160 , \33161 , \33162 , \33163 , \33164 , \33165 , \33166 ,
         \33167 , \33168 , \33169 , \33170 , \33171 , \33172 , \33173 , \33174 , \33175 , \33176 ,
         \33177 , \33178 , \33179 , \33180 , \33181_nG9bae , \33182 , \33183 , \33184 , \33185 , \33186 ,
         \33187 , \33188 , \33189 , \33190 , \33191 , \33192 , \33193 , \33194 , \33195 , \33196 ,
         \33197 , \33198 , \33199 , \33200 , \33201 , \33202 , \33203 , \33204 , \33205 , \33206 ,
         \33207 , \33208 , \33209 , \33210 , \33211 , \33212 , \33213 , \33214 , \33215 , \33216 ,
         \33217 , \33218 , \33219 , \33220 , \33221 , \33222 , \33223 , \33224 , \33225 , \33226 ,
         \33227 , \33228 , \33229 , \33230 , \33231 , \33232 , \33233 , \33234 , \33235 , \33236 ,
         \33237 , \33238 , \33239 , \33240 , \33241 , \33242 , \33243 , \33244 , \33245 , \33246 ,
         \33247 , \33248 , \33249 , \33250 , \33251 , \33252 , \33253 , \33254 , \33255 , \33256 ,
         \33257 , \33258 , \33259 , \33260 , \33261 , \33262 , \33263 , \33264 , \33265 , \33266 ,
         \33267 , \33268 , \33269 , \33270 , \33271 , \33272 , \33273 , \33274 , \33275 , \33276 ,
         \33277 , \33278 , \33279 , \33280 , \33281 , \33282 , \33283 , \33284 , \33285 , \33286 ,
         \33287 , \33288 , \33289 , \33290 , \33291 , \33292 , \33293 , \33294 , \33295 , \33296 ,
         \33297 , \33298 , \33299 , \33300 , \33301 , \33302 , \33303 , \33304 , \33305 , \33306 ,
         \33307 , \33308 , \33309 , \33310 , \33311 , \33312 , \33313 , \33314 , \33315 , \33316 ,
         \33317 , \33318 , \33319 , \33320 , \33321 , \33322 , \33323 , \33324 , \33325 , \33326 ,
         \33327 , \33328 , \33329 , \33330 , \33331 , \33332 , \33333 , \33334 , \33335 , \33336 ,
         \33337 , \33338 , \33339 , \33340 , \33341 , \33342 , \33343 , \33344 , \33345 , \33346 ,
         \33347 , \33348 , \33349 , \33350 , \33351 , \33352 , \33353 , \33354 , \33355 , \33356 ,
         \33357 , \33358 , \33359 , \33360 , \33361 , \33362 , \33363 , \33364 , \33365 , \33366 ,
         \33367 , \33368 , \33369 , \33370 , \33371 , \33372 , \33373 , \33374 , \33375 , \33376 ,
         \33377 , \33378 , \33379 , \33380 , \33381 , \33382 , \33383 , \33384 , \33385 , \33386 ,
         \33387 , \33388 , \33389 , \33390 , \33391 , \33392 , \33393 , \33394 , \33395 , \33396 ,
         \33397 , \33398 , \33399 , \33400 , \33401 , \33402 , \33403 , \33404 , \33405 , \33406 ,
         \33407 , \33408 , \33409 , \33410 , \33411 , \33412 , \33413 , \33414 , \33415 , \33416 ,
         \33417 , \33418 , \33419 , \33420 , \33421 , \33422 , \33423 , \33424 , \33425 , \33426 ,
         \33427 , \33428 , \33429 , \33430 , \33431 , \33432 , \33433 , \33434 , \33435 , \33436 ,
         \33437 , \33438 , \33439 , \33440 , \33441 , \33442 , \33443 , \33444 , \33445 , \33446 ,
         \33447 , \33448 , \33449 , \33450 , \33451 , \33452 , \33453 , \33454 , \33455 , \33456 ,
         \33457 , \33458 , \33459 , \33460 , \33461 , \33462 , \33463 , \33464 , \33465 , \33466 ,
         \33467 , \33468 , \33469 , \33470 , \33471 , \33472 , \33473 , \33474 , \33475 , \33476 ,
         \33477 , \33478 , \33479 , \33480 , \33481 , \33482 , \33483 , \33484 , \33485 , \33486 ,
         \33487 , \33488 , \33489 , \33490 , \33491 , \33492 , \33493 , \33494 , \33495 , \33496 ,
         \33497 , \33498 , \33499 , \33500 , \33501 , \33502 , \33503 , \33504 , \33505 , \33506 ,
         \33507 , \33508 , \33509 , \33510 , \33511 , \33512 , \33513 , \33514 , \33515 , \33516 ,
         \33517 , \33518 , \33519 , \33520 , \33521 , \33522 , \33523 , \33524 , \33525 , \33526 ,
         \33527 , \33528 , \33529 , \33530 , \33531 , \33532 , \33533 , \33534 , \33535 , \33536 ,
         \33537 , \33538 , \33539 , \33540 , \33541 , \33542 , \33543 , \33544 , \33545 , \33546 ,
         \33547 , \33548 , \33549 , \33550 , \33551 , \33552 , \33553 , \33554 , \33555 , \33556 ,
         \33557 , \33558 , \33559 , \33560 , \33561 , \33562 , \33563 , \33564 , \33565 , \33566 ,
         \33567 , \33568 , \33569 , \33570 , \33571 , \33572 , \33573 , \33574 , \33575 , \33576 ,
         \33577 , \33578 , \33579 , \33580 , \33581 , \33582 , \33583 , \33584 , \33585 , \33586 ,
         \33587 , \33588 , \33589 , \33590 , \33591 , \33592 , \33593 , \33594 , \33595 , \33596 ,
         \33597 , \33598 , \33599 , \33600 , \33601 , \33602 , \33603 , \33604 , \33605 , \33606 ,
         \33607 , \33608 , \33609 , \33610 , \33611 , \33612 , \33613_nG9bab , \33614 , \33615 , \33616 ,
         \33617 , \33618 , \33619 , \33620 , \33621 , \33622 , \33623 , \33624 , \33625 , \33626 ,
         \33627 , \33628 , \33629 , \33630 , \33631 , \33632 , \33633 , \33634 , \33635 , \33636 ,
         \33637 , \33638 , \33639 , \33640 , \33641 , \33642 , \33643 , \33644 , \33645 , \33646 ,
         \33647 , \33648 , \33649 , \33650 , \33651 , \33652 , \33653 , \33654 , \33655 , \33656 ,
         \33657 , \33658 , \33659 , \33660 , \33661 , \33662 , \33663 , \33664 , \33665 , \33666 ,
         \33667 , \33668 , \33669 , \33670 , \33671 , \33672 , \33673 , \33674 , \33675 , \33676 ,
         \33677 , \33678 , \33679 , \33680 , \33681 , \33682 , \33683 , \33684 , \33685 , \33686 ,
         \33687 , \33688 , \33689 , \33690 , \33691 , \33692 , \33693 , \33694 , \33695 , \33696 ,
         \33697 , \33698 , \33699 , \33700 , \33701 , \33702 , \33703 , \33704 , \33705 , \33706 ,
         \33707 , \33708 , \33709 , \33710 , \33711 , \33712 , \33713 , \33714 , \33715 , \33716 ,
         \33717 , \33718 , \33719 , \33720 , \33721 , \33722 , \33723 , \33724 , \33725 , \33726 ,
         \33727 , \33728 , \33729 , \33730 , \33731 , \33732 , \33733 , \33734 , \33735 , \33736 ,
         \33737 , \33738 , \33739 , \33740 , \33741 , \33742 , \33743 , \33744 , \33745 , \33746 ,
         \33747 , \33748 , \33749 , \33750 , \33751 , \33752 , \33753 , \33754 , \33755 , \33756 ,
         \33757 , \33758 , \33759 , \33760 , \33761 , \33762 , \33763 , \33764 , \33765 , \33766 ,
         \33767 , \33768 , \33769 , \33770 , \33771 , \33772 , \33773 , \33774 , \33775 , \33776 ,
         \33777 , \33778 , \33779 , \33780 , \33781 , \33782 , \33783 , \33784 , \33785 , \33786 ,
         \33787 , \33788 , \33789 , \33790 , \33791 , \33792 , \33793 , \33794 , \33795 , \33796 ,
         \33797 , \33798 , \33799 , \33800 , \33801 , \33802 , \33803 , \33804 , \33805 , \33806 ,
         \33807 , \33808 , \33809 , \33810 , \33811 , \33812 , \33813 , \33814 , \33815 , \33816 ,
         \33817 , \33818 , \33819 , \33820 , \33821 , \33822 , \33823 , \33824 , \33825 , \33826 ,
         \33827 , \33828 , \33829 , \33830 , \33831 , \33832 , \33833 , \33834 , \33835 , \33836 ,
         \33837 , \33838 , \33839 , \33840 , \33841 , \33842 , \33843 , \33844 , \33845 , \33846 ,
         \33847 , \33848 , \33849 , \33850 , \33851 , \33852 , \33853 , \33854 , \33855 , \33856 ,
         \33857 , \33858 , \33859 , \33860 , \33861 , \33862 , \33863 , \33864 , \33865 , \33866 ,
         \33867 , \33868 , \33869 , \33870 , \33871 , \33872 , \33873 , \33874 , \33875 , \33876 ,
         \33877 , \33878 , \33879 , \33880 , \33881 , \33882 , \33883 , \33884 , \33885 , \33886 ,
         \33887 , \33888 , \33889 , \33890 , \33891 , \33892 , \33893 , \33894 , \33895 , \33896 ,
         \33897 , \33898 , \33899 , \33900 , \33901 , \33902 , \33903 , \33904 , \33905 , \33906 ,
         \33907 , \33908 , \33909 , \33910 , \33911 , \33912 , \33913 , \33914 , \33915 , \33916 ,
         \33917 , \33918 , \33919 , \33920 , \33921 , \33922 , \33923 , \33924 , \33925 , \33926 ,
         \33927 , \33928 , \33929 , \33930 , \33931 , \33932 , \33933 , \33934 , \33935 , \33936 ,
         \33937 , \33938 , \33939 , \33940 , \33941 , \33942 , \33943 , \33944 , \33945 , \33946 ,
         \33947 , \33948 , \33949 , \33950 , \33951 , \33952 , \33953 , \33954 , \33955 , \33956 ,
         \33957 , \33958 , \33959 , \33960 , \33961 , \33962 , \33963 , \33964 , \33965 , \33966 ,
         \33967 , \33968 , \33969 , \33970 , \33971 , \33972 , \33973 , \33974 , \33975 , \33976 ,
         \33977 , \33978 , \33979 , \33980 , \33981 , \33982 , \33983 , \33984 , \33985 , \33986 ,
         \33987 , \33988 , \33989 , \33990 , \33991 , \33992 , \33993 , \33994 , \33995 , \33996 ,
         \33997 , \33998 , \33999 , \34000 , \34001 , \34002 , \34003 , \34004 , \34005 , \34006 ,
         \34007 , \34008 , \34009 , \34010 , \34011 , \34012 , \34013 , \34014 , \34015 , \34016 ,
         \34017 , \34018 , \34019 , \34020 , \34021 , \34022 , \34023 , \34024 , \34025 , \34026 ,
         \34027 , \34028 , \34029 , \34030 , \34031 , \34032 , \34033 , \34034 , \34035 , \34036 ,
         \34037 , \34038 , \34039 , \34040 , \34041_nG9ba8 , \34042 , \34043 , \34044 , \34045 , \34046 ,
         \34047 , \34048 , \34049 , \34050 , \34051 , \34052 , \34053 , \34054 , \34055 , \34056 ,
         \34057 , \34058 , \34059 , \34060 , \34061 , \34062 , \34063 , \34064 , \34065 , \34066 ,
         \34067 , \34068 , \34069 , \34070 , \34071 , \34072 , \34073 , \34074 , \34075 , \34076 ,
         \34077 , \34078 , \34079 , \34080 , \34081 , \34082 , \34083 , \34084 , \34085 , \34086 ,
         \34087 , \34088 , \34089 , \34090 , \34091 , \34092 , \34093 , \34094 , \34095 , \34096 ,
         \34097 , \34098 , \34099 , \34100 , \34101 , \34102 , \34103 , \34104 , \34105 , \34106 ,
         \34107 , \34108 , \34109 , \34110 , \34111 , \34112 , \34113 , \34114 , \34115 , \34116 ,
         \34117 , \34118 , \34119 , \34120 , \34121 , \34122 , \34123 , \34124 , \34125 , \34126 ,
         \34127 , \34128 , \34129 , \34130 , \34131 , \34132 , \34133 , \34134 , \34135 , \34136 ,
         \34137 , \34138 , \34139 , \34140 , \34141 , \34142 , \34143 , \34144 , \34145 , \34146 ,
         \34147 , \34148 , \34149 , \34150 , \34151 , \34152 , \34153 , \34154 , \34155 , \34156 ,
         \34157 , \34158 , \34159 , \34160 , \34161 , \34162 , \34163 , \34164 , \34165 , \34166 ,
         \34167 , \34168 , \34169 , \34170 , \34171 , \34172 , \34173 , \34174 , \34175 , \34176 ,
         \34177 , \34178 , \34179 , \34180 , \34181 , \34182 , \34183 , \34184 , \34185 , \34186 ,
         \34187 , \34188 , \34189 , \34190 , \34191 , \34192 , \34193 , \34194 , \34195 , \34196 ,
         \34197 , \34198 , \34199 , \34200 , \34201 , \34202 , \34203 , \34204 , \34205 , \34206 ,
         \34207 , \34208 , \34209 , \34210 , \34211 , \34212 , \34213 , \34214 , \34215 , \34216 ,
         \34217 , \34218 , \34219 , \34220 , \34221 , \34222 , \34223 , \34224 , \34225 , \34226 ,
         \34227 , \34228 , \34229 , \34230 , \34231 , \34232 , \34233 , \34234 , \34235 , \34236 ,
         \34237 , \34238 , \34239 , \34240 , \34241 , \34242 , \34243 , \34244 , \34245 , \34246 ,
         \34247 , \34248 , \34249 , \34250 , \34251 , \34252 , \34253 , \34254 , \34255 , \34256 ,
         \34257 , \34258 , \34259 , \34260 , \34261 , \34262 , \34263 , \34264 , \34265 , \34266 ,
         \34267 , \34268 , \34269 , \34270 , \34271 , \34272 , \34273 , \34274 , \34275 , \34276 ,
         \34277 , \34278 , \34279 , \34280 , \34281 , \34282 , \34283 , \34284 , \34285 , \34286 ,
         \34287 , \34288 , \34289 , \34290 , \34291 , \34292 , \34293 , \34294_nG9ba5 , \34295 , \34296 ,
         \34297 , \34298 , \34299 , \34300 , \34301 , \34302 , \34303 , \34304 , \34305 , \34306 ,
         \34307 , \34308 , \34309 , \34310 , \34311 , \34312 , \34313 , \34314 , \34315 , \34316 ,
         \34317 , \34318 , \34319 , \34320 , \34321 , \34322 , \34323 , \34324 , \34325 , \34326 ,
         \34327 , \34328 , \34329 , \34330 , \34331 , \34332 , \34333 , \34334 , \34335 , \34336 ,
         \34337 , \34338 , \34339 , \34340 , \34341 , \34342 , \34343 , \34344 , \34345 , \34346 ,
         \34347 , \34348 , \34349 , \34350 , \34351 , \34352 , \34353 , \34354 , \34355 , \34356 ,
         \34357 , \34358 , \34359 , \34360 , \34361 , \34362 , \34363 , \34364 , \34365 , \34366 ,
         \34367 , \34368 , \34369 , \34370 , \34371 , \34372 , \34373 , \34374 , \34375 , \34376 ,
         \34377 , \34378 , \34379 , \34380 , \34381 , \34382 , \34383 , \34384 , \34385 , \34386 ,
         \34387 , \34388 , \34389 , \34390 , \34391 , \34392 , \34393 , \34394 , \34395 , \34396 ,
         \34397 , \34398 , \34399 , \34400 , \34401 , \34402 , \34403 , \34404 , \34405 , \34406 ,
         \34407 , \34408 , \34409 , \34410 , \34411 , \34412 , \34413 , \34414 , \34415 , \34416 ,
         \34417 , \34418 , \34419 , \34420 , \34421 , \34422 , \34423 , \34424 , \34425 , \34426 ,
         \34427 , \34428 , \34429 , \34430 , \34431 , \34432 , \34433 , \34434 , \34435 , \34436 ,
         \34437 , \34438 , \34439 , \34440 , \34441 , \34442 , \34443 , \34444 , \34445 , \34446 ,
         \34447 , \34448 , \34449 , \34450 , \34451 , \34452 , \34453 , \34454 , \34455 , \34456 ,
         \34457 , \34458 , \34459 , \34460 , \34461 , \34462 , \34463 , \34464 , \34465 , \34466 ,
         \34467 , \34468 , \34469 , \34470 , \34471 , \34472 , \34473 , \34474 , \34475 , \34476 ,
         \34477 , \34478 , \34479 , \34480 , \34481 , \34482 , \34483 , \34484 , \34485 , \34486 ,
         \34487 , \34488 , \34489 , \34490 , \34491 , \34492 , \34493 , \34494 , \34495 , \34496 ,
         \34497 , \34498 , \34499 , \34500 , \34501 , \34502 , \34503 , \34504 , \34505 , \34506 ,
         \34507 , \34508 , \34509 , \34510 , \34511 , \34512 , \34513 , \34514 , \34515 , \34516 ,
         \34517 , \34518 , \34519 , \34520 , \34521 , \34522 , \34523 , \34524 , \34525 , \34526 ,
         \34527 , \34528 , \34529 , \34530 , \34531 , \34532 , \34533 , \34534 , \34535 , \34536 ,
         \34537 , \34538 , \34539 , \34540 , \34541 , \34542 , \34543 , \34544 , \34545 , \34546 ,
         \34547 , \34548 , \34549 , \34550 , \34551 , \34552 , \34553 , \34554 , \34555 , \34556 ,
         \34557 , \34558 , \34559 , \34560 , \34561 , \34562 , \34563 , \34564 , \34565 , \34566 ,
         \34567 , \34568 , \34569 , \34570 , \34571 , \34572 , \34573 , \34574 , \34575 , \34576 ,
         \34577 , \34578 , \34579 , \34580 , \34581 , \34582 , \34583 , \34584 , \34585 , \34586 ,
         \34587 , \34588 , \34589 , \34590 , \34591 , \34592 , \34593 , \34594 , \34595 , \34596 ,
         \34597 , \34598 , \34599 , \34600 , \34601 , \34602 , \34603 , \34604 , \34605 , \34606 ,
         \34607 , \34608 , \34609 , \34610 , \34611 , \34612 , \34613 , \34614 , \34615 , \34616 ,
         \34617 , \34618 , \34619 , \34620 , \34621 , \34622 , \34623 , \34624 , \34625 , \34626 ,
         \34627 , \34628 , \34629 , \34630 , \34631 , \34632 , \34633 , \34634 , \34635 , \34636 ,
         \34637 , \34638 , \34639 , \34640 , \34641 , \34642 , \34643_nG9ba2 , \34644 , \34645 , \34646 ,
         \34647 , \34648 , \34649 , \34650 , \34651 , \34652 , \34653 , \34654 , \34655 , \34656 ,
         \34657 , \34658 , \34659 , \34660 , \34661 , \34662 , \34663 , \34664 , \34665 , \34666 ,
         \34667 , \34668 , \34669 , \34670 , \34671 , \34672 , \34673 , \34674 , \34675 , \34676 ,
         \34677 , \34678 , \34679 , \34680 , \34681 , \34682 , \34683 , \34684 , \34685 , \34686 ,
         \34687 , \34688 , \34689 , \34690 , \34691 , \34692 , \34693 , \34694 , \34695 , \34696 ,
         \34697 , \34698 , \34699 , \34700 , \34701 , \34702 , \34703 , \34704 , \34705 , \34706 ,
         \34707 , \34708 , \34709 , \34710 , \34711 , \34712 , \34713 , \34714 , \34715 , \34716 ,
         \34717 , \34718 , \34719 , \34720 , \34721 , \34722 , \34723 , \34724 , \34725 , \34726 ,
         \34727 , \34728 , \34729 , \34730 , \34731 , \34732 , \34733 , \34734 , \34735 , \34736 ,
         \34737 , \34738 , \34739 , \34740 , \34741 , \34742 , \34743 , \34744 , \34745 , \34746 ,
         \34747 , \34748 , \34749 , \34750 , \34751 , \34752 , \34753 , \34754 , \34755 , \34756 ,
         \34757 , \34758 , \34759 , \34760 , \34761 , \34762 , \34763 , \34764 , \34765 , \34766 ,
         \34767 , \34768 , \34769 , \34770 , \34771 , \34772 , \34773 , \34774 , \34775 , \34776 ,
         \34777 , \34778 , \34779 , \34780 , \34781 , \34782 , \34783 , \34784 , \34785 , \34786 ,
         \34787 , \34788 , \34789 , \34790 , \34791 , \34792 , \34793 , \34794 , \34795 , \34796 ,
         \34797 , \34798 , \34799 , \34800 , \34801 , \34802 , \34803 , \34804 , \34805 , \34806 ,
         \34807 , \34808 , \34809 , \34810 , \34811 , \34812 , \34813 , \34814 , \34815 , \34816 ,
         \34817 , \34818 , \34819 , \34820 , \34821 , \34822 , \34823 , \34824 , \34825 , \34826 ,
         \34827 , \34828 , \34829 , \34830 , \34831 , \34832 , \34833 , \34834 , \34835 , \34836 ,
         \34837 , \34838 , \34839 , \34840 , \34841 , \34842 , \34843 , \34844 , \34845 , \34846 ,
         \34847 , \34848 , \34849 , \34850 , \34851 , \34852 , \34853 , \34854 , \34855 , \34856 ,
         \34857 , \34858 , \34859 , \34860 , \34861 , \34862 , \34863 , \34864 , \34865 , \34866 ,
         \34867 , \34868 , \34869 , \34870 , \34871 , \34872 , \34873 , \34874 , \34875 , \34876 ,
         \34877 , \34878 , \34879 , \34880 , \34881 , \34882 , \34883 , \34884 , \34885 , \34886 ,
         \34887 , \34888 , \34889 , \34890 , \34891 , \34892 , \34893 , \34894 , \34895 , \34896 ,
         \34897 , \34898 , \34899 , \34900 , \34901 , \34902 , \34903 , \34904 , \34905 , \34906 ,
         \34907 , \34908 , \34909 , \34910 , \34911 , \34912 , \34913 , \34914 , \34915 , \34916 ,
         \34917 , \34918 , \34919 , \34920 , \34921 , \34922 , \34923 , \34924 , \34925 , \34926 ,
         \34927 , \34928 , \34929 , \34930 , \34931 , \34932 , \34933 , \34934 , \34935 , \34936 ,
         \34937 , \34938 , \34939 , \34940 , \34941 , \34942 , \34943 , \34944 , \34945 , \34946 ,
         \34947 , \34948 , \34949 , \34950 , \34951 , \34952 , \34953 , \34954 , \34955 , \34956 ,
         \34957 , \34958 , \34959 , \34960 , \34961 , \34962 , \34963 , \34964 , \34965 , \34966 ,
         \34967 , \34968 , \34969 , \34970 , \34971 , \34972 , \34973 , \34974 , \34975 , \34976 ,
         \34977 , \34978 , \34979 , \34980 , \34981 , \34982 , \34983 , \34984 , \34985 , \34986 ,
         \34987 , \34988 , \34989 , \34990 , \34991 , \34992 , \34993 , \34994 , \34995 , \34996 ,
         \34997 , \34998 , \34999 , \35000 , \35001 , \35002 , \35003 , \35004 , \35005 , \35006 ,
         \35007 , \35008 , \35009 , \35010 , \35011 , \35012 , \35013 , \35014 , \35015 , \35016 ,
         \35017 , \35018 , \35019 , \35020 , \35021 , \35022 , \35023 , \35024 , \35025 , \35026 ,
         \35027 , \35028 , \35029 , \35030 , \35031 , \35032 , \35033 , \35034 , \35035 , \35036 ,
         \35037 , \35038 , \35039 , \35040 , \35041 , \35042 , \35043 , \35044 , \35045 , \35046 ,
         \35047 , \35048 , \35049 , \35050 , \35051 , \35052 , \35053 , \35054 , \35055 , \35056 ,
         \35057 , \35058 , \35059 , \35060 , \35061 , \35062 , \35063 , \35064 , \35065 , \35066 ,
         \35067 , \35068 , \35069 , \35070 , \35071 , \35072 , \35073 , \35074 , \35075 , \35076 ,
         \35077 , \35078 , \35079 , \35080 , \35081 , \35082 , \35083 , \35084 , \35085 , \35086 ,
         \35087 , \35088 , \35089 , \35090 , \35091 , \35092 , \35093 , \35094_nG9b9f , \35095 , \35096 ,
         \35097 , \35098 , \35099 , \35100 , \35101 , \35102 , \35103 , \35104 , \35105 , \35106 ,
         \35107 , \35108 , \35109 , \35110 , \35111 , \35112 , \35113 , \35114 , \35115 , \35116 ,
         \35117 , \35118 , \35119 , \35120 , \35121 , \35122 , \35123 , \35124 , \35125 , \35126 ,
         \35127 , \35128 , \35129 , \35130 , \35131 , \35132 , \35133 , \35134 , \35135 , \35136 ,
         \35137 , \35138 , \35139 , \35140 , \35141 , \35142 , \35143 , \35144 , \35145 , \35146 ,
         \35147 , \35148 , \35149 , \35150 , \35151 , \35152 , \35153 , \35154 , \35155 , \35156 ,
         \35157 , \35158 , \35159 , \35160 , \35161 , \35162 , \35163 , \35164 , \35165 , \35166 ,
         \35167 , \35168 , \35169 , \35170 , \35171 , \35172 , \35173 , \35174 , \35175 , \35176 ,
         \35177 , \35178 , \35179 , \35180 , \35181 , \35182 , \35183 , \35184 , \35185 , \35186 ,
         \35187 , \35188 , \35189 , \35190 , \35191 , \35192 , \35193 , \35194 , \35195 , \35196 ,
         \35197 , \35198 , \35199 , \35200 , \35201 , \35202 , \35203 , \35204 , \35205 , \35206 ,
         \35207 , \35208 , \35209 , \35210 , \35211 , \35212 , \35213 , \35214 , \35215 , \35216 ,
         \35217 , \35218 , \35219 , \35220 , \35221 , \35222 , \35223 , \35224 , \35225 , \35226 ,
         \35227 , \35228 , \35229 , \35230 , \35231 , \35232 , \35233 , \35234 , \35235 , \35236 ,
         \35237 , \35238 , \35239 , \35240 , \35241 , \35242 , \35243 , \35244 , \35245 , \35246 ,
         \35247 , \35248 , \35249 , \35250 , \35251 , \35252 , \35253 , \35254 , \35255 , \35256 ,
         \35257 , \35258 , \35259 , \35260 , \35261 , \35262 , \35263 , \35264 , \35265 , \35266 ,
         \35267 , \35268 , \35269 , \35270 , \35271 , \35272 , \35273 , \35274 , \35275 , \35276 ,
         \35277 , \35278 , \35279 , \35280 , \35281 , \35282 , \35283 , \35284 , \35285 , \35286 ,
         \35287 , \35288 , \35289 , \35290 , \35291 , \35292 , \35293 , \35294 , \35295 , \35296 ,
         \35297 , \35298 , \35299 , \35300 , \35301 , \35302 , \35303 , \35304 , \35305 , \35306 ,
         \35307 , \35308 , \35309 , \35310 , \35311 , \35312 , \35313 , \35314 , \35315 , \35316 ,
         \35317 , \35318 , \35319 , \35320 , \35321 , \35322 , \35323 , \35324 , \35325 , \35326 ,
         \35327 , \35328 , \35329 , \35330 , \35331 , \35332 , \35333 , \35334 , \35335 , \35336 ,
         \35337 , \35338 , \35339 , \35340 , \35341 , \35342 , \35343 , \35344 , \35345 , \35346 ,
         \35347 , \35348 , \35349 , \35350 , \35351 , \35352 , \35353 , \35354 , \35355 , \35356 ,
         \35357 , \35358 , \35359 , \35360 , \35361 , \35362 , \35363 , \35364 , \35365 , \35366 ,
         \35367 , \35368 , \35369 , \35370 , \35371 , \35372 , \35373 , \35374 , \35375 , \35376 ,
         \35377 , \35378 , \35379 , \35380 , \35381 , \35382 , \35383 , \35384 , \35385 , \35386 ,
         \35387 , \35388 , \35389 , \35390 , \35391 , \35392 , \35393 , \35394 , \35395 , \35396 ,
         \35397 , \35398 , \35399 , \35400 , \35401 , \35402 , \35403 , \35404 , \35405 , \35406 ,
         \35407 , \35408 , \35409 , \35410 , \35411 , \35412 , \35413 , \35414 , \35415 , \35416 ,
         \35417 , \35418 , \35419 , \35420 , \35421 , \35422 , \35423 , \35424 , \35425 , \35426 ,
         \35427 , \35428 , \35429 , \35430 , \35431 , \35432 , \35433 , \35434 , \35435 , \35436 ,
         \35437 , \35438 , \35439 , \35440 , \35441 , \35442 , \35443 , \35444 , \35445 , \35446 ,
         \35447 , \35448 , \35449 , \35450 , \35451 , \35452 , \35453 , \35454 , \35455 , \35456 ,
         \35457 , \35458 , \35459 , \35460 , \35461 , \35462 , \35463 , \35464 , \35465 , \35466 ,
         \35467 , \35468 , \35469 , \35470 , \35471 , \35472 , \35473 , \35474 , \35475 , \35476 ,
         \35477 , \35478 , \35479 , \35480 , \35481 , \35482 , \35483 , \35484 , \35485 , \35486 ,
         \35487 , \35488 , \35489 , \35490 , \35491 , \35492 , \35493 , \35494 , \35495 , \35496 ,
         \35497 , \35498 , \35499 , \35500 , \35501 , \35502 , \35503 , \35504 , \35505 , \35506 ,
         \35507 , \35508 , \35509 , \35510 , \35511 , \35512 , \35513 , \35514 , \35515 , \35516 ,
         \35517 , \35518 , \35519 , \35520 , \35521 , \35522 , \35523 , \35524 , \35525 , \35526 ,
         \35527 , \35528 , \35529 , \35530 , \35531 , \35532 , \35533 , \35534 , \35535 , \35536 ,
         \35537 , \35538 , \35539 , \35540 , \35541 , \35542 , \35543 , \35544 , \35545 , \35546 ,
         \35547 , \35548 , \35549 , \35550 , \35551 , \35552 , \35553 , \35554 , \35555 , \35556 ,
         \35557 , \35558 , \35559 , \35560 , \35561 , \35562 , \35563 , \35564 , \35565 , \35566 ,
         \35567 , \35568 , \35569 , \35570_nG9b9c , \35571 , \35572 , \35573 , \35574 , \35575 , \35576 ,
         \35577 , \35578 , \35579 , \35580 , \35581 , \35582 , \35583 , \35584 , \35585 , \35586 ,
         \35587 , \35588 , \35589 , \35590 , \35591 , \35592 , \35593 , \35594 , \35595 , \35596 ,
         \35597 , \35598 , \35599 , \35600 , \35601 , \35602 , \35603 , \35604 , \35605 , \35606 ,
         \35607 , \35608 , \35609 , \35610 , \35611 , \35612 , \35613 , \35614 , \35615 , \35616 ,
         \35617 , \35618 , \35619 , \35620 , \35621 , \35622 , \35623 , \35624 , \35625 , \35626 ,
         \35627 , \35628 , \35629 , \35630 , \35631 , \35632 , \35633 , \35634 , \35635 , \35636 ,
         \35637 , \35638 , \35639 , \35640 , \35641 , \35642 , \35643 , \35644 , \35645 , \35646 ,
         \35647 , \35648 , \35649 , \35650 , \35651 , \35652 , \35653 , \35654 , \35655 , \35656 ,
         \35657 , \35658 , \35659 , \35660 , \35661 , \35662 , \35663 , \35664 , \35665 , \35666 ,
         \35667 , \35668 , \35669 , \35670 , \35671 , \35672 , \35673 , \35674 , \35675 , \35676 ,
         \35677 , \35678 , \35679 , \35680 , \35681 , \35682 , \35683 , \35684 , \35685 , \35686 ,
         \35687 , \35688 , \35689 , \35690 , \35691 , \35692 , \35693 , \35694 , \35695 , \35696 ,
         \35697 , \35698 , \35699 , \35700 , \35701 , \35702 , \35703 , \35704 , \35705 , \35706 ,
         \35707 , \35708 , \35709 , \35710 , \35711 , \35712 , \35713 , \35714 , \35715 , \35716 ,
         \35717 , \35718 , \35719 , \35720 , \35721 , \35722 , \35723 , \35724 , \35725 , \35726 ,
         \35727 , \35728 , \35729 , \35730 , \35731 , \35732 , \35733 , \35734 , \35735 , \35736 ,
         \35737 , \35738 , \35739 , \35740 , \35741 , \35742 , \35743 , \35744 , \35745 , \35746 ,
         \35747 , \35748 , \35749 , \35750 , \35751 , \35752 , \35753 , \35754 , \35755 , \35756 ,
         \35757 , \35758 , \35759 , \35760 , \35761 , \35762 , \35763 , \35764 , \35765 , \35766 ,
         \35767 , \35768 , \35769 , \35770 , \35771 , \35772 , \35773 , \35774 , \35775 , \35776 ,
         \35777 , \35778 , \35779 , \35780 , \35781 , \35782 , \35783 , \35784 , \35785 , \35786 ,
         \35787 , \35788 , \35789 , \35790 , \35791 , \35792 , \35793 , \35794 , \35795 , \35796 ,
         \35797 , \35798 , \35799 , \35800 , \35801_nG9b99 , \35802 , \35803 , \35804 , \35805 , \35806 ,
         \35807 , \35808 , \35809 , \35810 , \35811 , \35812 , \35813 , \35814 , \35815 , \35816 ,
         \35817 , \35818 , \35819 , \35820 , \35821 , \35822 , \35823 , \35824 , \35825 , \35826 ,
         \35827 , \35828 , \35829 , \35830 , \35831 , \35832 , \35833 , \35834 , \35835 , \35836 ,
         \35837 , \35838 , \35839 , \35840 , \35841 , \35842 , \35843 , \35844 , \35845 , \35846 ,
         \35847 , \35848 , \35849 , \35850 , \35851 , \35852 , \35853 , \35854 , \35855 , \35856 ,
         \35857 , \35858 , \35859 , \35860 , \35861 , \35862 , \35863 , \35864 , \35865 , \35866 ,
         \35867 , \35868 , \35869 , \35870 , \35871 , \35872 , \35873 , \35874 , \35875 , \35876 ,
         \35877 , \35878 , \35879 , \35880 , \35881 , \35882 , \35883 , \35884 , \35885 , \35886 ,
         \35887 , \35888 , \35889 , \35890 , \35891 , \35892 , \35893 , \35894 , \35895 , \35896 ,
         \35897 , \35898 , \35899 , \35900 , \35901 , \35902 , \35903 , \35904 , \35905 , \35906 ,
         \35907 , \35908 , \35909 , \35910 , \35911 , \35912 , \35913 , \35914 , \35915 , \35916 ,
         \35917 , \35918 , \35919 , \35920 , \35921 , \35922 , \35923 , \35924 , \35925 , \35926 ,
         \35927 , \35928 , \35929 , \35930 , \35931 , \35932 , \35933 , \35934 , \35935 , \35936 ,
         \35937 , \35938 , \35939 , \35940 , \35941 , \35942 , \35943 , \35944 , \35945 , \35946 ,
         \35947 , \35948 , \35949 , \35950 , \35951 , \35952 , \35953 , \35954 , \35955 , \35956 ,
         \35957 , \35958 , \35959 , \35960 , \35961 , \35962 , \35963 , \35964 , \35965 , \35966 ,
         \35967 , \35968 , \35969 , \35970 , \35971 , \35972 , \35973 , \35974 , \35975 , \35976 ,
         \35977 , \35978 , \35979 , \35980 , \35981 , \35982 , \35983 , \35984 , \35985 , \35986 ,
         \35987 , \35988 , \35989 , \35990 , \35991 , \35992 , \35993 , \35994 , \35995 , \35996 ,
         \35997 , \35998 , \35999 , \36000 , \36001 , \36002 , \36003 , \36004 , \36005 , \36006 ,
         \36007 , \36008 , \36009 , \36010 , \36011 , \36012 , \36013 , \36014 , \36015 , \36016 ,
         \36017 , \36018 , \36019 , \36020 , \36021 , \36022 , \36023 , \36024 , \36025 , \36026 ,
         \36027 , \36028 , \36029 , \36030 , \36031 , \36032 , \36033 , \36034 , \36035 , \36036 ,
         \36037 , \36038 , \36039 , \36040 , \36041 , \36042 , \36043 , \36044 , \36045 , \36046 ,
         \36047 , \36048 , \36049 , \36050 , \36051 , \36052 , \36053 , \36054 , \36055 , \36056 ,
         \36057 , \36058 , \36059 , \36060 , \36061 , \36062 , \36063 , \36064 , \36065 , \36066 ,
         \36067 , \36068 , \36069 , \36070 , \36071 , \36072 , \36073 , \36074 , \36075 , \36076 ,
         \36077 , \36078 , \36079 , \36080 , \36081 , \36082 , \36083 , \36084 , \36085 , \36086 ,
         \36087 , \36088 , \36089 , \36090 , \36091 , \36092 , \36093 , \36094 , \36095 , \36096 ,
         \36097 , \36098 , \36099 , \36100 , \36101 , \36102 , \36103 , \36104 , \36105 , \36106 ,
         \36107 , \36108 , \36109 , \36110 , \36111 , \36112 , \36113 , \36114 , \36115 , \36116 ,
         \36117 , \36118 , \36119 , \36120 , \36121 , \36122 , \36123 , \36124 , \36125 , \36126 ,
         \36127 , \36128 , \36129 , \36130 , \36131 , \36132 , \36133 , \36134 , \36135 , \36136 ,
         \36137 , \36138 , \36139 , \36140 , \36141 , \36142 , \36143 , \36144 , \36145 , \36146 ,
         \36147 , \36148 , \36149 , \36150 , \36151 , \36152 , \36153 , \36154 , \36155 , \36156 ,
         \36157 , \36158 , \36159 , \36160 , \36161 , \36162 , \36163 , \36164 , \36165 , \36166 ,
         \36167 , \36168 , \36169 , \36170 , \36171 , \36172_nG9b96 , \36173 , \36174 , \36175 , \36176 ,
         \36177 , \36178 , \36179 , \36180 , \36181 , \36182 , \36183 , \36184 , \36185 , \36186 ,
         \36187 , \36188 , \36189 , \36190 , \36191 , \36192 , \36193 , \36194 , \36195 , \36196 ,
         \36197 , \36198 , \36199 , \36200 , \36201 , \36202 , \36203 , \36204 , \36205 , \36206 ,
         \36207 , \36208 , \36209 , \36210 , \36211 , \36212 , \36213 , \36214 , \36215 , \36216 ,
         \36217 , \36218 , \36219 , \36220 , \36221 , \36222 , \36223 , \36224 , \36225 , \36226 ,
         \36227 , \36228 , \36229 , \36230 , \36231 , \36232 , \36233 , \36234 , \36235 , \36236 ,
         \36237 , \36238 , \36239 , \36240 , \36241 , \36242 , \36243 , \36244 , \36245 , \36246 ,
         \36247 , \36248 , \36249 , \36250 , \36251 , \36252 , \36253 , \36254 , \36255 , \36256 ,
         \36257 , \36258 , \36259 , \36260 , \36261 , \36262 , \36263 , \36264 , \36265 , \36266 ,
         \36267 , \36268 , \36269 , \36270 , \36271 , \36272 , \36273 , \36274 , \36275 , \36276 ,
         \36277 , \36278 , \36279 , \36280 , \36281 , \36282 , \36283 , \36284 , \36285 , \36286 ,
         \36287 , \36288 , \36289 , \36290 , \36291 , \36292 , \36293 , \36294 , \36295 , \36296 ,
         \36297 , \36298 , \36299 , \36300 , \36301 , \36302 , \36303 , \36304 , \36305 , \36306 ,
         \36307 , \36308 , \36309 , \36310 , \36311 , \36312 , \36313 , \36314 , \36315 , \36316 ,
         \36317 , \36318 , \36319 , \36320 , \36321 , \36322 , \36323 , \36324 , \36325 , \36326 ,
         \36327 , \36328 , \36329 , \36330 , \36331 , \36332 , \36333 , \36334 , \36335 , \36336 ,
         \36337 , \36338 , \36339 , \36340 , \36341 , \36342 , \36343 , \36344 , \36345 , \36346 ,
         \36347 , \36348 , \36349 , \36350 , \36351 , \36352 , \36353 , \36354 , \36355 , \36356 ,
         \36357 , \36358 , \36359 , \36360 , \36361 , \36362 , \36363 , \36364 , \36365 , \36366 ,
         \36367 , \36368 , \36369 , \36370 , \36371 , \36372 , \36373 , \36374 , \36375 , \36376 ,
         \36377 , \36378 , \36379 , \36380 , \36381 , \36382 , \36383 , \36384 , \36385 , \36386 ,
         \36387 , \36388 , \36389 , \36390 , \36391 , \36392 , \36393 , \36394 , \36395 , \36396 ,
         \36397 , \36398 , \36399 , \36400 , \36401 , \36402 , \36403 , \36404 , \36405 , \36406 ,
         \36407 , \36408 , \36409 , \36410 , \36411 , \36412 , \36413 , \36414 , \36415 , \36416 ,
         \36417 , \36418 , \36419 , \36420 , \36421 , \36422 , \36423 , \36424 , \36425 , \36426 ,
         \36427 , \36428 , \36429 , \36430 , \36431 , \36432 , \36433 , \36434 , \36435 , \36436 ,
         \36437 , \36438 , \36439 , \36440 , \36441 , \36442 , \36443 , \36444 , \36445 , \36446 ,
         \36447 , \36448 , \36449 , \36450 , \36451 , \36452 , \36453 , \36454 , \36455 , \36456 ,
         \36457 , \36458 , \36459 , \36460 , \36461 , \36462 , \36463 , \36464 , \36465 , \36466 ,
         \36467 , \36468 , \36469 , \36470 , \36471 , \36472 , \36473 , \36474 , \36475 , \36476 ,
         \36477 , \36478 , \36479 , \36480 , \36481 , \36482 , \36483 , \36484 , \36485 , \36486 ,
         \36487 , \36488 , \36489 , \36490 , \36491 , \36492 , \36493 , \36494 , \36495 , \36496 ,
         \36497 , \36498 , \36499 , \36500 , \36501 , \36502 , \36503 , \36504 , \36505 , \36506 ,
         \36507 , \36508 , \36509 , \36510 , \36511 , \36512 , \36513 , \36514 , \36515 , \36516 ,
         \36517 , \36518 , \36519 , \36520 , \36521 , \36522 , \36523 , \36524 , \36525 , \36526 ,
         \36527 , \36528 , \36529 , \36530 , \36531 , \36532 , \36533 , \36534 , \36535 , \36536 ,
         \36537 , \36538 , \36539 , \36540 , \36541 , \36542 , \36543 , \36544 , \36545 , \36546 ,
         \36547 , \36548 , \36549 , \36550 , \36551 , \36552 , \36553 , \36554 , \36555 , \36556 ,
         \36557 , \36558 , \36559 , \36560 , \36561 , \36562 , \36563 , \36564 , \36565 , \36566 ,
         \36567 , \36568 , \36569 , \36570 , \36571 , \36572 , \36573 , \36574 , \36575 , \36576 ,
         \36577 , \36578 , \36579 , \36580 , \36581 , \36582 , \36583 , \36584 , \36585 , \36586 ,
         \36587 , \36588 , \36589_nG9b93 , \36590 , \36591 , \36592 , \36593 , \36594 , \36595 , \36596 ,
         \36597 , \36598 , \36599 , \36600 , \36601 , \36602 , \36603 , \36604 , \36605 , \36606 ,
         \36607 , \36608 , \36609 , \36610 , \36611 , \36612 , \36613 , \36614 , \36615 , \36616 ,
         \36617 , \36618 , \36619 , \36620 , \36621 , \36622 , \36623 , \36624 , \36625 , \36626 ,
         \36627 , \36628 , \36629 , \36630 , \36631 , \36632 , \36633 , \36634 , \36635 , \36636 ,
         \36637 , \36638 , \36639 , \36640 , \36641 , \36642 , \36643 , \36644 , \36645 , \36646 ,
         \36647 , \36648 , \36649 , \36650 , \36651 , \36652 , \36653 , \36654 , \36655 , \36656 ,
         \36657 , \36658 , \36659 , \36660 , \36661 , \36662 , \36663 , \36664 , \36665 , \36666 ,
         \36667 , \36668 , \36669 , \36670 , \36671 , \36672 , \36673 , \36674 , \36675 , \36676 ,
         \36677 , \36678 , \36679 , \36680 , \36681 , \36682 , \36683 , \36684 , \36685 , \36686 ,
         \36687 , \36688 , \36689 , \36690 , \36691 , \36692 , \36693 , \36694 , \36695 , \36696 ,
         \36697 , \36698 , \36699 , \36700 , \36701 , \36702 , \36703 , \36704 , \36705 , \36706 ,
         \36707 , \36708 , \36709 , \36710 , \36711 , \36712 , \36713 , \36714 , \36715 , \36716 ,
         \36717 , \36718 , \36719 , \36720 , \36721 , \36722 , \36723 , \36724 , \36725 , \36726 ,
         \36727 , \36728 , \36729 , \36730 , \36731 , \36732 , \36733 , \36734 , \36735 , \36736 ,
         \36737 , \36738 , \36739 , \36740 , \36741 , \36742 , \36743 , \36744 , \36745 , \36746 ,
         \36747 , \36748 , \36749 , \36750 , \36751 , \36752 , \36753 , \36754 , \36755 , \36756 ,
         \36757 , \36758 , \36759 , \36760 , \36761 , \36762 , \36763 , \36764 , \36765 , \36766 ,
         \36767 , \36768 , \36769 , \36770 , \36771 , \36772 , \36773 , \36774 , \36775 , \36776 ,
         \36777 , \36778 , \36779 , \36780 , \36781 , \36782 , \36783 , \36784 , \36785 , \36786 ,
         \36787 , \36788 , \36789 , \36790 , \36791 , \36792 , \36793 , \36794 , \36795 , \36796 ,
         \36797 , \36798 , \36799 , \36800 , \36801 , \36802 , \36803 , \36804 , \36805 , \36806 ,
         \36807 , \36808 , \36809 , \36810 , \36811 , \36812 , \36813 , \36814 , \36815 , \36816 ,
         \36817 , \36818 , \36819 , \36820 , \36821 , \36822 , \36823 , \36824 , \36825 , \36826 ,
         \36827 , \36828 , \36829 , \36830 , \36831 , \36832 , \36833 , \36834 , \36835 , \36836 ,
         \36837 , \36838 , \36839 , \36840 , \36841 , \36842 , \36843 , \36844 , \36845 , \36846 ,
         \36847 , \36848 , \36849 , \36850 , \36851 , \36852 , \36853 , \36854 , \36855 , \36856 ,
         \36857 , \36858 , \36859 , \36860 , \36861 , \36862 , \36863 , \36864 , \36865 , \36866 ,
         \36867 , \36868 , \36869 , \36870 , \36871 , \36872 , \36873 , \36874 , \36875 , \36876 ,
         \36877 , \36878 , \36879 , \36880 , \36881 , \36882 , \36883 , \36884 , \36885 , \36886 ,
         \36887 , \36888 , \36889 , \36890 , \36891 , \36892 , \36893 , \36894 , \36895 , \36896 ,
         \36897 , \36898 , \36899 , \36900 , \36901 , \36902 , \36903 , \36904 , \36905 , \36906 ,
         \36907 , \36908 , \36909 , \36910 , \36911 , \36912 , \36913 , \36914 , \36915 , \36916 ,
         \36917 , \36918 , \36919 , \36920 , \36921 , \36922 , \36923 , \36924 , \36925 , \36926 ,
         \36927 , \36928 , \36929 , \36930 , \36931 , \36932 , \36933 , \36934 , \36935 , \36936 ,
         \36937 , \36938 , \36939 , \36940 , \36941 , \36942 , \36943 , \36944 , \36945 , \36946 ,
         \36947 , \36948 , \36949 , \36950 , \36951 , \36952 , \36953 , \36954 , \36955 , \36956 ,
         \36957 , \36958 , \36959 , \36960 , \36961 , \36962 , \36963 , \36964 , \36965 , \36966 ,
         \36967 , \36968 , \36969 , \36970 , \36971 , \36972 , \36973 , \36974 , \36975 , \36976 ,
         \36977 , \36978 , \36979 , \36980 , \36981 , \36982 , \36983 , \36984 , \36985 , \36986_nG9b90 ,
         \36987 , \36988 , \36989 , \36990 , \36991 , \36992 , \36993 , \36994 , \36995 , \36996 ,
         \36997 , \36998 , \36999 , \37000 , \37001 , \37002 , \37003 , \37004 , \37005 , \37006 ,
         \37007 , \37008 , \37009 , \37010 , \37011 , \37012 , \37013 , \37014 , \37015 , \37016 ,
         \37017 , \37018 , \37019 , \37020 , \37021 , \37022 , \37023 , \37024 , \37025 , \37026 ,
         \37027 , \37028 , \37029 , \37030 , \37031 , \37032 , \37033 , \37034 , \37035 , \37036 ,
         \37037 , \37038 , \37039 , \37040 , \37041 , \37042 , \37043 , \37044 , \37045 , \37046 ,
         \37047 , \37048 , \37049 , \37050 , \37051 , \37052 , \37053 , \37054 , \37055 , \37056 ,
         \37057 , \37058 , \37059 , \37060 , \37061 , \37062 , \37063 , \37064 , \37065 , \37066 ,
         \37067 , \37068 , \37069 , \37070 , \37071 , \37072 , \37073 , \37074 , \37075 , \37076 ,
         \37077 , \37078 , \37079 , \37080 , \37081 , \37082 , \37083 , \37084 , \37085 , \37086 ,
         \37087 , \37088 , \37089 , \37090 , \37091 , \37092 , \37093 , \37094 , \37095 , \37096 ,
         \37097 , \37098 , \37099 , \37100 , \37101 , \37102 , \37103 , \37104 , \37105 , \37106 ,
         \37107 , \37108 , \37109 , \37110 , \37111 , \37112 , \37113 , \37114 , \37115 , \37116 ,
         \37117 , \37118 , \37119 , \37120 , \37121 , \37122 , \37123 , \37124 , \37125 , \37126 ,
         \37127 , \37128 , \37129 , \37130 , \37131 , \37132 , \37133 , \37134 , \37135 , \37136 ,
         \37137 , \37138 , \37139 , \37140 , \37141 , \37142 , \37143 , \37144 , \37145 , \37146 ,
         \37147 , \37148 , \37149 , \37150 , \37151 , \37152 , \37153 , \37154 , \37155 , \37156 ,
         \37157 , \37158 , \37159 , \37160 , \37161 , \37162 , \37163 , \37164 , \37165 , \37166 ,
         \37167 , \37168 , \37169 , \37170 , \37171 , \37172 , \37173 , \37174 , \37175 , \37176 ,
         \37177 , \37178 , \37179 , \37180 , \37181 , \37182 , \37183 , \37184 , \37185 , \37186 ,
         \37187 , \37188 , \37189 , \37190 , \37191 , \37192 , \37193 , \37194 , \37195 , \37196 ,
         \37197 , \37198 , \37199 , \37200 , \37201 , \37202 , \37203 , \37204 , \37205 , \37206 ,
         \37207 , \37208 , \37209 , \37210 , \37211 , \37212 , \37213 , \37214 , \37215 , \37216 ,
         \37217 , \37218 , \37219 , \37220 , \37221 , \37222 , \37223 , \37224 , \37225 , \37226 ,
         \37227 , \37228 , \37229 , \37230 , \37231 , \37232 , \37233 , \37234 , \37235 , \37236 ,
         \37237 , \37238 , \37239 , \37240 , \37241 , \37242 , \37243 , \37244 , \37245 , \37246 ,
         \37247 , \37248 , \37249 , \37250_nG9b8d , \37251 , \37252 , \37253 , \37254 , \37255 , \37256 ,
         \37257 , \37258 , \37259 , \37260 , \37261 , \37262 , \37263 , \37264 , \37265 , \37266 ,
         \37267 , \37268 , \37269 , \37270 , \37271 , \37272 , \37273 , \37274 , \37275 , \37276 ,
         \37277 , \37278 , \37279 , \37280 , \37281 , \37282 , \37283 , \37284 , \37285 , \37286 ,
         \37287 , \37288 , \37289 , \37290 , \37291 , \37292 , \37293 , \37294 , \37295 , \37296 ,
         \37297 , \37298 , \37299 , \37300 , \37301 , \37302 , \37303 , \37304 , \37305 , \37306 ,
         \37307 , \37308 , \37309 , \37310 , \37311 , \37312 , \37313 , \37314 , \37315 , \37316 ,
         \37317 , \37318 , \37319 , \37320 , \37321 , \37322 , \37323 , \37324 , \37325 , \37326 ,
         \37327 , \37328 , \37329 , \37330 , \37331 , \37332 , \37333 , \37334 , \37335 , \37336 ,
         \37337 , \37338 , \37339 , \37340 , \37341 , \37342 , \37343 , \37344 , \37345 , \37346 ,
         \37347 , \37348 , \37349 , \37350 , \37351 , \37352 , \37353 , \37354 , \37355 , \37356 ,
         \37357 , \37358 , \37359 , \37360 , \37361 , \37362 , \37363 , \37364 , \37365 , \37366 ,
         \37367 , \37368 , \37369 , \37370 , \37371 , \37372 , \37373 , \37374 , \37375 , \37376 ,
         \37377 , \37378 , \37379 , \37380 , \37381 , \37382 , \37383 , \37384 , \37385 , \37386 ,
         \37387 , \37388 , \37389 , \37390 , \37391 , \37392 , \37393 , \37394 , \37395 , \37396 ,
         \37397 , \37398 , \37399 , \37400 , \37401 , \37402 , \37403 , \37404 , \37405 , \37406 ,
         \37407 , \37408 , \37409 , \37410 , \37411 , \37412 , \37413 , \37414 , \37415 , \37416 ,
         \37417 , \37418 , \37419 , \37420 , \37421 , \37422 , \37423 , \37424 , \37425 , \37426 ,
         \37427 , \37428 , \37429 , \37430 , \37431 , \37432 , \37433 , \37434 , \37435 , \37436 ,
         \37437 , \37438 , \37439 , \37440 , \37441 , \37442 , \37443 , \37444 , \37445 , \37446 ,
         \37447 , \37448 , \37449 , \37450 , \37451 , \37452 , \37453 , \37454 , \37455 , \37456 ,
         \37457 , \37458 , \37459 , \37460 , \37461 , \37462 , \37463 , \37464 , \37465 , \37466 ,
         \37467 , \37468 , \37469 , \37470 , \37471 , \37472 , \37473 , \37474 , \37475 , \37476 ,
         \37477 , \37478 , \37479 , \37480 , \37481 , \37482 , \37483 , \37484 , \37485 , \37486 ,
         \37487 , \37488 , \37489 , \37490 , \37491 , \37492 , \37493 , \37494 , \37495 , \37496 ,
         \37497 , \37498 , \37499 , \37500 , \37501 , \37502 , \37503 , \37504 , \37505 , \37506 ,
         \37507 , \37508 , \37509 , \37510 , \37511 , \37512 , \37513 , \37514 , \37515 , \37516 ,
         \37517 , \37518 , \37519 , \37520 , \37521 , \37522 , \37523 , \37524 , \37525 , \37526 ,
         \37527 , \37528 , \37529 , \37530 , \37531 , \37532 , \37533 , \37534 , \37535 , \37536 ,
         \37537 , \37538 , \37539 , \37540 , \37541 , \37542 , \37543 , \37544 , \37545 , \37546 ,
         \37547 , \37548 , \37549 , \37550 , \37551 , \37552 , \37553 , \37554 , \37555 , \37556 ,
         \37557 , \37558 , \37559 , \37560 , \37561 , \37562 , \37563 , \37564 , \37565 , \37566 ,
         \37567 , \37568 , \37569 , \37570 , \37571 , \37572 , \37573 , \37574 , \37575 , \37576 ,
         \37577 , \37578 , \37579 , \37580 , \37581 , \37582 , \37583 , \37584 , \37585 , \37586 ,
         \37587 , \37588 , \37589 , \37590 , \37591 , \37592 , \37593 , \37594 , \37595 , \37596 ,
         \37597 , \37598 , \37599 , \37600 , \37601 , \37602 , \37603 , \37604 , \37605 , \37606 ,
         \37607_nG9b8a , \37608 , \37609 , \37610 , \37611 , \37612 , \37613 , \37614 , \37615 , \37616 ,
         \37617 , \37618 , \37619 , \37620 , \37621 , \37622 , \37623 , \37624 , \37625 , \37626 ,
         \37627 , \37628 , \37629 , \37630 , \37631 , \37632 , \37633 , \37634 , \37635 , \37636 ,
         \37637 , \37638 , \37639 , \37640 , \37641 , \37642 , \37643 , \37644 , \37645 , \37646 ,
         \37647 , \37648 , \37649 , \37650 , \37651 , \37652 , \37653 , \37654 , \37655 , \37656 ,
         \37657 , \37658 , \37659 , \37660 , \37661 , \37662 , \37663 , \37664 , \37665 , \37666 ,
         \37667 , \37668 , \37669 , \37670 , \37671 , \37672 , \37673 , \37674 , \37675 , \37676 ,
         \37677 , \37678 , \37679 , \37680 , \37681 , \37682 , \37683 , \37684 , \37685 , \37686 ,
         \37687 , \37688 , \37689 , \37690 , \37691 , \37692 , \37693 , \37694 , \37695 , \37696 ,
         \37697 , \37698 , \37699 , \37700 , \37701 , \37702 , \37703 , \37704 , \37705 , \37706 ,
         \37707 , \37708 , \37709 , \37710 , \37711 , \37712 , \37713 , \37714 , \37715 , \37716 ,
         \37717 , \37718 , \37719 , \37720 , \37721 , \37722 , \37723 , \37724 , \37725 , \37726 ,
         \37727 , \37728 , \37729 , \37730 , \37731 , \37732 , \37733 , \37734 , \37735 , \37736 ,
         \37737 , \37738 , \37739 , \37740 , \37741 , \37742 , \37743 , \37744 , \37745 , \37746 ,
         \37747 , \37748 , \37749 , \37750 , \37751 , \37752 , \37753 , \37754 , \37755 , \37756 ,
         \37757 , \37758 , \37759 , \37760 , \37761 , \37762 , \37763 , \37764 , \37765 , \37766 ,
         \37767 , \37768 , \37769 , \37770 , \37771 , \37772 , \37773 , \37774 , \37775 , \37776 ,
         \37777 , \37778 , \37779 , \37780 , \37781 , \37782 , \37783 , \37784 , \37785 , \37786 ,
         \37787 , \37788 , \37789 , \37790 , \37791 , \37792 , \37793 , \37794 , \37795 , \37796 ,
         \37797 , \37798 , \37799 , \37800 , \37801 , \37802 , \37803 , \37804 , \37805 , \37806 ,
         \37807 , \37808 , \37809 , \37810 , \37811 , \37812 , \37813 , \37814 , \37815 , \37816 ,
         \37817 , \37818 , \37819 , \37820 , \37821 , \37822 , \37823 , \37824 , \37825 , \37826 ,
         \37827 , \37828 , \37829 , \37830 , \37831 , \37832 , \37833 , \37834 , \37835 , \37836 ,
         \37837 , \37838 , \37839 , \37840 , \37841 , \37842 , \37843 , \37844 , \37845 , \37846 ,
         \37847 , \37848 , \37849 , \37850 , \37851 , \37852 , \37853 , \37854 , \37855 , \37856 ,
         \37857 , \37858 , \37859 , \37860 , \37861 , \37862 , \37863 , \37864 , \37865 , \37866 ,
         \37867 , \37868 , \37869 , \37870 , \37871 , \37872 , \37873 , \37874 , \37875 , \37876 ,
         \37877 , \37878 , \37879 , \37880 , \37881 , \37882 , \37883 , \37884 , \37885 , \37886 ,
         \37887 , \37888 , \37889 , \37890 , \37891 , \37892 , \37893 , \37894 , \37895 , \37896 ,
         \37897 , \37898 , \37899 , \37900 , \37901 , \37902 , \37903 , \37904 , \37905 , \37906 ,
         \37907 , \37908 , \37909 , \37910 , \37911 , \37912 , \37913 , \37914 , \37915 , \37916 ,
         \37917 , \37918 , \37919 , \37920 , \37921 , \37922 , \37923 , \37924 , \37925 , \37926 ,
         \37927 , \37928 , \37929 , \37930 , \37931 , \37932 , \37933 , \37934 , \37935 , \37936 ,
         \37937 , \37938 , \37939 , \37940 , \37941 , \37942 , \37943 , \37944 , \37945 , \37946 ,
         \37947 , \37948 , \37949 , \37950 , \37951 , \37952 , \37953 , \37954 , \37955 , \37956 ,
         \37957 , \37958 , \37959 , \37960 , \37961 , \37962 , \37963 , \37964 , \37965 , \37966 ,
         \37967 , \37968 , \37969 , \37970 , \37971 , \37972 , \37973 , \37974_nG9b87 , \37975 , \37976 ,
         \37977 , \37978 , \37979 , \37980 , \37981 , \37982 , \37983 , \37984 , \37985 , \37986 ,
         \37987 , \37988 , \37989 , \37990 , \37991 , \37992 , \37993 , \37994 , \37995 , \37996 ,
         \37997 , \37998 , \37999 , \38000 , \38001 , \38002 , \38003 , \38004 , \38005 , \38006 ,
         \38007 , \38008 , \38009 , \38010 , \38011 , \38012 , \38013 , \38014 , \38015 , \38016 ,
         \38017 , \38018 , \38019 , \38020 , \38021 , \38022 , \38023 , \38024 , \38025 , \38026 ,
         \38027 , \38028 , \38029 , \38030 , \38031 , \38032 , \38033 , \38034 , \38035 , \38036 ,
         \38037 , \38038 , \38039 , \38040 , \38041 , \38042 , \38043 , \38044 , \38045 , \38046 ,
         \38047 , \38048 , \38049 , \38050 , \38051 , \38052 , \38053 , \38054 , \38055 , \38056 ,
         \38057 , \38058 , \38059 , \38060 , \38061 , \38062 , \38063 , \38064 , \38065 , \38066 ,
         \38067 , \38068 , \38069 , \38070 , \38071 , \38072 , \38073 , \38074 , \38075 , \38076 ,
         \38077 , \38078 , \38079 , \38080 , \38081 , \38082 , \38083 , \38084 , \38085 , \38086 ,
         \38087 , \38088 , \38089 , \38090 , \38091 , \38092 , \38093 , \38094 , \38095 , \38096 ,
         \38097 , \38098 , \38099 , \38100 , \38101 , \38102 , \38103 , \38104 , \38105 , \38106 ,
         \38107 , \38108 , \38109 , \38110 , \38111 , \38112 , \38113 , \38114 , \38115 , \38116 ,
         \38117 , \38118 , \38119 , \38120 , \38121 , \38122 , \38123 , \38124 , \38125 , \38126 ,
         \38127 , \38128 , \38129 , \38130 , \38131 , \38132 , \38133 , \38134 , \38135 , \38136 ,
         \38137 , \38138 , \38139 , \38140 , \38141 , \38142 , \38143 , \38144 , \38145 , \38146 ,
         \38147 , \38148 , \38149 , \38150 , \38151 , \38152 , \38153 , \38154 , \38155 , \38156 ,
         \38157 , \38158 , \38159 , \38160 , \38161 , \38162 , \38163 , \38164 , \38165 , \38166 ,
         \38167 , \38168 , \38169 , \38170 , \38171 , \38172 , \38173 , \38174 , \38175 , \38176 ,
         \38177 , \38178 , \38179 , \38180 , \38181 , \38182 , \38183 , \38184 , \38185 , \38186 ,
         \38187 , \38188 , \38189 , \38190 , \38191 , \38192 , \38193 , \38194 , \38195 , \38196 ,
         \38197 , \38198 , \38199 , \38200 , \38201 , \38202 , \38203 , \38204 , \38205 , \38206 ,
         \38207 , \38208 , \38209 , \38210 , \38211 , \38212 , \38213 , \38214 , \38215 , \38216 ,
         \38217 , \38218 , \38219 , \38220 , \38221 , \38222 , \38223 , \38224 , \38225 , \38226 ,
         \38227 , \38228 , \38229 , \38230 , \38231 , \38232 , \38233 , \38234 , \38235 , \38236 ,
         \38237 , \38238 , \38239 , \38240 , \38241 , \38242 , \38243 , \38244 , \38245 , \38246 ,
         \38247 , \38248 , \38249 , \38250 , \38251 , \38252 , \38253 , \38254 , \38255 , \38256 ,
         \38257 , \38258 , \38259 , \38260 , \38261 , \38262 , \38263 , \38264 , \38265 , \38266 ,
         \38267 , \38268 , \38269 , \38270 , \38271 , \38272 , \38273 , \38274 , \38275 , \38276 ,
         \38277 , \38278 , \38279 , \38280 , \38281 , \38282 , \38283 , \38284 , \38285 , \38286 ,
         \38287 , \38288 , \38289 , \38290 , \38291 , \38292 , \38293 , \38294 , \38295 , \38296 ,
         \38297 , \38298 , \38299 , \38300 , \38301 , \38302 , \38303 , \38304 , \38305 , \38306 ,
         \38307 , \38308 , \38309 , \38310 , \38311 , \38312 , \38313 , \38314 , \38315 , \38316 ,
         \38317 , \38318 , \38319 , \38320 , \38321 , \38322 , \38323 , \38324 , \38325 , \38326 ,
         \38327 , \38328 , \38329 , \38330 , \38331 , \38332 , \38333 , \38334 , \38335 , \38336 ,
         \38337_nG9b84 , \38338 , \38339 , \38340 , \38341 , \38342 , \38343 , \38344 , \38345 , \38346 ,
         \38347 , \38348 , \38349 , \38350 , \38351 , \38352 , \38353 , \38354 , \38355 , \38356 ,
         \38357 , \38358 , \38359 , \38360 , \38361 , \38362 , \38363 , \38364 , \38365 , \38366 ,
         \38367 , \38368 , \38369 , \38370 , \38371 , \38372 , \38373 , \38374 , \38375 , \38376 ,
         \38377 , \38378 , \38379 , \38380 , \38381 , \38382 , \38383 , \38384 , \38385 , \38386 ,
         \38387 , \38388 , \38389 , \38390 , \38391 , \38392 , \38393 , \38394 , \38395 , \38396 ,
         \38397 , \38398 , \38399 , \38400 , \38401 , \38402 , \38403 , \38404 , \38405 , \38406 ,
         \38407 , \38408 , \38409 , \38410 , \38411 , \38412 , \38413 , \38414 , \38415 , \38416 ,
         \38417 , \38418 , \38419 , \38420 , \38421 , \38422 , \38423 , \38424 , \38425 , \38426 ,
         \38427 , \38428 , \38429 , \38430 , \38431 , \38432 , \38433 , \38434 , \38435 , \38436 ,
         \38437 , \38438 , \38439 , \38440 , \38441 , \38442 , \38443 , \38444 , \38445 , \38446 ,
         \38447 , \38448 , \38449 , \38450 , \38451 , \38452 , \38453 , \38454 , \38455 , \38456 ,
         \38457 , \38458 , \38459 , \38460 , \38461 , \38462 , \38463 , \38464 , \38465 , \38466 ,
         \38467 , \38468 , \38469 , \38470 , \38471 , \38472 , \38473 , \38474 , \38475 , \38476 ,
         \38477 , \38478 , \38479 , \38480 , \38481 , \38482 , \38483 , \38484 , \38485 , \38486 ,
         \38487 , \38488 , \38489 , \38490 , \38491 , \38492 , \38493 , \38494 , \38495 , \38496 ,
         \38497 , \38498 , \38499 , \38500 , \38501 , \38502 , \38503 , \38504 , \38505 , \38506 ,
         \38507 , \38508 , \38509 , \38510 , \38511 , \38512 , \38513 , \38514 , \38515 , \38516 ,
         \38517 , \38518 , \38519 , \38520 , \38521 , \38522 , \38523 , \38524 , \38525 , \38526 ,
         \38527 , \38528 , \38529 , \38530 , \38531 , \38532 , \38533 , \38534 , \38535 , \38536 ,
         \38537 , \38538 , \38539 , \38540 , \38541 , \38542 , \38543 , \38544 , \38545 , \38546 ,
         \38547 , \38548 , \38549 , \38550 , \38551 , \38552 , \38553 , \38554 , \38555 , \38556 ,
         \38557 , \38558 , \38559 , \38560 , \38561 , \38562 , \38563 , \38564 , \38565 , \38566 ,
         \38567 , \38568 , \38569 , \38570 , \38571 , \38572 , \38573 , \38574 , \38575 , \38576 ,
         \38577 , \38578 , \38579 , \38580 , \38581 , \38582 , \38583 , \38584 , \38585 , \38586 ,
         \38587 , \38588 , \38589 , \38590 , \38591 , \38592 , \38593 , \38594 , \38595 , \38596 ,
         \38597 , \38598 , \38599 , \38600 , \38601 , \38602 , \38603 , \38604 , \38605 , \38606 ,
         \38607 , \38608 , \38609 , \38610 , \38611 , \38612 , \38613 , \38614 , \38615 , \38616 ,
         \38617 , \38618 , \38619 , \38620 , \38621 , \38622 , \38623 , \38624 , \38625 , \38626 ,
         \38627 , \38628 , \38629 , \38630 , \38631 , \38632 , \38633 , \38634 , \38635 , \38636 ,
         \38637 , \38638 , \38639 , \38640 , \38641 , \38642 , \38643 , \38644 , \38645 , \38646 ,
         \38647 , \38648 , \38649 , \38650 , \38651 , \38652 , \38653 , \38654 , \38655 , \38656 ,
         \38657 , \38658 , \38659 , \38660 , \38661 , \38662 , \38663_nG9b81 , \38664 , \38665 , \38666 ,
         \38667 , \38668 , \38669 , \38670 , \38671 , \38672 , \38673 , \38674 , \38675 , \38676 ,
         \38677 , \38678 , \38679 , \38680 , \38681 , \38682 , \38683 , \38684 , \38685 , \38686 ,
         \38687 , \38688 , \38689 , \38690 , \38691 , \38692 , \38693 , \38694 , \38695 , \38696 ,
         \38697 , \38698 , \38699 , \38700 , \38701 , \38702 , \38703 , \38704 , \38705 , \38706 ,
         \38707 , \38708 , \38709 , \38710 , \38711 , \38712 , \38713 , \38714 , \38715 , \38716 ,
         \38717 , \38718 , \38719 , \38720 , \38721 , \38722 , \38723 , \38724 , \38725 , \38726 ,
         \38727 , \38728 , \38729 , \38730 , \38731 , \38732 , \38733 , \38734 , \38735 , \38736 ,
         \38737 , \38738 , \38739 , \38740 , \38741 , \38742 , \38743 , \38744 , \38745 , \38746 ,
         \38747 , \38748 , \38749 , \38750 , \38751 , \38752 , \38753 , \38754 , \38755 , \38756 ,
         \38757 , \38758 , \38759 , \38760 , \38761 , \38762 , \38763 , \38764 , \38765 , \38766 ,
         \38767 , \38768 , \38769 , \38770 , \38771 , \38772 , \38773 , \38774 , \38775 , \38776 ,
         \38777 , \38778 , \38779 , \38780 , \38781 , \38782 , \38783 , \38784 , \38785 , \38786 ,
         \38787 , \38788 , \38789 , \38790 , \38791 , \38792 , \38793 , \38794 , \38795 , \38796 ,
         \38797 , \38798 , \38799 , \38800 , \38801 , \38802 , \38803 , \38804 , \38805 , \38806 ,
         \38807 , \38808 , \38809 , \38810 , \38811 , \38812 , \38813 , \38814 , \38815 , \38816 ,
         \38817 , \38818 , \38819 , \38820 , \38821 , \38822 , \38823 , \38824 , \38825 , \38826 ,
         \38827 , \38828 , \38829 , \38830 , \38831 , \38832 , \38833 , \38834 , \38835 , \38836 ,
         \38837 , \38838 , \38839 , \38840 , \38841 , \38842 , \38843 , \38844 , \38845 , \38846 ,
         \38847 , \38848 , \38849 , \38850 , \38851 , \38852 , \38853 , \38854 , \38855 , \38856 ,
         \38857 , \38858 , \38859 , \38860 , \38861 , \38862 , \38863 , \38864 , \38865 , \38866 ,
         \38867 , \38868 , \38869 , \38870 , \38871 , \38872 , \38873 , \38874 , \38875 , \38876 ,
         \38877 , \38878 , \38879 , \38880 , \38881 , \38882 , \38883 , \38884 , \38885 , \38886 ,
         \38887 , \38888 , \38889 , \38890 , \38891 , \38892 , \38893 , \38894 , \38895 , \38896 ,
         \38897 , \38898 , \38899 , \38900 , \38901 , \38902 , \38903 , \38904 , \38905 , \38906 ,
         \38907 , \38908 , \38909 , \38910 , \38911 , \38912 , \38913 , \38914 , \38915 , \38916 ,
         \38917 , \38918 , \38919 , \38920 , \38921 , \38922 , \38923 , \38924 , \38925 , \38926 ,
         \38927 , \38928 , \38929 , \38930 , \38931 , \38932 , \38933 , \38934 , \38935 , \38936 ,
         \38937 , \38938 , \38939 , \38940 , \38941 , \38942 , \38943 , \38944 , \38945 , \38946 ,
         \38947 , \38948 , \38949 , \38950 , \38951 , \38952 , \38953 , \38954 , \38955 , \38956 ,
         \38957 , \38958 , \38959 , \38960 , \38961 , \38962 , \38963 , \38964 , \38965 , \38966 ,
         \38967 , \38968_nG9b7e , \38969 , \38970 , \38971 , \38972 , \38973 , \38974 , \38975 , \38976 ,
         \38977 , \38978 , \38979 , \38980 , \38981 , \38982 , \38983 , \38984 , \38985 , \38986 ,
         \38987 , \38988 , \38989 , \38990 , \38991 , \38992 , \38993 , \38994 , \38995 , \38996 ,
         \38997 , \38998 , \38999 , \39000 , \39001 , \39002 , \39003 , \39004 , \39005 , \39006 ,
         \39007 , \39008 , \39009 , \39010 , \39011 , \39012 , \39013 , \39014 , \39015 , \39016 ,
         \39017 , \39018 , \39019 , \39020 , \39021 , \39022 , \39023 , \39024 , \39025 , \39026 ,
         \39027 , \39028 , \39029 , \39030 , \39031 , \39032 , \39033 , \39034 , \39035 , \39036 ,
         \39037 , \39038 , \39039 , \39040 , \39041 , \39042 , \39043 , \39044 , \39045 , \39046 ,
         \39047 , \39048 , \39049 , \39050 , \39051 , \39052 , \39053 , \39054 , \39055 , \39056 ,
         \39057 , \39058 , \39059 , \39060 , \39061 , \39062 , \39063 , \39064 , \39065 , \39066 ,
         \39067 , \39068 , \39069 , \39070 , \39071 , \39072 , \39073 , \39074 , \39075 , \39076 ,
         \39077 , \39078 , \39079 , \39080 , \39081 , \39082 , \39083 , \39084 , \39085 , \39086 ,
         \39087 , \39088 , \39089 , \39090 , \39091 , \39092 , \39093 , \39094 , \39095 , \39096 ,
         \39097 , \39098 , \39099 , \39100 , \39101 , \39102 , \39103 , \39104 , \39105 , \39106 ,
         \39107 , \39108 , \39109 , \39110 , \39111 , \39112 , \39113 , \39114 , \39115 , \39116 ,
         \39117 , \39118 , \39119 , \39120 , \39121 , \39122 , \39123 , \39124 , \39125 , \39126 ,
         \39127 , \39128 , \39129 , \39130 , \39131 , \39132 , \39133 , \39134 , \39135 , \39136 ,
         \39137 , \39138 , \39139 , \39140 , \39141 , \39142 , \39143 , \39144 , \39145 , \39146 ,
         \39147 , \39148 , \39149 , \39150 , \39151 , \39152 , \39153 , \39154 , \39155 , \39156 ,
         \39157 , \39158 , \39159 , \39160 , \39161 , \39162 , \39163 , \39164 , \39165 , \39166 ,
         \39167 , \39168 , \39169 , \39170 , \39171 , \39172 , \39173 , \39174 , \39175 , \39176 ,
         \39177 , \39178 , \39179 , \39180 , \39181 , \39182 , \39183 , \39184 , \39185 , \39186 ,
         \39187 , \39188 , \39189 , \39190 , \39191 , \39192 , \39193 , \39194 , \39195 , \39196 ,
         \39197 , \39198 , \39199 , \39200 , \39201 , \39202 , \39203 , \39204 , \39205 , \39206 ,
         \39207 , \39208 , \39209 , \39210 , \39211 , \39212 , \39213 , \39214 , \39215 , \39216 ,
         \39217 , \39218 , \39219 , \39220 , \39221 , \39222 , \39223 , \39224 , \39225 , \39226 ,
         \39227 , \39228 , \39229 , \39230 , \39231 , \39232 , \39233 , \39234 , \39235 , \39236 ,
         \39237 , \39238 , \39239 , \39240 , \39241 , \39242 , \39243 , \39244 , \39245 , \39246 ,
         \39247 , \39248 , \39249 , \39250 , \39251 , \39252 , \39253 , \39254 , \39255 , \39256 ,
         \39257 , \39258 , \39259 , \39260 , \39261 , \39262 , \39263 , \39264 , \39265 , \39266 ,
         \39267 , \39268 , \39269 , \39270 , \39271 , \39272 , \39273 , \39274 , \39275 , \39276 ,
         \39277 , \39278 , \39279 , \39280 , \39281 , \39282 , \39283 , \39284 , \39285 , \39286 ,
         \39287 , \39288 , \39289 , \39290 , \39291 , \39292 , \39293 , \39294 , \39295 , \39296 ,
         \39297 , \39298 , \39299 , \39300 , \39301 , \39302 , \39303 , \39304 , \39305 , \39306 ,
         \39307 , \39308 , \39309 , \39310 , \39311 , \39312 , \39313 , \39314 , \39315 , \39316 ,
         \39317 , \39318 , \39319 , \39320 , \39321 , \39322 , \39323 , \39324 , \39325 , \39326 ,
         \39327 , \39328 , \39329 , \39330 , \39331 , \39332 , \39333 , \39334_nG9b7b , \39335 , \39336 ,
         \39337 , \39338 , \39339 , \39340 , \39341 , \39342 , \39343 , \39344 , \39345 , \39346 ,
         \39347 , \39348 , \39349 , \39350 , \39351 , \39352 , \39353 , \39354 , \39355 , \39356 ,
         \39357 , \39358 , \39359 , \39360 , \39361 , \39362 , \39363 , \39364 , \39365 , \39366 ,
         \39367 , \39368 , \39369 , \39370 , \39371 , \39372 , \39373 , \39374 , \39375 , \39376 ,
         \39377 , \39378 , \39379 , \39380 , \39381 , \39382 , \39383 , \39384 , \39385 , \39386 ,
         \39387 , \39388 , \39389 , \39390 , \39391 , \39392 , \39393 , \39394 , \39395 , \39396 ,
         \39397 , \39398 , \39399 , \39400 , \39401 , \39402 , \39403 , \39404 , \39405 , \39406 ,
         \39407 , \39408 , \39409 , \39410 , \39411 , \39412 , \39413 , \39414 , \39415 , \39416 ,
         \39417 , \39418 , \39419 , \39420 , \39421 , \39422 , \39423 , \39424 , \39425 , \39426 ,
         \39427 , \39428 , \39429 , \39430 , \39431 , \39432 , \39433 , \39434 , \39435 , \39436 ,
         \39437 , \39438 , \39439 , \39440 , \39441 , \39442 , \39443 , \39444 , \39445 , \39446 ,
         \39447 , \39448 , \39449 , \39450 , \39451 , \39452 , \39453 , \39454 , \39455 , \39456 ,
         \39457 , \39458 , \39459 , \39460 , \39461 , \39462 , \39463 , \39464 , \39465 , \39466 ,
         \39467 , \39468 , \39469 , \39470 , \39471 , \39472 , \39473 , \39474 , \39475 , \39476 ,
         \39477 , \39478 , \39479 , \39480 , \39481 , \39482 , \39483 , \39484 , \39485 , \39486 ,
         \39487 , \39488 , \39489 , \39490 , \39491 , \39492 , \39493 , \39494 , \39495 , \39496 ,
         \39497 , \39498 , \39499 , \39500 , \39501 , \39502 , \39503 , \39504 , \39505 , \39506 ,
         \39507 , \39508 , \39509 , \39510 , \39511 , \39512 , \39513 , \39514 , \39515 , \39516 ,
         \39517 , \39518 , \39519 , \39520 , \39521 , \39522 , \39523 , \39524 , \39525 , \39526 ,
         \39527 , \39528 , \39529 , \39530 , \39531 , \39532 , \39533 , \39534 , \39535 , \39536 ,
         \39537 , \39538 , \39539 , \39540 , \39541 , \39542 , \39543 , \39544 , \39545 , \39546 ,
         \39547 , \39548 , \39549 , \39550 , \39551 , \39552 , \39553 , \39554 , \39555 , \39556 ,
         \39557 , \39558 , \39559 , \39560 , \39561 , \39562 , \39563 , \39564 , \39565 , \39566 ,
         \39567 , \39568 , \39569 , \39570 , \39571 , \39572 , \39573 , \39574 , \39575 , \39576 ,
         \39577 , \39578 , \39579 , \39580 , \39581 , \39582 , \39583 , \39584 , \39585 , \39586 ,
         \39587 , \39588 , \39589 , \39590 , \39591_nG9b78 , \39592 , \39593 , \39594 , \39595 , \39596 ,
         \39597 , \39598 , \39599 , \39600 , \39601 , \39602 , \39603 , \39604 , \39605 , \39606 ,
         \39607 , \39608 , \39609 , \39610 , \39611 , \39612 , \39613 , \39614 , \39615 , \39616 ,
         \39617 , \39618 , \39619 , \39620 , \39621 , \39622 , \39623 , \39624 , \39625 , \39626 ,
         \39627 , \39628 , \39629 , \39630 , \39631 , \39632 , \39633 , \39634 , \39635 , \39636 ,
         \39637 , \39638 , \39639 , \39640 , \39641 , \39642 , \39643 , \39644 , \39645 , \39646 ,
         \39647 , \39648 , \39649 , \39650 , \39651 , \39652 , \39653 , \39654 , \39655 , \39656 ,
         \39657 , \39658 , \39659 , \39660 , \39661 , \39662 , \39663 , \39664 , \39665 , \39666 ,
         \39667 , \39668 , \39669 , \39670 , \39671 , \39672 , \39673 , \39674 , \39675 , \39676 ,
         \39677 , \39678 , \39679 , \39680 , \39681 , \39682 , \39683 , \39684 , \39685 , \39686 ,
         \39687 , \39688 , \39689 , \39690 , \39691 , \39692 , \39693 , \39694 , \39695 , \39696 ,
         \39697 , \39698 , \39699 , \39700 , \39701 , \39702 , \39703 , \39704 , \39705 , \39706 ,
         \39707 , \39708 , \39709 , \39710 , \39711 , \39712 , \39713 , \39714 , \39715 , \39716 ,
         \39717 , \39718 , \39719 , \39720 , \39721 , \39722 , \39723 , \39724 , \39725 , \39726 ,
         \39727 , \39728 , \39729 , \39730 , \39731 , \39732 , \39733 , \39734 , \39735 , \39736 ,
         \39737 , \39738 , \39739 , \39740 , \39741 , \39742 , \39743 , \39744 , \39745 , \39746 ,
         \39747 , \39748 , \39749 , \39750 , \39751 , \39752 , \39753 , \39754 , \39755 , \39756 ,
         \39757 , \39758 , \39759 , \39760 , \39761 , \39762 , \39763 , \39764 , \39765 , \39766 ,
         \39767 , \39768 , \39769 , \39770 , \39771 , \39772 , \39773 , \39774 , \39775 , \39776 ,
         \39777 , \39778 , \39779 , \39780 , \39781 , \39782 , \39783 , \39784 , \39785 , \39786 ,
         \39787 , \39788 , \39789 , \39790 , \39791 , \39792 , \39793 , \39794 , \39795 , \39796 ,
         \39797 , \39798 , \39799 , \39800 , \39801 , \39802 , \39803 , \39804 , \39805 , \39806 ,
         \39807 , \39808 , \39809 , \39810 , \39811 , \39812 , \39813 , \39814 , \39815 , \39816 ,
         \39817 , \39818 , \39819 , \39820 , \39821 , \39822 , \39823 , \39824 , \39825 , \39826 ,
         \39827 , \39828 , \39829 , \39830 , \39831 , \39832 , \39833 , \39834 , \39835 , \39836 ,
         \39837 , \39838 , \39839 , \39840 , \39841 , \39842 , \39843 , \39844 , \39845 , \39846 ,
         \39847 , \39848 , \39849 , \39850 , \39851 , \39852 , \39853 , \39854 , \39855 , \39856 ,
         \39857 , \39858 , \39859 , \39860 , \39861 , \39862 , \39863 , \39864 , \39865 , \39866 ,
         \39867 , \39868 , \39869 , \39870 , \39871 , \39872 , \39873 , \39874 , \39875 , \39876 ,
         \39877 , \39878 , \39879 , \39880 , \39881 , \39882 , \39883 , \39884 , \39885 , \39886 ,
         \39887 , \39888 , \39889 , \39890 , \39891 , \39892 , \39893 , \39894 , \39895 , \39896 ,
         \39897 , \39898 , \39899 , \39900 , \39901 , \39902 , \39903 , \39904 , \39905 , \39906 ,
         \39907 , \39908 , \39909 , \39910 , \39911 , \39912 , \39913 , \39914 , \39915 , \39916 ,
         \39917 , \39918 , \39919 , \39920 , \39921 , \39922 , \39923 , \39924 , \39925 , \39926 ,
         \39927 , \39928 , \39929 , \39930 , \39931 , \39932 , \39933 , \39934 , \39935 , \39936 ,
         \39937 , \39938 , \39939 , \39940 , \39941 , \39942 , \39943 , \39944 , \39945 , \39946 ,
         \39947 , \39948 , \39949 , \39950 , \39951 , \39952 , \39953 , \39954 , \39955 , \39956 ,
         \39957 , \39958 , \39959 , \39960 , \39961 , \39962 , \39963_nG9b75 , \39964 , \39965 , \39966 ,
         \39967 , \39968 , \39969 , \39970 , \39971 , \39972 , \39973 , \39974 , \39975 , \39976 ,
         \39977 , \39978 , \39979 , \39980 , \39981 , \39982 , \39983 , \39984 , \39985 , \39986 ,
         \39987 , \39988 , \39989 , \39990 , \39991 , \39992 , \39993 , \39994 , \39995 , \39996 ,
         \39997 , \39998 , \39999 , \40000 , \40001 , \40002 , \40003 , \40004 , \40005 , \40006 ,
         \40007 , \40008 , \40009 , \40010 , \40011 , \40012 , \40013 , \40014 , \40015 , \40016 ,
         \40017 , \40018 , \40019 , \40020 , \40021 , \40022 , \40023 , \40024 , \40025 , \40026 ,
         \40027 , \40028 , \40029 , \40030 , \40031 , \40032 , \40033 , \40034 , \40035 , \40036 ,
         \40037 , \40038 , \40039 , \40040 , \40041 , \40042 , \40043 , \40044 , \40045 , \40046 ,
         \40047 , \40048 , \40049 , \40050 , \40051 , \40052 , \40053 , \40054 , \40055 , \40056 ,
         \40057 , \40058 , \40059 , \40060 , \40061 , \40062 , \40063 , \40064 , \40065 , \40066 ,
         \40067 , \40068 , \40069 , \40070 , \40071 , \40072 , \40073 , \40074 , \40075 , \40076 ,
         \40077 , \40078 , \40079 , \40080 , \40081 , \40082 , \40083 , \40084 , \40085 , \40086 ,
         \40087 , \40088 , \40089 , \40090 , \40091 , \40092 , \40093 , \40094 , \40095 , \40096 ,
         \40097 , \40098 , \40099 , \40100 , \40101 , \40102 , \40103 , \40104 , \40105 , \40106 ,
         \40107 , \40108 , \40109 , \40110 , \40111 , \40112 , \40113 , \40114 , \40115 , \40116 ,
         \40117 , \40118 , \40119 , \40120 , \40121 , \40122 , \40123 , \40124 , \40125 , \40126 ,
         \40127 , \40128 , \40129 , \40130 , \40131 , \40132 , \40133 , \40134 , \40135 , \40136 ,
         \40137 , \40138 , \40139 , \40140 , \40141 , \40142 , \40143 , \40144 , \40145 , \40146 ,
         \40147 , \40148 , \40149 , \40150 , \40151 , \40152 , \40153 , \40154 , \40155 , \40156 ,
         \40157 , \40158 , \40159 , \40160 , \40161 , \40162 , \40163 , \40164 , \40165 , \40166 ,
         \40167 , \40168 , \40169 , \40170 , \40171 , \40172 , \40173 , \40174 , \40175 , \40176 ,
         \40177 , \40178 , \40179 , \40180 , \40181 , \40182 , \40183 , \40184 , \40185 , \40186 ,
         \40187 , \40188 , \40189 , \40190 , \40191 , \40192 , \40193 , \40194 , \40195 , \40196 ,
         \40197 , \40198 , \40199 , \40200 , \40201 , \40202 , \40203 , \40204_nG9b72 , \40205 , \40206 ,
         \40207 , \40208 , \40209 , \40210 , \40211 , \40212 , \40213 , \40214 , \40215 , \40216 ,
         \40217 , \40218 , \40219 , \40220 , \40221 , \40222 , \40223 , \40224 , \40225 , \40226 ,
         \40227 , \40228 , \40229 , \40230 , \40231 , \40232 , \40233 , \40234 , \40235 , \40236 ,
         \40237 , \40238 , \40239 , \40240 , \40241 , \40242 , \40243 , \40244 , \40245 , \40246 ,
         \40247 , \40248 , \40249 , \40250 , \40251 , \40252 , \40253 , \40254 , \40255 , \40256 ,
         \40257 , \40258 , \40259 , \40260 , \40261 , \40262 , \40263 , \40264 , \40265 , \40266 ,
         \40267 , \40268 , \40269 , \40270 , \40271 , \40272 , \40273 , \40274 , \40275 , \40276 ,
         \40277 , \40278 , \40279 , \40280 , \40281 , \40282 , \40283 , \40284 , \40285 , \40286 ,
         \40287 , \40288 , \40289 , \40290 , \40291 , \40292 , \40293 , \40294 , \40295 , \40296 ,
         \40297 , \40298 , \40299 , \40300 , \40301 , \40302 , \40303 , \40304 , \40305 , \40306 ,
         \40307 , \40308 , \40309 , \40310 , \40311 , \40312 , \40313 , \40314 , \40315 , \40316 ,
         \40317 , \40318 , \40319 , \40320 , \40321 , \40322 , \40323 , \40324 , \40325 , \40326 ,
         \40327 , \40328 , \40329 , \40330 , \40331 , \40332 , \40333 , \40334 , \40335 , \40336 ,
         \40337 , \40338 , \40339 , \40340 , \40341 , \40342 , \40343 , \40344 , \40345 , \40346 ,
         \40347 , \40348 , \40349 , \40350 , \40351 , \40352 , \40353 , \40354 , \40355 , \40356 ,
         \40357 , \40358 , \40359 , \40360 , \40361 , \40362 , \40363 , \40364 , \40365 , \40366 ,
         \40367 , \40368 , \40369 , \40370 , \40371 , \40372 , \40373 , \40374 , \40375 , \40376 ,
         \40377 , \40378 , \40379 , \40380 , \40381 , \40382 , \40383 , \40384 , \40385 , \40386 ,
         \40387 , \40388 , \40389 , \40390 , \40391 , \40392 , \40393 , \40394 , \40395 , \40396 ,
         \40397 , \40398 , \40399 , \40400 , \40401 , \40402 , \40403 , \40404 , \40405 , \40406 ,
         \40407 , \40408 , \40409 , \40410 , \40411 , \40412 , \40413 , \40414 , \40415 , \40416 ,
         \40417 , \40418 , \40419 , \40420 , \40421 , \40422 , \40423 , \40424 , \40425 , \40426 ,
         \40427 , \40428 , \40429 , \40430 , \40431 , \40432 , \40433 , \40434 , \40435 , \40436 ,
         \40437 , \40438 , \40439 , \40440 , \40441 , \40442 , \40443 , \40444 , \40445 , \40446 ,
         \40447 , \40448 , \40449 , \40450 , \40451 , \40452_nG9b6f , \40453 , \40454 , \40455 , \40456 ,
         \40457 , \40458 , \40459 , \40460 , \40461 , \40462 , \40463 , \40464 , \40465 , \40466 ,
         \40467 , \40468 , \40469 , \40470 , \40471 , \40472 , \40473 , \40474 , \40475 , \40476 ,
         \40477 , \40478 , \40479 , \40480 , \40481 , \40482 , \40483 , \40484 , \40485 , \40486 ,
         \40487 , \40488 , \40489 , \40490 , \40491 , \40492 , \40493 , \40494 , \40495 , \40496 ,
         \40497 , \40498 , \40499 , \40500 , \40501 , \40502 , \40503 , \40504 , \40505 , \40506 ,
         \40507 , \40508 , \40509 , \40510 , \40511 , \40512 , \40513 , \40514 , \40515 , \40516 ,
         \40517 , \40518 , \40519 , \40520 , \40521 , \40522 , \40523 , \40524 , \40525 , \40526 ,
         \40527 , \40528 , \40529 , \40530 , \40531 , \40532 , \40533 , \40534 , \40535 , \40536 ,
         \40537 , \40538 , \40539 , \40540 , \40541 , \40542 , \40543 , \40544 , \40545 , \40546 ,
         \40547 , \40548 , \40549 , \40550 , \40551 , \40552 , \40553 , \40554 , \40555 , \40556 ,
         \40557 , \40558 , \40559 , \40560 , \40561 , \40562 , \40563 , \40564 , \40565 , \40566 ,
         \40567 , \40568 , \40569 , \40570 , \40571 , \40572 , \40573 , \40574 , \40575 , \40576 ,
         \40577 , \40578 , \40579 , \40580 , \40581 , \40582 , \40583 , \40584 , \40585 , \40586 ,
         \40587 , \40588 , \40589 , \40590 , \40591 , \40592 , \40593 , \40594 , \40595 , \40596 ,
         \40597 , \40598 , \40599 , \40600 , \40601 , \40602 , \40603 , \40604 , \40605 , \40606 ,
         \40607 , \40608 , \40609 , \40610 , \40611 , \40612 , \40613 , \40614 , \40615 , \40616 ,
         \40617 , \40618 , \40619 , \40620 , \40621 , \40622 , \40623 , \40624 , \40625 , \40626 ,
         \40627 , \40628 , \40629 , \40630 , \40631 , \40632 , \40633 , \40634 , \40635 , \40636 ,
         \40637 , \40638 , \40639 , \40640 , \40641 , \40642 , \40643 , \40644 , \40645 , \40646 ,
         \40647 , \40648 , \40649 , \40650 , \40651 , \40652 , \40653 , \40654 , \40655 , \40656 ,
         \40657 , \40658 , \40659 , \40660 , \40661 , \40662 , \40663 , \40664 , \40665 , \40666 ,
         \40667 , \40668 , \40669 , \40670 , \40671 , \40672 , \40673 , \40674 , \40675 , \40676 ,
         \40677 , \40678 , \40679 , \40680 , \40681 , \40682 , \40683 , \40684 , \40685 , \40686 ,
         \40687 , \40688 , \40689 , \40690 , \40691 , \40692 , \40693 , \40694 , \40695 , \40696 ,
         \40697 , \40698 , \40699 , \40700 , \40701 , \40702 , \40703 , \40704 , \40705 , \40706 ,
         \40707 , \40708 , \40709 , \40710 , \40711 , \40712 , \40713 , \40714 , \40715 , \40716 ,
         \40717 , \40718 , \40719 , \40720 , \40721 , \40722 , \40723 , \40724 , \40725 , \40726 ,
         \40727 , \40728 , \40729 , \40730 , \40731 , \40732 , \40733 , \40734 , \40735 , \40736 ,
         \40737 , \40738 , \40739 , \40740 , \40741 , \40742 , \40743 , \40744 , \40745 , \40746 ,
         \40747 , \40748 , \40749 , \40750 , \40751 , \40752 , \40753 , \40754 , \40755 , \40756 ,
         \40757 , \40758 , \40759 , \40760 , \40761 , \40762 , \40763 , \40764 , \40765 , \40766 ,
         \40767 , \40768 , \40769 , \40770 , \40771 , \40772 , \40773 , \40774 , \40775 , \40776 ,
         \40777 , \40778 , \40779 , \40780 , \40781 , \40782 , \40783 , \40784 , \40785 , \40786 ,
         \40787 , \40788 , \40789 , \40790 , \40791 , \40792 , \40793 , \40794 , \40795 , \40796 ,
         \40797 , \40798 , \40799 , \40800 , \40801 , \40802 , \40803 , \40804 , \40805 , \40806 ,
         \40807 , \40808 , \40809 , \40810 , \40811 , \40812 , \40813 , \40814 , \40815 , \40816 ,
         \40817 , \40818 , \40819 , \40820 , \40821 , \40822 , \40823 , \40824 , \40825 , \40826 ,
         \40827 , \40828 , \40829 , \40830 , \40831 , \40832 , \40833 , \40834 , \40835 , \40836 ,
         \40837 , \40838 , \40839 , \40840 , \40841 , \40842 , \40843_nG9b6c , \40844 , \40845 , \40846 ,
         \40847 , \40848 , \40849 , \40850 , \40851 , \40852 , \40853 , \40854 , \40855 , \40856 ,
         \40857 , \40858 , \40859 , \40860 , \40861 , \40862 , \40863 , \40864 , \40865 , \40866 ,
         \40867 , \40868 , \40869 , \40870 , \40871 , \40872 , \40873 , \40874 , \40875 , \40876 ,
         \40877 , \40878 , \40879 , \40880 , \40881 , \40882 , \40883 , \40884 , \40885 , \40886 ,
         \40887 , \40888 , \40889 , \40890 , \40891 , \40892 , \40893 , \40894 , \40895 , \40896 ,
         \40897 , \40898 , \40899 , \40900 , \40901 , \40902 , \40903 , \40904 , \40905 , \40906 ,
         \40907 , \40908 , \40909 , \40910 , \40911 , \40912 , \40913 , \40914 , \40915 , \40916 ,
         \40917 , \40918 , \40919 , \40920 , \40921 , \40922 , \40923 , \40924 , \40925 , \40926 ,
         \40927 , \40928 , \40929 , \40930 , \40931 , \40932 , \40933 , \40934 , \40935 , \40936 ,
         \40937 , \40938 , \40939 , \40940 , \40941 , \40942 , \40943 , \40944 , \40945 , \40946 ,
         \40947 , \40948 , \40949 , \40950 , \40951 , \40952 , \40953 , \40954 , \40955 , \40956 ,
         \40957 , \40958 , \40959 , \40960 , \40961 , \40962 , \40963 , \40964 , \40965 , \40966 ,
         \40967 , \40968 , \40969 , \40970 , \40971 , \40972 , \40973 , \40974 , \40975 , \40976 ,
         \40977 , \40978 , \40979 , \40980 , \40981 , \40982 , \40983 , \40984 , \40985 , \40986 ,
         \40987 , \40988 , \40989 , \40990 , \40991 , \40992 , \40993 , \40994 , \40995 , \40996 ,
         \40997 , \40998 , \40999 , \41000 , \41001 , \41002 , \41003 , \41004 , \41005 , \41006 ,
         \41007 , \41008 , \41009 , \41010 , \41011 , \41012 , \41013 , \41014 , \41015 , \41016 ,
         \41017 , \41018 , \41019 , \41020 , \41021 , \41022 , \41023 , \41024 , \41025 , \41026 ,
         \41027 , \41028 , \41029 , \41030 , \41031 , \41032 , \41033 , \41034 , \41035 , \41036 ,
         \41037 , \41038 , \41039 , \41040_nG9b69 , \41041 , \41042 , \41043 , \41044 , \41045 , \41046 ,
         \41047 , \41048 , \41049 , \41050 , \41051 , \41052 , \41053 , \41054 , \41055 , \41056 ,
         \41057 , \41058 , \41059 , \41060 , \41061 , \41062 , \41063 , \41064 , \41065 , \41066 ,
         \41067 , \41068 , \41069 , \41070 , \41071 , \41072 , \41073 , \41074 , \41075 , \41076 ,
         \41077 , \41078 , \41079 , \41080 , \41081 , \41082 , \41083 , \41084 , \41085 , \41086 ,
         \41087 , \41088 , \41089 , \41090 , \41091 , \41092 , \41093 , \41094 , \41095 , \41096 ,
         \41097 , \41098 , \41099 , \41100 , \41101 , \41102 , \41103 , \41104 , \41105 , \41106 ,
         \41107 , \41108 , \41109 , \41110 , \41111 , \41112 , \41113 , \41114 , \41115 , \41116 ,
         \41117 , \41118 , \41119 , \41120 , \41121 , \41122 , \41123 , \41124 , \41125 , \41126 ,
         \41127 , \41128 , \41129 , \41130 , \41131 , \41132 , \41133 , \41134 , \41135 , \41136 ,
         \41137 , \41138 , \41139 , \41140 , \41141 , \41142 , \41143 , \41144 , \41145 , \41146 ,
         \41147 , \41148 , \41149 , \41150 , \41151 , \41152 , \41153 , \41154 , \41155 , \41156 ,
         \41157 , \41158 , \41159 , \41160 , \41161 , \41162 , \41163 , \41164 , \41165 , \41166 ,
         \41167 , \41168 , \41169 , \41170 , \41171 , \41172 , \41173 , \41174 , \41175 , \41176 ,
         \41177 , \41178 , \41179 , \41180 , \41181 , \41182 , \41183 , \41184 , \41185 , \41186 ,
         \41187 , \41188 , \41189 , \41190 , \41191 , \41192 , \41193 , \41194 , \41195 , \41196 ,
         \41197 , \41198 , \41199 , \41200 , \41201 , \41202 , \41203 , \41204 , \41205 , \41206 ,
         \41207 , \41208 , \41209 , \41210 , \41211 , \41212 , \41213 , \41214 , \41215 , \41216 ,
         \41217 , \41218 , \41219 , \41220 , \41221 , \41222 , \41223 , \41224 , \41225 , \41226 ,
         \41227 , \41228 , \41229 , \41230 , \41231 , \41232 , \41233 , \41234 , \41235 , \41236 ,
         \41237 , \41238 , \41239 , \41240 , \41241 , \41242 , \41243 , \41244 , \41245 , \41246 ,
         \41247 , \41248 , \41249 , \41250 , \41251 , \41252 , \41253 , \41254 , \41255 , \41256 ,
         \41257 , \41258 , \41259 , \41260 , \41261 , \41262 , \41263 , \41264 , \41265 , \41266 ,
         \41267 , \41268 , \41269 , \41270 , \41271 , \41272 , \41273 , \41274 , \41275 , \41276 ,
         \41277 , \41278 , \41279 , \41280 , \41281 , \41282 , \41283 , \41284 , \41285 , \41286 ,
         \41287 , \41288 , \41289 , \41290 , \41291 , \41292 , \41293 , \41294 , \41295 , \41296 ,
         \41297 , \41298 , \41299 , \41300 , \41301 , \41302 , \41303 , \41304 , \41305 , \41306 ,
         \41307 , \41308 , \41309 , \41310 , \41311 , \41312 , \41313 , \41314 , \41315 , \41316 ,
         \41317 , \41318 , \41319 , \41320 , \41321 , \41322 , \41323 , \41324 , \41325 , \41326 ,
         \41327 , \41328 , \41329 , \41330 , \41331 , \41332 , \41333 , \41334 , \41335 , \41336 ,
         \41337 , \41338 , \41339 , \41340 , \41341 , \41342 , \41343 , \41344 , \41345 , \41346 ,
         \41347 , \41348 , \41349 , \41350 , \41351 , \41352 , \41353 , \41354 , \41355 , \41356 ,
         \41357 , \41358 , \41359 , \41360 , \41361 , \41362 , \41363 , \41364 , \41365 , \41366 ,
         \41367 , \41368 , \41369 , \41370 , \41371 , \41372 , \41373 , \41374 , \41375 , \41376 ,
         \41377 , \41378 , \41379 , \41380 , \41381_nG9b66 , \41382 , \41383 , \41384 , \41385 , \41386 ,
         \41387 , \41388 , \41389 , \41390 , \41391 , \41392 , \41393 , \41394 , \41395 , \41396 ,
         \41397 , \41398 , \41399 , \41400 , \41401 , \41402 , \41403 , \41404 , \41405 , \41406 ,
         \41407 , \41408 , \41409 , \41410 , \41411 , \41412 , \41413 , \41414 , \41415 , \41416 ,
         \41417 , \41418 , \41419 , \41420 , \41421 , \41422 , \41423 , \41424 , \41425 , \41426 ,
         \41427 , \41428 , \41429 , \41430 , \41431 , \41432 , \41433 , \41434 , \41435 , \41436 ,
         \41437 , \41438 , \41439 , \41440 , \41441 , \41442 , \41443 , \41444 , \41445 , \41446 ,
         \41447 , \41448 , \41449 , \41450 , \41451 , \41452 , \41453 , \41454 , \41455 , \41456 ,
         \41457 , \41458 , \41459 , \41460 , \41461 , \41462 , \41463 , \41464 , \41465 , \41466 ,
         \41467 , \41468 , \41469 , \41470 , \41471 , \41472 , \41473 , \41474 , \41475 , \41476 ,
         \41477 , \41478 , \41479 , \41480 , \41481 , \41482 , \41483 , \41484 , \41485 , \41486 ,
         \41487 , \41488 , \41489 , \41490 , \41491 , \41492 , \41493 , \41494 , \41495 , \41496 ,
         \41497 , \41498 , \41499 , \41500 , \41501 , \41502 , \41503 , \41504 , \41505 , \41506 ,
         \41507 , \41508 , \41509 , \41510 , \41511 , \41512 , \41513 , \41514 , \41515 , \41516 ,
         \41517 , \41518 , \41519 , \41520 , \41521 , \41522 , \41523 , \41524 , \41525 , \41526 ,
         \41527 , \41528 , \41529 , \41530 , \41531 , \41532 , \41533 , \41534 , \41535 , \41536 ,
         \41537 , \41538 , \41539 , \41540 , \41541 , \41542 , \41543 , \41544 , \41545 , \41546 ,
         \41547 , \41548 , \41549 , \41550 , \41551 , \41552 , \41553 , \41554 , \41555 , \41556 ,
         \41557 , \41558 , \41559 , \41560 , \41561 , \41562 , \41563 , \41564 , \41565 , \41566 ,
         \41567 , \41568 , \41569 , \41570 , \41571 , \41572 , \41573 , \41574 , \41575 , \41576 ,
         \41577 , \41578 , \41579 , \41580 , \41581 , \41582 , \41583 , \41584 , \41585 , \41586 ,
         \41587 , \41588 , \41589 , \41590 , \41591 , \41592 , \41593 , \41594 , \41595 , \41596 ,
         \41597 , \41598 , \41599 , \41600 , \41601 , \41602 , \41603 , \41604 , \41605 , \41606 ,
         \41607 , \41608 , \41609 , \41610 , \41611 , \41612 , \41613 , \41614 , \41615 , \41616 ,
         \41617 , \41618 , \41619 , \41620 , \41621 , \41622 , \41623 , \41624 , \41625 , \41626 ,
         \41627 , \41628 , \41629 , \41630 , \41631 , \41632 , \41633 , \41634 , \41635 , \41636 ,
         \41637 , \41638 , \41639 , \41640 , \41641 , \41642 , \41643 , \41644 , \41645 , \41646 ,
         \41647 , \41648 , \41649 , \41650 , \41651 , \41652 , \41653 , \41654 , \41655 , \41656 ,
         \41657 , \41658 , \41659 , \41660 , \41661 , \41662 , \41663 , \41664 , \41665 , \41666 ,
         \41667 , \41668 , \41669 , \41670 , \41671 , \41672 , \41673 , \41674 , \41675 , \41676 ,
         \41677 , \41678 , \41679 , \41680 , \41681 , \41682 , \41683 , \41684 , \41685_nG9b63 , \41686 ,
         \41687 , \41688 , \41689 , \41690 , \41691 , \41692 , \41693 , \41694 , \41695 , \41696 ,
         \41697 , \41698 , \41699 , \41700 , \41701 , \41702 , \41703 , \41704 , \41705 , \41706 ,
         \41707 , \41708 , \41709 , \41710 , \41711 , \41712 , \41713 , \41714 , \41715 , \41716 ,
         \41717 , \41718 , \41719 , \41720 , \41721 , \41722 , \41723 , \41724 , \41725 , \41726 ,
         \41727 , \41728 , \41729 , \41730 , \41731 , \41732 , \41733 , \41734 , \41735 , \41736 ,
         \41737 , \41738 , \41739 , \41740 , \41741 , \41742 , \41743 , \41744 , \41745 , \41746 ,
         \41747 , \41748 , \41749 , \41750 , \41751 , \41752 , \41753 , \41754 , \41755 , \41756 ,
         \41757 , \41758 , \41759 , \41760 , \41761 , \41762 , \41763 , \41764 , \41765 , \41766 ,
         \41767 , \41768 , \41769 , \41770 , \41771 , \41772 , \41773 , \41774 , \41775 , \41776 ,
         \41777 , \41778 , \41779 , \41780 , \41781 , \41782 , \41783 , \41784 , \41785 , \41786 ,
         \41787 , \41788 , \41789 , \41790 , \41791 , \41792 , \41793 , \41794 , \41795 , \41796 ,
         \41797 , \41798 , \41799 , \41800 , \41801 , \41802 , \41803 , \41804 , \41805 , \41806 ,
         \41807 , \41808 , \41809 , \41810 , \41811 , \41812 , \41813 , \41814 , \41815 , \41816 ,
         \41817 , \41818 , \41819 , \41820 , \41821 , \41822 , \41823 , \41824 , \41825 , \41826 ,
         \41827 , \41828 , \41829 , \41830 , \41831 , \41832 , \41833 , \41834 , \41835 , \41836 ,
         \41837 , \41838 , \41839 , \41840 , \41841 , \41842 , \41843 , \41844 , \41845 , \41846 ,
         \41847 , \41848 , \41849 , \41850 , \41851 , \41852 , \41853 , \41854 , \41855 , \41856 ,
         \41857 , \41858 , \41859 , \41860 , \41861 , \41862 , \41863 , \41864 , \41865 , \41866 ,
         \41867 , \41868 , \41869 , \41870 , \41871 , \41872 , \41873 , \41874 , \41875 , \41876 ,
         \41877 , \41878 , \41879 , \41880 , \41881 , \41882 , \41883 , \41884 , \41885 , \41886 ,
         \41887 , \41888 , \41889 , \41890 , \41891 , \41892 , \41893 , \41894 , \41895 , \41896 ,
         \41897 , \41898 , \41899 , \41900 , \41901 , \41902 , \41903 , \41904 , \41905 , \41906 ,
         \41907 , \41908 , \41909 , \41910 , \41911 , \41912 , \41913 , \41914 , \41915 , \41916 ,
         \41917 , \41918 , \41919 , \41920 , \41921 , \41922 , \41923 , \41924 , \41925 , \41926 ,
         \41927 , \41928 , \41929 , \41930 , \41931 , \41932 , \41933 , \41934 , \41935 , \41936 ,
         \41937 , \41938 , \41939 , \41940 , \41941 , \41942 , \41943 , \41944 , \41945 , \41946 ,
         \41947 , \41948 , \41949 , \41950 , \41951 , \41952 , \41953 , \41954 , \41955 , \41956 ,
         \41957 , \41958 , \41959 , \41960 , \41961 , \41962 , \41963_nG9b60 , \41964 , \41965 , \41966 ,
         \41967 , \41968 , \41969 , \41970 , \41971 , \41972 , \41973 , \41974 , \41975 , \41976 ,
         \41977 , \41978 , \41979 , \41980 , \41981 , \41982 , \41983 , \41984 , \41985 , \41986 ,
         \41987 , \41988 , \41989 , \41990 , \41991 , \41992 , \41993 , \41994 , \41995 , \41996 ,
         \41997 , \41998 , \41999 , \42000 , \42001 , \42002 , \42003 , \42004 , \42005 , \42006 ,
         \42007 , \42008 , \42009 , \42010 , \42011 , \42012 , \42013 , \42014 , \42015 , \42016 ,
         \42017 , \42018 , \42019 , \42020 , \42021 , \42022 , \42023 , \42024 , \42025 , \42026 ,
         \42027 , \42028 , \42029 , \42030 , \42031 , \42032 , \42033 , \42034 , \42035 , \42036 ,
         \42037 , \42038 , \42039 , \42040 , \42041 , \42042 , \42043 , \42044 , \42045 , \42046 ,
         \42047 , \42048 , \42049 , \42050 , \42051 , \42052 , \42053 , \42054 , \42055 , \42056 ,
         \42057 , \42058 , \42059 , \42060 , \42061 , \42062 , \42063 , \42064 , \42065 , \42066 ,
         \42067 , \42068 , \42069 , \42070 , \42071 , \42072 , \42073 , \42074 , \42075 , \42076 ,
         \42077 , \42078 , \42079 , \42080 , \42081 , \42082 , \42083 , \42084 , \42085 , \42086 ,
         \42087 , \42088 , \42089 , \42090 , \42091 , \42092 , \42093 , \42094 , \42095 , \42096 ,
         \42097 , \42098 , \42099 , \42100 , \42101 , \42102 , \42103 , \42104 , \42105 , \42106 ,
         \42107 , \42108 , \42109 , \42110 , \42111 , \42112 , \42113 , \42114 , \42115 , \42116 ,
         \42117 , \42118 , \42119 , \42120 , \42121 , \42122 , \42123 , \42124 , \42125 , \42126 ,
         \42127 , \42128 , \42129 , \42130 , \42131 , \42132 , \42133 , \42134 , \42135 , \42136 ,
         \42137 , \42138 , \42139 , \42140 , \42141 , \42142 , \42143 , \42144 , \42145 , \42146 ,
         \42147 , \42148 , \42149 , \42150 , \42151 , \42152 , \42153 , \42154 , \42155 , \42156 ,
         \42157 , \42158 , \42159 , \42160 , \42161 , \42162 , \42163 , \42164 , \42165 , \42166 ,
         \42167 , \42168 , \42169 , \42170 , \42171 , \42172 , \42173 , \42174 , \42175 , \42176 ,
         \42177 , \42178 , \42179 , \42180 , \42181 , \42182 , \42183 , \42184 , \42185 , \42186 ,
         \42187 , \42188 , \42189 , \42190 , \42191 , \42192 , \42193 , \42194 , \42195 , \42196 ,
         \42197 , \42198 , \42199 , \42200 , \42201_nG9b5d , \42202 , \42203 , \42204 , \42205 , \42206 ,
         \42207 , \42208 , \42209 , \42210 , \42211 , \42212 , \42213 , \42214 , \42215 , \42216 ,
         \42217 , \42218 , \42219 , \42220 , \42221 , \42222 , \42223 , \42224 , \42225 , \42226 ,
         \42227 , \42228 , \42229 , \42230 , \42231 , \42232 , \42233 , \42234 , \42235 , \42236 ,
         \42237 , \42238 , \42239 , \42240 , \42241 , \42242 , \42243 , \42244 , \42245 , \42246 ,
         \42247 , \42248 , \42249 , \42250 , \42251 , \42252 , \42253 , \42254 , \42255 , \42256 ,
         \42257 , \42258 , \42259 , \42260 , \42261 , \42262 , \42263 , \42264 , \42265 , \42266 ,
         \42267 , \42268 , \42269 , \42270 , \42271 , \42272 , \42273 , \42274 , \42275 , \42276 ,
         \42277 , \42278 , \42279 , \42280 , \42281 , \42282 , \42283 , \42284 , \42285 , \42286 ,
         \42287 , \42288 , \42289 , \42290 , \42291 , \42292 , \42293 , \42294 , \42295 , \42296 ,
         \42297 , \42298 , \42299 , \42300 , \42301 , \42302 , \42303 , \42304 , \42305 , \42306 ,
         \42307 , \42308 , \42309 , \42310 , \42311 , \42312 , \42313 , \42314 , \42315 , \42316 ,
         \42317 , \42318 , \42319 , \42320 , \42321 , \42322 , \42323 , \42324 , \42325 , \42326 ,
         \42327 , \42328 , \42329 , \42330 , \42331 , \42332 , \42333 , \42334 , \42335 , \42336 ,
         \42337 , \42338 , \42339 , \42340 , \42341 , \42342 , \42343 , \42344 , \42345 , \42346 ,
         \42347 , \42348 , \42349 , \42350 , \42351 , \42352 , \42353 , \42354 , \42355 , \42356 ,
         \42357 , \42358 , \42359 , \42360 , \42361 , \42362 , \42363 , \42364 , \42365 , \42366 ,
         \42367 , \42368 , \42369 , \42370 , \42371 , \42372 , \42373 , \42374 , \42375 , \42376 ,
         \42377 , \42378 , \42379 , \42380 , \42381 , \42382 , \42383 , \42384 , \42385 , \42386 ,
         \42387 , \42388 , \42389 , \42390 , \42391 , \42392 , \42393 , \42394 , \42395 , \42396 ,
         \42397 , \42398 , \42399 , \42400 , \42401 , \42402 , \42403 , \42404 , \42405 , \42406 ,
         \42407 , \42408 , \42409 , \42410 , \42411 , \42412 , \42413 , \42414 , \42415 , \42416 ,
         \42417 , \42418 , \42419 , \42420 , \42421 , \42422 , \42423 , \42424 , \42425 , \42426 ,
         \42427 , \42428 , \42429 , \42430 , \42431 , \42432 , \42433_nG9b5a , \42434 , \42435 , \42436 ,
         \42437 , \42438 , \42439 , \42440 , \42441 , \42442 , \42443 , \42444 , \42445 , \42446 ,
         \42447 , \42448 , \42449 , \42450 , \42451 , \42452 , \42453 , \42454 , \42455 , \42456 ,
         \42457 , \42458 , \42459 , \42460 , \42461 , \42462 , \42463 , \42464 , \42465 , \42466 ,
         \42467 , \42468 , \42469 , \42470 , \42471 , \42472 , \42473 , \42474 , \42475 , \42476 ,
         \42477 , \42478 , \42479 , \42480 , \42481 , \42482 , \42483 , \42484 , \42485 , \42486 ,
         \42487 , \42488 , \42489 , \42490 , \42491 , \42492 , \42493 , \42494 , \42495 , \42496 ,
         \42497 , \42498 , \42499 , \42500 , \42501 , \42502 , \42503 , \42504 , \42505 , \42506 ,
         \42507 , \42508 , \42509 , \42510 , \42511 , \42512 , \42513 , \42514 , \42515 , \42516 ,
         \42517 , \42518 , \42519 , \42520 , \42521 , \42522 , \42523 , \42524 , \42525 , \42526 ,
         \42527 , \42528 , \42529 , \42530 , \42531 , \42532 , \42533 , \42534 , \42535 , \42536 ,
         \42537 , \42538 , \42539 , \42540 , \42541 , \42542 , \42543 , \42544 , \42545 , \42546 ,
         \42547 , \42548 , \42549 , \42550 , \42551 , \42552 , \42553 , \42554 , \42555 , \42556 ,
         \42557 , \42558 , \42559 , \42560 , \42561 , \42562 , \42563 , \42564 , \42565 , \42566 ,
         \42567 , \42568 , \42569 , \42570 , \42571 , \42572 , \42573 , \42574 , \42575 , \42576 ,
         \42577 , \42578 , \42579 , \42580 , \42581 , \42582 , \42583 , \42584 , \42585 , \42586 ,
         \42587 , \42588 , \42589 , \42590 , \42591 , \42592 , \42593 , \42594 , \42595 , \42596 ,
         \42597 , \42598 , \42599 , \42600 , \42601 , \42602 , \42603 , \42604 , \42605 , \42606 ,
         \42607 , \42608 , \42609 , \42610 , \42611 , \42612 , \42613 , \42614 , \42615 , \42616 ,
         \42617 , \42618 , \42619 , \42620 , \42621 , \42622 , \42623 , \42624 , \42625 , \42626 ,
         \42627 , \42628 , \42629 , \42630 , \42631 , \42632 , \42633 , \42634 , \42635 , \42636 ,
         \42637 , \42638 , \42639 , \42640 , \42641 , \42642 , \42643 , \42644 , \42645 , \42646 ,
         \42647 , \42648 , \42649 , \42650 , \42651 , \42652 , \42653 , \42654 , \42655 , \42656 ,
         \42657 , \42658 , \42659 , \42660 , \42661 , \42662 , \42663 , \42664 , \42665 , \42666 ,
         \42667 , \42668 , \42669 , \42670 , \42671 , \42672 , \42673 , \42674 , \42675 , \42676 ,
         \42677 , \42678 , \42679 , \42680 , \42681 , \42682 , \42683 , \42684 , \42685 , \42686 ,
         \42687 , \42688 , \42689 , \42690 , \42691 , \42692 , \42693 , \42694 , \42695 , \42696 ,
         \42697 , \42698 , \42699 , \42700 , \42701 , \42702 , \42703 , \42704 , \42705 , \42706 ,
         \42707 , \42708 , \42709 , \42710 , \42711 , \42712 , \42713 , \42714 , \42715 , \42716 ,
         \42717 , \42718 , \42719 , \42720 , \42721 , \42722 , \42723 , \42724 , \42725 , \42726 ,
         \42727 , \42728 , \42729 , \42730 , \42731 , \42732 , \42733 , \42734 , \42735 , \42736 ,
         \42737 , \42738 , \42739 , \42740 , \42741 , \42742 , \42743 , \42744 , \42745 , \42746 ,
         \42747 , \42748 , \42749 , \42750 , \42751 , \42752 , \42753 , \42754 , \42755 , \42756 ,
         \42757 , \42758 , \42759 , \42760 , \42761 , \42762 , \42763 , \42764 , \42765 , \42766_nG9b57 ,
         \42767 , \42768 , \42769 , \42770 , \42771 , \42772 , \42773 , \42774 , \42775 , \42776 ,
         \42777 , \42778 , \42779 , \42780 , \42781 , \42782 , \42783 , \42784 , \42785 , \42786 ,
         \42787 , \42788 , \42789 , \42790 , \42791 , \42792 , \42793 , \42794 , \42795 , \42796 ,
         \42797 , \42798 , \42799 , \42800 , \42801 , \42802 , \42803 , \42804 , \42805 , \42806 ,
         \42807 , \42808 , \42809 , \42810 , \42811 , \42812 , \42813 , \42814 , \42815 , \42816 ,
         \42817 , \42818 , \42819 , \42820 , \42821 , \42822 , \42823 , \42824 , \42825 , \42826 ,
         \42827 , \42828 , \42829 , \42830 , \42831 , \42832 , \42833 , \42834 , \42835 , \42836 ,
         \42837 , \42838 , \42839 , \42840 , \42841 , \42842 , \42843 , \42844 , \42845 , \42846 ,
         \42847 , \42848_nG9b54 , \42849 , \42850 , \42851 , \42852 , \42853 , \42854 , \42855 , \42856 ,
         \42857 , \42858 , \42859 , \42860 , \42861 , \42862 , \42863 , \42864 , \42865 , \42866 ,
         \42867 , \42868 , \42869 , \42870 , \42871 , \42872 , \42873 , \42874 , \42875 , \42876 ,
         \42877 , \42878 , \42879 , \42880 , \42881 , \42882 , \42883 , \42884 , \42885 , \42886 ,
         \42887 , \42888 , \42889 , \42890 , \42891 , \42892 , \42893 , \42894 , \42895 , \42896 ,
         \42897 , \42898 , \42899 , \42900 , \42901 , \42902 , \42903 , \42904 , \42905 , \42906 ,
         \42907 , \42908 , \42909 , \42910 , \42911 , \42912 , \42913 , \42914 , \42915 , \42916 ,
         \42917 , \42918 , \42919 , \42920 , \42921 , \42922 , \42923 , \42924 , \42925 , \42926 ,
         \42927 , \42928 , \42929 , \42930 , \42931 , \42932 , \42933 , \42934 , \42935 , \42936 ,
         \42937 , \42938 , \42939 , \42940 , \42941 , \42942 , \42943 , \42944 , \42945 , \42946 ,
         \42947 , \42948 , \42949 , \42950 , \42951 , \42952 , \42953 , \42954 , \42955 , \42956 ,
         \42957 , \42958 , \42959 , \42960 , \42961 , \42962 , \42963 , \42964 , \42965 , \42966 ,
         \42967 , \42968 , \42969 , \42970 , \42971 , \42972 , \42973 , \42974 , \42975 , \42976 ,
         \42977 , \42978 , \42979 , \42980 , \42981 , \42982 , \42983 , \42984 , \42985 , \42986 ,
         \42987 , \42988 , \42989 , \42990 , \42991 , \42992 , \42993 , \42994 , \42995 , \42996 ,
         \42997 , \42998 , \42999 , \43000 , \43001 , \43002 , \43003 , \43004 , \43005 , \43006 ,
         \43007 , \43008 , \43009 , \43010 , \43011 , \43012 , \43013 , \43014 , \43015 , \43016 ,
         \43017 , \43018 , \43019 , \43020 , \43021 , \43022 , \43023 , \43024 , \43025 , \43026 ,
         \43027 , \43028 , \43029 , \43030 , \43031 , \43032 , \43033 , \43034 , \43035 , \43036 ,
         \43037 , \43038 , \43039 , \43040 , \43041 , \43042 , \43043 , \43044 , \43045 , \43046 ,
         \43047 , \43048 , \43049 , \43050 , \43051 , \43052 , \43053 , \43054 , \43055 , \43056 ,
         \43057 , \43058 , \43059 , \43060 , \43061 , \43062 , \43063 , \43064 , \43065 , \43066 ,
         \43067 , \43068 , \43069 , \43070 , \43071 , \43072 , \43073 , \43074 , \43075 , \43076 ,
         \43077 , \43078 , \43079 , \43080 , \43081 , \43082 , \43083 , \43084 , \43085 , \43086 ,
         \43087 , \43088 , \43089 , \43090 , \43091 , \43092 , \43093 , \43094 , \43095 , \43096 ,
         \43097 , \43098 , \43099 , \43100 , \43101 , \43102 , \43103 , \43104 , \43105 , \43106 ,
         \43107 , \43108 , \43109 , \43110 , \43111 , \43112 , \43113 , \43114 , \43115 , \43116 ,
         \43117 , \43118 , \43119 , \43120 , \43121 , \43122 , \43123 , \43124 , \43125 , \43126 ,
         \43127 , \43128 , \43129 , \43130 , \43131 , \43132 , \43133 , \43134 , \43135 , \43136 ,
         \43137 , \43138 , \43139 , \43140 , \43141 , \43142 , \43143 , \43144 , \43145 , \43146 ,
         \43147 , \43148 , \43149 , \43150 , \43151 , \43152 , \43153 , \43154 , \43155 , \43156 ,
         \43157 , \43158 , \43159 , \43160 , \43161 , \43162 , \43163 , \43164 , \43165 , \43166 ,
         \43167 , \43168 , \43169 , \43170 , \43171 , \43172 , \43173 , \43174 , \43175 , \43176 ,
         \43177 , \43178 , \43179_nG9b51 , \43180 , \43181 , \43182 , \43183 , \43184 , \43185 , \43186 ,
         \43187 , \43188 , \43189 , \43190 , \43191 , \43192 , \43193 , \43194 , \43195 , \43196 ,
         \43197 , \43198 , \43199 , \43200 , \43201 , \43202 , \43203 , \43204 , \43205 , \43206 ,
         \43207 , \43208 , \43209 , \43210 , \43211 , \43212 , \43213 , \43214 , \43215 , \43216 ,
         \43217 , \43218 , \43219 , \43220 , \43221 , \43222 , \43223 , \43224 , \43225 , \43226 ,
         \43227 , \43228 , \43229 , \43230 , \43231 , \43232 , \43233 , \43234 , \43235 , \43236 ,
         \43237 , \43238 , \43239 , \43240 , \43241 , \43242 , \43243 , \43244 , \43245 , \43246 ,
         \43247 , \43248 , \43249 , \43250 , \43251 , \43252 , \43253 , \43254 , \43255 , \43256 ,
         \43257 , \43258 , \43259 , \43260 , \43261 , \43262 , \43263 , \43264 , \43265 , \43266 ,
         \43267 , \43268 , \43269 , \43270 , \43271 , \43272 , \43273 , \43274 , \43275 , \43276 ,
         \43277 , \43278 , \43279 , \43280 , \43281 , \43282 , \43283 , \43284 , \43285 , \43286 ,
         \43287 , \43288 , \43289 , \43290 , \43291 , \43292 , \43293 , \43294 , \43295 , \43296 ,
         \43297 , \43298 , \43299 , \43300 , \43301 , \43302 , \43303 , \43304 , \43305 , \43306 ,
         \43307 , \43308 , \43309 , \43310 , \43311 , \43312 , \43313 , \43314 , \43315 , \43316 ,
         \43317 , \43318 , \43319 , \43320 , \43321 , \43322 , \43323 , \43324 , \43325 , \43326 ,
         \43327 , \43328 , \43329 , \43330 , \43331 , \43332 , \43333 , \43334 , \43335 , \43336 ,
         \43337 , \43338 , \43339 , \43340 , \43341 , \43342 , \43343 , \43344 , \43345 , \43346 ,
         \43347 , \43348 , \43349 , \43350 , \43351 , \43352 , \43353 , \43354 , \43355 , \43356 ,
         \43357 , \43358 , \43359 , \43360 , \43361 , \43362 , \43363 , \43364 , \43365 , \43366 ,
         \43367 , \43368 , \43369 , \43370 , \43371 , \43372 , \43373 , \43374 , \43375 , \43376 ,
         \43377 , \43378 , \43379 , \43380 , \43381 , \43382 , \43383 , \43384 , \43385 , \43386 ,
         \43387 , \43388 , \43389 , \43390 , \43391 , \43392 , \43393 , \43394 , \43395 , \43396 ,
         \43397 , \43398 , \43399 , \43400 , \43401 , \43402 , \43403 , \43404 , \43405 , \43406 ,
         \43407 , \43408 , \43409 , \43410 , \43411 , \43412 , \43413 , \43414 , \43415 , \43416 ,
         \43417 , \43418 , \43419 , \43420 , \43421 , \43422 , \43423 , \43424 , \43425 , \43426 ,
         \43427 , \43428 , \43429 , \43430 , \43431 , \43432 , \43433 , \43434 , \43435 , \43436 ,
         \43437 , \43438 , \43439 , \43440 , \43441 , \43442 , \43443 , \43444 , \43445 , \43446 ,
         \43447 , \43448 , \43449 , \43450 , \43451 , \43452 , \43453 , \43454 , \43455 , \43456 ,
         \43457 , \43458 , \43459 , \43460 , \43461 , \43462 , \43463 , \43464 , \43465 , \43466 ,
         \43467 , \43468 , \43469 , \43470 , \43471 , \43472 , \43473 , \43474 , \43475 , \43476 ,
         \43477 , \43478 , \43479 , \43480 , \43481 , \43482 , \43483 , \43484 , \43485 , \43486 ,
         \43487 , \43488 , \43489 , \43490 , \43491 , \43492 , \43493 , \43494 , \43495 , \43496 ,
         \43497 , \43498 , \43499 , \43500 , \43501 , \43502 , \43503 , \43504 , \43505 , \43506 ,
         \43507 , \43508 , \43509 , \43510 , \43511 , \43512 , \43513 , \43514 , \43515 , \43516 ,
         \43517 , \43518 , \43519 , \43520 , \43521 , \43522 , \43523 , \43524 , \43525 , \43526 ,
         \43527 , \43528 , \43529 , \43530 , \43531 , \43532 , \43533 , \43534 , \43535 , \43536 ,
         \43537 , \43538 , \43539 , \43540 , \43541 , \43542 , \43543 , \43544 , \43545 , \43546 ,
         \43547 , \43548 , \43549 , \43550 , \43551 , \43552 , \43553 , \43554 , \43555 , \43556 ,
         \43557 , \43558 , \43559 , \43560 , \43561 , \43562 , \43563 , \43564 , \43565 , \43566 ,
         \43567 , \43568 , \43569 , \43570 , \43571 , \43572 , \43573 , \43574 , \43575 , \43576 ,
         \43577 , \43578 , \43579 , \43580 , \43581 , \43582 , \43583 , \43584 , \43585 , \43586 ,
         \43587 , \43588 , \43589 , \43590 , \43591 , \43592 , \43593 , \43594 , \43595 , \43596 ,
         \43597 , \43598 , \43599 , \43600 , \43601 , \43602 , \43603 , \43604 , \43605 , \43606 ,
         \43607 , \43608 , \43609 , \43610 , \43611 , \43612 , \43613 , \43614 , \43615 , \43616 ,
         \43617 , \43618 , \43619 , \43620 , \43621 , \43622 , \43623 , \43624 , \43625 , \43626 ,
         \43627 , \43628 , \43629 , \43630 , \43631 , \43632 , \43633 , \43634 , \43635 , \43636 ,
         \43637 , \43638 , \43639 , \43640 , \43641 , \43642 , \43643 , \43644 , \43645 , \43646 ,
         \43647 , \43648 , \43649 , \43650 , \43651 , \43652 , \43653 , \43654 , \43655 , \43656 ,
         \43657 , \43658 , \43659 , \43660 , \43661 , \43662 , \43663 , \43664 , \43665 , \43666 ,
         \43667 , \43668 , \43669 , \43670 , \43671 , \43672 , \43673 , \43674 , \43675 , \43676 ,
         \43677 , \43678 , \43679 , \43680 , \43681 , \43682 , \43683 , \43684 , \43685 , \43686 ,
         \43687 , \43688 , \43689 , \43690 , \43691 , \43692 , \43693 , \43694 , \43695 , \43696 ,
         \43697 , \43698 , \43699 , \43700 , \43701 , \43702 , \43703 , \43704 , \43705 , \43706 ,
         \43707 , \43708 , \43709 , \43710 , \43711 , \43712 , \43713 , \43714 , \43715 , \43716 ,
         \43717 , \43718 , \43719 , \43720 , \43721 , \43722 , \43723 , \43724 , \43725 , \43726 ,
         \43727 , \43728 , \43729 , \43730 , \43731 , \43732 , \43733 , \43734 , \43735 , \43736 ,
         \43737 , \43738 , \43739 , \43740 , \43741 , \43742 , \43743 , \43744 , \43745 , \43746 ,
         \43747 , \43748 , \43749 , \43750 , \43751 , \43752 , \43753 , \43754 , \43755 , \43756 ,
         \43757 , \43758 , \43759 , \43760 , \43761 , \43762 , \43763 , \43764 , \43765 , \43766 ,
         \43767 , \43768 , \43769 , \43770 , \43771 , \43772 , \43773 , \43774 , \43775 , \43776 ,
         \43777 , \43778 , \43779 , \43780 , \43781 , \43782 , \43783 , \43784 , \43785 , \43786 ,
         \43787 , \43788 , \43789 , \43790 , \43791 , \43792 , \43793 , \43794 , \43795 , \43796 ,
         \43797 , \43798 , \43799 , \43800 , \43801 , \43802 , \43803 , \43804 , \43805 , \43806 ,
         \43807 , \43808 , \43809 , \43810 , \43811 , \43812 , \43813 , \43814 , \43815 , \43816 ,
         \43817 , \43818 , \43819 , \43820 , \43821 , \43822 , \43823 , \43824 , \43825 , \43826 ,
         \43827 , \43828 , \43829 , \43830 , \43831 , \43832 , \43833 , \43834 , \43835 , \43836 ,
         \43837 , \43838 , \43839 , \43840 , \43841 , \43842 , \43843 , \43844 , \43845 , \43846 ,
         \43847 , \43848 , \43849 , \43850 , \43851 , \43852 , \43853 , \43854 , \43855 , \43856 ,
         \43857 , \43858 , \43859 , \43860 , \43861 , \43862 , \43863 , \43864 , \43865 , \43866 ,
         \43867 , \43868 , \43869 , \43870 , \43871 , \43872 , \43873 , \43874 , \43875 , \43876 ,
         \43877 , \43878 , \43879 , \43880 , \43881 , \43882 , \43883 , \43884 , \43885 , \43886 ,
         \43887 , \43888 , \43889 , \43890 , \43891 , \43892 , \43893 , \43894 , \43895 , \43896 ,
         \43897 , \43898 , \43899 , \43900 , \43901 , \43902 , \43903 , \43904 , \43905 , \43906 ,
         \43907 , \43908 , \43909 , \43910 , \43911 , \43912 , \43913 , \43914 , \43915 , \43916 ,
         \43917 , \43918 , \43919 , \43920 , \43921 , \43922 , \43923 , \43924 , \43925 , \43926 ,
         \43927 , \43928 , \43929 , \43930 , \43931 , \43932 , \43933 , \43934 , \43935 , \43936 ,
         \43937 , \43938 , \43939 , \43940 , \43941 , \43942 , \43943 , \43944 , \43945 , \43946 ,
         \43947 , \43948 , \43949 , \43950 , \43951 , \43952 , \43953 , \43954 , \43955 , \43956 ,
         \43957 , \43958 , \43959 , \43960 , \43961 , \43962 , \43963 , \43964 , \43965 , \43966 ,
         \43967 , \43968 , \43969 , \43970 , \43971 , \43972 , \43973 , \43974 , \43975 , \43976 ,
         \43977 , \43978 , \43979 , \43980 , \43981 , \43982 , \43983 , \43984 , \43985 , \43986 ,
         \43987 , \43988 , \43989 , \43990 , \43991 , \43992 , \43993 , \43994 , \43995 , \43996 ,
         \43997 , \43998 , \43999 , \44000 , \44001 , \44002 , \44003 , \44004 , \44005 , \44006 ,
         \44007 , \44008 , \44009 , \44010 , \44011 , \44012 , \44013 , \44014 , \44015 , \44016 ,
         \44017 , \44018 , \44019 , \44020 , \44021 , \44022 , \44023 , \44024 , \44025 , \44026 ,
         \44027 , \44028 , \44029 , \44030 , \44031 , \44032 , \44033 , \44034 , \44035 , \44036 ,
         \44037 , \44038 , \44039 , \44040 , \44041 , \44042 , \44043 , \44044 , \44045 , \44046 ,
         \44047 , \44048 , \44049 , \44050 , \44051 , \44052 , \44053 , \44054 , \44055 , \44056 ,
         \44057 , \44058 , \44059 , \44060 , \44061 , \44062 , \44063 , \44064 , \44065 , \44066 ,
         \44067 , \44068 , \44069 , \44070 , \44071 , \44072 , \44073 , \44074 , \44075 , \44076 ,
         \44077 , \44078 , \44079 , \44080 , \44081 , \44082 , \44083 , \44084 , \44085 , \44086 ,
         \44087 , \44088 , \44089 , \44090 , \44091 , \44092 , \44093 , \44094 , \44095 , \44096 ,
         \44097 , \44098 , \44099 , \44100 , \44101 , \44102 , \44103 , \44104 , \44105 , \44106 ,
         \44107 , \44108 , \44109 , \44110 , \44111 , \44112 , \44113 , \44114 , \44115 , \44116 ,
         \44117 , \44118 , \44119 , \44120 , \44121 , \44122 , \44123 , \44124 , \44125 , \44126 ,
         \44127 , \44128 , \44129 , \44130 , \44131 , \44132 , \44133 , \44134 , \44135 , \44136 ,
         \44137 , \44138 , \44139 , \44140 , \44141 , \44142 , \44143 , \44144 , \44145 , \44146 ,
         \44147 , \44148 , \44149 , \44150 , \44151 , \44152 , \44153 , \44154 , \44155 , \44156 ,
         \44157 , \44158 , \44159 , \44160 , \44161 , \44162 , \44163 , \44164 , \44165 , \44166 ,
         \44167 , \44168 , \44169 , \44170 , \44171 , \44172 , \44173 , \44174 , \44175 , \44176 ,
         \44177 , \44178 , \44179 , \44180 , \44181 , \44182 , \44183 , \44184 , \44185 , \44186 ,
         \44187 , \44188 , \44189 , \44190 , \44191 , \44192 , \44193 , \44194 , \44195 , \44196 ,
         \44197 , \44198 , \44199 , \44200 , \44201 , \44202 , \44203 , \44204 , \44205 , \44206 ,
         \44207 , \44208 , \44209 , \44210 , \44211 , \44212 , \44213 , \44214 , \44215 , \44216 ,
         \44217 , \44218 , \44219 , \44220 , \44221 , \44222 , \44223 , \44224 , \44225 , \44226 ,
         \44227 , \44228 , \44229 , \44230 , \44231 , \44232 , \44233 , \44234 , \44235 , \44236 ,
         \44237 , \44238 , \44239 , \44240 , \44241 , \44242 , \44243 , \44244 , \44245 , \44246 ,
         \44247 , \44248 , \44249 , \44250 , \44251 , \44252 , \44253 , \44254 , \44255 , \44256 ,
         \44257 , \44258 , \44259 , \44260 , \44261 , \44262 , \44263 , \44264 , \44265 , \44266 ,
         \44267 , \44268 , \44269 , \44270 , \44271 , \44272 , \44273 , \44274 , \44275 , \44276 ,
         \44277 , \44278 , \44279 , \44280 , \44281 , \44282 , \44283 , \44284 , \44285 , \44286 ,
         \44287 , \44288 , \44289 , \44290 , \44291 , \44292 , \44293 , \44294 , \44295 , \44296 ,
         \44297 , \44298 , \44299 , \44300 , \44301 , \44302 , \44303 , \44304 , \44305 , \44306 ,
         \44307 , \44308 , \44309 , \44310 , \44311 , \44312 , \44313 , \44314 , \44315 , \44316 ,
         \44317 , \44318 , \44319 , \44320 , \44321 , \44322 , \44323 , \44324 , \44325 , \44326 ,
         \44327 , \44328 , \44329 , \44330 , \44331 , \44332 , \44333 , \44334 , \44335 , \44336 ,
         \44337 , \44338 , \44339 , \44340 , \44341 , \44342 , \44343 , \44344 , \44345 , \44346 ,
         \44347 , \44348 , \44349 , \44350 , \44351 , \44352 , \44353 , \44354 , \44355 , \44356 ,
         \44357 , \44358 , \44359 , \44360 , \44361 , \44362 , \44363 , \44364 , \44365 , \44366 ,
         \44367 , \44368 , \44369 , \44370 , \44371 , \44372 , \44373 , \44374 , \44375 , \44376 ,
         \44377 , \44378 , \44379 , \44380 , \44381 , \44382 , \44383 , \44384 , \44385 , \44386 ,
         \44387 , \44388 , \44389 , \44390 , \44391 , \44392 , \44393 , \44394 , \44395 , \44396 ,
         \44397 , \44398 , \44399 , \44400 , \44401 , \44402 , \44403 , \44404 , \44405 , \44406 ,
         \44407 , \44408 , \44409 , \44410 , \44411 , \44412 , \44413 , \44414 , \44415 , \44416 ,
         \44417 , \44418 , \44419 , \44420 , \44421 , \44422 , \44423 , \44424 , \44425 , \44426 ,
         \44427 , \44428 , \44429 , \44430 , \44431 , \44432 , \44433 , \44434 , \44435 , \44436 ,
         \44437 , \44438 , \44439 , \44440 , \44441 , \44442 , \44443 , \44444 , \44445 , \44446 ,
         \44447 , \44448 , \44449 , \44450 , \44451 , \44452 , \44453 , \44454 , \44455 , \44456 ,
         \44457 , \44458 , \44459 , \44460 , \44461 , \44462 , \44463 , \44464 , \44465 , \44466 ,
         \44467 , \44468 , \44469 , \44470 , \44471 , \44472 , \44473 , \44474 , \44475 , \44476 ,
         \44477 , \44478 , \44479 , \44480 , \44481 , \44482 , \44483 , \44484 , \44485 , \44486 ,
         \44487 , \44488 , \44489 , \44490 , \44491 , \44492 , \44493 , \44494 , \44495 , \44496 ,
         \44497 , \44498 , \44499 , \44500 , \44501 , \44502 , \44503 , \44504 , \44505 , \44506 ,
         \44507 , \44508 , \44509 , \44510 , \44511 , \44512 , \44513 , \44514 , \44515 , \44516 ,
         \44517 , \44518 , \44519 , \44520 , \44521 , \44522 , \44523 , \44524 , \44525 , \44526 ,
         \44527 , \44528 , \44529 , \44530 , \44531 , \44532 , \44533 , \44534 , \44535 , \44536 ,
         \44537 , \44538 , \44539 , \44540 , \44541 , \44542 , \44543 , \44544 , \44545 , \44546 ,
         \44547 , \44548 , \44549 , \44550 , \44551 , \44552 , \44553 , \44554 , \44555 , \44556 ,
         \44557 , \44558 , \44559 , \44560 , \44561 , \44562 , \44563 , \44564 , \44565 , \44566 ,
         \44567 , \44568 , \44569 , \44570 , \44571 , \44572 , \44573 , \44574 , \44575 , \44576 ,
         \44577 , \44578 , \44579 , \44580 , \44581 , \44582 , \44583 , \44584 , \44585 , \44586 ,
         \44587 , \44588 , \44589 , \44590 , \44591 , \44592 , \44593 , \44594 , \44595 , \44596 ,
         \44597 , \44598 , \44599 , \44600 , \44601 , \44602 , \44603 , \44604 , \44605 , \44606 ,
         \44607 , \44608 , \44609 , \44610 , \44611 , \44612 , \44613 , \44614 , \44615 , \44616 ,
         \44617 , \44618 , \44619 , \44620 , \44621 , \44622 , \44623 , \44624 , \44625 , \44626 ,
         \44627 , \44628 , \44629 , \44630 , \44631 , \44632 , \44633 , \44634 , \44635 , \44636 ,
         \44637 , \44638 , \44639 , \44640 , \44641 , \44642 , \44643 , \44644 , \44645 , \44646 ,
         \44647 , \44648 , \44649 , \44650 , \44651 , \44652 , \44653 , \44654 , \44655 , \44656 ,
         \44657 , \44658 , \44659 , \44660 , \44661 , \44662 , \44663 , \44664 , \44665 , \44666 ,
         \44667 , \44668 , \44669 , \44670 , \44671 , \44672 , \44673 , \44674 , \44675 , \44676 ,
         \44677 , \44678 , \44679 , \44680 , \44681 , \44682 , \44683 , \44684 , \44685 , \44686 ,
         \44687 , \44688 , \44689 , \44690 , \44691 , \44692 , \44693 , \44694 , \44695 , \44696 ,
         \44697 , \44698 , \44699 , \44700 , \44701 , \44702 , \44703 , \44704 , \44705 , \44706 ,
         \44707 , \44708 , \44709 , \44710 , \44711 , \44712 , \44713 , \44714 , \44715 , \44716 ,
         \44717 , \44718 , \44719 , \44720 , \44721 , \44722 , \44723 , \44724 , \44725 , \44726 ,
         \44727 , \44728 , \44729 , \44730 , \44731 , \44732 , \44733 , \44734 , \44735 , \44736 ,
         \44737 , \44738 , \44739 , \44740 , \44741 , \44742 , \44743 , \44744 , \44745 , \44746 ,
         \44747 , \44748 , \44749 , \44750 , \44751 , \44752 , \44753 , \44754 , \44755 , \44756 ,
         \44757 , \44758 , \44759 , \44760 , \44761 , \44762 , \44763 , \44764 , \44765 , \44766 ,
         \44767 , \44768 , \44769 , \44770 , \44771 , \44772 , \44773 , \44774 , \44775 , \44776 ,
         \44777 , \44778 , \44779 , \44780 , \44781 , \44782 , \44783 , \44784 , \44785 , \44786 ,
         \44787 , \44788 , \44789 , \44790 , \44791 , \44792 , \44793 , \44794 , \44795 , \44796 ,
         \44797 , \44798 , \44799 , \44800 , \44801 , \44802 , \44803 , \44804 , \44805 , \44806 ,
         \44807 , \44808 , \44809 , \44810 , \44811 , \44812 , \44813 , \44814 , \44815 , \44816 ,
         \44817 , \44818 , \44819 , \44820 , \44821 , \44822 , \44823 , \44824 , \44825 , \44826 ,
         \44827 , \44828 , \44829 , \44830 , \44831 , \44832 , \44833 , \44834 , \44835 , \44836 ,
         \44837 , \44838 , \44839 , \44840 , \44841 , \44842 , \44843 , \44844 , \44845 , \44846 ,
         \44847 , \44848 , \44849 , \44850 , \44851 , \44852 , \44853 , \44854 , \44855 , \44856 ,
         \44857 , \44858 , \44859 , \44860 , \44861 , \44862 , \44863 , \44864 , \44865 , \44866 ,
         \44867 , \44868 , \44869 , \44870 , \44871 , \44872 , \44873 , \44874 , \44875 , \44876 ,
         \44877 , \44878 , \44879 , \44880 , \44881 , \44882 , \44883 , \44884 , \44885 , \44886 ,
         \44887 , \44888 , \44889 , \44890 , \44891 , \44892 , \44893 , \44894 , \44895 , \44896 ,
         \44897 , \44898 , \44899 , \44900 , \44901 , \44902 , \44903 , \44904 , \44905 , \44906 ,
         \44907 , \44908 , \44909 , \44910 , \44911 , \44912 , \44913 , \44914 , \44915 , \44916 ,
         \44917 , \44918 , \44919 , \44920 , \44921 , \44922 , \44923 , \44924 , \44925 , \44926 ,
         \44927 , \44928 , \44929 , \44930 , \44931 , \44932 , \44933 , \44934 , \44935 , \44936 ,
         \44937 , \44938 , \44939 , \44940 , \44941 , \44942 , \44943 , \44944 , \44945 , \44946 ,
         \44947 , \44948 , \44949 , \44950 , \44951 , \44952 , \44953 , \44954 , \44955 , \44956 ,
         \44957 , \44958 , \44959 , \44960 , \44961 , \44962 , \44963 , \44964 , \44965 , \44966 ,
         \44967 , \44968 , \44969 , \44970 , \44971 , \44972 , \44973 , \44974 , \44975 , \44976 ,
         \44977 , \44978 , \44979 , \44980 , \44981 , \44982 , \44983 , \44984 , \44985 , \44986 ,
         \44987 , \44988 , \44989 , \44990 , \44991 , \44992 , \44993 , \44994 , \44995 , \44996 ,
         \44997 , \44998 , \44999 , \45000 , \45001 , \45002 , \45003 , \45004 , \45005 , \45006 ,
         \45007 , \45008 , \45009 , \45010 , \45011 , \45012 , \45013 , \45014 , \45015 , \45016 ,
         \45017 , \45018 , \45019 , \45020 , \45021 , \45022 , \45023 , \45024 , \45025 , \45026 ,
         \45027 , \45028 , \45029 , \45030 , \45031 , \45032 , \45033 , \45034 , \45035 , \45036 ,
         \45037 , \45038 , \45039 , \45040 , \45041 , \45042 , \45043 , \45044 , \45045 , \45046 ,
         \45047 , \45048 , \45049 , \45050 , \45051 , \45052 , \45053 , \45054 , \45055 , \45056 ,
         \45057 , \45058 , \45059 , \45060 , \45061 , \45062 , \45063 , \45064 , \45065 , \45066 ,
         \45067 , \45068 , \45069 , \45070 , \45071 , \45072 , \45073 , \45074 , \45075 , \45076 ,
         \45077 , \45078 , \45079 , \45080 , \45081 , \45082 , \45083 , \45084 , \45085 , \45086 ,
         \45087 , \45088 , \45089 , \45090 , \45091 , \45092 , \45093 , \45094 , \45095 , \45096 ,
         \45097 , \45098 , \45099 , \45100 , \45101 , \45102 , \45103 , \45104 , \45105 , \45106 ,
         \45107 , \45108 , \45109 , \45110 , \45111 , \45112 , \45113 , \45114 , \45115 , \45116 ,
         \45117 , \45118 , \45119 , \45120 , \45121 , \45122 , \45123 , \45124 , \45125 , \45126 ,
         \45127 , \45128 , \45129 , \45130 , \45131 , \45132 , \45133 , \45134 , \45135 , \45136 ,
         \45137 , \45138 , \45139 , \45140 , \45141 , \45142 , \45143 , \45144 , \45145 , \45146 ,
         \45147 , \45148 , \45149 , \45150 , \45151 , \45152 , \45153 , \45154 , \45155 , \45156 ,
         \45157 , \45158 , \45159 , \45160 , \45161 , \45162 , \45163 , \45164 , \45165 , \45166 ,
         \45167 , \45168 , \45169 , \45170 , \45171 , \45172 , \45173 , \45174 , \45175 , \45176 ,
         \45177 , \45178 , \45179 , \45180 , \45181 , \45182 , \45183 , \45184 , \45185 , \45186 ,
         \45187 , \45188 , \45189 , \45190 , \45191 , \45192 , \45193 , \45194 , \45195 , \45196 ,
         \45197 , \45198 , \45199 , \45200 , \45201 , \45202 , \45203 , \45204 , \45205 , \45206 ,
         \45207 , \45208 , \45209 , \45210 , \45211 , \45212 , \45213 , \45214 , \45215 , \45216 ,
         \45217 , \45218 , \45219 , \45220 , \45221 , \45222 , \45223 , \45224 , \45225 , \45226 ,
         \45227 , \45228 , \45229 , \45230 , \45231 , \45232 , \45233 , \45234 , \45235 , \45236 ,
         \45237 , \45238 , \45239 , \45240 , \45241 , \45242 , \45243 , \45244 , \45245 , \45246 ,
         \45247 , \45248 , \45249 , \45250 , \45251 , \45252 , \45253 , \45254 , \45255 , \45256 ,
         \45257 , \45258 , \45259 , \45260 , \45261 , \45262 , \45263 , \45264 , \45265 , \45266 ,
         \45267 , \45268 , \45269 , \45270 , \45271 , \45272 , \45273 , \45274 , \45275 , \45276 ,
         \45277 , \45278 , \45279 , \45280 , \45281 , \45282 , \45283 , \45284 , \45285 , \45286 ,
         \45287 , \45288 , \45289 , \45290 , \45291 , \45292 , \45293 , \45294 , \45295 , \45296 ,
         \45297 , \45298 , \45299 , \45300 , \45301 , \45302 , \45303 , \45304 , \45305 , \45306 ,
         \45307 , \45308 , \45309 , \45310 , \45311 , \45312 , \45313 , \45314 , \45315 , \45316 ,
         \45317 , \45318 , \45319 , \45320 , \45321 , \45322 , \45323 , \45324 , \45325 , \45326 ,
         \45327 , \45328 , \45329 , \45330 , \45331 , \45332 , \45333 , \45334 , \45335 , \45336 ,
         \45337 , \45338 , \45339 , \45340 , \45341 , \45342 , \45343 , \45344 , \45345 , \45346 ,
         \45347 , \45348 , \45349 , \45350 , \45351 , \45352 , \45353 , \45354 , \45355 , \45356 ,
         \45357 , \45358 , \45359 , \45360 , \45361 , \45362 , \45363 , \45364 , \45365 , \45366 ,
         \45367 , \45368 , \45369 , \45370 , \45371 , \45372 , \45373 , \45374 , \45375 , \45376 ,
         \45377 , \45378 , \45379 , \45380 , \45381 , \45382 , \45383 , \45384 , \45385 , \45386 ,
         \45387 , \45388 , \45389 , \45390 , \45391 , \45392 , \45393 , \45394 , \45395 , \45396 ,
         \45397 , \45398 , \45399 , \45400 , \45401 , \45402 , \45403 , \45404 , \45405 , \45406 ,
         \45407 , \45408 , \45409 , \45410 , \45411 , \45412 , \45413 , \45414 , \45415 , \45416 ,
         \45417 , \45418 , \45419 , \45420 , \45421 , \45422 , \45423 , \45424 , \45425 , \45426 ,
         \45427 , \45428 , \45429 , \45430 , \45431 , \45432 , \45433 , \45434 , \45435 , \45436 ,
         \45437 , \45438 , \45439 , \45440 , \45441 , \45442 , \45443 , \45444 , \45445 , \45446 ,
         \45447 , \45448 , \45449 , \45450 , \45451 , \45452 , \45453 , \45454 , \45455 , \45456 ,
         \45457 , \45458 , \45459 , \45460 , \45461 , \45462 , \45463 , \45464 , \45465 , \45466 ,
         \45467 , \45468 , \45469 , \45470 , \45471 , \45472 , \45473 , \45474 , \45475 , \45476 ,
         \45477 , \45478 , \45479 , \45480 , \45481 , \45482 , \45483 , \45484 , \45485 , \45486 ,
         \45487 , \45488 , \45489 , \45490 , \45491 , \45492 , \45493 , \45494 , \45495 , \45496 ,
         \45497 , \45498 , \45499 , \45500 , \45501 , \45502 , \45503 , \45504 , \45505 , \45506 ,
         \45507 , \45508 , \45509 , \45510 , \45511 , \45512 , \45513 , \45514 , \45515 , \45516 ,
         \45517 , \45518 , \45519 , \45520 , \45521 , \45522 , \45523 , \45524 , \45525 , \45526 ,
         \45527 , \45528 , \45529 , \45530 , \45531 , \45532 , \45533 , \45534 , \45535 , \45536 ,
         \45537 , \45538 , \45539 , \45540 , \45541 , \45542 , \45543 , \45544 , \45545 , \45546 ,
         \45547 , \45548 , \45549 , \45550 , \45551 , \45552 , \45553 , \45554 , \45555 , \45556 ,
         \45557 , \45558 , \45559 , \45560 , \45561 , \45562 , \45563 , \45564 , \45565 , \45566 ,
         \45567 , \45568 , \45569 , \45570 , \45571 , \45572 , \45573 , \45574 , \45575 , \45576 ,
         \45577 , \45578 , \45579 , \45580 , \45581 , \45582 , \45583 , \45584 , \45585 , \45586 ,
         \45587 , \45588 , \45589 , \45590 , \45591 , \45592 , \45593 , \45594 , \45595 , \45596 ,
         \45597 , \45598 , \45599 , \45600 , \45601 , \45602 , \45603 , \45604 , \45605 , \45606 ,
         \45607 , \45608 , \45609 , \45610 , \45611 , \45612 , \45613 , \45614 , \45615 , \45616 ,
         \45617 , \45618 , \45619 , \45620 , \45621 , \45622 , \45623 , \45624 , \45625 , \45626 ,
         \45627 , \45628 , \45629 , \45630 , \45631 , \45632 , \45633 , \45634 , \45635 , \45636 ,
         \45637 , \45638 , \45639 , \45640 , \45641 , \45642 , \45643 , \45644 , \45645 , \45646 ,
         \45647 , \45648 , \45649 , \45650 , \45651 , \45652 , \45653 , \45654 , \45655 , \45656 ,
         \45657 , \45658 , \45659 , \45660 , \45661 , \45662 , \45663 , \45664 , \45665 , \45666 ,
         \45667 , \45668 , \45669 , \45670 , \45671 , \45672 , \45673 , \45674 , \45675 , \45676 ,
         \45677 , \45678 , \45679 , \45680 , \45681 , \45682 , \45683 , \45684 , \45685 , \45686 ,
         \45687 , \45688 , \45689 , \45690 , \45691 , \45692 , \45693 , \45694 , \45695 , \45696 ,
         \45697 , \45698 , \45699 , \45700 , \45701 , \45702 , \45703 , \45704 , \45705 , \45706 ,
         \45707 , \45708 , \45709 , \45710 , \45711 , \45712 , \45713 , \45714 , \45715 , \45716 ,
         \45717 , \45718 , \45719 , \45720 , \45721 , \45722 , \45723 , \45724 , \45725 , \45726 ,
         \45727 , \45728 , \45729 , \45730 , \45731 , \45732 , \45733 , \45734 , \45735 , \45736 ,
         \45737 , \45738 , \45739 , \45740 , \45741 , \45742 , \45743 , \45744 , \45745 , \45746 ,
         \45747 , \45748 , \45749 , \45750 , \45751 , \45752 , \45753 , \45754 , \45755 , \45756 ,
         \45757 , \45758 , \45759 , \45760 , \45761 , \45762 , \45763 , \45764 , \45765 , \45766 ,
         \45767 , \45768 , \45769 , \45770 , \45771 , \45772 , \45773 , \45774 , \45775 , \45776 ,
         \45777 , \45778 , \45779 , \45780 , \45781 , \45782 , \45783 , \45784 , \45785 , \45786 ,
         \45787 , \45788 , \45789 , \45790 , \45791 , \45792 , \45793 , \45794 , \45795 , \45796 ,
         \45797 , \45798 , \45799 , \45800 , \45801 , \45802 , \45803 , \45804 , \45805 , \45806 ,
         \45807 , \45808 , \45809 , \45810 , \45811 , \45812 , \45813 , \45814 , \45815 , \45816 ,
         \45817 , \45818 , \45819 , \45820 , \45821 , \45822 , \45823 , \45824 , \45825 , \45826 ,
         \45827 , \45828 , \45829 , \45830 , \45831 , \45832 , \45833 , \45834 , \45835 , \45836 ,
         \45837 , \45838 , \45839 , \45840 , \45841 , \45842 , \45843 , \45844 , \45845 , \45846 ,
         \45847 , \45848 , \45849 , \45850 , \45851 , \45852 , \45853 , \45854 , \45855 , \45856 ,
         \45857 , \45858 , \45859 , \45860 , \45861 , \45862 , \45863 , \45864 , \45865 , \45866 ,
         \45867 , \45868 , \45869 , \45870 , \45871 , \45872 , \45873 , \45874 , \45875 , \45876 ,
         \45877 , \45878 , \45879 , \45880 , \45881 , \45882 , \45883 , \45884 , \45885 , \45886 ,
         \45887 , \45888 , \45889 , \45890 , \45891 , \45892 , \45893 , \45894 , \45895 , \45896 ,
         \45897 , \45898 , \45899 , \45900 , \45901 , \45902 , \45903 , \45904 , \45905 , \45906 ,
         \45907 , \45908 , \45909 , \45910 , \45911 , \45912 , \45913 , \45914 , \45915 , \45916 ,
         \45917 , \45918 , \45919 , \45920 , \45921 , \45922 , \45923 , \45924 , \45925 , \45926 ,
         \45927 , \45928 , \45929 , \45930 , \45931 , \45932 , \45933 , \45934 , \45935 , \45936 ,
         \45937 , \45938 , \45939 , \45940 , \45941 , \45942 , \45943 , \45944 , \45945 , \45946 ,
         \45947 , \45948 , \45949 , \45950 , \45951 , \45952 , \45953 , \45954 , \45955 , \45956 ,
         \45957 , \45958 , \45959 , \45960 , \45961 , \45962 , \45963 , \45964 , \45965 , \45966 ,
         \45967 , \45968 , \45969 , \45970 , \45971 , \45972 , \45973 , \45974 , \45975 , \45976 ,
         \45977 , \45978 , \45979 , \45980 , \45981 , \45982 , \45983 , \45984 , \45985 , \45986 ,
         \45987 , \45988 , \45989 , \45990 , \45991 , \45992 , \45993 , \45994 , \45995 , \45996 ,
         \45997 , \45998 , \45999 , \46000 , \46001 , \46002 , \46003 , \46004 , \46005 , \46006 ,
         \46007 , \46008 , \46009 , \46010 , \46011 , \46012 , \46013 , \46014 , \46015 , \46016 ,
         \46017 , \46018 , \46019 , \46020 , \46021 , \46022 , \46023 , \46024 , \46025 , \46026 ,
         \46027 , \46028 , \46029 , \46030 , \46031 , \46032 , \46033 , \46034 , \46035 , \46036 ,
         \46037 , \46038 , \46039 , \46040 , \46041 , \46042 , \46043 , \46044 , \46045 , \46046 ,
         \46047 , \46048 , \46049 , \46050 , \46051 , \46052 , \46053 , \46054 , \46055 , \46056 ,
         \46057 , \46058 , \46059 , \46060 , \46061 , \46062 , \46063 , \46064 , \46065 , \46066 ,
         \46067 , \46068 , \46069 , \46070 , \46071 , \46072 , \46073 , \46074 , \46075 , \46076 ,
         \46077 , \46078 , \46079 , \46080 , \46081 , \46082 , \46083 , \46084 , \46085 , \46086 ,
         \46087 , \46088 , \46089 , \46090 , \46091 , \46092 , \46093 , \46094 , \46095 , \46096 ,
         \46097 , \46098 , \46099 , \46100 , \46101 , \46102 , \46103 , \46104 , \46105 , \46106 ,
         \46107 , \46108 , \46109 , \46110 , \46111 , \46112 , \46113 , \46114 , \46115 , \46116 ,
         \46117 , \46118 , \46119 , \46120 , \46121 , \46122 , \46123 , \46124 , \46125 , \46126 ,
         \46127 , \46128 , \46129 , \46130 , \46131 , \46132 , \46133 , \46134 , \46135 , \46136 ,
         \46137 , \46138 , \46139 , \46140 , \46141 , \46142 , \46143 , \46144 , \46145 , \46146 ,
         \46147 , \46148 , \46149 , \46150 , \46151 , \46152 , \46153 , \46154 , \46155 , \46156 ,
         \46157 , \46158 , \46159 , \46160 , \46161 , \46162 , \46163 , \46164 , \46165 , \46166 ,
         \46167 , \46168 , \46169 , \46170 , \46171 , \46172 , \46173 , \46174 , \46175 , \46176 ,
         \46177 , \46178 , \46179 , \46180 , \46181 , \46182 , \46183 , \46184 , \46185 , \46186 ,
         \46187 , \46188 , \46189 , \46190 , \46191 , \46192 , \46193 , \46194 , \46195 , \46196 ,
         \46197 , \46198 , \46199 , \46200 , \46201 , \46202 , \46203 , \46204 , \46205 , \46206 ,
         \46207 , \46208 , \46209 , \46210 , \46211 , \46212 , \46213 , \46214 , \46215 , \46216 ,
         \46217 , \46218 , \46219 , \46220 , \46221 , \46222 , \46223 , \46224 , \46225 , \46226 ,
         \46227 , \46228 , \46229 , \46230 , \46231 , \46232 , \46233 , \46234 , \46235 , \46236 ,
         \46237 , \46238 , \46239 , \46240 , \46241 , \46242 , \46243 , \46244 , \46245 , \46246 ,
         \46247 , \46248 , \46249 , \46250 , \46251 , \46252 , \46253 , \46254 , \46255 , \46256 ,
         \46257 , \46258 , \46259 , \46260 , \46261 , \46262 , \46263 , \46264 , \46265 , \46266 ,
         \46267 , \46268 , \46269 , \46270 , \46271 , \46272 , \46273 , \46274 , \46275 , \46276 ,
         \46277 , \46278 , \46279 , \46280 , \46281 , \46282 , \46283 , \46284 , \46285 , \46286 ,
         \46287 , \46288 , \46289 , \46290 , \46291 , \46292 , \46293 , \46294 , \46295 , \46296 ,
         \46297 , \46298 , \46299 , \46300 , \46301 , \46302 , \46303 , \46304 , \46305 , \46306 ,
         \46307 , \46308 , \46309 , \46310 , \46311 , \46312 , \46313 , \46314 , \46315 , \46316 ,
         \46317 , \46318 , \46319 , \46320 , \46321 , \46322 , \46323 , \46324 , \46325 , \46326 ,
         \46327 , \46328 , \46329 , \46330 , \46331 , \46332 , \46333 , \46334 , \46335 , \46336 ,
         \46337 , \46338 , \46339 , \46340 , \46341 , \46342 , \46343 , \46344 , \46345 , \46346 ,
         \46347 , \46348 , \46349 , \46350 , \46351 , \46352 , \46353 , \46354 , \46355 , \46356 ,
         \46357 , \46358 , \46359 , \46360 , \46361 , \46362 , \46363 , \46364 , \46365 , \46366 ,
         \46367 , \46368 , \46369 , \46370 , \46371 , \46372 , \46373 , \46374 , \46375 , \46376 ,
         \46377 , \46378 , \46379 , \46380 , \46381 , \46382 , \46383 , \46384 , \46385 , \46386 ,
         \46387 , \46388 , \46389 , \46390 , \46391 , \46392 , \46393 , \46394 , \46395 , \46396 ,
         \46397 , \46398 , \46399 , \46400 , \46401 , \46402 , \46403 , \46404 , \46405 , \46406 ,
         \46407 , \46408 , \46409 , \46410 , \46411 , \46412 , \46413 , \46414 , \46415 , \46416 ,
         \46417 , \46418 , \46419 , \46420 , \46421 , \46422 , \46423 , \46424 , \46425 , \46426 ,
         \46427 , \46428 , \46429 , \46430 , \46431 , \46432 , \46433 , \46434 , \46435 , \46436 ,
         \46437 , \46438 , \46439 , \46440 , \46441 , \46442 , \46443 , \46444 , \46445 , \46446 ,
         \46447 , \46448 , \46449 , \46450 , \46451 , \46452 , \46453 , \46454 , \46455 , \46456 ,
         \46457 , \46458 , \46459 , \46460 , \46461 , \46462 , \46463 , \46464 , \46465 , \46466 ,
         \46467 , \46468 , \46469 , \46470 , \46471 , \46472 , \46473 , \46474 , \46475 , \46476 ,
         \46477 , \46478 , \46479 , \46480 , \46481 , \46482 , \46483 , \46484 , \46485 , \46486 ,
         \46487 , \46488 , \46489 , \46490 , \46491 , \46492 , \46493 , \46494 , \46495 , \46496 ,
         \46497 , \46498 , \46499 , \46500 , \46501 , \46502 , \46503 , \46504 , \46505 , \46506 ,
         \46507 , \46508 , \46509 , \46510 , \46511 , \46512 , \46513 , \46514 , \46515 , \46516 ,
         \46517 , \46518 , \46519 , \46520 , \46521 , \46522 , \46523 , \46524 , \46525 , \46526 ,
         \46527 , \46528 , \46529 , \46530 , \46531 , \46532 , \46533 , \46534 , \46535 , \46536 ,
         \46537 , \46538 , \46539 , \46540 , \46541 , \46542 , \46543 , \46544 , \46545 , \46546 ,
         \46547 , \46548 , \46549 , \46550 , \46551 , \46552 , \46553 , \46554 , \46555 , \46556 ,
         \46557 , \46558 , \46559 , \46560 , \46561 , \46562 , \46563 , \46564 , \46565 , \46566 ,
         \46567 , \46568 , \46569 , \46570 , \46571 , \46572 , \46573 , \46574 , \46575 , \46576 ,
         \46577 , \46578 , \46579 , \46580 , \46581 , \46582 , \46583 , \46584 , \46585 , \46586 ,
         \46587 , \46588 , \46589 , \46590 , \46591 , \46592 , \46593 , \46594 , \46595 , \46596 ,
         \46597 , \46598 , \46599 , \46600 , \46601 , \46602 , \46603 , \46604 , \46605 , \46606 ,
         \46607 , \46608 , \46609 , \46610 , \46611 , \46612 , \46613 , \46614 , \46615 , \46616 ,
         \46617 , \46618 , \46619 , \46620 , \46621 , \46622 , \46623 , \46624 , \46625 , \46626 ,
         \46627 , \46628 , \46629 , \46630 , \46631 , \46632 , \46633 , \46634 , \46635 , \46636 ,
         \46637 , \46638 , \46639 , \46640 , \46641 , \46642 , \46643 , \46644 , \46645 , \46646 ,
         \46647 , \46648 , \46649 , \46650 , \46651 , \46652 , \46653 , \46654 , \46655 , \46656 ,
         \46657 , \46658 , \46659 , \46660 , \46661 , \46662 , \46663 , \46664 , \46665 , \46666 ,
         \46667 , \46668 , \46669 , \46670 , \46671 , \46672 , \46673 , \46674 , \46675 , \46676 ,
         \46677 , \46678 , \46679 , \46680 , \46681 , \46682 , \46683 , \46684 , \46685 , \46686 ,
         \46687 , \46688 , \46689 , \46690 , \46691 , \46692 , \46693 , \46694 , \46695 , \46696 ,
         \46697 , \46698 , \46699 , \46700 , \46701 , \46702 , \46703 , \46704 , \46705 , \46706 ,
         \46707 , \46708 , \46709 , \46710 , \46711 , \46712 , \46713 , \46714 , \46715 , \46716 ,
         \46717 , \46718 , \46719 , \46720 , \46721 , \46722 , \46723 , \46724 , \46725 , \46726 ,
         \46727 , \46728 , \46729 , \46730 , \46731 , \46732 , \46733 , \46734 , \46735 , \46736 ,
         \46737 , \46738 , \46739 , \46740 , \46741 , \46742 , \46743 , \46744 , \46745 , \46746 ,
         \46747 , \46748 , \46749 , \46750 , \46751 , \46752 , \46753 , \46754 , \46755 , \46756 ,
         \46757 , \46758 , \46759 , \46760 , \46761 , \46762 , \46763 , \46764 , \46765 , \46766 ,
         \46767 , \46768 , \46769 , \46770 , \46771 , \46772 , \46773 , \46774 , \46775 , \46776 ,
         \46777 , \46778 , \46779 , \46780 , \46781 , \46782 , \46783 , \46784 , \46785 , \46786 ,
         \46787 , \46788 , \46789 , \46790 , \46791 , \46792 , \46793 , \46794 , \46795 , \46796 ,
         \46797 , \46798 , \46799 , \46800 , \46801 , \46802 , \46803 , \46804 , \46805 , \46806 ,
         \46807 , \46808 , \46809 , \46810 , \46811 , \46812 , \46813 , \46814 , \46815 , \46816 ,
         \46817 , \46818 , \46819 , \46820 , \46821 , \46822 , \46823 , \46824 , \46825 , \46826 ,
         \46827 , \46828 , \46829 , \46830 , \46831 , \46832 , \46833 , \46834 , \46835 , \46836 ,
         \46837 , \46838 , \46839 , \46840 , \46841 , \46842 , \46843 , \46844 , \46845 , \46846 ,
         \46847 , \46848 , \46849 , \46850 , \46851 , \46852 , \46853 , \46854 , \46855 , \46856 ,
         \46857 , \46858 , \46859 , \46860 , \46861 , \46862 , \46863 , \46864 , \46865 , \46866 ,
         \46867 , \46868 , \46869 , \46870 , \46871 , \46872 , \46873 , \46874 , \46875 , \46876 ,
         \46877 , \46878 , \46879 , \46880 , \46881 , \46882 , \46883 , \46884 , \46885 , \46886 ,
         \46887 , \46888 , \46889 , \46890 , \46891 , \46892 , \46893 , \46894 , \46895 , \46896 ,
         \46897 , \46898 , \46899 , \46900 , \46901 , \46902 , \46903 , \46904 , \46905 , \46906 ,
         \46907 , \46908 , \46909 , \46910 , \46911 , \46912 , \46913 , \46914 , \46915 , \46916 ,
         \46917 , \46918 , \46919 , \46920 , \46921 , \46922 , \46923 , \46924 , \46925 , \46926 ,
         \46927 , \46928 , \46929 , \46930 , \46931 , \46932 , \46933 , \46934 , \46935 , \46936 ,
         \46937 , \46938 , \46939 , \46940 , \46941 , \46942 , \46943 , \46944 , \46945 , \46946 ,
         \46947 , \46948 , \46949 , \46950 , \46951 , \46952 , \46953 , \46954 , \46955 , \46956 ,
         \46957 , \46958 , \46959 , \46960 , \46961 , \46962 , \46963 , \46964 , \46965 , \46966 ,
         \46967 , \46968 , \46969 , \46970 , \46971 , \46972 , \46973 , \46974 , \46975 , \46976 ,
         \46977 , \46978 , \46979 , \46980 , \46981 , \46982 , \46983 , \46984 , \46985 , \46986 ,
         \46987 , \46988 , \46989 , \46990 , \46991 , \46992 , \46993 , \46994 , \46995 , \46996 ,
         \46997 , \46998 , \46999 , \47000 , \47001 , \47002 , \47003 , \47004 , \47005 , \47006 ,
         \47007 , \47008 , \47009 , \47010 , \47011 , \47012 , \47013 , \47014 , \47015 , \47016 ,
         \47017 , \47018 , \47019 , \47020 , \47021 , \47022 , \47023 , \47024 , \47025 , \47026 ,
         \47027 , \47028 , \47029 , \47030 , \47031 , \47032 , \47033 , \47034 , \47035 , \47036 ,
         \47037 , \47038 , \47039 , \47040 , \47041 , \47042 , \47043 , \47044 , \47045 , \47046 ,
         \47047 , \47048 , \47049 , \47050 , \47051 , \47052 , \47053 , \47054 , \47055 , \47056 ,
         \47057 , \47058 , \47059 , \47060 , \47061 , \47062 , \47063 , \47064 , \47065 , \47066 ,
         \47067 , \47068 , \47069 , \47070 , \47071 , \47072 , \47073 , \47074 , \47075 , \47076 ,
         \47077 , \47078 , \47079 , \47080 , \47081 , \47082 , \47083 , \47084 , \47085 , \47086 ,
         \47087 , \47088 , \47089 , \47090 , \47091 , \47092 , \47093 , \47094 , \47095 , \47096 ,
         \47097 , \47098 , \47099 , \47100 , \47101 , \47102 , \47103 , \47104 , \47105 , \47106 ,
         \47107 , \47108 , \47109 , \47110 , \47111 , \47112 , \47113 , \47114 , \47115 , \47116 ,
         \47117 , \47118 , \47119 , \47120 , \47121 , \47122 , \47123 , \47124 , \47125 , \47126 ,
         \47127 , \47128 , \47129 , \47130 , \47131 , \47132 , \47133 , \47134 , \47135 , \47136 ,
         \47137 , \47138 , \47139 , \47140 , \47141 , \47142 , \47143 , \47144 , \47145 , \47146 ,
         \47147 , \47148 , \47149 , \47150 , \47151 , \47152 , \47153 , \47154 , \47155 , \47156 ,
         \47157 , \47158 , \47159 , \47160 , \47161 , \47162 , \47163 , \47164 , \47165 , \47166 ,
         \47167 , \47168 , \47169 , \47170 , \47171 , \47172 , \47173 , \47174 , \47175 , \47176 ,
         \47177 , \47178 , \47179 , \47180 , \47181 , \47182 , \47183 , \47184 , \47185 , \47186 ,
         \47187 , \47188 , \47189 , \47190 , \47191 , \47192 , \47193 , \47194 , \47195 , \47196 ,
         \47197 , \47198 , \47199 , \47200 , \47201 , \47202 , \47203 , \47204 , \47205 , \47206 ,
         \47207 , \47208 , \47209 , \47210 , \47211 , \47212 , \47213 , \47214 , \47215 , \47216 ,
         \47217 , \47218 , \47219 , \47220 , \47221 , \47222 , \47223 , \47224 , \47225 , \47226 ,
         \47227 , \47228 , \47229 , \47230 , \47231 , \47232 , \47233 , \47234 , \47235 , \47236 ,
         \47237 , \47238 , \47239 , \47240 , \47241 , \47242 , \47243 , \47244 , \47245 , \47246 ,
         \47247 , \47248 , \47249 , \47250 , \47251 , \47252 , \47253 , \47254 , \47255 , \47256 ,
         \47257 , \47258 , \47259 , \47260 , \47261 , \47262 , \47263 , \47264 , \47265 , \47266 ,
         \47267 , \47268 , \47269 , \47270 , \47271 , \47272 , \47273 , \47274 , \47275 , \47276 ,
         \47277 , \47278 , \47279 , \47280 , \47281 , \47282 , \47283 , \47284 , \47285 , \47286 ,
         \47287 , \47288 , \47289 , \47290 , \47291 , \47292 , \47293 , \47294 , \47295 , \47296 ,
         \47297 , \47298 , \47299 , \47300 , \47301 , \47302 , \47303 , \47304 , \47305 , \47306 ,
         \47307 , \47308 , \47309 , \47310 , \47311 , \47312 , \47313 , \47314 , \47315 , \47316 ,
         \47317 , \47318 , \47319 , \47320 , \47321 , \47322 , \47323 , \47324 , \47325 , \47326 ,
         \47327 , \47328 , \47329 , \47330 , \47331 , \47332 , \47333 , \47334 , \47335 , \47336 ,
         \47337 , \47338 , \47339 , \47340 , \47341 , \47342 , \47343 , \47344 , \47345 , \47346 ,
         \47347 , \47348 , \47349 , \47350 , \47351 , \47352 , \47353 , \47354 , \47355 , \47356 ,
         \47357 , \47358 , \47359 , \47360 , \47361 , \47362 , \47363 , \47364 , \47365 , \47366 ,
         \47367 , \47368 , \47369 , \47370 , \47371 , \47372 , \47373 , \47374 , \47375 , \47376 ,
         \47377 , \47378 , \47379 , \47380 , \47381 , \47382 , \47383 , \47384 , \47385 , \47386 ,
         \47387 , \47388 , \47389 , \47390 , \47391 , \47392 , \47393 , \47394 , \47395 , \47396 ,
         \47397 , \47398 , \47399 , \47400 , \47401 , \47402 , \47403 , \47404 , \47405 , \47406 ,
         \47407 , \47408 , \47409 , \47410 , \47411 , \47412 , \47413 , \47414 , \47415 , \47416 ,
         \47417 , \47418 , \47419 , \47420 , \47421 , \47422 , \47423 , \47424 , \47425 , \47426 ,
         \47427 , \47428 , \47429 , \47430 , \47431 , \47432 , \47433 , \47434 , \47435 , \47436 ,
         \47437 , \47438 , \47439 , \47440 , \47441 , \47442 , \47443 , \47444 , \47445 , \47446 ,
         \47447 , \47448 , \47449 , \47450 , \47451 , \47452 , \47453 , \47454 , \47455 , \47456 ,
         \47457 , \47458 , \47459 , \47460 , \47461 , \47462 , \47463 , \47464 , \47465 , \47466 ,
         \47467 , \47468 , \47469 , \47470 , \47471 , \47472 , \47473 , \47474 , \47475 , \47476 ,
         \47477 , \47478 , \47479 , \47480 , \47481 , \47482 , \47483 , \47484 , \47485 , \47486 ,
         \47487 , \47488 , \47489 , \47490 , \47491 , \47492 , \47493 , \47494 , \47495 , \47496 ,
         \47497 , \47498 , \47499 , \47500 , \47501 , \47502 , \47503 , \47504 , \47505 , \47506 ,
         \47507 , \47508 , \47509 , \47510 , \47511 , \47512 , \47513 , \47514 , \47515 , \47516 ,
         \47517 , \47518 , \47519 , \47520 , \47521 , \47522 , \47523 , \47524 , \47525 , \47526 ,
         \47527 , \47528 , \47529 , \47530 , \47531 , \47532 , \47533 , \47534 , \47535 , \47536 ,
         \47537 , \47538 , \47539 , \47540 , \47541 , \47542 , \47543 , \47544 , \47545 , \47546 ,
         \47547 , \47548 , \47549 , \47550 , \47551 , \47552 , \47553 , \47554 , \47555 , \47556 ,
         \47557 , \47558 , \47559 , \47560 , \47561 , \47562 , \47563 , \47564 , \47565 , \47566 ,
         \47567 , \47568 , \47569 , \47570 , \47571 , \47572 , \47573 , \47574 , \47575 , \47576 ,
         \47577 , \47578 , \47579 , \47580 , \47581 , \47582 , \47583 , \47584 , \47585 , \47586 ,
         \47587 , \47588 , \47589 , \47590 , \47591 , \47592 , \47593 , \47594 , \47595 , \47596 ,
         \47597 , \47598 , \47599 , \47600 , \47601 , \47602 , \47603 , \47604 , \47605 , \47606 ,
         \47607 , \47608_nGdf4e , \47609 , \47610 , \47611 , \47612_nGdf51 , \47613 , \47614 , \47615_nGdf53 , \47616 ,
         \47617 , \47618_nGdf55 , \47619 , \47620 , \47621_nGdf57 , \47622 , \47623 , \47624_nGdf59 , \47625 , \47626 ,
         \47627_nGdf5b , \47628 , \47629 , \47630_nGdf5d , \47631 , \47632 , \47633_nGdf5f , \47634 , \47635 , \47636_nGdf61 ,
         \47637 , \47638 , \47639_nGdf63 , \47640 , \47641 , \47642_nGdf65 , \47643 , \47644 , \47645_nGdf67 , \47646 ,
         \47647 , \47648_nGdf69 , \47649 , \47650 , \47651_nGdf6b , \47652 , \47653 , \47654_nGdf6d , \47655 , \47656 ,
         \47657_nGdf6f , \47658 , \47659 , \47660_nGdf71 , \47661 , \47662 , \47663_nGdf73 , \47664 , \47665 , \47666_nGdf75 ,
         \47667 , \47668 , \47669_nGdf77 , \47670 , \47671 , \47672_nGdf79 , \47673 , \47674 , \47675_nGdf7b , \47676 ,
         \47677 , \47678_nGdf7d , \47679 , \47680 , \47681_nGdf7f , \47682 , \47683 , \47684_nGdf81 , \47685 , \47686 ,
         \47687_nGdf83 , \47688 , \47689 , \47690_nGdf85 , \47691 , \47692 , \47693_nGdf87 , \47694 , \47695 , \47696_nGdf89 ,
         \47697 , \47698 , \47699_nGdf8b , \47700 , \47701 , \47702_nGdf8d , \47703 , \47704 , \47705_nGdf8f , \47706 ,
         \47707 , \47708_nGdf91 , \47709 , \47710 , \47711_nGdf93 , \47712 , \47713 , \47714_nGdf95 , \47715 , \47716 ,
         \47717_nGdf97 , \47718 , \47719 , \47720_nGdf99 , \47721 , \47722 , \47723_nGdf9b , \47724 , \47725 , \47726_nGdf9d ,
         \47727 , \47728 , \47729_nGdf9f , \47730 , \47731 , \47732_nGdfa1 , \47733 , \47734 , \47735_nGdfa3 , \47736 ,
         \47737 , \47738_nGdfa5 , \47739 , \47740 , \47741_nGdfa7 , \47742 , \47743 , \47744_nGdfa9 , \47745 , \47746 ,
         \47747_nGdfab , \47748 , \47749 , \47750_nGdfad , \47751 , \47752 , \47753_nGdfaf , \47754 , \47755 , \47756_nGdfb1 ,
         \47757 , \47758 , \47759_nGdfb3 , \47760 , \47761 , \47762_nGdfb5 , \47763 , \47764 , \47765_nGdfb7 , \47766 ,
         \47767 , \47768_nGdfb9 , \47769 , \47770 , \47771_nGdfbb , \47772 , \47773 , \47774_nGdfbd , \47775 , \47776 ,
         \47777_nGdfbf , \47778 , \47779 , \47780_nGdfc1 , \47781 , \47782 , \47783_nGdfc3 , \47784 , \47785 , \47786_nGdfc5 ,
         \47787 , \47788 , \47789_nGdfc7 , \47790 , \47791 , \47792 , \47793_nGdfca , \47794 , \47795 , \47796 ,
         \47797_nGdfcd , \47798 , \47799 , \47800 , \47801_nGdfd0 , \47802 , \47803 , \47804_nGdfd2 , \47805 , \47806 ,
         \47807 , \47808_nGdfd5 , \47809 , \47810 , \47811_nGdfd7 , \47812 , \47813 , \47814 , \47815_nGdfda , \47816 ,
         \47817 , \47818_nGdfdc , \47819 , \47820 , \47821 , \47822_nGdfdf , \47823 , \47824 , \47825_nGdfe1 , \47826 ,
         \47827 , \47828 , \47829_nGdfe4 , \47830 , \47831 , \47832_nGdfe6 , \47833 , \47834 , \47835 , \47836_nGdfe9 ,
         \47837 , \47838 , \47839_nGdfeb , \47840 , \47841 , \47842 , \47843_nGdfee , \47844 , \47845 , \47846_nGdff0 ,
         \47847 , \47848 , \47849 , \47850_nGdff3 , \47851 , \47852 , \47853_nGdff5 , \47854 , \47855 , \47856 ,
         \47857_nGdff8 , \47858 , \47859 , \47860_nGdffa , \47861 , \47862 , \47863 , \47864_nGdffd , \47865 , \47866 ,
         \47867_nGdfff , \47868 , \47869 , \47870 , \47871_nGe002 , \47872 , \47873 , \47874_nGe004 , \47875 , \47876 ,
         \47877 , \47878_nGe007 , \47879 , \47880 , \47881_nGe009 , \47882 , \47883 , \47884 , \47885_nGe00c , \47886 ,
         \47887 , \47888_nGe00e , \47889 , \47890 , \47891 , \47892_nGe011 , \47893 , \47894 , \47895_nGe013 , \47896 ,
         \47897 , \47898 , \47899_nGe016 , \47900 , \47901 , \47902_nGe018 , \47903 ;
buf \U$labaj5628 ( R_58_102f1b78, \47609 );
buf \U$labaj5629 ( R_59_be1fc68, \47613 );
buf \U$labaj5630 ( R_5a_10279198, \47616 );
buf \U$labaj5631 ( R_5b_102299e8, \47619 );
buf \U$labaj5632 ( R_5c_101d0448, \47622 );
buf \U$labaj5633 ( R_5d_f7f82f0, \47625 );
buf \U$labaj5634 ( R_5e_be21600, \47628 );
buf \U$labaj5635 ( R_5f_f7fa5b8, \47631 );
buf \U$labaj5636 ( R_60_1027d530, \47634 );
buf \U$labaj5637 ( R_61_10205ae8, \47637 );
buf \U$labaj5638 ( R_62_10283510, \47640 );
buf \U$labaj5639 ( R_63_f82b578, \47643 );
buf \U$labaj5640 ( R_64_ace4e68, \47646 );
buf \U$labaj5641 ( R_65_f8204e0, \47649 );
buf \U$labaj5642 ( R_66_1027a0b0, \47652 );
buf \U$labaj5643 ( R_67_1022dc30, \47655 );
buf \U$labaj5644 ( R_68_102478a8, \47658 );
buf \U$labaj5645 ( R_69_10286f78, \47661 );
buf \U$labaj5646 ( R_6a_f7edd80, \47664 );
buf \U$labaj5647 ( R_6b_101c3628, \47667 );
buf \U$labaj5648 ( R_6c_f7fbe00, \47670 );
buf \U$labaj5649 ( R_6d_f7ce9f8, \47673 );
buf \U$labaj5650 ( R_6e_f7c8830, \47676 );
buf \U$labaj5651 ( R_6f_101ffc68, \47679 );
buf \U$labaj5652 ( R_70_f7d4000, \47682 );
buf \U$labaj5653 ( R_71_acee958, \47685 );
buf \U$labaj5654 ( R_72_94046c0, \47688 );
buf \U$labaj5655 ( R_73_101ee420, \47691 );
buf \U$labaj5656 ( R_74_102eb268, \47694 );
buf \U$labaj5657 ( R_75_b320c50, \47697 );
buf \U$labaj5658 ( R_76_ad80a90, \47700 );
buf \U$labaj5659 ( R_77_1027fd48, \47703 );
buf \U$labaj5660 ( R_78_f7ce4b8, \47706 );
buf \U$labaj5661 ( R_79_ad77048, \47709 );
buf \U$labaj5662 ( R_7a_102a6ae0, \47712 );
buf \U$labaj5663 ( R_7b_f7e4c78, \47715 );
buf \U$labaj5664 ( R_7c_e2a6ce0, \47718 );
buf \U$labaj5665 ( R_7d_101e86e0, \47721 );
buf \U$labaj5666 ( R_7e_e2a9cc8, \47724 );
buf \U$labaj5667 ( R_7f_10292be0, \47727 );
buf \U$labaj5668 ( R_80_b33cde8, \47730 );
buf \U$labaj5669 ( R_81_101e2908, \47733 );
buf \U$labaj5670 ( R_82_102e9780, \47736 );
buf \U$labaj5671 ( R_83_f8157a0, \47739 );
buf \U$labaj5672 ( R_84_f819358, \47742 );
buf \U$labaj5673 ( R_85_ace8b70, \47745 );
buf \U$labaj5674 ( R_86_be142b0, \47748 );
buf \U$labaj5675 ( R_87_f81b770, \47751 );
buf \U$labaj5676 ( R_88_b330278, \47754 );
buf \U$labaj5677 ( R_89_f7fe9f8, \47757 );
buf \U$labaj5678 ( R_8a_101cf488, \47760 );
buf \U$labaj5679 ( R_8b_f8225c0, \47763 );
buf \U$labaj5680 ( R_8c_101d4738, \47766 );
buf \U$labaj5681 ( R_8d_101c4000, \47769 );
buf \U$labaj5682 ( R_8e_101fe960, \47772 );
buf \U$labaj5683 ( R_8f_102a0330, \47775 );
buf \U$labaj5684 ( R_90_f7f4bd0, \47778 );
buf \U$labaj5685 ( R_91_1023e5a8, \47781 );
buf \U$labaj5686 ( R_92_10248da8, \47784 );
buf \U$labaj5687 ( R_93_be2c938, \47787 );
buf \U$labaj5688 ( R_94_f7f5458, \47790 );
buf \U$labaj5689 ( R_95_f7c6808, \47794 );
buf \U$labaj5690 ( R_96_be316a8, \47798 );
buf \U$labaj5691 ( R_97_e2a0328, \47802 );
buf \U$labaj5692 ( R_98_be2d850, \47805 );
buf \U$labaj5693 ( R_99_10217db0, \47809 );
buf \U$labaj5694 ( R_9a_f7ec340, \47812 );
buf \U$labaj5695 ( R_9b_be23ec0, \47816 );
buf \U$labaj5696 ( R_9c_101d4540, \47819 );
buf \U$labaj5697 ( R_9d_f800828, \47823 );
buf \U$labaj5698 ( R_9e_102970c8, \47826 );
buf \U$labaj5699 ( R_9f_10221de0, \47830 );
buf \U$labaj5700 ( R_a0_ad8d568, \47833 );
buf \U$labaj5701 ( R_a1_be4eb58, \47837 );
buf \U$labaj5702 ( R_a2_f7c5500, \47840 );
buf \U$labaj5703 ( R_a3_ad88f30, \47844 );
buf \U$labaj5704 ( R_a4_f82f088, \47847 );
buf \U$labaj5705 ( R_a5_f7dcbc8, \47851 );
buf \U$labaj5706 ( R_a6_10292940, \47854 );
buf \U$labaj5707 ( R_a7_be138d8, \47858 );
buf \U$labaj5708 ( R_a8_acee418, \47861 );
buf \U$labaj5709 ( R_a9_ad84450, \47865 );
buf \U$labaj5710 ( R_aa_be10838, \47868 );
buf \U$labaj5711 ( R_ab_be31fd8, \47872 );
buf \U$labaj5712 ( R_ac_acdaef0, \47875 );
buf \U$labaj5713 ( R_ad_acea908, \47879 );
buf \U$labaj5714 ( R_ae_101f8830, \47882 );
buf \U$labaj5715 ( R_af_f7dec98, \47886 );
buf \U$labaj5716 ( R_b0_101e2c50, \47889 );
buf \U$labaj5717 ( R_b1_f801b30, \47893 );
buf \U$labaj5718 ( R_b2_be16e00, \47896 );
buf \U$labaj5719 ( R_b3_102e3cf0, \47900 );
buf \U$labaj5720 ( R_b4_10291788, \47903 );
not \U$1 ( \9052 , RIbc62af0_23);
not \U$2 ( \9053 , RIbc62a78_22);
not \U$3 ( \9054 , RIbc62a00_21);
not \U$4 ( \9055 , RIbc62988_20);
not \U$5 ( \9056 , RIbc62910_19);
not \U$6 ( \9057 , RIbc62898_18);
not \U$7 ( \9058 , RIbc62820_17);
nor \U$8 ( \9059 , \9052 , \9053 , \9054 , \9055 , \9056 , \9057 , \9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$9 ( \9060 , RIdec64b8_720, \9059 );
nor \U$10 ( \9061 , RIbc62af0_23, \9053 , \9054 , \9055 , \9056 , \9057 , \9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$11 ( \9062 , RIdec37b8_688, \9061 );
nor \U$12 ( \9063 , \9052 , RIbc62a78_22, \9054 , \9055 , \9056 , \9057 , \9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$13 ( \9064 , RIfc8daa0_6634, \9063 );
nor \U$14 ( \9065 , RIbc62af0_23, RIbc62a78_22, \9054 , \9055 , \9056 , \9057 , \9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$15 ( \9066 , RIdec0ab8_656, \9065 );
nor \U$16 ( \9067 , \9052 , \9053 , RIbc62a00_21, \9055 , \9056 , \9057 , \9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$17 ( \9068 , RIfc56348_6003, \9067 );
nor \U$18 ( \9069 , RIbc62af0_23, \9053 , RIbc62a00_21, \9055 , \9056 , \9057 , \9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$19 ( \9070 , RIdebddb8_624, \9069 );
nor \U$20 ( \9071 , \9052 , RIbc62a78_22, RIbc62a00_21, \9055 , \9056 , \9057 , \9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$21 ( \9072 , RIdebb0b8_592, \9071 );
nor \U$22 ( \9073 , RIbc62af0_23, RIbc62a78_22, RIbc62a00_21, \9055 , \9056 , \9057 , \9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$23 ( \9074 , RIdeb83b8_560, \9073 );
nor \U$24 ( \9075 , \9052 , \9053 , \9054 , RIbc62988_20, \9056 , \9057 , \9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$25 ( \9076 , RIfc98798_6757, \9075 );
nor \U$26 ( \9077 , RIbc62af0_23, \9053 , \9054 , RIbc62988_20, \9056 , \9057 , \9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$27 ( \9078 , RIdeb29b8_496, \9077 );
nor \U$28 ( \9079 , \9052 , RIbc62a78_22, \9054 , RIbc62988_20, \9056 , \9057 , \9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$29 ( \9080 , RIfcbd098_7173, \9079 );
nor \U$30 ( \9081 , RIbc62af0_23, RIbc62a78_22, \9054 , RIbc62988_20, \9056 , \9057 , \9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$31 ( \9082 , RIdeafcb8_464, \9081 );
nor \U$32 ( \9083 , \9052 , \9053 , RIbc62a00_21, RIbc62988_20, \9056 , \9057 , \9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$33 ( \9084 , RIfc8dc08_6635, \9083 );
nor \U$34 ( \9085 , RIbc62af0_23, \9053 , RIbc62a00_21, RIbc62988_20, \9056 , \9057 , \9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$35 ( \9086 , RIdeacb80_432, \9085 );
nor \U$36 ( \9087 , \9052 , RIbc62a78_22, RIbc62a00_21, RIbc62988_20, \9056 , \9057 , \9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$37 ( \9088 , RIdea6280_400, \9087 );
nor \U$38 ( \9089 , RIbc62af0_23, RIbc62a78_22, RIbc62a00_21, RIbc62988_20, \9056 , \9057 , \9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$39 ( \9090 , RIde9f980_368, \9089 );
nor \U$40 ( \9091 , \9052 , \9053 , \9054 , \9055 , RIbc62910_19, \9057 , \9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$41 ( \9092 , RIfcd6868_7463, \9091 );
nor \U$42 ( \9093 , RIbc62af0_23, \9053 , \9054 , \9055 , RIbc62910_19, \9057 , \9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$43 ( \9094 , RIfc8ded8_6637, \9093 );
nor \U$44 ( \9095 , \9052 , RIbc62a78_22, \9054 , \9055 , RIbc62910_19, \9057 , \9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$45 ( \9096 , RIfc7dd80_6454, \9095 );
nor \U$46 ( \9097 , RIbc62af0_23, RIbc62a78_22, \9054 , \9055 , RIbc62910_19, \9057 , \9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$47 ( \9098 , RIfc56618_6005, \9097 );
nor \U$48 ( \9099 , \9052 , \9053 , RIbc62a00_21, \9055 , RIbc62910_19, \9057 , \9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$49 ( \9100 , RIde92e10_306, \9099 );
nor \U$50 ( \9101 , RIbc62af0_23, \9053 , RIbc62a00_21, \9055 , RIbc62910_19, \9057 , \9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$51 ( \9102 , RIde8f300_288, \9101 );
nor \U$52 ( \9103 , \9052 , RIbc62a78_22, RIbc62a00_21, \9055 , RIbc62910_19, \9057 , \9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$53 ( \9104 , RIde8b160_268, \9103 );
nor \U$54 ( \9105 , RIbc62af0_23, RIbc62a78_22, RIbc62a00_21, \9055 , RIbc62910_19, \9057 , \9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$55 ( \9106 , RIde86fc0_248, \9105 );
nor \U$56 ( \9107 , \9052 , \9053 , \9054 , RIbc62988_20, RIbc62910_19, \9057 , \9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$57 ( \9108 , RIde82ad8_227, \9107 );
nor \U$58 ( \9109 , RIbc62af0_23, \9053 , \9054 , RIbc62988_20, RIbc62910_19, \9057 , \9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$59 ( \9110 , RIfc8e040_6638, \9109 );
nor \U$60 ( \9111 , \9052 , RIbc62a78_22, \9054 , RIbc62988_20, RIbc62910_19, \9057 , \9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$61 ( \9112 , RIfcd96d0_7496, \9111 );
nor \U$62 ( \9113 , RIbc62af0_23, RIbc62a78_22, \9054 , RIbc62988_20, RIbc62910_19, \9057 , \9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$63 ( \9114 , RIfca1e10_6864, \9113 );
nor \U$64 ( \9115 , \9052 , \9053 , RIbc62a00_21, RIbc62988_20, RIbc62910_19, \9057 , \9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$65 ( \9116 , RIfcbd200_7174, \9115 );
nor \U$66 ( \9117 , RIbc62af0_23, \9053 , RIbc62a00_21, RIbc62988_20, RIbc62910_19, \9057 , \9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$67 ( \9118 , RIe16c5c0_2610, \9117 );
nor \U$68 ( \9119 , \9052 , RIbc62a78_22, RIbc62a00_21, RIbc62988_20, RIbc62910_19, \9057 , \9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$69 ( \9120 , RIe16a298_2585, \9119 );
nor \U$70 ( \9121 , RIbc62af0_23, RIbc62a78_22, RIbc62a00_21, RIbc62988_20, RIbc62910_19, \9057 , \9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$71 ( \9122 , RIe168ab0_2568, \9121 );
nor \U$72 ( \9123 , \9052 , \9053 , \9054 , \9055 , \9056 , RIbc62898_18, \9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$73 ( \9124 , RIe1664b8_2541, \9123 );
nor \U$74 ( \9125 , RIbc62af0_23, \9053 , \9054 , \9055 , \9056 , RIbc62898_18, \9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$75 ( \9126 , RIe1637b8_2509, \9125 );
nor \U$76 ( \9127 , \9052 , RIbc62a78_22, \9054 , \9055 , \9056 , RIbc62898_18, \9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$77 ( \9128 , RIee37f00_5095, \9127 );
nor \U$78 ( \9129 , RIbc62af0_23, RIbc62a78_22, \9054 , \9055 , \9056 , RIbc62898_18, \9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$79 ( \9130 , RIe160ab8_2477, \9129 );
nor \U$80 ( \9131 , \9052 , \9053 , RIbc62a00_21, \9055 , \9056 , RIbc62898_18, \9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$81 ( \9132 , RIfc8ea18_6645, \9131 );
nor \U$82 ( \9133 , RIbc62af0_23, \9053 , RIbc62a00_21, \9055 , \9056 , RIbc62898_18, \9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$83 ( \9134 , RIe15ddb8_2445, \9133 );
nor \U$84 ( \9135 , \9052 , RIbc62a78_22, RIbc62a00_21, \9055 , \9056 , RIbc62898_18, \9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$85 ( \9136 , RIe1583b8_2381, \9135 );
nor \U$86 ( \9137 , RIbc62af0_23, RIbc62a78_22, RIbc62a00_21, \9055 , \9056 , RIbc62898_18, \9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$87 ( \9138 , RIe1556b8_2349, \9137 );
nor \U$88 ( \9139 , \9052 , \9053 , \9054 , RIbc62988_20, \9056 , RIbc62898_18, \9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$89 ( \9140 , RIfe9f828_8159, \9139 );
nor \U$90 ( \9141 , RIbc62af0_23, \9053 , \9054 , RIbc62988_20, \9056 , RIbc62898_18, \9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$91 ( \9142 , RIe1529b8_2317, \9141 );
nor \U$92 ( \9143 , \9052 , RIbc62a78_22, \9054 , RIbc62988_20, \9056 , RIbc62898_18, \9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$93 ( \9144 , RIfe9f990_8160, \9143 );
nor \U$94 ( \9145 , RIbc62af0_23, RIbc62a78_22, \9054 , RIbc62988_20, \9056 , RIbc62898_18, \9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$95 ( \9146 , RIe14fcb8_2285, \9145 );
nor \U$96 ( \9147 , \9052 , \9053 , RIbc62a00_21, RIbc62988_20, \9056 , RIbc62898_18, \9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$97 ( \9148 , RIfcbd368_7175, \9147 );
nor \U$98 ( \9149 , RIbc62af0_23, \9053 , RIbc62a00_21, RIbc62988_20, \9056 , RIbc62898_18, \9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$99 ( \9150 , RIe14cfb8_2253, \9149 );
nor \U$100 ( \9151 , \9052 , RIbc62a78_22, RIbc62a00_21, RIbc62988_20, \9056 , RIbc62898_18, \9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$101 ( \9152 , RIe14a2b8_2221, \9151 );
nor \U$102 ( \9153 , RIbc62af0_23, RIbc62a78_22, RIbc62a00_21, RIbc62988_20, \9056 , RIbc62898_18, \9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$103 ( \9154 , RIe1475b8_2189, \9153 );
nor \U$104 ( \9155 , \9052 , \9053 , \9054 , \9055 , RIbc62910_19, RIbc62898_18, \9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$105 ( \9156 , RIfc8ee50_6648, \9155 );
nor \U$106 ( \9157 , RIbc62af0_23, \9053 , \9054 , \9055 , RIbc62910_19, RIbc62898_18, \9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$107 ( \9158 , RIfc45278_5809, \9157 );
nor \U$108 ( \9159 , \9052 , RIbc62a78_22, \9054 , \9055 , RIbc62910_19, RIbc62898_18, \9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$109 ( \9160 , RIfc98360_6754, \9159 );
nor \U$110 ( \9161 , RIbc62af0_23, RIbc62a78_22, \9054 , \9055 , RIbc62910_19, RIbc62898_18, \9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$111 ( \9162 , RIfca2248_6867, \9161 );
nor \U$112 ( \9163 , \9052 , \9053 , RIbc62a00_21, \9055 , RIbc62910_19, RIbc62898_18, \9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$113 ( \9164 , RIe141d20_2126, \9163 );
nor \U$114 ( \9165 , RIbc62af0_23, \9053 , RIbc62a00_21, \9055 , RIbc62910_19, RIbc62898_18, \9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$115 ( \9166 , RIe13f9f8_2101, \9165 );
nor \U$116 ( \9167 , \9052 , RIbc62a78_22, RIbc62a00_21, \9055 , RIbc62910_19, RIbc62898_18, \9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$117 ( \9168 , RIdf3d900_2077, \9167 );
nor \U$118 ( \9169 , RIbc62af0_23, RIbc62a78_22, RIbc62a00_21, \9055 , RIbc62910_19, RIbc62898_18, \9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$119 ( \9170 , RIdf3b470_2051, \9169 );
nor \U$120 ( \9171 , \9052 , \9053 , \9054 , RIbc62988_20, RIbc62910_19, RIbc62898_18, \9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$121 ( \9172 , RIfcd6ca0_7466, \9171 );
nor \U$122 ( \9173 , RIbc62af0_23, \9053 , \9054 , RIbc62988_20, RIbc62910_19, RIbc62898_18, \9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$123 ( \9174 , RIee2ff08_5004, \9173 );
nor \U$124 ( \9175 , \9052 , RIbc62a78_22, \9054 , RIbc62988_20, RIbc62910_19, RIbc62898_18, \9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$125 ( \9176 , RIfc8ece8_6647, \9175 );
nor \U$126 ( \9177 , RIbc62af0_23, RIbc62a78_22, \9054 , RIbc62988_20, RIbc62910_19, RIbc62898_18, \9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$127 ( \9178 , RIee2dd48_4980, \9177 );
nor \U$128 ( \9179 , \9052 , \9053 , RIbc62a00_21, RIbc62988_20, RIbc62910_19, RIbc62898_18, \9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$129 ( \9180 , RIdf36718_1996, \9179 );
nor \U$130 ( \9181 , RIbc62af0_23, \9053 , RIbc62a00_21, RIbc62988_20, RIbc62910_19, RIbc62898_18, \9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$131 ( \9182 , RIdf34120_1969, \9181 );
nor \U$132 ( \9183 , \9052 , RIbc62a78_22, RIbc62a00_21, RIbc62988_20, RIbc62910_19, RIbc62898_18, \9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$133 ( \9184 , RIdf31f60_1945, \9183 );
nor \U$134 ( \9185 , RIbc62af0_23, RIbc62a78_22, RIbc62a00_21, RIbc62988_20, RIbc62910_19, RIbc62898_18, \9058 , RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$135 ( \9186 , RIfe9f6c0_8158, \9185 );
or \U$136 ( \9187 , \9060 , \9062 , \9064 , \9066 , \9068 , \9070 , \9072 , \9074 , \9076 , \9078 , \9080 , \9082 , \9084 , \9086 , \9088 , \9090 , \9092 , \9094 , \9096 , \9098 , \9100 , \9102 , \9104 , \9106 , \9108 , \9110 , \9112 , \9114 , \9116 , \9118 , \9120 , \9122 , \9124 , \9126 , \9128 , \9130 , \9132 , \9134 , \9136 , \9138 , \9140 , \9142 , \9144 , \9146 , \9148 , \9150 , \9152 , \9154 , \9156 , \9158 , \9160 , \9162 , \9164 , \9166 , \9168 , \9170 , \9172 , \9174 , \9176 , \9178 , \9180 , \9182 , \9184 , \9186 );
nor \U$137 ( \9188 , \9052 , \9053 , \9054 , \9055 , \9056 , \9057 , RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$138 ( \9189 , RIfcb4560_7074, \9188 );
nor \U$139 ( \9190 , RIbc62af0_23, \9053 , \9054 , \9055 , \9056 , \9057 , RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$140 ( \9191 , RIfc45db8_5817, \9190 );
nor \U$141 ( \9192 , \9052 , RIbc62a78_22, \9054 , \9055 , \9056 , \9057 , RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$142 ( \9193 , RIfc8e1a8_6639, \9192 );
nor \U$143 ( \9194 , RIbc62af0_23, RIbc62a78_22, \9054 , \9055 , \9056 , \9057 , RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$144 ( \9195 , RIfc7d678_6449, \9194 );
nor \U$145 ( \9196 , \9052 , \9053 , RIbc62a00_21, \9055 , \9056 , \9057 , RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$146 ( \9197 , RIdf2aee0_1865, \9196 );
nor \U$147 ( \9198 , RIbc62af0_23, \9053 , RIbc62a00_21, \9055 , \9056 , \9057 , RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$148 ( \9199 , RIdf28ff0_1843, \9198 );
nor \U$149 ( \9200 , \9052 , RIbc62a78_22, RIbc62a00_21, \9055 , \9056 , \9057 , RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$150 ( \9201 , RIdf26e30_1819, \9200 );
nor \U$151 ( \9202 , RIbc62af0_23, RIbc62a78_22, RIbc62a00_21, \9055 , \9056 , \9057 , RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$152 ( \9203 , RIdf25378_1800, \9202 );
nor \U$153 ( \9204 , \9052 , \9053 , \9054 , RIbc62988_20, \9056 , \9057 , RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$154 ( \9205 , RIfcb43f8_7073, \9204 );
nor \U$155 ( \9206 , RIbc62af0_23, \9053 , \9054 , RIbc62988_20, \9056 , \9057 , RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$156 ( \9207 , RIfc8e748_6643, \9206 );
nor \U$157 ( \9208 , \9052 , RIbc62a78_22, \9054 , RIbc62988_20, \9056 , \9057 , RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$158 ( \9209 , RIdf23488_1778, \9208 );
nor \U$159 ( \9210 , RIbc62af0_23, RIbc62a78_22, \9054 , RIbc62988_20, \9056 , \9057 , RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$160 ( \9211 , RIfcc2c00_7238, \9210 );
nor \U$161 ( \9212 , \9052 , \9053 , RIbc62a00_21, RIbc62988_20, \9056 , \9057 , RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$162 ( \9213 , RIdf21e08_1762, \9212 );
nor \U$163 ( \9214 , RIbc62af0_23, \9053 , RIbc62a00_21, RIbc62988_20, \9056 , \9057 , RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$164 ( \9215 , RIdf20788_1746, \9214 );
nor \U$165 ( \9216 , \9052 , RIbc62a78_22, RIbc62a00_21, RIbc62988_20, \9056 , \9057 , RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$166 ( \9217 , RIdf1b760_1689, \9216 );
nor \U$167 ( \9218 , RIbc62af0_23, RIbc62a78_22, RIbc62a00_21, RIbc62988_20, \9056 , \9057 , RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$168 ( \9219 , RIdf1a248_1674, \9218 );
nor \U$169 ( \9220 , \9052 , \9053 , \9054 , \9055 , RIbc62910_19, \9057 , RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$170 ( \9221 , RIdf18088_1650, \9220 );
nor \U$171 ( \9222 , RIbc62af0_23, \9053 , \9054 , \9055 , RIbc62910_19, \9057 , RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$172 ( \9223 , RIdf15388_1618, \9222 );
nor \U$173 ( \9224 , \9052 , RIbc62a78_22, \9054 , \9055 , RIbc62910_19, \9057 , RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$174 ( \9225 , RIdf12688_1586, \9224 );
nor \U$175 ( \9226 , RIbc62af0_23, RIbc62a78_22, \9054 , \9055 , RIbc62910_19, \9057 , RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$176 ( \9227 , RIdf0f988_1554, \9226 );
nor \U$177 ( \9228 , \9052 , \9053 , RIbc62a00_21, \9055 , RIbc62910_19, \9057 , RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$178 ( \9229 , RIdf0cc88_1522, \9228 );
nor \U$179 ( \9230 , RIbc62af0_23, \9053 , RIbc62a00_21, \9055 , RIbc62910_19, \9057 , RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$180 ( \9231 , RIdf09f88_1490, \9230 );
nor \U$181 ( \9232 , \9052 , RIbc62a78_22, RIbc62a00_21, \9055 , RIbc62910_19, \9057 , RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$182 ( \9233 , RIdf07288_1458, \9232 );
nor \U$183 ( \9234 , RIbc62af0_23, RIbc62a78_22, RIbc62a00_21, \9055 , RIbc62910_19, \9057 , RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$184 ( \9235 , RIdf04588_1426, \9234 );
nor \U$185 ( \9236 , \9052 , \9053 , \9054 , RIbc62988_20, RIbc62910_19, \9057 , RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$186 ( \9237 , RIdefeb88_1362, \9236 );
nor \U$187 ( \9238 , RIbc62af0_23, \9053 , \9054 , RIbc62988_20, RIbc62910_19, \9057 , RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$188 ( \9239 , RIdefbe88_1330, \9238 );
nor \U$189 ( \9240 , \9052 , RIbc62a78_22, \9054 , RIbc62988_20, RIbc62910_19, \9057 , RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$190 ( \9241 , RIdef9188_1298, \9240 );
nor \U$191 ( \9242 , RIbc62af0_23, RIbc62a78_22, \9054 , RIbc62988_20, RIbc62910_19, \9057 , RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$192 ( \9243 , RIdef6488_1266, \9242 );
nor \U$193 ( \9244 , \9052 , \9053 , RIbc62a00_21, RIbc62988_20, RIbc62910_19, \9057 , RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$194 ( \9245 , RIdef3788_1234, \9244 );
nor \U$195 ( \9246 , RIbc62af0_23, \9053 , RIbc62a00_21, RIbc62988_20, RIbc62910_19, \9057 , RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$196 ( \9247 , RIdef0a88_1202, \9246 );
nor \U$197 ( \9248 , \9052 , RIbc62a78_22, RIbc62a00_21, RIbc62988_20, RIbc62910_19, \9057 , RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$198 ( \9249 , RIdeedd88_1170, \9248 );
nor \U$199 ( \9250 , RIbc62af0_23, RIbc62a78_22, RIbc62a00_21, RIbc62988_20, RIbc62910_19, \9057 , RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$200 ( \9251 , RIdeeb088_1138, \9250 );
nor \U$201 ( \9252 , \9052 , \9053 , \9054 , \9055 , \9056 , RIbc62898_18, RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$202 ( \9253 , RIfc8efb8_6649, \9252 );
nor \U$203 ( \9254 , RIbc62af0_23, \9053 , \9054 , \9055 , \9056 , RIbc62898_18, RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$204 ( \9255 , RIfc44e40_5806, \9254 );
nor \U$205 ( \9256 , \9052 , RIbc62a78_22, \9054 , \9055 , \9056 , RIbc62898_18, RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$206 ( \9257 , RIfc57860_6018, \9256 );
nor \U$207 ( \9258 , RIbc62af0_23, RIbc62a78_22, \9054 , \9055 , \9056 , RIbc62898_18, RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$208 ( \9259 , RIfca23b0_6868, \9258 );
nor \U$209 ( \9260 , \9052 , \9053 , RIbc62a00_21, \9055 , \9056 , RIbc62898_18, RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$210 ( \9261 , RIfe9faf8_8161, \9260 );
nor \U$211 ( \9262 , RIbc62af0_23, \9053 , RIbc62a00_21, \9055 , \9056 , RIbc62898_18, RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$212 ( \9263 , RIdee3900_1053, \9262 );
nor \U$213 ( \9264 , \9052 , RIbc62a78_22, RIbc62a00_21, \9055 , \9056 , RIbc62898_18, RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$214 ( \9265 , RIdee1740_1029, \9264 );
nor \U$215 ( \9266 , RIbc62af0_23, RIbc62a78_22, RIbc62a00_21, \9055 , \9056 , RIbc62898_18, RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$216 ( \9267 , RIdedf6e8_1006, \9266 );
nor \U$217 ( \9268 , \9052 , \9053 , \9054 , RIbc62988_20, \9056 , RIbc62898_18, RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$218 ( \9269 , RIfcbd4d0_7176, \9268 );
nor \U$219 ( \9270 , RIbc62af0_23, \9053 , \9054 , RIbc62988_20, \9056 , RIbc62898_18, RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$220 ( \9271 , RIee22678_4850, \9270 );
nor \U$221 ( \9272 , \9052 , RIbc62a78_22, \9054 , RIbc62988_20, \9056 , RIbc62898_18, RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$222 ( \9273 , RIfc98090_6752, \9272 );
nor \U$223 ( \9274 , RIbc62af0_23, RIbc62a78_22, \9054 , RIbc62988_20, \9056 , RIbc62898_18, RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$224 ( \9275 , RIee21598_4838, \9274 );
nor \U$225 ( \9276 , \9052 , \9053 , RIbc62a00_21, RIbc62988_20, \9056 , RIbc62898_18, RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$226 ( \9277 , RIfe9fc60_8162, \9276 );
nor \U$227 ( \9278 , RIbc62af0_23, \9053 , RIbc62a00_21, RIbc62988_20, \9056 , RIbc62898_18, RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$228 ( \9279 , RIded80c8_922, \9278 );
nor \U$229 ( \9280 , \9052 , RIbc62a78_22, RIbc62a00_21, RIbc62988_20, \9056 , RIbc62898_18, RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$230 ( \9281 , RIfe9fdc8_8163, \9280 );
nor \U$231 ( \9282 , RIbc62af0_23, RIbc62a78_22, RIbc62a00_21, RIbc62988_20, \9056 , RIbc62898_18, RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$232 ( \9283 , RIded3be0_873, \9282 );
nor \U$233 ( \9284 , \9052 , \9053 , \9054 , \9055 , RIbc62910_19, RIbc62898_18, RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$234 ( \9285 , RIded18b8_848, \9284 );
nor \U$235 ( \9286 , RIbc62af0_23, \9053 , \9054 , \9055 , RIbc62910_19, RIbc62898_18, RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$236 ( \9287 , RIdecebb8_816, \9286 );
nor \U$237 ( \9288 , \9052 , RIbc62a78_22, \9054 , \9055 , RIbc62910_19, RIbc62898_18, RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$238 ( \9289 , RIdecbeb8_784, \9288 );
nor \U$239 ( \9290 , RIbc62af0_23, RIbc62a78_22, \9054 , \9055 , RIbc62910_19, RIbc62898_18, RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$240 ( \9291 , RIdec91b8_752, \9290 );
nor \U$241 ( \9292 , \9052 , \9053 , RIbc62a00_21, \9055 , RIbc62910_19, RIbc62898_18, RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$242 ( \9293 , RIdeb56b8_528, \9292 );
nor \U$243 ( \9294 , RIbc62af0_23, \9053 , RIbc62a00_21, \9055 , RIbc62910_19, RIbc62898_18, RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$244 ( \9295 , RIde99080_336, \9294 );
nor \U$245 ( \9296 , \9052 , RIbc62a78_22, RIbc62a00_21, \9055 , RIbc62910_19, RIbc62898_18, RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$246 ( \9297 , RIe16f2c0_2642, \9296 );
nor \U$247 ( \9298 , RIbc62af0_23, RIbc62a78_22, RIbc62a00_21, \9055 , RIbc62910_19, RIbc62898_18, RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$248 ( \9299 , RIe15b0b8_2413, \9298 );
nor \U$249 ( \9300 , \9052 , \9053 , \9054 , RIbc62988_20, RIbc62910_19, RIbc62898_18, RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$250 ( \9301 , RIe1448b8_2157, \9300 );
nor \U$251 ( \9302 , RIbc62af0_23, \9053 , \9054 , RIbc62988_20, RIbc62910_19, RIbc62898_18, RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$252 ( \9303 , RIdf392b0_2027, \9302 );
nor \U$253 ( \9304 , \9052 , RIbc62a78_22, \9054 , RIbc62988_20, RIbc62910_19, RIbc62898_18, RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$254 ( \9305 , RIdf2d910_1895, \9304 );
nor \U$255 ( \9306 , RIbc62af0_23, RIbc62a78_22, \9054 , RIbc62988_20, RIbc62910_19, RIbc62898_18, RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$256 ( \9307 , RIdf1e190_1719, \9306 );
nor \U$257 ( \9308 , \9052 , \9053 , RIbc62a00_21, RIbc62988_20, RIbc62910_19, RIbc62898_18, RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$258 ( \9309 , RIdf01888_1394, \9308 );
nor \U$259 ( \9310 , RIbc62af0_23, \9053 , RIbc62a00_21, RIbc62988_20, RIbc62910_19, RIbc62898_18, RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$260 ( \9311 , RIdee8388_1106, \9310 );
nor \U$261 ( \9312 , \9052 , RIbc62a78_22, RIbc62a00_21, RIbc62988_20, RIbc62910_19, RIbc62898_18, RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$262 ( \9313 , RIdedd0f0_979, \9312 );
nor \U$263 ( \9314 , RIbc62af0_23, RIbc62a78_22, RIbc62a00_21, RIbc62988_20, RIbc62910_19, RIbc62898_18, RIbc62820_17, RIbc627a8_16, RIbc62730_15, RIbc626b8_14, RIbc62640_13);
and \U$264 ( \9315 , RIde7efc8_209, \9314 );
or \U$265 ( \9316 , \9189 , \9191 , \9193 , \9195 , \9197 , \9199 , \9201 , \9203 , \9205 , \9207 , \9209 , \9211 , \9213 , \9215 , \9217 , \9219 , \9221 , \9223 , \9225 , \9227 , \9229 , \9231 , \9233 , \9235 , \9237 , \9239 , \9241 , \9243 , \9245 , \9247 , \9249 , \9251 , \9253 , \9255 , \9257 , \9259 , \9261 , \9263 , \9265 , \9267 , \9269 , \9271 , \9273 , \9275 , \9277 , \9279 , \9281 , \9283 , \9285 , \9287 , \9289 , \9291 , \9293 , \9295 , \9297 , \9299 , \9301 , \9303 , \9305 , \9307 , \9309 , \9311 , \9313 , \9315 );
or \U$266 ( \9317 , \9187 , \9316 );
buf \U$267 ( \9318 , RIbc627a8_16);
buf \U$268 ( \9319 , RIbc62730_15);
buf \U$269 ( \9320 , RIbc626b8_14);
buf \U$270 ( \9321 , RIbc62640_13);
or \U$271 ( \9322 , \9318 , \9319 , \9320 , \9321 );
buf \U$272 ( \9323 , \9322 );
_DC g30c1 ( \9324_nG30c1 , \9317 , \9323 );
buf \U$273 ( \9325 , \9324_nG30c1 );
not \U$274 ( \9326 , RIbc625c8_12);
not \U$275 ( \9327 , RIbc62550_11);
not \U$276 ( \9328 , RIbc624d8_10);
not \U$277 ( \9329 , RIbc62460_9);
not \U$278 ( \9330 , RIbc623e8_8);
not \U$279 ( \9331 , RIbc62370_7);
not \U$280 ( \9332 , RIbc622f8_6);
nor \U$281 ( \9333 , \9326 , \9327 , \9328 , \9329 , \9330 , \9331 , \9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$282 ( \9334 , RIe19e750_3180, \9333 );
nor \U$283 ( \9335 , RIbc625c8_12, \9327 , \9328 , \9329 , \9330 , \9331 , \9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$284 ( \9336 , RIe19ba50_3148, \9335 );
nor \U$285 ( \9337 , \9326 , RIbc62550_11, \9328 , \9329 , \9330 , \9331 , \9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$286 ( \9338 , RIfc479d8_5837, \9337 );
nor \U$287 ( \9339 , RIbc625c8_12, RIbc62550_11, \9328 , \9329 , \9330 , \9331 , \9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$288 ( \9340 , RIe198d50_3116, \9339 );
nor \U$289 ( \9341 , \9326 , \9327 , RIbc624d8_10, \9329 , \9330 , \9331 , \9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$290 ( \9342 , RIfe9f558_8157, \9341 );
nor \U$291 ( \9343 , RIbc625c8_12, \9327 , RIbc624d8_10, \9329 , \9330 , \9331 , \9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$292 ( \9344 , RIe196050_3084, \9343 );
nor \U$293 ( \9345 , \9326 , RIbc62550_11, RIbc624d8_10, \9329 , \9330 , \9331 , \9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$294 ( \9346 , RIe193350_3052, \9345 );
nor \U$295 ( \9347 , RIbc625c8_12, RIbc62550_11, RIbc624d8_10, \9329 , \9330 , \9331 , \9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$296 ( \9348 , RIe190650_3020, \9347 );
nor \U$297 ( \9349 , \9326 , \9327 , \9328 , RIbc62460_9, \9330 , \9331 , \9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$298 ( \9350 , RIe18ac50_2956, \9349 );
nor \U$299 ( \9351 , RIbc625c8_12, \9327 , \9328 , RIbc62460_9, \9330 , \9331 , \9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$300 ( \9352 , RIe187f50_2924, \9351 );
nor \U$301 ( \9353 , \9326 , RIbc62550_11, \9328 , RIbc62460_9, \9330 , \9331 , \9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$302 ( \9354 , RIfc47870_5836, \9353 );
nor \U$303 ( \9355 , RIbc625c8_12, RIbc62550_11, \9328 , RIbc62460_9, \9330 , \9331 , \9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$304 ( \9356 , RIe185250_2892, \9355 );
nor \U$305 ( \9357 , \9326 , \9327 , RIbc624d8_10, RIbc62460_9, \9330 , \9331 , \9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$306 ( \9358 , RIf142ef8_5221, \9357 );
nor \U$307 ( \9359 , RIbc625c8_12, \9327 , RIbc624d8_10, RIbc62460_9, \9330 , \9331 , \9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$308 ( \9360 , RIe182550_2860, \9359 );
nor \U$309 ( \9361 , \9326 , RIbc62550_11, RIbc624d8_10, RIbc62460_9, \9330 , \9331 , \9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$310 ( \9362 , RIe17f850_2828, \9361 );
nor \U$311 ( \9363 , RIbc625c8_12, RIbc62550_11, RIbc624d8_10, RIbc62460_9, \9330 , \9331 , \9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$312 ( \9364 , RIe17cb50_2796, \9363 );
nor \U$313 ( \9365 , \9326 , \9327 , \9328 , \9329 , RIbc623e8_8, \9331 , \9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$314 ( \9366 , RIfcb5208_7083, \9365 );
nor \U$315 ( \9367 , RIbc625c8_12, \9327 , \9328 , \9329 , RIbc623e8_8, \9331 , \9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$316 ( \9368 , RIfcbc6c0_7166, \9367 );
nor \U$317 ( \9369 , \9326 , RIbc62550_11, \9328 , \9329 , RIbc623e8_8, \9331 , \9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$318 ( \9370 , RIe177588_2735, \9369 );
nor \U$319 ( \9371 , RIbc625c8_12, RIbc62550_11, \9328 , \9329 , RIbc623e8_8, \9331 , \9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$320 ( \9372 , RIe176610_2724, \9371 );
nor \U$321 ( \9373 , \9326 , \9327 , RIbc624d8_10, \9329 , RIbc623e8_8, \9331 , \9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$322 ( \9374 , RIf13fdc0_5186, \9373 );
nor \U$323 ( \9375 , RIbc625c8_12, \9327 , RIbc624d8_10, \9329 , RIbc623e8_8, \9331 , \9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$324 ( \9376 , RIfe9f3f0_8156, \9375 );
nor \U$325 ( \9377 , \9326 , RIbc62550_11, RIbc624d8_10, \9329 , RIbc623e8_8, \9331 , \9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$326 ( \9378 , RIfce40f8_7617, \9377 );
nor \U$327 ( \9379 , RIbc625c8_12, RIbc62550_11, RIbc624d8_10, \9329 , RIbc623e8_8, \9331 , \9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$328 ( \9380 , RIfc47708_5835, \9379 );
nor \U$329 ( \9381 , \9326 , \9327 , \9328 , RIbc62460_9, RIbc623e8_8, \9331 , \9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$330 ( \9382 , RIfc47438_5833, \9381 );
nor \U$331 ( \9383 , RIbc625c8_12, \9327 , \9328 , RIbc62460_9, RIbc623e8_8, \9331 , \9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$332 ( \9384 , RIfca15a0_6858, \9383 );
nor \U$333 ( \9385 , \9326 , RIbc62550_11, \9328 , RIbc62460_9, RIbc623e8_8, \9331 , \9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$334 ( \9386 , RIfc99170_6764, \9385 );
nor \U$335 ( \9387 , RIbc625c8_12, RIbc62550_11, \9328 , RIbc62460_9, RIbc623e8_8, \9331 , \9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$336 ( \9388 , RIe1745b8_2701, \9387 );
nor \U$337 ( \9389 , \9326 , \9327 , RIbc624d8_10, RIbc62460_9, RIbc623e8_8, \9331 , \9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$338 ( \9390 , RIfc8cc90_6624, \9389 );
nor \U$339 ( \9391 , RIbc625c8_12, \9327 , RIbc624d8_10, RIbc62460_9, RIbc623e8_8, \9331 , \9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$340 ( \9392 , RIfc556a0_5994, \9391 );
nor \U$341 ( \9393 , \9326 , RIbc62550_11, RIbc624d8_10, RIbc62460_9, RIbc623e8_8, \9331 , \9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$342 ( \9394 , RIfc7ee60_6466, \9393 );
nor \U$343 ( \9395 , RIbc625c8_12, RIbc62550_11, RIbc624d8_10, RIbc62460_9, RIbc623e8_8, \9331 , \9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$344 ( \9396 , RIfce8e50_7672, \9395 );
nor \U$345 ( \9397 , \9326 , \9327 , \9328 , \9329 , \9330 , RIbc62370_7, \9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$346 ( \9398 , RIfe9f288_8155, \9397 );
nor \U$347 ( \9399 , RIbc625c8_12, \9327 , \9328 , \9329 , \9330 , RIbc62370_7, \9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$348 ( \9400 , RIe224aa8_4707, \9399 );
nor \U$349 ( \9401 , \9326 , RIbc62550_11, \9328 , \9329 , \9330 , RIbc62370_7, \9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$350 ( \9402 , RIfc55808_5995, \9401 );
nor \U$351 ( \9403 , RIbc625c8_12, RIbc62550_11, \9328 , \9329 , \9330 , RIbc62370_7, \9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$352 ( \9404 , RIe221da8_4675, \9403 );
nor \U$353 ( \9405 , \9326 , \9327 , RIbc624d8_10, \9329 , \9330 , RIbc62370_7, \9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$354 ( \9406 , RIfcb50a0_7082, \9405 );
nor \U$355 ( \9407 , RIbc625c8_12, \9327 , RIbc624d8_10, \9329 , \9330 , RIbc62370_7, \9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$356 ( \9408 , RIe21f0a8_4643, \9407 );
nor \U$357 ( \9409 , \9326 , RIbc62550_11, RIbc624d8_10, \9329 , \9330 , RIbc62370_7, \9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$358 ( \9410 , RIe2196a8_4579, \9409 );
nor \U$359 ( \9411 , RIbc625c8_12, RIbc62550_11, RIbc624d8_10, \9329 , \9330 , RIbc62370_7, \9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$360 ( \9412 , RIe2169a8_4547, \9411 );
nor \U$361 ( \9413 , \9326 , \9327 , \9328 , RIbc62460_9, \9330 , RIbc62370_7, \9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$362 ( \9414 , RIfcbc828_7167, \9413 );
nor \U$363 ( \9415 , RIbc625c8_12, \9327 , \9328 , RIbc62460_9, \9330 , RIbc62370_7, \9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$364 ( \9416 , RIe213ca8_4515, \9415 );
nor \U$365 ( \9417 , \9326 , RIbc62550_11, \9328 , RIbc62460_9, \9330 , RIbc62370_7, \9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$366 ( \9418 , RIfc47000_5830, \9417 );
nor \U$367 ( \9419 , RIbc625c8_12, RIbc62550_11, \9328 , RIbc62460_9, \9330 , RIbc62370_7, \9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$368 ( \9420 , RIe210fa8_4483, \9419 );
nor \U$369 ( \9421 , \9326 , \9327 , RIbc624d8_10, RIbc62460_9, \9330 , RIbc62370_7, \9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$370 ( \9422 , RIfcbc990_7168, \9421 );
nor \U$371 ( \9423 , RIbc625c8_12, \9327 , RIbc624d8_10, RIbc62460_9, \9330 , RIbc62370_7, \9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$372 ( \9424 , RIe20e2a8_4451, \9423 );
nor \U$373 ( \9425 , \9326 , RIbc62550_11, RIbc624d8_10, RIbc62460_9, \9330 , RIbc62370_7, \9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$374 ( \9426 , RIe20b5a8_4419, \9425 );
nor \U$375 ( \9427 , RIbc625c8_12, RIbc62550_11, RIbc624d8_10, RIbc62460_9, \9330 , RIbc62370_7, \9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$376 ( \9428 , RIe2088a8_4387, \9427 );
nor \U$377 ( \9429 , \9326 , \9327 , \9328 , \9329 , RIbc623e8_8, RIbc62370_7, \9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$378 ( \9430 , RIfc46bc8_5827, \9429 );
nor \U$379 ( \9431 , RIbc625c8_12, \9327 , \9328 , \9329 , RIbc623e8_8, RIbc62370_7, \9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$380 ( \9432 , RIfcd6598_7461, \9431 );
nor \U$381 ( \9433 , \9326 , RIbc62550_11, \9328 , \9329 , RIbc623e8_8, RIbc62370_7, \9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$382 ( \9434 , RIe2032e0_4326, \9433 );
nor \U$383 ( \9435 , RIbc625c8_12, RIbc62550_11, \9328 , \9329 , RIbc623e8_8, RIbc62370_7, \9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$384 ( \9436 , RIe2016c0_4306, \9435 );
nor \U$385 ( \9437 , \9326 , \9327 , RIbc624d8_10, \9329 , RIbc623e8_8, RIbc62370_7, \9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$386 ( \9438 , RIfc98ea0_6762, \9437 );
nor \U$387 ( \9439 , RIbc625c8_12, \9327 , RIbc624d8_10, \9329 , RIbc623e8_8, RIbc62370_7, \9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$388 ( \9440 , RIfc7eb90_6464, \9439 );
nor \U$389 ( \9441 , \9326 , RIbc62550_11, RIbc624d8_10, \9329 , RIbc623e8_8, RIbc62370_7, \9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$390 ( \9442 , RIfce0318_7573, \9441 );
nor \U$391 ( \9443 , RIbc625c8_12, RIbc62550_11, RIbc624d8_10, \9329 , RIbc623e8_8, RIbc62370_7, \9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$392 ( \9444 , RIfcbcaf8_7169, \9443 );
nor \U$393 ( \9445 , \9326 , \9327 , \9328 , RIbc62460_9, RIbc623e8_8, RIbc62370_7, \9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$394 ( \9446 , RIfc8cf60_6626, \9445 );
nor \U$395 ( \9447 , RIbc625c8_12, \9327 , \9328 , RIbc62460_9, RIbc623e8_8, RIbc62370_7, \9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$396 ( \9448 , RIfcb4dd0_7080, \9447 );
nor \U$397 ( \9449 , \9326 , RIbc62550_11, \9328 , RIbc62460_9, RIbc623e8_8, RIbc62370_7, \9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$398 ( \9450 , RIe1fd340_4258, \9449 );
nor \U$399 ( \9451 , RIbc625c8_12, RIbc62550_11, \9328 , RIbc62460_9, RIbc623e8_8, RIbc62370_7, \9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$400 ( \9452 , RIe1fc260_4246, \9451 );
nor \U$401 ( \9453 , \9326 , \9327 , RIbc624d8_10, RIbc62460_9, RIbc623e8_8, RIbc62370_7, \9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$402 ( \9454 , RIf15cf38_5517, \9453 );
nor \U$403 ( \9455 , RIbc625c8_12, \9327 , RIbc624d8_10, RIbc62460_9, RIbc623e8_8, RIbc62370_7, \9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$404 ( \9456 , RIfe9f120_8154, \9455 );
nor \U$405 ( \9457 , \9326 , RIbc62550_11, RIbc624d8_10, RIbc62460_9, RIbc623e8_8, RIbc62370_7, \9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$406 ( \9458 , RIfc7ea28_6463, \9457 );
nor \U$407 ( \9459 , RIbc625c8_12, RIbc62550_11, RIbc624d8_10, RIbc62460_9, RIbc623e8_8, RIbc62370_7, \9332 , RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$408 ( \9460 , RIfc8d0c8_6627, \9459 );
or \U$409 ( \9461 , \9334 , \9336 , \9338 , \9340 , \9342 , \9344 , \9346 , \9348 , \9350 , \9352 , \9354 , \9356 , \9358 , \9360 , \9362 , \9364 , \9366 , \9368 , \9370 , \9372 , \9374 , \9376 , \9378 , \9380 , \9382 , \9384 , \9386 , \9388 , \9390 , \9392 , \9394 , \9396 , \9398 , \9400 , \9402 , \9404 , \9406 , \9408 , \9410 , \9412 , \9414 , \9416 , \9418 , \9420 , \9422 , \9424 , \9426 , \9428 , \9430 , \9432 , \9434 , \9436 , \9438 , \9440 , \9442 , \9444 , \9446 , \9448 , \9450 , \9452 , \9454 , \9456 , \9458 , \9460 );
nor \U$410 ( \9462 , \9326 , \9327 , \9328 , \9329 , \9330 , \9331 , RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$411 ( \9463 , RIfcbcc60_7170, \9462 );
nor \U$412 ( \9464 , RIbc625c8_12, \9327 , \9328 , \9329 , \9330 , \9331 , RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$413 ( \9465 , RIfc98bd0_6760, \9464 );
nor \U$414 ( \9466 , \9326 , RIbc62550_11, \9328 , \9329 , \9330 , \9331 , RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$415 ( \9467 , RIfce2d48_7603, \9466 );
nor \U$416 ( \9468 , RIbc625c8_12, RIbc62550_11, \9328 , \9329 , \9330 , \9331 , RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$417 ( \9469 , RIe1fb018_4233, \9468 );
nor \U$418 ( \9470 , \9326 , \9327 , RIbc624d8_10, \9329 , \9330 , \9331 , RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$419 ( \9471 , RIfc55f10_6000, \9470 );
nor \U$420 ( \9472 , RIbc625c8_12, \9327 , RIbc624d8_10, \9329 , \9330 , \9331 , RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$421 ( \9473 , RIfc7e8c0_6462, \9472 );
nor \U$422 ( \9474 , \9326 , RIbc62550_11, RIbc624d8_10, \9329 , \9330 , \9331 , RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$423 ( \9475 , RIfc8d230_6628, \9474 );
nor \U$424 ( \9476 , RIbc625c8_12, RIbc62550_11, RIbc624d8_10, \9329 , \9330 , \9331 , RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$425 ( \9477 , RIe1f6590_4180, \9476 );
nor \U$426 ( \9478 , \9326 , \9327 , \9328 , RIbc62460_9, \9330 , \9331 , RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$427 ( \9479 , RIfce58e0_7634, \9478 );
nor \U$428 ( \9480 , RIbc625c8_12, \9327 , \9328 , RIbc62460_9, \9330 , \9331 , RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$429 ( \9481 , RIfc468f8_5825, \9480 );
nor \U$430 ( \9482 , \9326 , RIbc62550_11, \9328 , RIbc62460_9, \9330 , \9331 , RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$431 ( \9483 , RIfcc2ed0_7240, \9482 );
nor \U$432 ( \9484 , RIbc625c8_12, RIbc62550_11, \9328 , RIbc62460_9, \9330 , \9331 , RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$433 ( \9485 , RIe1f4100_4154, \9484 );
nor \U$434 ( \9486 , \9326 , \9327 , RIbc624d8_10, RIbc62460_9, \9330 , \9331 , RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$435 ( \9487 , RIfceedf0_7740, \9486 );
nor \U$436 ( \9488 , RIbc625c8_12, \9327 , RIbc624d8_10, RIbc62460_9, \9330 , \9331 , RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$437 ( \9489 , RIfc8d398_6629, \9488 );
nor \U$438 ( \9490 , \9326 , RIbc62550_11, RIbc624d8_10, RIbc62460_9, \9330 , \9331 , RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$439 ( \9491 , RIfc8d500_6630, \9490 );
nor \U$440 ( \9492 , RIbc625c8_12, RIbc62550_11, RIbc624d8_10, RIbc62460_9, \9330 , \9331 , RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$441 ( \9493 , RIe1eef70_4096, \9492 );
nor \U$442 ( \9494 , \9326 , \9327 , \9328 , \9329 , RIbc623e8_8, \9331 , RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$443 ( \9495 , RIe1ec810_4068, \9494 );
nor \U$444 ( \9496 , RIbc625c8_12, \9327 , \9328 , \9329 , RIbc623e8_8, \9331 , RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$445 ( \9497 , RIe1e9b10_4036, \9496 );
nor \U$446 ( \9498 , \9326 , RIbc62550_11, \9328 , \9329 , RIbc623e8_8, \9331 , RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$447 ( \9499 , RIe1e6e10_4004, \9498 );
nor \U$448 ( \9500 , RIbc625c8_12, RIbc62550_11, \9328 , \9329 , RIbc623e8_8, \9331 , RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$449 ( \9501 , RIe1e4110_3972, \9500 );
nor \U$450 ( \9502 , \9326 , \9327 , RIbc624d8_10, \9329 , RIbc623e8_8, \9331 , RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$451 ( \9503 , RIe1e1410_3940, \9502 );
nor \U$452 ( \9504 , RIbc625c8_12, \9327 , RIbc624d8_10, \9329 , RIbc623e8_8, \9331 , RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$453 ( \9505 , RIe1de710_3908, \9504 );
nor \U$454 ( \9506 , \9326 , RIbc62550_11, RIbc624d8_10, \9329 , RIbc623e8_8, \9331 , RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$455 ( \9507 , RIe1dba10_3876, \9506 );
nor \U$456 ( \9508 , RIbc625c8_12, RIbc62550_11, RIbc624d8_10, \9329 , RIbc623e8_8, \9331 , RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$457 ( \9509 , RIe1d8d10_3844, \9508 );
nor \U$458 ( \9510 , \9326 , \9327 , \9328 , RIbc62460_9, RIbc623e8_8, \9331 , RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$459 ( \9511 , RIe1d3310_3780, \9510 );
nor \U$460 ( \9512 , RIbc625c8_12, \9327 , \9328 , RIbc62460_9, RIbc623e8_8, \9331 , RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$461 ( \9513 , RIe1d0610_3748, \9512 );
nor \U$462 ( \9514 , \9326 , RIbc62550_11, \9328 , RIbc62460_9, RIbc623e8_8, \9331 , RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$463 ( \9515 , RIe1cd910_3716, \9514 );
nor \U$464 ( \9516 , RIbc625c8_12, RIbc62550_11, \9328 , RIbc62460_9, RIbc623e8_8, \9331 , RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$465 ( \9517 , RIe1cac10_3684, \9516 );
nor \U$466 ( \9518 , \9326 , \9327 , RIbc624d8_10, RIbc62460_9, RIbc623e8_8, \9331 , RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$467 ( \9519 , RIe1c7f10_3652, \9518 );
nor \U$468 ( \9520 , RIbc625c8_12, \9327 , RIbc624d8_10, RIbc62460_9, RIbc623e8_8, \9331 , RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$469 ( \9521 , RIe1c5210_3620, \9520 );
nor \U$470 ( \9522 , \9326 , RIbc62550_11, RIbc624d8_10, RIbc62460_9, RIbc623e8_8, \9331 , RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$471 ( \9523 , RIe1c2510_3588, \9522 );
nor \U$472 ( \9524 , RIbc625c8_12, RIbc62550_11, RIbc624d8_10, RIbc62460_9, RIbc623e8_8, \9331 , RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$473 ( \9525 , RIe1bf810_3556, \9524 );
nor \U$474 ( \9526 , \9326 , \9327 , \9328 , \9329 , \9330 , RIbc62370_7, RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$475 ( \9527 , RIf14d0b0_5336, \9526 );
nor \U$476 ( \9528 , RIbc625c8_12, \9327 , \9328 , \9329 , \9330 , RIbc62370_7, RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$477 ( \9529 , RIfe9efb8_8153, \9528 );
nor \U$478 ( \9530 , \9326 , RIbc62550_11, \9328 , \9329 , \9330 , RIbc62370_7, RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$479 ( \9531 , RIe1ba248_3495, \9530 );
nor \U$480 ( \9532 , RIbc625c8_12, RIbc62550_11, \9328 , \9329 , \9330 , RIbc62370_7, RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$481 ( \9533 , RIe1b8088_3471, \9532 );
nor \U$482 ( \9534 , \9326 , \9327 , RIbc624d8_10, \9329 , \9330 , RIbc62370_7, RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$483 ( \9535 , RIfec4dd0_8360, \9534 );
nor \U$484 ( \9536 , RIbc625c8_12, \9327 , RIbc624d8_10, \9329 , \9330 , RIbc62370_7, RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$485 ( \9537 , RIfec50a0_8362, \9536 );
nor \U$486 ( \9538 , \9326 , RIbc62550_11, RIbc624d8_10, \9329 , \9330 , RIbc62370_7, RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$487 ( \9539 , RIe1b5ec8_3447, \9538 );
nor \U$488 ( \9540 , RIbc625c8_12, RIbc62550_11, RIbc624d8_10, \9329 , \9330 , RIbc62370_7, RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$489 ( \9541 , RIe1b46e0_3430, \9540 );
nor \U$490 ( \9542 , \9326 , \9327 , \9328 , RIbc62460_9, \9330 , RIbc62370_7, RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$491 ( \9543 , RIfcb4998_7077, \9542 );
nor \U$492 ( \9544 , RIbc625c8_12, \9327 , \9328 , RIbc62460_9, \9330 , RIbc62370_7, RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$493 ( \9545 , RIfcb4c68_7079, \9544 );
nor \U$494 ( \9546 , \9326 , RIbc62550_11, \9328 , RIbc62460_9, \9330 , RIbc62370_7, RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$495 ( \9547 , RIfec5370_8364, \9546 );
nor \U$496 ( \9548 , RIbc625c8_12, RIbc62550_11, \9328 , RIbc62460_9, \9330 , RIbc62370_7, RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$497 ( \9549 , RIfe9ee50_8152, \9548 );
nor \U$498 ( \9550 , \9326 , \9327 , RIbc624d8_10, RIbc62460_9, \9330 , RIbc62370_7, RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$499 ( \9551 , RIfcbcdc8_7171, \9550 );
nor \U$500 ( \9552 , RIbc625c8_12, \9327 , RIbc624d8_10, RIbc62460_9, \9330 , RIbc62370_7, RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$501 ( \9553 , RIfc46358_5821, \9552 );
nor \U$502 ( \9554 , \9326 , RIbc62550_11, RIbc624d8_10, RIbc62460_9, \9330 , RIbc62370_7, RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$503 ( \9555 , RIfec5208_8363, \9554 );
nor \U$504 ( \9556 , RIbc625c8_12, RIbc62550_11, RIbc624d8_10, RIbc62460_9, \9330 , RIbc62370_7, RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$505 ( \9557 , RIfec4f38_8361, \9556 );
nor \U$506 ( \9558 , \9326 , \9327 , \9328 , \9329 , RIbc623e8_8, RIbc62370_7, RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$507 ( \9559 , RIe1a9b50_3308, \9558 );
nor \U$508 ( \9560 , RIbc625c8_12, \9327 , \9328 , \9329 , RIbc623e8_8, RIbc62370_7, RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$509 ( \9561 , RIe1a6e50_3276, \9560 );
nor \U$510 ( \9562 , \9326 , RIbc62550_11, \9328 , \9329 , RIbc623e8_8, RIbc62370_7, RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$511 ( \9563 , RIe1a4150_3244, \9562 );
nor \U$512 ( \9564 , RIbc625c8_12, RIbc62550_11, \9328 , \9329 , RIbc623e8_8, RIbc62370_7, RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$513 ( \9565 , RIe1a1450_3212, \9564 );
nor \U$514 ( \9566 , \9326 , \9327 , RIbc624d8_10, \9329 , RIbc623e8_8, RIbc62370_7, RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$515 ( \9567 , RIe18d950_2988, \9566 );
nor \U$516 ( \9568 , RIbc625c8_12, \9327 , RIbc624d8_10, \9329 , RIbc623e8_8, RIbc62370_7, RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$517 ( \9569 , RIe179e50_2764, \9568 );
nor \U$518 ( \9570 , \9326 , RIbc62550_11, RIbc624d8_10, \9329 , RIbc623e8_8, RIbc62370_7, RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$519 ( \9571 , RIe2277a8_4739, \9570 );
nor \U$520 ( \9572 , RIbc625c8_12, RIbc62550_11, RIbc624d8_10, \9329 , RIbc623e8_8, RIbc62370_7, RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$521 ( \9573 , RIe21c3a8_4611, \9572 );
nor \U$522 ( \9574 , \9326 , \9327 , \9328 , RIbc62460_9, RIbc623e8_8, RIbc62370_7, RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$523 ( \9575 , RIe205ba8_4355, \9574 );
nor \U$524 ( \9576 , RIbc625c8_12, \9327 , \9328 , RIbc62460_9, RIbc623e8_8, RIbc62370_7, RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$525 ( \9577 , RIe1ffc08_4287, \9576 );
nor \U$526 ( \9578 , \9326 , RIbc62550_11, \9328 , RIbc62460_9, RIbc623e8_8, RIbc62370_7, RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$527 ( \9579 , RIe1f8fc0_4210, \9578 );
nor \U$528 ( \9580 , RIbc625c8_12, RIbc62550_11, \9328 , RIbc62460_9, RIbc623e8_8, RIbc62370_7, RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$529 ( \9581 , RIe1f1b08_4127, \9580 );
nor \U$530 ( \9582 , \9326 , \9327 , RIbc624d8_10, RIbc62460_9, RIbc623e8_8, RIbc62370_7, RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$531 ( \9583 , RIe1d6010_3812, \9582 );
nor \U$532 ( \9584 , RIbc625c8_12, \9327 , RIbc624d8_10, RIbc62460_9, RIbc623e8_8, RIbc62370_7, RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$533 ( \9585 , RIe1bcb10_3524, \9584 );
nor \U$534 ( \9586 , \9326 , RIbc62550_11, RIbc624d8_10, RIbc62460_9, RIbc623e8_8, RIbc62370_7, RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$535 ( \9587 , RIe1af988_3375, \9586 );
nor \U$536 ( \9588 , RIbc625c8_12, RIbc62550_11, RIbc624d8_10, RIbc62460_9, RIbc623e8_8, RIbc62370_7, RIbc622f8_6, RIbc62280_5, RIbc62208_4, RIbc62190_3, RIbc62118_2);
and \U$537 ( \9589 , RIe171fc0_2674, \9588 );
or \U$538 ( \9590 , \9463 , \9465 , \9467 , \9469 , \9471 , \9473 , \9475 , \9477 , \9479 , \9481 , \9483 , \9485 , \9487 , \9489 , \9491 , \9493 , \9495 , \9497 , \9499 , \9501 , \9503 , \9505 , \9507 , \9509 , \9511 , \9513 , \9515 , \9517 , \9519 , \9521 , \9523 , \9525 , \9527 , \9529 , \9531 , \9533 , \9535 , \9537 , \9539 , \9541 , \9543 , \9545 , \9547 , \9549 , \9551 , \9553 , \9555 , \9557 , \9559 , \9561 , \9563 , \9565 , \9567 , \9569 , \9571 , \9573 , \9575 , \9577 , \9579 , \9581 , \9583 , \9585 , \9587 , \9589 );
or \U$539 ( \9591 , \9461 , \9590 );
buf \U$540 ( \9592 , RIbc62280_5);
buf \U$541 ( \9593 , RIbc62208_4);
buf \U$542 ( \9594 , RIbc62190_3);
buf \U$543 ( \9595 , RIbc62118_2);
or \U$544 ( \9596 , \9592 , \9593 , \9594 , \9595 );
buf \U$545 ( \9597 , \9596 );
_DC g41ee ( \9598_nG41ee , \9591 , \9597 );
buf \U$546 ( \9599 , \9598_nG41ee );
xor \U$547 ( \9600 , \9325 , \9599 );
and \U$548 ( \9601 , RIdec6080_717, \9059 );
and \U$549 ( \9602 , RIdec3380_685, \9061 );
and \U$550 ( \9603 , RIee204b8_4826, \9063 );
and \U$551 ( \9604 , RIdec0680_653, \9065 );
and \U$552 ( \9605 , RIfcd70d8_7469, \9067 );
and \U$553 ( \9606 , RIdebd980_621, \9069 );
and \U$554 ( \9607 , RIdebac80_589, \9071 );
and \U$555 ( \9608 , RIdeb7f80_557, \9073 );
and \U$556 ( \9609 , RIfcbe448_7187, \9075 );
and \U$557 ( \9610 , RIdeb2580_493, \9077 );
and \U$558 ( \9611 , RIfcb3480_7062, \9079 );
and \U$559 ( \9612 , RIdeaf880_461, \9081 );
and \U$560 ( \9613 , RIfc43928_5791, \9083 );
and \U$561 ( \9614 , RIdeac1a8_429, \9085 );
and \U$562 ( \9615 , RIdea58a8_397, \9087 );
and \U$563 ( \9616 , RIde9efa8_365, \9089 );
and \U$564 ( \9617 , RIfcd88c0_7486, \9091 );
and \U$565 ( \9618 , RIee1c408_4780, \9093 );
and \U$566 ( \9619 , RIfcc77f0_7292, \9095 );
and \U$567 ( \9620 , RIfea04d0_8168, \9097 );
and \U$568 ( \9621 , RIde92438_303, \9099 );
and \U$569 ( \9622 , RIde8ec70_286, \9101 );
and \U$570 ( \9623 , RIde8aad0_266, \9103 );
and \U$571 ( \9624 , RIde86930_246, \9105 );
and \U$572 ( \9625 , RIfca31c0_6878, \9107 );
and \U$573 ( \9626 , RIfc59a20_6042, \9109 );
and \U$574 ( \9627 , RIfcd1de0_7410, \9111 );
and \U$575 ( \9628 , RIfc91448_6675, \9113 );
and \U$576 ( \9629 , RIfc97280_6742, \9115 );
and \U$577 ( \9630 , RIe16c188_2607, \9117 );
and \U$578 ( \9631 , RIfc97118_6741, \9119 );
and \U$579 ( \9632 , RIe168948_2567, \9121 );
and \U$580 ( \9633 , RIe166080_2538, \9123 );
and \U$581 ( \9634 , RIe163380_2506, \9125 );
and \U$582 ( \9635 , RIee37ac8_5092, \9127 );
and \U$583 ( \9636 , RIe160680_2474, \9129 );
and \U$584 ( \9637 , RIfcd1c78_7409, \9131 );
and \U$585 ( \9638 , RIe15d980_2442, \9133 );
and \U$586 ( \9639 , RIe157f80_2378, \9135 );
and \U$587 ( \9640 , RIe155280_2346, \9137 );
and \U$588 ( \9641 , RIfc3f530_5746, \9139 );
and \U$589 ( \9642 , RIe152580_2314, \9141 );
and \U$590 ( \9643 , RIee35368_5064, \9143 );
and \U$591 ( \9644 , RIe14f880_2282, \9145 );
and \U$592 ( \9645 , RIfc7a3d8_6413, \9147 );
and \U$593 ( \9646 , RIe14cb80_2250, \9149 );
and \U$594 ( \9647 , RIe149e80_2218, \9151 );
and \U$595 ( \9648 , RIe147180_2186, \9153 );
and \U$596 ( \9649 , RIfc42b18_5781, \9155 );
and \U$597 ( \9650 , RIfc7a270_6412, \9157 );
and \U$598 ( \9651 , RIfc5a560_6050, \9159 );
and \U$599 ( \9652 , RIfc96b78_6737, \9161 );
and \U$600 ( \9653 , RIfea6fb0_8216, \9163 );
and \U$601 ( \9654 , RIe13f5c0_2098, \9165 );
and \U$602 ( \9655 , RIdf3d4c8_2074, \9167 );
and \U$603 ( \9656 , RIdf3b038_2048, \9169 );
and \U$604 ( \9657 , RIfce5bb0_7636, \9171 );
and \U$605 ( \9658 , RIee2fc38_5002, \9173 );
and \U$606 ( \9659 , RIfc91cb8_6681, \9175 );
and \U$607 ( \9660 , RIee2d910_4977, \9177 );
and \U$608 ( \9661 , RIdf362e0_1993, \9179 );
and \U$609 ( \9662 , RIdf33e50_1967, \9181 );
and \U$610 ( \9663 , RIdf31c90_1943, \9183 );
and \U$611 ( \9664 , RIdf2fda0_1921, \9185 );
or \U$612 ( \9665 , \9601 , \9602 , \9603 , \9604 , \9605 , \9606 , \9607 , \9608 , \9609 , \9610 , \9611 , \9612 , \9613 , \9614 , \9615 , \9616 , \9617 , \9618 , \9619 , \9620 , \9621 , \9622 , \9623 , \9624 , \9625 , \9626 , \9627 , \9628 , \9629 , \9630 , \9631 , \9632 , \9633 , \9634 , \9635 , \9636 , \9637 , \9638 , \9639 , \9640 , \9641 , \9642 , \9643 , \9644 , \9645 , \9646 , \9647 , \9648 , \9649 , \9650 , \9651 , \9652 , \9653 , \9654 , \9655 , \9656 , \9657 , \9658 , \9659 , \9660 , \9661 , \9662 , \9663 , \9664 );
and \U$613 ( \9666 , RIfc43658_5789, \9188 );
and \U$614 ( \9667 , RIfc59e58_6045, \9190 );
and \U$615 ( \9668 , RIfc96fb0_6740, \9192 );
and \U$616 ( \9669 , RIfc7ac48_6419, \9194 );
and \U$617 ( \9670 , RIfea0368_8167, \9196 );
and \U$618 ( \9671 , RIdf28bb8_1840, \9198 );
and \U$619 ( \9672 , RIdf26cc8_1818, \9200 );
and \U$620 ( \9673 , RIdf25210_1799, \9202 );
and \U$621 ( \9674 , RIfc91718_6677, \9204 );
and \U$622 ( \9675 , RIfcb3318_7061, \9206 );
and \U$623 ( \9676 , RIfc919e8_6679, \9208 );
and \U$624 ( \9677 , RIfc91880_6678, \9210 );
and \U$625 ( \9678 , RIfc430b8_5785, \9212 );
and \U$626 ( \9679 , RIdf20350_1743, \9214 );
and \U$627 ( \9680 , RIfc7a978_6417, \9216 );
and \U$628 ( \9681 , RIdf19e10_1671, \9218 );
and \U$629 ( \9682 , RIdf17c50_1647, \9220 );
and \U$630 ( \9683 , RIdf14f50_1615, \9222 );
and \U$631 ( \9684 , RIdf12250_1583, \9224 );
and \U$632 ( \9685 , RIdf0f550_1551, \9226 );
and \U$633 ( \9686 , RIdf0c850_1519, \9228 );
and \U$634 ( \9687 , RIdf09b50_1487, \9230 );
and \U$635 ( \9688 , RIdf06e50_1455, \9232 );
and \U$636 ( \9689 , RIdf04150_1423, \9234 );
and \U$637 ( \9690 , RIdefe750_1359, \9236 );
and \U$638 ( \9691 , RIdefba50_1327, \9238 );
and \U$639 ( \9692 , RIdef8d50_1295, \9240 );
and \U$640 ( \9693 , RIdef6050_1263, \9242 );
and \U$641 ( \9694 , RIdef3350_1231, \9244 );
and \U$642 ( \9695 , RIdef0650_1199, \9246 );
and \U$643 ( \9696 , RIdeed950_1167, \9248 );
and \U$644 ( \9697 , RIdeeac50_1135, \9250 );
and \U$645 ( \9698 , RIfcd1b10_7408, \9252 );
and \U$646 ( \9699 , RIfc968a8_6735, \9254 );
and \U$647 ( \9700 , RIfc91f88_6683, \9256 );
and \U$648 ( \9701 , RIfcdfc10_7568, \9258 );
and \U$649 ( \9702 , RIfea99e0_8246, \9260 );
and \U$650 ( \9703 , RIdee3630_1051, \9262 );
and \U$651 ( \9704 , RIdee1308_1026, \9264 );
and \U$652 ( \9705 , RIdedf2b0_1003, \9266 );
and \U$653 ( \9706 , RIfcc7d90_7296, \9268 );
and \U$654 ( \9707 , RIfcd85f0_7484, \9270 );
and \U$655 ( \9708 , RIfce3888_7611, \9272 );
and \U$656 ( \9709 , RIfc5a830_6052, \9274 );
and \U$657 ( \9710 , RIdeda3f0_947, \9276 );
and \U$658 ( \9711 , RIfea9878_8245, \9278 );
and \U$659 ( \9712 , RIded5f08_898, \9280 );
and \U$660 ( \9713 , RIded37a8_870, \9282 );
and \U$661 ( \9714 , RIded1480_845, \9284 );
and \U$662 ( \9715 , RIdece780_813, \9286 );
and \U$663 ( \9716 , RIdecba80_781, \9288 );
and \U$664 ( \9717 , RIdec8d80_749, \9290 );
and \U$665 ( \9718 , RIdeb5280_525, \9292 );
and \U$666 ( \9719 , RIde986a8_333, \9294 );
and \U$667 ( \9720 , RIe16ee88_2639, \9296 );
and \U$668 ( \9721 , RIe15ac80_2410, \9298 );
and \U$669 ( \9722 , RIe144480_2154, \9300 );
and \U$670 ( \9723 , RIdf38e78_2024, \9302 );
and \U$671 ( \9724 , RIdf2d4d8_1892, \9304 );
and \U$672 ( \9725 , RIdf1dd58_1716, \9306 );
and \U$673 ( \9726 , RIdf01450_1391, \9308 );
and \U$674 ( \9727 , RIdee7f50_1103, \9310 );
and \U$675 ( \9728 , RIdedccb8_976, \9312 );
and \U$676 ( \9729 , RIde7e5f0_206, \9314 );
or \U$677 ( \9730 , \9666 , \9667 , \9668 , \9669 , \9670 , \9671 , \9672 , \9673 , \9674 , \9675 , \9676 , \9677 , \9678 , \9679 , \9680 , \9681 , \9682 , \9683 , \9684 , \9685 , \9686 , \9687 , \9688 , \9689 , \9690 , \9691 , \9692 , \9693 , \9694 , \9695 , \9696 , \9697 , \9698 , \9699 , \9700 , \9701 , \9702 , \9703 , \9704 , \9705 , \9706 , \9707 , \9708 , \9709 , \9710 , \9711 , \9712 , \9713 , \9714 , \9715 , \9716 , \9717 , \9718 , \9719 , \9720 , \9721 , \9722 , \9723 , \9724 , \9725 , \9726 , \9727 , \9728 , \9729 );
or \U$678 ( \9731 , \9665 , \9730 );
_DC g3146 ( \9732_nG3146 , \9731 , \9323 );
buf \U$679 ( \9733 , \9732_nG3146 );
and \U$680 ( \9734 , RIe19e318_3177, \9333 );
and \U$681 ( \9735 , RIe19b618_3145, \9335 );
and \U$682 ( \9736 , RIfc8f3f0_6652, \9337 );
and \U$683 ( \9737 , RIe198918_3113, \9339 );
and \U$684 ( \9738 , RIf144b18_5241, \9341 );
and \U$685 ( \9739 , RIe195c18_3081, \9343 );
and \U$686 ( \9740 , RIe192f18_3049, \9345 );
and \U$687 ( \9741 , RIe190218_3017, \9347 );
and \U$688 ( \9742 , RIe18a818_2953, \9349 );
and \U$689 ( \9743 , RIe187b18_2921, \9351 );
and \U$690 ( \9744 , RIf143d08_5231, \9353 );
and \U$691 ( \9745 , RIe184e18_2889, \9355 );
and \U$692 ( \9746 , RIfcb3cf0_7068, \9357 );
and \U$693 ( \9747 , RIe182118_2857, \9359 );
and \U$694 ( \9748 , RIe17f418_2825, \9361 );
and \U$695 ( \9749 , RIe17c718_2793, \9363 );
and \U$696 ( \9750 , RIfc448a0_5802, \9365 );
and \U$697 ( \9751 , RIf141170_5200, \9367 );
and \U$698 ( \9752 , RIfc7c9d0_6440, \9369 );
and \U$699 ( \9753 , RIfea0098_8165, \9371 );
and \U$700 ( \9754 , RIfc57e00_6022, \9373 );
and \U$701 ( \9755 , RIf13f550_5180, \9375 );
and \U$702 ( \9756 , RIfcd6e08_7467, \9377 );
and \U$703 ( \9757 , RIee3d900_5159, \9379 );
and \U$704 ( \9758 , RIfc8f6c0_6654, \9381 );
and \U$705 ( \9759 , RIfce0048_7571, \9383 );
and \U$706 ( \9760 , RIfca27e8_6871, \9385 );
and \U$707 ( \9761 , RIe1742e8_2699, \9387 );
and \U$708 ( \9762 , RIfc7c700_6438, \9389 );
and \U$709 ( \9763 , RIfc8f990_6656, \9391 );
and \U$710 ( \9764 , RIfce9828_7679, \9393 );
and \U$711 ( \9765 , RIfc583a0_6026, \9395 );
and \U$712 ( \9766 , RIf16cdc0_5698, \9397 );
and \U$713 ( \9767 , RIe224670_4704, \9399 );
and \U$714 ( \9768 , RIf16c118_5689, \9401 );
and \U$715 ( \9769 , RIe221970_4672, \9403 );
and \U$716 ( \9770 , RIfc58508_6027, \9405 );
and \U$717 ( \9771 , RIe21ec70_4640, \9407 );
and \U$718 ( \9772 , RIe219270_4576, \9409 );
and \U$719 ( \9773 , RIe216570_4544, \9411 );
and \U$720 ( \9774 , RIfc3ff08_5753, \9413 );
and \U$721 ( \9775 , RIe213870_4512, \9415 );
and \U$722 ( \9776 , RIf1696e8_5659, \9417 );
and \U$723 ( \9777 , RIe210b70_4480, \9419 );
and \U$724 ( \9778 , RIfc58940_6030, \9421 );
and \U$725 ( \9779 , RIe20de70_4448, \9423 );
and \U$726 ( \9780 , RIe20b170_4416, \9425 );
and \U$727 ( \9781 , RIe208470_4384, \9427 );
and \U$728 ( \9782 , RIfc8fc60_6658, \9429 );
and \U$729 ( \9783 , RIfc97820_6746, \9431 );
and \U$730 ( \9784 , RIe202ea8_4323, \9433 );
and \U$731 ( \9785 , RIe201288_4303, \9435 );
and \U$732 ( \9786 , RIfcc27c8_7235, \9437 );
and \U$733 ( \9787 , RIfcdfee0_7570, \9439 );
and \U$734 ( \9788 , RIfc44198_5797, \9441 );
and \U$735 ( \9789 , RIfc58670_6028, \9443 );
and \U$736 ( \9790 , RIf1608e0_5558, \9445 );
and \U$737 ( \9791 , RIf15e9f0_5536, \9447 );
and \U$738 ( \9792 , RIfe9ff30_8164, \9449 );
and \U$739 ( \9793 , RIe1fc0f8_4245, \9451 );
and \U$740 ( \9794 , RIfc7be90_6432, \9453 );
and \U$741 ( \9795 , RIf15bb88_5503, \9455 );
and \U$742 ( \9796 , RIfcd8cf8_7489, \9457 );
and \U$743 ( \9797 , RIfcd8e60_7490, \9459 );
or \U$744 ( \9798 , \9734 , \9735 , \9736 , \9737 , \9738 , \9739 , \9740 , \9741 , \9742 , \9743 , \9744 , \9745 , \9746 , \9747 , \9748 , \9749 , \9750 , \9751 , \9752 , \9753 , \9754 , \9755 , \9756 , \9757 , \9758 , \9759 , \9760 , \9761 , \9762 , \9763 , \9764 , \9765 , \9766 , \9767 , \9768 , \9769 , \9770 , \9771 , \9772 , \9773 , \9774 , \9775 , \9776 , \9777 , \9778 , \9779 , \9780 , \9781 , \9782 , \9783 , \9784 , \9785 , \9786 , \9787 , \9788 , \9789 , \9790 , \9791 , \9792 , \9793 , \9794 , \9795 , \9796 , \9797 );
and \U$745 ( \9799 , RIfca2d88_6875, \9462 );
and \U$746 ( \9800 , RIfcbdea8_7183, \9464 );
and \U$747 ( \9801 , RIfcb3a20_7066, \9466 );
and \U$748 ( \9802 , RIe1fabe0_4230, \9468 );
and \U$749 ( \9803 , RIfc90098_6661, \9470 );
and \U$750 ( \9804 , RIfc90200_6662, \9472 );
and \U$751 ( \9805 , RIfcd20b0_7412, \9474 );
and \U$752 ( \9806 , RIe1f6158_4177, \9476 );
and \U$753 ( \9807 , RIfc904d0_6664, \9478 );
and \U$754 ( \9808 , RIfca2ef0_6876, \9480 );
and \U$755 ( \9809 , RIfc97550_6744, \9482 );
and \U$756 ( \9810 , RIe1f3e30_4152, \9484 );
and \U$757 ( \9811 , RIfc59048_6035, \9486 );
and \U$758 ( \9812 , RIfc907a0_6666, \9488 );
and \U$759 ( \9813 , RIfc90638_6665, \9490 );
and \U$760 ( \9814 , RIe1eeb38_4093, \9492 );
and \U$761 ( \9815 , RIe1ec3d8_4065, \9494 );
and \U$762 ( \9816 , RIe1e96d8_4033, \9496 );
and \U$763 ( \9817 , RIe1e69d8_4001, \9498 );
and \U$764 ( \9818 , RIe1e3cd8_3969, \9500 );
and \U$765 ( \9819 , RIe1e0fd8_3937, \9502 );
and \U$766 ( \9820 , RIe1de2d8_3905, \9504 );
and \U$767 ( \9821 , RIe1db5d8_3873, \9506 );
and \U$768 ( \9822 , RIe1d88d8_3841, \9508 );
and \U$769 ( \9823 , RIe1d2ed8_3777, \9510 );
and \U$770 ( \9824 , RIe1d01d8_3745, \9512 );
and \U$771 ( \9825 , RIe1cd4d8_3713, \9514 );
and \U$772 ( \9826 , RIe1ca7d8_3681, \9516 );
and \U$773 ( \9827 , RIe1c7ad8_3649, \9518 );
and \U$774 ( \9828 , RIe1c4dd8_3617, \9520 );
and \U$775 ( \9829 , RIe1c20d8_3585, \9522 );
and \U$776 ( \9830 , RIe1bf3d8_3553, \9524 );
and \U$777 ( \9831 , RIfcc73b8_7289, \9526 );
and \U$778 ( \9832 , RIfce3cc0_7614, \9528 );
and \U$779 ( \9833 , RIe1b9e10_3492, \9530 );
and \U$780 ( \9834 , RIe1b7c50_3468, \9532 );
and \U$781 ( \9835 , RIfcd6f70_7468, \9534 );
and \U$782 ( \9836 , RIf149e10_5300, \9536 );
and \U$783 ( \9837 , RIe1b5a90_3444, \9538 );
and \U$784 ( \9838 , RIfea0200_8166, \9540 );
and \U$785 ( \9839 , RIfc90bd8_6669, \9542 );
and \U$786 ( \9840 , RIfcdfd78_7569, \9544 );
and \U$787 ( \9841 , RIe1b2ef8_3413, \9546 );
and \U$788 ( \9842 , RIe1b15a8_3395, \9548 );
and \U$789 ( \9843 , RIfc973e8_6743, \9550 );
and \U$790 ( \9844 , RIfcc7520_7290, \9552 );
and \U$791 ( \9845 , RIe1acdf0_3344, \9554 );
and \U$792 ( \9846 , RIe1ab608_3327, \9556 );
and \U$793 ( \9847 , RIe1a9718_3305, \9558 );
and \U$794 ( \9848 , RIe1a6a18_3273, \9560 );
and \U$795 ( \9849 , RIe1a3d18_3241, \9562 );
and \U$796 ( \9850 , RIe1a1018_3209, \9564 );
and \U$797 ( \9851 , RIe18d518_2985, \9566 );
and \U$798 ( \9852 , RIe179a18_2761, \9568 );
and \U$799 ( \9853 , RIe227370_4736, \9570 );
and \U$800 ( \9854 , RIe21bf70_4608, \9572 );
and \U$801 ( \9855 , RIe205770_4352, \9574 );
and \U$802 ( \9856 , RIe1ff7d0_4284, \9576 );
and \U$803 ( \9857 , RIe1f8b88_4207, \9578 );
and \U$804 ( \9858 , RIe1f16d0_4124, \9580 );
and \U$805 ( \9859 , RIe1d5bd8_3809, \9582 );
and \U$806 ( \9860 , RIe1bc6d8_3521, \9584 );
and \U$807 ( \9861 , RIe1af550_3372, \9586 );
and \U$808 ( \9862 , RIe171b88_2671, \9588 );
or \U$809 ( \9863 , \9799 , \9800 , \9801 , \9802 , \9803 , \9804 , \9805 , \9806 , \9807 , \9808 , \9809 , \9810 , \9811 , \9812 , \9813 , \9814 , \9815 , \9816 , \9817 , \9818 , \9819 , \9820 , \9821 , \9822 , \9823 , \9824 , \9825 , \9826 , \9827 , \9828 , \9829 , \9830 , \9831 , \9832 , \9833 , \9834 , \9835 , \9836 , \9837 , \9838 , \9839 , \9840 , \9841 , \9842 , \9843 , \9844 , \9845 , \9846 , \9847 , \9848 , \9849 , \9850 , \9851 , \9852 , \9853 , \9854 , \9855 , \9856 , \9857 , \9858 , \9859 , \9860 , \9861 , \9862 );
or \U$810 ( \9864 , \9798 , \9863 );
_DC g4273 ( \9865_nG4273 , \9864 , \9597 );
buf \U$811 ( \9866 , \9865_nG4273 );
and \U$812 ( \9867 , \9733 , \9866 );
and \U$813 ( \9868 , RIdec5108_706, \9059 );
and \U$814 ( \9869 , RIdec2408_674, \9061 );
and \U$815 ( \9870 , RIfc93608_6699, \9063 );
and \U$816 ( \9871 , RIdebf708_642, \9065 );
and \U$817 ( \9872 , RIfc934a0_6698, \9067 );
and \U$818 ( \9873 , RIdebca08_610, \9069 );
and \U$819 ( \9874 , RIdeb9d08_578, \9071 );
and \U$820 ( \9875 , RIdeb7008_546, \9073 );
and \U$821 ( \9876 , RIfcdf7d8_7565, \9075 );
and \U$822 ( \9877 , RIdeb1608_482, \9077 );
and \U$823 ( \9878 , RIfc78218_6389, \9079 );
and \U$824 ( \9879 , RIdeae908_450, \9081 );
and \U$825 ( \9880 , RIfcc8498_7301, \9083 );
and \U$826 ( \9881 , RIdea9d90_418, \9085 );
and \U$827 ( \9882 , RIdea3490_386, \9087 );
and \U$828 ( \9883 , RIde9cb90_354, \9089 );
and \U$829 ( \9884 , RIee1cc78_4786, \9091 );
and \U$830 ( \9885 , RIee1bb98_4774, \9093 );
and \U$831 ( \9886 , RIee1b328_4768, \9095 );
and \U$832 ( \9887 , RIee1aab8_4762, \9097 );
and \U$833 ( \9888 , RIde909f8_295, \9099 );
and \U$834 ( \9889 , RIde8d578_279, \9101 );
and \U$835 ( \9890 , RIfea8ea0_8238, \9103 );
and \U$836 ( \9891 , RIde85238_239, \9105 );
and \U$837 ( \9892 , RIde813e0_220, \9107 );
and \U$838 ( \9893 , RIfc938d8_6701, \9109 );
and \U$839 ( \9894 , RIfce5e80_7638, \9111 );
and \U$840 ( \9895 , RIfcbfd98_7205, \9113 );
and \U$841 ( \9896 , RIfce8ce8_7671, \9115 );
and \U$842 ( \9897 , RIe16b4e0_2598, \9117 );
and \U$843 ( \9898 , RIfea8d38_8237, \9119 );
and \U$844 ( \9899 , RIfea9f80_8250, \9121 );
and \U$845 ( \9900 , RIe165108_2527, \9123 );
and \U$846 ( \9901 , RIe162408_2495, \9125 );
and \U$847 ( \9902 , RIfc779a8_6383, \9127 );
and \U$848 ( \9903 , RIe15f708_2463, \9129 );
and \U$849 ( \9904 , RIfe9dc08_8139, \9131 );
and \U$850 ( \9905 , RIe15ca08_2431, \9133 );
and \U$851 ( \9906 , RIe157008_2367, \9135 );
and \U$852 ( \9907 , RIe154308_2335, \9137 );
and \U$853 ( \9908 , RIfea7550_8220, \9139 );
and \U$854 ( \9909 , RIe151608_2303, \9141 );
and \U$855 ( \9910 , RIfcd6160_7458, \9143 );
and \U$856 ( \9911 , RIe14e908_2271, \9145 );
and \U$857 ( \9912 , RIfcd1408_7403, \9147 );
and \U$858 ( \9913 , RIe14bc08_2239, \9149 );
and \U$859 ( \9914 , RIe148f08_2207, \9151 );
and \U$860 ( \9915 , RIe146208_2175, \9153 );
and \U$861 ( \9916 , RIfceb718_7701, \9155 );
and \U$862 ( \9917 , RIfcb19c8_7043, \9157 );
and \U$863 ( \9918 , RIfc93e78_6705, \9159 );
and \U$864 ( \9919 , RIfce7938_7657, \9161 );
and \U$865 ( \9920 , RIe140da8_2115, \9163 );
and \U$866 ( \9921 , RIdf3ecb0_2091, \9165 );
and \U$867 ( \9922 , RIdf3c988_2066, \9167 );
and \U$868 ( \9923 , RIfe9daa0_8138, \9169 );
and \U$869 ( \9924 , RIfce8478_7665, \9171 );
and \U$870 ( \9925 , RIfcdbf98_7525, \9173 );
and \U$871 ( \9926 , RIfc776d8_6381, \9175 );
and \U$872 ( \9927 , RIfc93fe0_6706, \9177 );
and \U$873 ( \9928 , RIdf354d0_1983, \9179 );
and \U$874 ( \9929 , RIdf33040_1957, \9181 );
and \U$875 ( \9930 , RIdf30fe8_1934, \9183 );
and \U$876 ( \9931 , RIdf2ee28_1910, \9185 );
or \U$877 ( \9932 , \9868 , \9869 , \9870 , \9871 , \9872 , \9873 , \9874 , \9875 , \9876 , \9877 , \9878 , \9879 , \9880 , \9881 , \9882 , \9883 , \9884 , \9885 , \9886 , \9887 , \9888 , \9889 , \9890 , \9891 , \9892 , \9893 , \9894 , \9895 , \9896 , \9897 , \9898 , \9899 , \9900 , \9901 , \9902 , \9903 , \9904 , \9905 , \9906 , \9907 , \9908 , \9909 , \9910 , \9911 , \9912 , \9913 , \9914 , \9915 , \9916 , \9917 , \9918 , \9919 , \9920 , \9921 , \9922 , \9923 , \9924 , \9925 , \9926 , \9927 , \9928 , \9929 , \9930 , \9931 );
and \U$878 ( \9933 , RIee2ba20_4955, \9188 );
and \U$879 ( \9934 , RIfc93ba8_6703, \9190 );
and \U$880 ( \9935 , RIfc77de0_6386, \9192 );
and \U$881 ( \9936 , RIee27ad8_4910, \9194 );
and \U$882 ( \9937 , RIfe9d668_8135, \9196 );
and \U$883 ( \9938 , RIfea8bd0_8236, \9198 );
and \U$884 ( \9939 , RIdf26458_1812, \9200 );
and \U$885 ( \9940 , RIfe9d7d0_8136, \9202 );
and \U$886 ( \9941 , RIfcb1c98_7045, \9204 );
and \U$887 ( \9942 , RIee26cc8_4900, \9206 );
and \U$888 ( \9943 , RIdf22ab0_1771, \9208 );
and \U$889 ( \9944 , RIfcc0068_7207, \9210 );
and \U$890 ( \9945 , RIdf21598_1756, \9212 );
and \U$891 ( \9946 , RIdf1f6a8_1734, \9214 );
and \U$892 ( \9947 , RIdf1aef0_1683, \9216 );
and \U$893 ( \9948 , RIfe9d938_8137, \9218 );
and \U$894 ( \9949 , RIdf16cd8_1636, \9220 );
and \U$895 ( \9950 , RIdf13fd8_1604, \9222 );
and \U$896 ( \9951 , RIdf112d8_1572, \9224 );
and \U$897 ( \9952 , RIdf0e5d8_1540, \9226 );
and \U$898 ( \9953 , RIdf0b8d8_1508, \9228 );
and \U$899 ( \9954 , RIdf08bd8_1476, \9230 );
and \U$900 ( \9955 , RIdf05ed8_1444, \9232 );
and \U$901 ( \9956 , RIdf031d8_1412, \9234 );
and \U$902 ( \9957 , RIdefd7d8_1348, \9236 );
and \U$903 ( \9958 , RIdefaad8_1316, \9238 );
and \U$904 ( \9959 , RIdef7dd8_1284, \9240 );
and \U$905 ( \9960 , RIdef50d8_1252, \9242 );
and \U$906 ( \9961 , RIdef23d8_1220, \9244 );
and \U$907 ( \9962 , RIdeef6d8_1188, \9246 );
and \U$908 ( \9963 , RIdeec9d8_1156, \9248 );
and \U$909 ( \9964 , RIdee9cd8_1124, \9250 );
and \U$910 ( \9965 , RIfc942b0_6708, \9252 );
and \U$911 ( \9966 , RIfcde6f8_7553, \9254 );
and \U$912 ( \9967 , RIfcd1138_7401, \9256 );
and \U$913 ( \9968 , RIfcde860_7554, \9258 );
and \U$914 ( \9969 , RIdee4878_1064, \9260 );
and \U$915 ( \9970 , RIdee2af0_1043, \9262 );
and \U$916 ( \9971 , RIdee0a98_1020, \9264 );
and \U$917 ( \9972 , RIdede8d8_996, \9266 );
and \U$918 ( \9973 , RIfc5c9f0_6076, \9268 );
and \U$919 ( \9974 , RIee22240_4847, \9270 );
and \U$920 ( \9975 , RIfcc8768_7303, \9272 );
and \U$921 ( \9976 , RIee21160_4835, \9274 );
and \U$922 ( \9977 , RIded95e0_937, \9276 );
and \U$923 ( \9978 , RIded7150_911, \9278 );
and \U$924 ( \9979 , RIded5260_889, \9280 );
and \U$925 ( \9980 , RIfea76b8_8221, \9282 );
and \U$926 ( \9981 , RIded0508_834, \9284 );
and \U$927 ( \9982 , RIdecd808_802, \9286 );
and \U$928 ( \9983 , RIdecab08_770, \9288 );
and \U$929 ( \9984 , RIdec7e08_738, \9290 );
and \U$930 ( \9985 , RIdeb4308_514, \9292 );
and \U$931 ( \9986 , RIde96290_322, \9294 );
and \U$932 ( \9987 , RIe16df10_2628, \9296 );
and \U$933 ( \9988 , RIe159d08_2399, \9298 );
and \U$934 ( \9989 , RIe143508_2143, \9300 );
and \U$935 ( \9990 , RIdf37f00_2013, \9302 );
and \U$936 ( \9991 , RIdf2c560_1881, \9304 );
and \U$937 ( \9992 , RIdf1cde0_1705, \9306 );
and \U$938 ( \9993 , RIdf004d8_1380, \9308 );
and \U$939 ( \9994 , RIdee6fd8_1092, \9310 );
and \U$940 ( \9995 , RIdedbd40_965, \9312 );
and \U$941 ( \9996 , RIde7c1d8_195, \9314 );
or \U$942 ( \9997 , \9933 , \9934 , \9935 , \9936 , \9937 , \9938 , \9939 , \9940 , \9941 , \9942 , \9943 , \9944 , \9945 , \9946 , \9947 , \9948 , \9949 , \9950 , \9951 , \9952 , \9953 , \9954 , \9955 , \9956 , \9957 , \9958 , \9959 , \9960 , \9961 , \9962 , \9963 , \9964 , \9965 , \9966 , \9967 , \9968 , \9969 , \9970 , \9971 , \9972 , \9973 , \9974 , \9975 , \9976 , \9977 , \9978 , \9979 , \9980 , \9981 , \9982 , \9983 , \9984 , \9985 , \9986 , \9987 , \9988 , \9989 , \9990 , \9991 , \9992 , \9993 , \9994 , \9995 , \9996 );
or \U$943 ( \9998 , \9932 , \9997 );
_DC g31cb ( \9999_nG31cb , \9998 , \9323 );
buf \U$944 ( \10000 , \9999_nG31cb );
and \U$945 ( \10001 , RIe19d3a0_3166, \9333 );
and \U$946 ( \10002 , RIe19a6a0_3134, \9335 );
and \U$947 ( \10003 , RIfcb2c10_7056, \9337 );
and \U$948 ( \10004 , RIe1979a0_3102, \9339 );
and \U$949 ( \10005 , RIfc923c0_6686, \9341 );
and \U$950 ( \10006 , RIe194ca0_3070, \9343 );
and \U$951 ( \10007 , RIe191fa0_3038, \9345 );
and \U$952 ( \10008 , RIe18f2a0_3006, \9347 );
and \U$953 ( \10009 , RIe1898a0_2942, \9349 );
and \U$954 ( \10010 , RIe186ba0_2910, \9351 );
and \U$955 ( \10011 , RIfc422a8_5775, \9353 );
and \U$956 ( \10012 , RIe183ea0_2878, \9355 );
and \U$957 ( \10013 , RIfcbecb8_7193, \9357 );
and \U$958 ( \10014 , RIe1811a0_2846, \9359 );
and \U$959 ( \10015 , RIe17e4a0_2814, \9361 );
and \U$960 ( \10016 , RIe17b7a0_2782, \9363 );
and \U$961 ( \10017 , RIf142250_5212, \9365 );
and \U$962 ( \10018 , RIf140bd0_5196, \9367 );
and \U$963 ( \10019 , RIfec43f8_8353, \9369 );
and \U$964 ( \10020 , RIe175968_2715, \9371 );
and \U$965 ( \10021 , RIfc79b68_6407, \9373 );
and \U$966 ( \10022 , RIf13efb0_5176, \9375 );
and \U$967 ( \10023 , RIfc92528_6687, \9377 );
and \U$968 ( \10024 , RIfcb2aa8_7055, \9379 );
and \U$969 ( \10025 , RIfcd8320_7482, \9381 );
and \U$970 ( \10026 , RIfcea200_7686, \9383 );
and \U$971 ( \10027 , RIfc79898_6405, \9385 );
and \U$972 ( \10028 , RIe1734d8_2689, \9387 );
and \U$973 ( \10029 , RIfcd7948_7475, \9389 );
and \U$974 ( \10030 , RIfcd7678_7473, \9391 );
and \U$975 ( \10031 , RIf16e170_5712, \9393 );
and \U$976 ( \10032 , RIfc927f8_6689, \9395 );
and \U$977 ( \10033 , RIfc92960_6690, \9397 );
and \U$978 ( \10034 , RIe2236f8_4693, \9399 );
and \U$979 ( \10035 , RIfc795c8_6403, \9401 );
and \U$980 ( \10036 , RIe2209f8_4661, \9403 );
and \U$981 ( \10037 , RIf16ad68_5675, \9405 );
and \U$982 ( \10038 , RIe21dcf8_4629, \9407 );
and \U$983 ( \10039 , RIe2182f8_4565, \9409 );
and \U$984 ( \10040 , RIe2155f8_4533, \9411 );
and \U$985 ( \10041 , RIfe9d398_8133, \9413 );
and \U$986 ( \10042 , RIe2128f8_4501, \9415 );
and \U$987 ( \10043 , RIfcdb9f8_7521, \9417 );
and \U$988 ( \10044 , RIe20fbf8_4469, \9419 );
and \U$989 ( \10045 , RIfc41d08_5771, \9421 );
and \U$990 ( \10046 , RIe20cef8_4437, \9423 );
and \U$991 ( \10047 , RIe20a1f8_4405, \9425 );
and \U$992 ( \10048 , RIe2074f8_4373, \9427 );
and \U$993 ( \10049 , RIfcd7510_7472, \9429 );
and \U$994 ( \10050 , RIf166010_5620, \9431 );
and \U$995 ( \10051 , RIfe9d230_8132, \9433 );
and \U$996 ( \10052 , RIe2008b0_4296, \9435 );
and \U$997 ( \10053 , RIf165098_5609, \9437 );
and \U$998 ( \10054 , RIfc41ba0_5770, \9439 );
and \U$999 ( \10055 , RIfc41a38_5769, \9441 );
and \U$1000 ( \10056 , RIfc92c30_6692, \9443 );
and \U$1001 ( \10057 , RIfc418d0_5768, \9445 );
and \U$1002 ( \10058 , RIfc79190_6400, \9447 );
and \U$1003 ( \10059 , RIe1fcad0_4252, \9449 );
and \U$1004 ( \10060 , RIfec4560_8354, \9451 );
and \U$1005 ( \10061 , RIfc79028_6399, \9453 );
and \U$1006 ( \10062 , RIfcbf258_7197, \9455 );
and \U$1007 ( \10063 , RIfcc1df0_7228, \9457 );
and \U$1008 ( \10064 , RIfcd81b8_7481, \9459 );
or \U$1009 ( \10065 , \10001 , \10002 , \10003 , \10004 , \10005 , \10006 , \10007 , \10008 , \10009 , \10010 , \10011 , \10012 , \10013 , \10014 , \10015 , \10016 , \10017 , \10018 , \10019 , \10020 , \10021 , \10022 , \10023 , \10024 , \10025 , \10026 , \10027 , \10028 , \10029 , \10030 , \10031 , \10032 , \10033 , \10034 , \10035 , \10036 , \10037 , \10038 , \10039 , \10040 , \10041 , \10042 , \10043 , \10044 , \10045 , \10046 , \10047 , \10048 , \10049 , \10050 , \10051 , \10052 , \10053 , \10054 , \10055 , \10056 , \10057 , \10058 , \10059 , \10060 , \10061 , \10062 , \10063 , \10064 );
and \U$1010 ( \10066 , RIfc92d98_6693, \9462 );
and \U$1011 ( \10067 , RIfc5b4d8_6061, \9464 );
and \U$1012 ( \10068 , RIfcd77e0_7474, \9466 );
and \U$1013 ( \10069 , RIe1fa0a0_4222, \9468 );
and \U$1014 ( \10070 , RIf156188_5439, \9470 );
and \U$1015 ( \10071 , RIfe9d500_8134, \9472 );
and \U$1016 ( \10072 , RIf1546d0_5420, \9474 );
and \U$1017 ( \10073 , RIe1f5348_4167, \9476 );
and \U$1018 ( \10074 , RIfec4830_8356, \9478 );
and \U$1019 ( \10075 , RIfec46c8_8355, \9480 );
and \U$1020 ( \10076 , RIf1508f0_5376, \9482 );
and \U$1021 ( \10077 , RIe1f3020_4142, \9484 );
and \U$1022 ( \10078 , RIfce3180_7606, \9486 );
and \U$1023 ( \10079 , RIfce8fb8_7673, \9488 );
and \U$1024 ( \10080 , RIfcbf690_7200, \9490 );
and \U$1025 ( \10081 , RIe1edd28_4083, \9492 );
and \U$1026 ( \10082 , RIe1eb460_4054, \9494 );
and \U$1027 ( \10083 , RIe1e8760_4022, \9496 );
and \U$1028 ( \10084 , RIe1e5a60_3990, \9498 );
and \U$1029 ( \10085 , RIe1e2d60_3958, \9500 );
and \U$1030 ( \10086 , RIe1e0060_3926, \9502 );
and \U$1031 ( \10087 , RIe1dd360_3894, \9504 );
and \U$1032 ( \10088 , RIe1da660_3862, \9506 );
and \U$1033 ( \10089 , RIe1d7960_3830, \9508 );
and \U$1034 ( \10090 , RIe1d1f60_3766, \9510 );
and \U$1035 ( \10091 , RIe1cf260_3734, \9512 );
and \U$1036 ( \10092 , RIe1cc560_3702, \9514 );
and \U$1037 ( \10093 , RIe1c9860_3670, \9516 );
and \U$1038 ( \10094 , RIe1c6b60_3638, \9518 );
and \U$1039 ( \10095 , RIe1c3e60_3606, \9520 );
and \U$1040 ( \10096 , RIe1c1160_3574, \9522 );
and \U$1041 ( \10097 , RIe1be460_3542, \9524 );
and \U$1042 ( \10098 , RIfe9d0c8_8131, \9526 );
and \U$1043 ( \10099 , RIfe9cc90_8128, \9528 );
and \U$1044 ( \10100 , RIe1b9168_3483, \9530 );
and \U$1045 ( \10101 , RIe1b7110_3460, \9532 );
and \U$1046 ( \10102 , RIf14a3b0_5304, \9534 );
and \U$1047 ( \10103 , RIfe9cb28_8127, \9536 );
and \U$1048 ( \10104 , RIfe9cf60_8130, \9538 );
and \U$1049 ( \10105 , RIfe9c9c0_8126, \9540 );
and \U$1050 ( \10106 , RIfce2208_7595, \9542 );
and \U$1051 ( \10107 , RIfce9558_7677, \9544 );
and \U$1052 ( \10108 , RIfe9c858_8125, \9546 );
and \U$1053 ( \10109 , RIfe9cdf8_8129, \9548 );
and \U$1054 ( \10110 , RIf147110_5268, \9550 );
and \U$1055 ( \10111 , RIf146468_5259, \9552 );
and \U$1056 ( \10112 , RIe1ac2b0_3336, \9554 );
and \U$1057 ( \10113 , RIe1aaac8_3319, \9556 );
and \U$1058 ( \10114 , RIe1a87a0_3294, \9558 );
and \U$1059 ( \10115 , RIe1a5aa0_3262, \9560 );
and \U$1060 ( \10116 , RIe1a2da0_3230, \9562 );
and \U$1061 ( \10117 , RIe1a00a0_3198, \9564 );
and \U$1062 ( \10118 , RIe18c5a0_2974, \9566 );
and \U$1063 ( \10119 , RIe178aa0_2750, \9568 );
and \U$1064 ( \10120 , RIe2263f8_4725, \9570 );
and \U$1065 ( \10121 , RIe21aff8_4597, \9572 );
and \U$1066 ( \10122 , RIe2047f8_4341, \9574 );
and \U$1067 ( \10123 , RIe1fe858_4273, \9576 );
and \U$1068 ( \10124 , RIe1f7c10_4196, \9578 );
and \U$1069 ( \10125 , RIe1f0758_4113, \9580 );
and \U$1070 ( \10126 , RIe1d4c60_3798, \9582 );
and \U$1071 ( \10127 , RIe1bb760_3510, \9584 );
and \U$1072 ( \10128 , RIe1ae5d8_3361, \9586 );
and \U$1073 ( \10129 , RIe170c10_2660, \9588 );
or \U$1074 ( \10130 , \10066 , \10067 , \10068 , \10069 , \10070 , \10071 , \10072 , \10073 , \10074 , \10075 , \10076 , \10077 , \10078 , \10079 , \10080 , \10081 , \10082 , \10083 , \10084 , \10085 , \10086 , \10087 , \10088 , \10089 , \10090 , \10091 , \10092 , \10093 , \10094 , \10095 , \10096 , \10097 , \10098 , \10099 , \10100 , \10101 , \10102 , \10103 , \10104 , \10105 , \10106 , \10107 , \10108 , \10109 , \10110 , \10111 , \10112 , \10113 , \10114 , \10115 , \10116 , \10117 , \10118 , \10119 , \10120 , \10121 , \10122 , \10123 , \10124 , \10125 , \10126 , \10127 , \10128 , \10129 );
or \U$1075 ( \10131 , \10065 , \10130 );
_DC g42f8 ( \10132_nG42f8 , \10131 , \9597 );
buf \U$1076 ( \10133 , \10132_nG42f8 );
and \U$1077 ( \10134 , \10000 , \10133 );
and \U$1078 ( \10135 , RIdec4190_695, \9059 );
and \U$1079 ( \10136 , RIdec1490_663, \9061 );
and \U$1080 ( \10137 , RIfceaa70_7692, \9063 );
and \U$1081 ( \10138 , RIdebe790_631, \9065 );
and \U$1082 ( \10139 , RIfc954f8_6721, \9067 );
and \U$1083 ( \10140 , RIdebba90_599, \9069 );
and \U$1084 ( \10141 , RIdeb8d90_567, \9071 );
and \U$1085 ( \10142 , RIdeb6090_535, \9073 );
and \U$1086 ( \10143 , RIfcebb50_7704, \9075 );
and \U$1087 ( \10144 , RIdeb0690_471, \9077 );
and \U$1088 ( \10145 , RIee1e190_4801, \9079 );
and \U$1089 ( \10146 , RIdead990_439, \9081 );
and \U$1090 ( \10147 , RIfcdf0d0_7560, \9083 );
and \U$1091 ( \10148 , RIdea7978_407, \9085 );
and \U$1092 ( \10149 , RIdea1078_375, \9087 );
and \U$1093 ( \10150 , RIde9a778_343, \9089 );
and \U$1094 ( \10151 , RIee1c840_4783, \9091 );
and \U$1095 ( \10152 , RIfc957c8_6723, \9093 );
and \U$1096 ( \10153 , RIfcc8e70_7308, \9095 );
and \U$1097 ( \10154 , RIfc5e610_6096, \9097 );
and \U$1098 ( \10155 , RIfe9e8b0_8148, \9099 );
and \U$1099 ( \10156 , RIde8c1c8_273, \9101 );
and \U$1100 ( \10157 , RIde88028_253, \9103 );
and \U$1101 ( \10158 , RIde83b40_232, \9105 );
and \U$1102 ( \10159 , RIfcb0bb8_7033, \9107 );
and \U$1103 ( \10160 , RIfca4b10_6896, \9109 );
and \U$1104 ( \10161 , RIfc75d88_6363, \9111 );
and \U$1105 ( \10162 , RIfca4c78_6897, \9113 );
and \U$1106 ( \10163 , RIfc95390_6720, \9115 );
and \U$1107 ( \10164 , RIe16a9a0_2590, \9117 );
and \U$1108 ( \10165 , RIfcc8fd8_7309, \9119 );
and \U$1109 ( \10166 , RIe166e90_2548, \9121 );
and \U$1110 ( \10167 , RIe164190_2516, \9123 );
and \U$1111 ( \10168 , RIe161490_2484, \9125 );
and \U$1112 ( \10169 , RIfe9e748_8147, \9127 );
and \U$1113 ( \10170 , RIe15e790_2452, \9129 );
and \U$1114 ( \10171 , RIfc74f78_6353, \9131 );
and \U$1115 ( \10172 , RIe15ba90_2420, \9133 );
and \U$1116 ( \10173 , RIe156090_2356, \9135 );
and \U$1117 ( \10174 , RIe153390_2324, \9137 );
and \U$1118 ( \10175 , RIfc3ecc0_5740, \9139 );
and \U$1119 ( \10176 , RIe150690_2292, \9141 );
and \U$1120 ( \10177 , RIfce8b80_7670, \9143 );
and \U$1121 ( \10178 , RIe14d990_2260, \9145 );
and \U$1122 ( \10179 , RIfca6730_6916, \9147 );
and \U$1123 ( \10180 , RIe14ac90_2228, \9149 );
and \U$1124 ( \10181 , RIe147f90_2196, \9151 );
and \U$1125 ( \10182 , RIe145290_2164, \9153 );
and \U$1126 ( \10183 , RIfcee2b0_7732, \9155 );
and \U$1127 ( \10184 , RIfc5f2b8_6105, \9157 );
and \U$1128 ( \10185 , RIfc753b0_6356, \9159 );
and \U$1129 ( \10186 , RIfc74b40_6350, \9161 );
and \U$1130 ( \10187 , RIe140268_2107, \9163 );
and \U$1131 ( \10188 , RIdf3e170_2083, \9165 );
and \U$1132 ( \10189 , RIdf3be48_2058, \9167 );
and \U$1133 ( \10190 , RIdf39c88_2034, \9169 );
and \U$1134 ( \10191 , RIfcc1c88_7227, \9171 );
and \U$1135 ( \10192 , RIfcc1850_7224, \9173 );
and \U$1136 ( \10193 , RIfc965d8_6733, \9175 );
and \U$1137 ( \10194 , RIfc96038_6729, \9177 );
and \U$1138 ( \10195 , RIdf34828_1974, \9179 );
and \U$1139 ( \10196 , RIdf327d0_1951, \9181 );
and \U$1140 ( \10197 , RIdf301d8_1924, \9183 );
and \U$1141 ( \10198 , RIdf2e2e8_1902, \9185 );
or \U$1142 ( \10199 , \10135 , \10136 , \10137 , \10138 , \10139 , \10140 , \10141 , \10142 , \10143 , \10144 , \10145 , \10146 , \10147 , \10148 , \10149 , \10150 , \10151 , \10152 , \10153 , \10154 , \10155 , \10156 , \10157 , \10158 , \10159 , \10160 , \10161 , \10162 , \10163 , \10164 , \10165 , \10166 , \10167 , \10168 , \10169 , \10170 , \10171 , \10172 , \10173 , \10174 , \10175 , \10176 , \10177 , \10178 , \10179 , \10180 , \10181 , \10182 , \10183 , \10184 , \10185 , \10186 , \10187 , \10188 , \10189 , \10190 , \10191 , \10192 , \10193 , \10194 , \10195 , \10196 , \10197 , \10198 );
and \U$1143 ( \10200 , RIfc5e778_6097, \9188 );
and \U$1144 ( \10201 , RIfcd0328_7391, \9190 );
and \U$1145 ( \10202 , RIfc757e8_6359, \9192 );
and \U$1146 ( \10203 , RIfcee6e8_7735, \9194 );
and \U$1147 ( \10204 , RIdf296f8_1848, \9196 );
and \U$1148 ( \10205 , RIdf273d0_1823, \9198 );
and \U$1149 ( \10206 , RIdf257b0_1803, \9200 );
and \U$1150 ( \10207 , RIdf23b90_1783, \9202 );
and \U$1151 ( \10208 , RIfc95d68_6727, \9204 );
and \U$1152 ( \10209 , RIfceda40_7726, \9206 );
and \U$1153 ( \10210 , RIfe9eb80_8150, \9208 );
and \U$1154 ( \10211 , RIfc75518_6357, \9210 );
and \U$1155 ( \10212 , RIfcd01c0_7390, \9212 );
and \U$1156 ( \10213 , RIdf1eb68_1726, \9214 );
and \U$1157 ( \10214 , RIfe9ece8_8151, \9216 );
and \U$1158 ( \10215 , RIfe9ea18_8149, \9218 );
and \U$1159 ( \10216 , RIdf15d60_1625, \9220 );
and \U$1160 ( \10217 , RIdf13060_1593, \9222 );
and \U$1161 ( \10218 , RIdf10360_1561, \9224 );
and \U$1162 ( \10219 , RIdf0d660_1529, \9226 );
and \U$1163 ( \10220 , RIdf0a960_1497, \9228 );
and \U$1164 ( \10221 , RIdf07c60_1465, \9230 );
and \U$1165 ( \10222 , RIdf04f60_1433, \9232 );
and \U$1166 ( \10223 , RIdf02260_1401, \9234 );
and \U$1167 ( \10224 , RIdefc860_1337, \9236 );
and \U$1168 ( \10225 , RIdef9b60_1305, \9238 );
and \U$1169 ( \10226 , RIdef6e60_1273, \9240 );
and \U$1170 ( \10227 , RIdef4160_1241, \9242 );
and \U$1171 ( \10228 , RIdef1460_1209, \9244 );
and \U$1172 ( \10229 , RIdeee760_1177, \9246 );
and \U$1173 ( \10230 , RIdeeba60_1145, \9248 );
and \U$1174 ( \10231 , RIdee8d60_1113, \9250 );
and \U$1175 ( \10232 , RIfc961a0_6730, \9252 );
and \U$1176 ( \10233 , RIfc96308_6731, \9254 );
and \U$1177 ( \10234 , RIfc5ee80_6102, \9256 );
and \U$1178 ( \10235 , RIfce6150_7640, \9258 );
and \U$1179 ( \10236 , RIdee42d8_1060, \9260 );
and \U$1180 ( \10237 , RIdee1e48_1034, \9262 );
and \U$1181 ( \10238 , RIdee00c0_1013, \9264 );
and \U$1182 ( \10239 , RIdeddac8_986, \9266 );
and \U$1183 ( \10240 , RIfc96470_6732, \9268 );
and \U$1184 ( \10241 , RIfc75248_6355, \9270 );
and \U$1185 ( \10242 , RIfc74ca8_6351, \9272 );
and \U$1186 ( \10243 , RIfcb0618_7029, \9274 );
and \U$1187 ( \10244 , RIded8938_928, \9276 );
and \U$1188 ( \10245 , RIded6610_903, \9278 );
and \U$1189 ( \10246 , RIded4450_879, \9280 );
and \U$1190 ( \10247 , RIded2290_855, \9282 );
and \U$1191 ( \10248 , RIdecf590_823, \9284 );
and \U$1192 ( \10249 , RIdecc890_791, \9286 );
and \U$1193 ( \10250 , RIdec9b90_759, \9288 );
and \U$1194 ( \10251 , RIdec6e90_727, \9290 );
and \U$1195 ( \10252 , RIdeb3390_503, \9292 );
and \U$1196 ( \10253 , RIde93e78_311, \9294 );
and \U$1197 ( \10254 , RIe16cf98_2617, \9296 );
and \U$1198 ( \10255 , RIe158d90_2388, \9298 );
and \U$1199 ( \10256 , RIe142590_2132, \9300 );
and \U$1200 ( \10257 , RIdf36f88_2002, \9302 );
and \U$1201 ( \10258 , RIdf2b5e8_1870, \9304 );
and \U$1202 ( \10259 , RIdf1be68_1694, \9306 );
and \U$1203 ( \10260 , RIdeff560_1369, \9308 );
and \U$1204 ( \10261 , RIdee6060_1081, \9310 );
and \U$1205 ( \10262 , RIdedadc8_954, \9312 );
and \U$1206 ( \10263 , RIde79dc0_184, \9314 );
or \U$1207 ( \10264 , \10200 , \10201 , \10202 , \10203 , \10204 , \10205 , \10206 , \10207 , \10208 , \10209 , \10210 , \10211 , \10212 , \10213 , \10214 , \10215 , \10216 , \10217 , \10218 , \10219 , \10220 , \10221 , \10222 , \10223 , \10224 , \10225 , \10226 , \10227 , \10228 , \10229 , \10230 , \10231 , \10232 , \10233 , \10234 , \10235 , \10236 , \10237 , \10238 , \10239 , \10240 , \10241 , \10242 , \10243 , \10244 , \10245 , \10246 , \10247 , \10248 , \10249 , \10250 , \10251 , \10252 , \10253 , \10254 , \10255 , \10256 , \10257 , \10258 , \10259 , \10260 , \10261 , \10262 , \10263 );
or \U$1208 ( \10265 , \10199 , \10264 );
_DC g3250 ( \10266_nG3250 , \10265 , \9323 );
buf \U$1209 ( \10267 , \10266_nG3250 );
and \U$1210 ( \10268 , RIe19c428_3155, \9333 );
and \U$1211 ( \10269 , RIe199728_3123, \9335 );
and \U$1212 ( \10270 , RIfe9e310_8144, \9337 );
and \U$1213 ( \10271 , RIe196a28_3091, \9339 );
and \U$1214 ( \10272 , RIfcc04a0_7210, \9341 );
and \U$1215 ( \10273 , RIe193d28_3059, \9343 );
and \U$1216 ( \10274 , RIe191028_3027, \9345 );
and \U$1217 ( \10275 , RIe18e328_2995, \9347 );
and \U$1218 ( \10276 , RIe188928_2931, \9349 );
and \U$1219 ( \10277 , RIe185c28_2899, \9351 );
and \U$1220 ( \10278 , RIfce1830_7588, \9353 );
and \U$1221 ( \10279 , RIe182f28_2867, \9355 );
and \U$1222 ( \10280 , RIfe9e478_8145, \9357 );
and \U$1223 ( \10281 , RIe180228_2835, \9359 );
and \U$1224 ( \10282 , RIe17d528_2803, \9361 );
and \U$1225 ( \10283 , RIe17a828_2771, \9363 );
and \U$1226 ( \10284 , RIf141878_5205, \9365 );
and \U$1227 ( \10285 , RIfcb12c0_7038, \9367 );
and \U$1228 ( \10286 , RIfc94418_6709, \9369 );
and \U$1229 ( \10287 , RIe174f90_2708, \9371 );
and \U$1230 ( \10288 , RIfc77408_6379, \9373 );
and \U$1231 ( \10289 , RIf13ea10_5172, \9375 );
and \U$1232 ( \10290 , RIfcdc100_7526, \9377 );
and \U$1233 ( \10291 , RIfc94580_6710, \9379 );
and \U$1234 ( \10292 , RIfc946e8_6711, \9381 );
and \U$1235 ( \10293 , RIfced338_7721, \9383 );
and \U$1236 ( \10294 , RIfce5fe8_7639, \9385 );
and \U$1237 ( \10295 , RIe172998_2681, \9387 );
and \U$1238 ( \10296 , RIfcdc268_7527, \9389 );
and \U$1239 ( \10297 , RIfcddff0_7548, \9391 );
and \U$1240 ( \10298 , RIfcc0608_7211, \9393 );
and \U$1241 ( \10299 , RIfce7230_7652, \9395 );
and \U$1242 ( \10300 , RIfc40340_5756, \9397 );
and \U$1243 ( \10301 , RIe222780_4682, \9399 );
and \U$1244 ( \10302 , RIfcdd618_7541, \9401 );
and \U$1245 ( \10303 , RIe21fa80_4650, \9403 );
and \U$1246 ( \10304 , RIfcd0b98_7397, \9405 );
and \U$1247 ( \10305 , RIe21cd80_4618, \9407 );
and \U$1248 ( \10306 , RIe217380_4554, \9409 );
and \U$1249 ( \10307 , RIe214680_4522, \9411 );
and \U$1250 ( \10308 , RIfec4998_8357, \9413 );
and \U$1251 ( \10309 , RIe211980_4490, \9415 );
and \U$1252 ( \10310 , RIf168608_5647, \9417 );
and \U$1253 ( \10311 , RIe20ec80_4458, \9419 );
and \U$1254 ( \10312 , RIfcc0770_7212, \9421 );
and \U$1255 ( \10313 , RIe20bf80_4426, \9423 );
and \U$1256 ( \10314 , RIe209280_4394, \9425 );
and \U$1257 ( \10315 , RIe206580_4362, \9427 );
and \U$1258 ( \10316 , RIfce2370_7596, \9429 );
and \U$1259 ( \10317 , RIfcee580_7734, \9431 );
and \U$1260 ( \10318 , RIfec4c68_8359, \9433 );
and \U$1261 ( \10319 , RIfec4b00_8358, \9435 );
and \U$1262 ( \10320 , RIfc949b8_6713, \9437 );
and \U$1263 ( \10321 , RIfcebcb8_7705, \9439 );
and \U$1264 ( \10322 , RIf162938_5581, \9441 );
and \U$1265 ( \10323 , RIf1612b8_5565, \9443 );
and \U$1266 ( \10324 , RIfccd088_7355, \9445 );
and \U$1267 ( \10325 , RIfcc08d8_7213, \9447 );
and \U$1268 ( \10326 , RIfe9e040_8142, \9449 );
and \U$1269 ( \10327 , RIfe9e1a8_8143, \9451 );
and \U$1270 ( \10328 , RIfcead40_7694, \9453 );
and \U$1271 ( \10329 , RIf15ad78_5493, \9455 );
and \U$1272 ( \10330 , RIfc94c88_6715, \9457 );
and \U$1273 ( \10331 , RIfccc3e0_7346, \9459 );
or \U$1274 ( \10332 , \10268 , \10269 , \10270 , \10271 , \10272 , \10273 , \10274 , \10275 , \10276 , \10277 , \10278 , \10279 , \10280 , \10281 , \10282 , \10283 , \10284 , \10285 , \10286 , \10287 , \10288 , \10289 , \10290 , \10291 , \10292 , \10293 , \10294 , \10295 , \10296 , \10297 , \10298 , \10299 , \10300 , \10301 , \10302 , \10303 , \10304 , \10305 , \10306 , \10307 , \10308 , \10309 , \10310 , \10311 , \10312 , \10313 , \10314 , \10315 , \10316 , \10317 , \10318 , \10319 , \10320 , \10321 , \10322 , \10323 , \10324 , \10325 , \10326 , \10327 , \10328 , \10329 , \10330 , \10331 );
and \U$1275 ( \10333 , RIfc765f8_6369, \9462 );
and \U$1276 ( \10334 , RIfc94df0_6716, \9464 );
and \U$1277 ( \10335 , RIfcc0a40_7214, \9466 );
and \U$1278 ( \10336 , RIe1f9998_4217, \9468 );
and \U$1279 ( \10337 , RIfcc8d08_7307, \9470 );
and \U$1280 ( \10338 , RIfce8748_7667, \9472 );
and \U$1281 ( \10339 , RIfceb2e0_7698, \9474 );
and \U$1282 ( \10340 , RIe1f4970_4160, \9476 );
and \U$1283 ( \10341 , RIf152510_5396, \9478 );
and \U$1284 ( \10342 , RIf1512c8_5383, \9480 );
and \U$1285 ( \10343 , RIfcb0ff0_7036, \9482 );
and \U$1286 ( \10344 , RIe1f24e0_4134, \9484 );
and \U$1287 ( \10345 , RIfc761c0_6366, \9486 );
and \U$1288 ( \10346 , RIfc950c0_6718, \9488 );
and \U$1289 ( \10347 , RIfcc0e78_7217, \9490 );
and \U$1290 ( \10348 , RIe1ed1e8_4075, \9492 );
and \U$1291 ( \10349 , RIe1ea4e8_4043, \9494 );
and \U$1292 ( \10350 , RIe1e77e8_4011, \9496 );
and \U$1293 ( \10351 , RIe1e4ae8_3979, \9498 );
and \U$1294 ( \10352 , RIe1e1de8_3947, \9500 );
and \U$1295 ( \10353 , RIe1df0e8_3915, \9502 );
and \U$1296 ( \10354 , RIe1dc3e8_3883, \9504 );
and \U$1297 ( \10355 , RIe1d96e8_3851, \9506 );
and \U$1298 ( \10356 , RIe1d69e8_3819, \9508 );
and \U$1299 ( \10357 , RIe1d0fe8_3755, \9510 );
and \U$1300 ( \10358 , RIe1ce2e8_3723, \9512 );
and \U$1301 ( \10359 , RIe1cb5e8_3691, \9514 );
and \U$1302 ( \10360 , RIe1c88e8_3659, \9516 );
and \U$1303 ( \10361 , RIe1c5be8_3627, \9518 );
and \U$1304 ( \10362 , RIe1c2ee8_3595, \9520 );
and \U$1305 ( \10363 , RIe1c01e8_3563, \9522 );
and \U$1306 ( \10364 , RIe1bd4e8_3531, \9524 );
and \U$1307 ( \10365 , RIf14bfd0_5324, \9526 );
and \U$1308 ( \10366 , RIf14ac20_5310, \9528 );
and \U$1309 ( \10367 , RIfe9ded8_8141, \9530 );
and \U$1310 ( \10368 , RIe1b65d0_3452, \9532 );
and \U$1311 ( \10369 , RIfcecd98_7717, \9534 );
and \U$1312 ( \10370 , RIfc76490_6368, \9536 );
and \U$1313 ( \10371 , RIe1b4c80_3434, \9538 );
and \U$1314 ( \10372 , RIe1b38d0_3420, \9540 );
and \U$1315 ( \10373 , RIfcc0fe0_7218, \9542 );
and \U$1316 ( \10374 , RIfceaea8_7695, \9544 );
and \U$1317 ( \10375 , RIe1b1f80_3402, \9546 );
and \U$1318 ( \10376 , RIe1b0360_3382, \9548 );
and \U$1319 ( \10377 , RIfcd0760_7394, \9550 );
and \U$1320 ( \10378 , RIf145ec8_5255, \9552 );
and \U$1321 ( \10379 , RIfe9e5e0_8146, \9554 );
and \U$1322 ( \10380 , RIfe9dd70_8140, \9556 );
and \U$1323 ( \10381 , RIe1a7828_3283, \9558 );
and \U$1324 ( \10382 , RIe1a4b28_3251, \9560 );
and \U$1325 ( \10383 , RIe1a1e28_3219, \9562 );
and \U$1326 ( \10384 , RIe19f128_3187, \9564 );
and \U$1327 ( \10385 , RIe18b628_2963, \9566 );
and \U$1328 ( \10386 , RIe177b28_2739, \9568 );
and \U$1329 ( \10387 , RIe225480_4714, \9570 );
and \U$1330 ( \10388 , RIe21a080_4586, \9572 );
and \U$1331 ( \10389 , RIe203880_4330, \9574 );
and \U$1332 ( \10390 , RIe1fd8e0_4262, \9576 );
and \U$1333 ( \10391 , RIe1f6c98_4185, \9578 );
and \U$1334 ( \10392 , RIe1ef7e0_4102, \9580 );
and \U$1335 ( \10393 , RIe1d3ce8_3787, \9582 );
and \U$1336 ( \10394 , RIe1ba7e8_3499, \9584 );
and \U$1337 ( \10395 , RIe1ad660_3350, \9586 );
and \U$1338 ( \10396 , RIe16fc98_2649, \9588 );
or \U$1339 ( \10397 , \10333 , \10334 , \10335 , \10336 , \10337 , \10338 , \10339 , \10340 , \10341 , \10342 , \10343 , \10344 , \10345 , \10346 , \10347 , \10348 , \10349 , \10350 , \10351 , \10352 , \10353 , \10354 , \10355 , \10356 , \10357 , \10358 , \10359 , \10360 , \10361 , \10362 , \10363 , \10364 , \10365 , \10366 , \10367 , \10368 , \10369 , \10370 , \10371 , \10372 , \10373 , \10374 , \10375 , \10376 , \10377 , \10378 , \10379 , \10380 , \10381 , \10382 , \10383 , \10384 , \10385 , \10386 , \10387 , \10388 , \10389 , \10390 , \10391 , \10392 , \10393 , \10394 , \10395 , \10396 );
or \U$1340 ( \10398 , \10332 , \10397 );
_DC g437d ( \10399_nG437d , \10398 , \9597 );
buf \U$1341 ( \10400 , \10399_nG437d );
and \U$1342 ( \10401 , \10267 , \10400 );
and \U$1343 ( \10402 , \10133 , \10401 );
and \U$1344 ( \10403 , \10000 , \10401 );
or \U$1345 ( \10404 , \10134 , \10402 , \10403 );
and \U$1346 ( \10405 , \9866 , \10404 );
and \U$1347 ( \10406 , \9733 , \10404 );
or \U$1348 ( \10407 , \9867 , \10405 , \10406 );
xor \U$1349 ( \10408 , \9600 , \10407 );
buf g444e ( \10409_nG444e , \10408 );
xor \U$1350 ( \10410 , \9733 , \9866 );
xor \U$1351 ( \10411 , \10410 , \10404 );
buf g4451 ( \10412_nG4451 , \10411 );
xor \U$1352 ( \10413 , \10000 , \10133 );
xor \U$1353 ( \10414 , \10413 , \10401 );
buf g4454 ( \10415_nG4454 , \10414 );
nand \U$1354 ( \10416 , \10412_nG4451 , \10415_nG4454 );
and \U$1355 ( \10417 , \10409_nG444e , \10416 );
xor \U$1356 ( \10418 , \10412_nG4451 , \10415_nG4454 );
not \U$1357 ( \10419 , \10418 );
xor \U$1358 ( \10420 , \10409_nG444e , \10412_nG4451 );
and \U$1359 ( \10421 , \10419 , \10420 );
and \U$1362 ( \10422 , RIdec4190_695, \9333 );
and \U$1363 ( \10423 , RIdec1490_663, \9335 );
and \U$1364 ( \10424 , RIfceaa70_7692, \9337 );
and \U$1365 ( \10425 , RIdebe790_631, \9339 );
and \U$1366 ( \10426 , RIfc954f8_6721, \9341 );
and \U$1367 ( \10427 , RIdebba90_599, \9343 );
and \U$1368 ( \10428 , RIdeb8d90_567, \9345 );
and \U$1369 ( \10429 , RIdeb6090_535, \9347 );
and \U$1370 ( \10430 , RIfcebb50_7704, \9349 );
and \U$1371 ( \10431 , RIdeb0690_471, \9351 );
and \U$1372 ( \10432 , RIee1e190_4801, \9353 );
and \U$1373 ( \10433 , RIdead990_439, \9355 );
and \U$1374 ( \10434 , RIfcdf0d0_7560, \9357 );
and \U$1375 ( \10435 , RIdea7978_407, \9359 );
and \U$1376 ( \10436 , RIdea1078_375, \9361 );
and \U$1377 ( \10437 , RIde9a778_343, \9363 );
and \U$1378 ( \10438 , RIee1c840_4783, \9365 );
and \U$1379 ( \10439 , RIfc957c8_6723, \9367 );
and \U$1380 ( \10440 , RIfcc8e70_7308, \9369 );
and \U$1381 ( \10441 , RIfc5e610_6096, \9371 );
and \U$1382 ( \10442 , RIfe9e8b0_8148, \9373 );
and \U$1383 ( \10443 , RIde8c1c8_273, \9375 );
and \U$1384 ( \10444 , RIde88028_253, \9377 );
and \U$1385 ( \10445 , RIde83b40_232, \9379 );
and \U$1386 ( \10446 , RIfcb0bb8_7033, \9381 );
and \U$1387 ( \10447 , RIfca4b10_6896, \9383 );
and \U$1388 ( \10448 , RIfc75d88_6363, \9385 );
and \U$1389 ( \10449 , RIfca4c78_6897, \9387 );
and \U$1390 ( \10450 , RIfc95390_6720, \9389 );
and \U$1391 ( \10451 , RIe16a9a0_2590, \9391 );
and \U$1392 ( \10452 , RIfcc8fd8_7309, \9393 );
and \U$1393 ( \10453 , RIe166e90_2548, \9395 );
and \U$1394 ( \10454 , RIe164190_2516, \9397 );
and \U$1395 ( \10455 , RIe161490_2484, \9399 );
and \U$1396 ( \10456 , RIfe9e748_8147, \9401 );
and \U$1397 ( \10457 , RIe15e790_2452, \9403 );
and \U$1398 ( \10458 , RIfc74f78_6353, \9405 );
and \U$1399 ( \10459 , RIe15ba90_2420, \9407 );
and \U$1400 ( \10460 , RIe156090_2356, \9409 );
and \U$1401 ( \10461 , RIe153390_2324, \9411 );
and \U$1402 ( \10462 , RIfc3ecc0_5740, \9413 );
and \U$1403 ( \10463 , RIe150690_2292, \9415 );
and \U$1404 ( \10464 , RIfce8b80_7670, \9417 );
and \U$1405 ( \10465 , RIe14d990_2260, \9419 );
and \U$1406 ( \10466 , RIfca6730_6916, \9421 );
and \U$1407 ( \10467 , RIe14ac90_2228, \9423 );
and \U$1408 ( \10468 , RIe147f90_2196, \9425 );
and \U$1409 ( \10469 , RIe145290_2164, \9427 );
and \U$1410 ( \10470 , RIfcee2b0_7732, \9429 );
and \U$1411 ( \10471 , RIfc5f2b8_6105, \9431 );
and \U$1412 ( \10472 , RIfc753b0_6356, \9433 );
and \U$1413 ( \10473 , RIfc74b40_6350, \9435 );
and \U$1414 ( \10474 , RIe140268_2107, \9437 );
and \U$1415 ( \10475 , RIdf3e170_2083, \9439 );
and \U$1416 ( \10476 , RIdf3be48_2058, \9441 );
and \U$1417 ( \10477 , RIdf39c88_2034, \9443 );
and \U$1418 ( \10478 , RIfcc1c88_7227, \9445 );
and \U$1419 ( \10479 , RIfcc1850_7224, \9447 );
and \U$1420 ( \10480 , RIfc965d8_6733, \9449 );
and \U$1421 ( \10481 , RIfc96038_6729, \9451 );
and \U$1422 ( \10482 , RIdf34828_1974, \9453 );
and \U$1423 ( \10483 , RIdf327d0_1951, \9455 );
and \U$1424 ( \10484 , RIdf301d8_1924, \9457 );
and \U$1425 ( \10485 , RIdf2e2e8_1902, \9459 );
or \U$1426 ( \10486 , \10422 , \10423 , \10424 , \10425 , \10426 , \10427 , \10428 , \10429 , \10430 , \10431 , \10432 , \10433 , \10434 , \10435 , \10436 , \10437 , \10438 , \10439 , \10440 , \10441 , \10442 , \10443 , \10444 , \10445 , \10446 , \10447 , \10448 , \10449 , \10450 , \10451 , \10452 , \10453 , \10454 , \10455 , \10456 , \10457 , \10458 , \10459 , \10460 , \10461 , \10462 , \10463 , \10464 , \10465 , \10466 , \10467 , \10468 , \10469 , \10470 , \10471 , \10472 , \10473 , \10474 , \10475 , \10476 , \10477 , \10478 , \10479 , \10480 , \10481 , \10482 , \10483 , \10484 , \10485 );
and \U$1427 ( \10487 , RIfc5e778_6097, \9462 );
and \U$1428 ( \10488 , RIfcd0328_7391, \9464 );
and \U$1429 ( \10489 , RIfc757e8_6359, \9466 );
and \U$1430 ( \10490 , RIfcee6e8_7735, \9468 );
and \U$1431 ( \10491 , RIdf296f8_1848, \9470 );
and \U$1432 ( \10492 , RIdf273d0_1823, \9472 );
and \U$1433 ( \10493 , RIdf257b0_1803, \9474 );
and \U$1434 ( \10494 , RIdf23b90_1783, \9476 );
and \U$1435 ( \10495 , RIfc95d68_6727, \9478 );
and \U$1436 ( \10496 , RIfceda40_7726, \9480 );
and \U$1437 ( \10497 , RIfe9eb80_8150, \9482 );
and \U$1438 ( \10498 , RIfc75518_6357, \9484 );
and \U$1439 ( \10499 , RIfcd01c0_7390, \9486 );
and \U$1440 ( \10500 , RIdf1eb68_1726, \9488 );
and \U$1441 ( \10501 , RIfe9ece8_8151, \9490 );
and \U$1442 ( \10502 , RIfe9ea18_8149, \9492 );
and \U$1443 ( \10503 , RIdf15d60_1625, \9494 );
and \U$1444 ( \10504 , RIdf13060_1593, \9496 );
and \U$1445 ( \10505 , RIdf10360_1561, \9498 );
and \U$1446 ( \10506 , RIdf0d660_1529, \9500 );
and \U$1447 ( \10507 , RIdf0a960_1497, \9502 );
and \U$1448 ( \10508 , RIdf07c60_1465, \9504 );
and \U$1449 ( \10509 , RIdf04f60_1433, \9506 );
and \U$1450 ( \10510 , RIdf02260_1401, \9508 );
and \U$1451 ( \10511 , RIdefc860_1337, \9510 );
and \U$1452 ( \10512 , RIdef9b60_1305, \9512 );
and \U$1453 ( \10513 , RIdef6e60_1273, \9514 );
and \U$1454 ( \10514 , RIdef4160_1241, \9516 );
and \U$1455 ( \10515 , RIdef1460_1209, \9518 );
and \U$1456 ( \10516 , RIdeee760_1177, \9520 );
and \U$1457 ( \10517 , RIdeeba60_1145, \9522 );
and \U$1458 ( \10518 , RIdee8d60_1113, \9524 );
and \U$1459 ( \10519 , RIfc961a0_6730, \9526 );
and \U$1460 ( \10520 , RIfc96308_6731, \9528 );
and \U$1461 ( \10521 , RIfc5ee80_6102, \9530 );
and \U$1462 ( \10522 , RIfce6150_7640, \9532 );
and \U$1463 ( \10523 , RIdee42d8_1060, \9534 );
and \U$1464 ( \10524 , RIdee1e48_1034, \9536 );
and \U$1465 ( \10525 , RIdee00c0_1013, \9538 );
and \U$1466 ( \10526 , RIdeddac8_986, \9540 );
and \U$1467 ( \10527 , RIfc96470_6732, \9542 );
and \U$1468 ( \10528 , RIfc75248_6355, \9544 );
and \U$1469 ( \10529 , RIfc74ca8_6351, \9546 );
and \U$1470 ( \10530 , RIfcb0618_7029, \9548 );
and \U$1471 ( \10531 , RIded8938_928, \9550 );
and \U$1472 ( \10532 , RIded6610_903, \9552 );
and \U$1473 ( \10533 , RIded4450_879, \9554 );
and \U$1474 ( \10534 , RIded2290_855, \9556 );
and \U$1475 ( \10535 , RIdecf590_823, \9558 );
and \U$1476 ( \10536 , RIdecc890_791, \9560 );
and \U$1477 ( \10537 , RIdec9b90_759, \9562 );
and \U$1478 ( \10538 , RIdec6e90_727, \9564 );
and \U$1479 ( \10539 , RIdeb3390_503, \9566 );
and \U$1480 ( \10540 , RIde93e78_311, \9568 );
and \U$1481 ( \10541 , RIe16cf98_2617, \9570 );
and \U$1482 ( \10542 , RIe158d90_2388, \9572 );
and \U$1483 ( \10543 , RIe142590_2132, \9574 );
and \U$1484 ( \10544 , RIdf36f88_2002, \9576 );
and \U$1485 ( \10545 , RIdf2b5e8_1870, \9578 );
and \U$1486 ( \10546 , RIdf1be68_1694, \9580 );
and \U$1487 ( \10547 , RIdeff560_1369, \9582 );
and \U$1488 ( \10548 , RIdee6060_1081, \9584 );
and \U$1489 ( \10549 , RIdedadc8_954, \9586 );
and \U$1490 ( \10550 , RIde79dc0_184, \9588 );
or \U$1491 ( \10551 , \10487 , \10488 , \10489 , \10490 , \10491 , \10492 , \10493 , \10494 , \10495 , \10496 , \10497 , \10498 , \10499 , \10500 , \10501 , \10502 , \10503 , \10504 , \10505 , \10506 , \10507 , \10508 , \10509 , \10510 , \10511 , \10512 , \10513 , \10514 , \10515 , \10516 , \10517 , \10518 , \10519 , \10520 , \10521 , \10522 , \10523 , \10524 , \10525 , \10526 , \10527 , \10528 , \10529 , \10530 , \10531 , \10532 , \10533 , \10534 , \10535 , \10536 , \10537 , \10538 , \10539 , \10540 , \10541 , \10542 , \10543 , \10544 , \10545 , \10546 , \10547 , \10548 , \10549 , \10550 );
or \U$1492 ( \10552 , \10486 , \10551 );
_DC g6577 ( \10553_nG6577 , \10552 , \9597 );
and \U$1493 ( \10554 , RIe19c428_3155, \9059 );
and \U$1494 ( \10555 , RIe199728_3123, \9061 );
and \U$1495 ( \10556 , RIfe9e310_8144, \9063 );
and \U$1496 ( \10557 , RIe196a28_3091, \9065 );
and \U$1497 ( \10558 , RIfcc04a0_7210, \9067 );
and \U$1498 ( \10559 , RIe193d28_3059, \9069 );
and \U$1499 ( \10560 , RIe191028_3027, \9071 );
and \U$1500 ( \10561 , RIe18e328_2995, \9073 );
and \U$1501 ( \10562 , RIe188928_2931, \9075 );
and \U$1502 ( \10563 , RIe185c28_2899, \9077 );
and \U$1503 ( \10564 , RIfce1830_7588, \9079 );
and \U$1504 ( \10565 , RIe182f28_2867, \9081 );
and \U$1505 ( \10566 , RIfe9e478_8145, \9083 );
and \U$1506 ( \10567 , RIe180228_2835, \9085 );
and \U$1507 ( \10568 , RIe17d528_2803, \9087 );
and \U$1508 ( \10569 , RIe17a828_2771, \9089 );
and \U$1509 ( \10570 , RIf141878_5205, \9091 );
and \U$1510 ( \10571 , RIfcb12c0_7038, \9093 );
and \U$1511 ( \10572 , RIfc94418_6709, \9095 );
and \U$1512 ( \10573 , RIe174f90_2708, \9097 );
and \U$1513 ( \10574 , RIfc77408_6379, \9099 );
and \U$1514 ( \10575 , RIf13ea10_5172, \9101 );
and \U$1515 ( \10576 , RIfcdc100_7526, \9103 );
and \U$1516 ( \10577 , RIfc94580_6710, \9105 );
and \U$1517 ( \10578 , RIfc946e8_6711, \9107 );
and \U$1518 ( \10579 , RIfced338_7721, \9109 );
and \U$1519 ( \10580 , RIfce5fe8_7639, \9111 );
and \U$1520 ( \10581 , RIe172998_2681, \9113 );
and \U$1521 ( \10582 , RIfcdc268_7527, \9115 );
and \U$1522 ( \10583 , RIfcddff0_7548, \9117 );
and \U$1523 ( \10584 , RIfcc0608_7211, \9119 );
and \U$1524 ( \10585 , RIfce7230_7652, \9121 );
and \U$1525 ( \10586 , RIfc40340_5756, \9123 );
and \U$1526 ( \10587 , RIe222780_4682, \9125 );
and \U$1527 ( \10588 , RIfcdd618_7541, \9127 );
and \U$1528 ( \10589 , RIe21fa80_4650, \9129 );
and \U$1529 ( \10590 , RIfcd0b98_7397, \9131 );
and \U$1530 ( \10591 , RIe21cd80_4618, \9133 );
and \U$1531 ( \10592 , RIe217380_4554, \9135 );
and \U$1532 ( \10593 , RIe214680_4522, \9137 );
and \U$1533 ( \10594 , RIfec4998_8357, \9139 );
and \U$1534 ( \10595 , RIe211980_4490, \9141 );
and \U$1535 ( \10596 , RIf168608_5647, \9143 );
and \U$1536 ( \10597 , RIe20ec80_4458, \9145 );
and \U$1537 ( \10598 , RIfcc0770_7212, \9147 );
and \U$1538 ( \10599 , RIe20bf80_4426, \9149 );
and \U$1539 ( \10600 , RIe209280_4394, \9151 );
and \U$1540 ( \10601 , RIe206580_4362, \9153 );
and \U$1541 ( \10602 , RIfce2370_7596, \9155 );
and \U$1542 ( \10603 , RIfcee580_7734, \9157 );
and \U$1543 ( \10604 , RIfec4c68_8359, \9159 );
and \U$1544 ( \10605 , RIfec4b00_8358, \9161 );
and \U$1545 ( \10606 , RIfc949b8_6713, \9163 );
and \U$1546 ( \10607 , RIfcebcb8_7705, \9165 );
and \U$1547 ( \10608 , RIf162938_5581, \9167 );
and \U$1548 ( \10609 , RIf1612b8_5565, \9169 );
and \U$1549 ( \10610 , RIfccd088_7355, \9171 );
and \U$1550 ( \10611 , RIfcc08d8_7213, \9173 );
and \U$1551 ( \10612 , RIfe9e040_8142, \9175 );
and \U$1552 ( \10613 , RIfe9e1a8_8143, \9177 );
and \U$1553 ( \10614 , RIfcead40_7694, \9179 );
and \U$1554 ( \10615 , RIf15ad78_5493, \9181 );
and \U$1555 ( \10616 , RIfc94c88_6715, \9183 );
and \U$1556 ( \10617 , RIfccc3e0_7346, \9185 );
or \U$1557 ( \10618 , \10554 , \10555 , \10556 , \10557 , \10558 , \10559 , \10560 , \10561 , \10562 , \10563 , \10564 , \10565 , \10566 , \10567 , \10568 , \10569 , \10570 , \10571 , \10572 , \10573 , \10574 , \10575 , \10576 , \10577 , \10578 , \10579 , \10580 , \10581 , \10582 , \10583 , \10584 , \10585 , \10586 , \10587 , \10588 , \10589 , \10590 , \10591 , \10592 , \10593 , \10594 , \10595 , \10596 , \10597 , \10598 , \10599 , \10600 , \10601 , \10602 , \10603 , \10604 , \10605 , \10606 , \10607 , \10608 , \10609 , \10610 , \10611 , \10612 , \10613 , \10614 , \10615 , \10616 , \10617 );
and \U$1558 ( \10619 , RIfc765f8_6369, \9188 );
and \U$1559 ( \10620 , RIfc94df0_6716, \9190 );
and \U$1560 ( \10621 , RIfcc0a40_7214, \9192 );
and \U$1561 ( \10622 , RIe1f9998_4217, \9194 );
and \U$1562 ( \10623 , RIfcc8d08_7307, \9196 );
and \U$1563 ( \10624 , RIfce8748_7667, \9198 );
and \U$1564 ( \10625 , RIfceb2e0_7698, \9200 );
and \U$1565 ( \10626 , RIe1f4970_4160, \9202 );
and \U$1566 ( \10627 , RIf152510_5396, \9204 );
and \U$1567 ( \10628 , RIf1512c8_5383, \9206 );
and \U$1568 ( \10629 , RIfcb0ff0_7036, \9208 );
and \U$1569 ( \10630 , RIe1f24e0_4134, \9210 );
and \U$1570 ( \10631 , RIfc761c0_6366, \9212 );
and \U$1571 ( \10632 , RIfc950c0_6718, \9214 );
and \U$1572 ( \10633 , RIfcc0e78_7217, \9216 );
and \U$1573 ( \10634 , RIe1ed1e8_4075, \9218 );
and \U$1574 ( \10635 , RIe1ea4e8_4043, \9220 );
and \U$1575 ( \10636 , RIe1e77e8_4011, \9222 );
and \U$1576 ( \10637 , RIe1e4ae8_3979, \9224 );
and \U$1577 ( \10638 , RIe1e1de8_3947, \9226 );
and \U$1578 ( \10639 , RIe1df0e8_3915, \9228 );
and \U$1579 ( \10640 , RIe1dc3e8_3883, \9230 );
and \U$1580 ( \10641 , RIe1d96e8_3851, \9232 );
and \U$1581 ( \10642 , RIe1d69e8_3819, \9234 );
and \U$1582 ( \10643 , RIe1d0fe8_3755, \9236 );
and \U$1583 ( \10644 , RIe1ce2e8_3723, \9238 );
and \U$1584 ( \10645 , RIe1cb5e8_3691, \9240 );
and \U$1585 ( \10646 , RIe1c88e8_3659, \9242 );
and \U$1586 ( \10647 , RIe1c5be8_3627, \9244 );
and \U$1587 ( \10648 , RIe1c2ee8_3595, \9246 );
and \U$1588 ( \10649 , RIe1c01e8_3563, \9248 );
and \U$1589 ( \10650 , RIe1bd4e8_3531, \9250 );
and \U$1590 ( \10651 , RIf14bfd0_5324, \9252 );
and \U$1591 ( \10652 , RIf14ac20_5310, \9254 );
and \U$1592 ( \10653 , RIfe9ded8_8141, \9256 );
and \U$1593 ( \10654 , RIe1b65d0_3452, \9258 );
and \U$1594 ( \10655 , RIfcecd98_7717, \9260 );
and \U$1595 ( \10656 , RIfc76490_6368, \9262 );
and \U$1596 ( \10657 , RIe1b4c80_3434, \9264 );
and \U$1597 ( \10658 , RIe1b38d0_3420, \9266 );
and \U$1598 ( \10659 , RIfcc0fe0_7218, \9268 );
and \U$1599 ( \10660 , RIfceaea8_7695, \9270 );
and \U$1600 ( \10661 , RIe1b1f80_3402, \9272 );
and \U$1601 ( \10662 , RIe1b0360_3382, \9274 );
and \U$1602 ( \10663 , RIfcd0760_7394, \9276 );
and \U$1603 ( \10664 , RIf145ec8_5255, \9278 );
and \U$1604 ( \10665 , RIfe9e5e0_8146, \9280 );
and \U$1605 ( \10666 , RIfe9dd70_8140, \9282 );
and \U$1606 ( \10667 , RIe1a7828_3283, \9284 );
and \U$1607 ( \10668 , RIe1a4b28_3251, \9286 );
and \U$1608 ( \10669 , RIe1a1e28_3219, \9288 );
and \U$1609 ( \10670 , RIe19f128_3187, \9290 );
and \U$1610 ( \10671 , RIe18b628_2963, \9292 );
and \U$1611 ( \10672 , RIe177b28_2739, \9294 );
and \U$1612 ( \10673 , RIe225480_4714, \9296 );
and \U$1613 ( \10674 , RIe21a080_4586, \9298 );
and \U$1614 ( \10675 , RIe203880_4330, \9300 );
and \U$1615 ( \10676 , RIe1fd8e0_4262, \9302 );
and \U$1616 ( \10677 , RIe1f6c98_4185, \9304 );
and \U$1617 ( \10678 , RIe1ef7e0_4102, \9306 );
and \U$1618 ( \10679 , RIe1d3ce8_3787, \9308 );
and \U$1619 ( \10680 , RIe1ba7e8_3499, \9310 );
and \U$1620 ( \10681 , RIe1ad660_3350, \9312 );
and \U$1621 ( \10682 , RIe16fc98_2649, \9314 );
or \U$1622 ( \10683 , \10619 , \10620 , \10621 , \10622 , \10623 , \10624 , \10625 , \10626 , \10627 , \10628 , \10629 , \10630 , \10631 , \10632 , \10633 , \10634 , \10635 , \10636 , \10637 , \10638 , \10639 , \10640 , \10641 , \10642 , \10643 , \10644 , \10645 , \10646 , \10647 , \10648 , \10649 , \10650 , \10651 , \10652 , \10653 , \10654 , \10655 , \10656 , \10657 , \10658 , \10659 , \10660 , \10661 , \10662 , \10663 , \10664 , \10665 , \10666 , \10667 , \10668 , \10669 , \10670 , \10671 , \10672 , \10673 , \10674 , \10675 , \10676 , \10677 , \10678 , \10679 , \10680 , \10681 , \10682 );
or \U$1623 ( \10684 , \10618 , \10683 );
_DC g6578 ( \10685_nG6578 , \10684 , \9323 );
and g6579 ( \10686_nG6579 , \10553_nG6577 , \10685_nG6578 );
buf \U$1624 ( \10687 , \10686_nG6579 );
_DC g44da ( \10688_nG44da , \10552 , \9597 );
_DC g455e ( \10689_nG455e , \10684 , \9323 );
xor g455f ( \10690_nG455f , \10688_nG44da , \10689_nG455e );
buf \U$1625 ( \10691 , \10690_nG455f );
and \U$1626 ( \10692 , \10687 , \10691 );
buf \U$1627 ( \10693 , \10692 );
buf g9c0e ( \10694_nG9c0e , \10693 );
and \U$1628 ( \10695 , \10418 , \10694_nG9c0e );
or \U$1629 ( \10696 , 1'b0 , \10695 );
xor \U$1630 ( \10697 , \10417 , \10696 );
xor \U$1631 ( \10698 , \10417 , \10697 );
buf \U$1632 ( \10699 , \10698 );
buf \U$1633 ( \10700 , \10699 );
xor \U$1634 ( \10701 , \10267 , \10400 );
buf g4456 ( \10702_nG4456 , \10701 );
and \U$1637 ( \10703 , \10415_nG4454 , 1'b1 );
xor \U$1638 ( \10704 , \10702_nG4456 , 1'b0 );
not \U$1639 ( \10705 , \10704 );
xor \U$1640 ( \10706 , \10415_nG4454 , \10702_nG4456 );
and \U$1641 ( \10707 , \10705 , \10706 );
and \U$1643 ( \10708 , \10704 , \10694_nG9c0e );
or \U$1644 ( \10709 , 1'b0 , \10708 );
xor \U$1645 ( \10710 , \10703 , \10709 );
and \U$1646 ( \10711 , \10703 , \10710 );
buf \U$1647 ( \10712 , \10711 );
buf \U$1649 ( \10713 , \10712 );
and \U$1650 ( \10714 , \10707 , \10694_nG9c0e );
and \U$1651 ( \10715 , RIdec5108_706, \9333 );
and \U$1652 ( \10716 , RIdec2408_674, \9335 );
and \U$1653 ( \10717 , RIfc93608_6699, \9337 );
and \U$1654 ( \10718 , RIdebf708_642, \9339 );
and \U$1655 ( \10719 , RIfc934a0_6698, \9341 );
and \U$1656 ( \10720 , RIdebca08_610, \9343 );
and \U$1657 ( \10721 , RIdeb9d08_578, \9345 );
and \U$1658 ( \10722 , RIdeb7008_546, \9347 );
and \U$1659 ( \10723 , RIfcdf7d8_7565, \9349 );
and \U$1660 ( \10724 , RIdeb1608_482, \9351 );
and \U$1661 ( \10725 , RIfc78218_6389, \9353 );
and \U$1662 ( \10726 , RIdeae908_450, \9355 );
and \U$1663 ( \10727 , RIfcc8498_7301, \9357 );
and \U$1664 ( \10728 , RIdea9d90_418, \9359 );
and \U$1665 ( \10729 , RIdea3490_386, \9361 );
and \U$1666 ( \10730 , RIde9cb90_354, \9363 );
and \U$1667 ( \10731 , RIee1cc78_4786, \9365 );
and \U$1668 ( \10732 , RIee1bb98_4774, \9367 );
and \U$1669 ( \10733 , RIee1b328_4768, \9369 );
and \U$1670 ( \10734 , RIee1aab8_4762, \9371 );
and \U$1671 ( \10735 , RIde909f8_295, \9373 );
and \U$1672 ( \10736 , RIde8d578_279, \9375 );
and \U$1673 ( \10737 , RIfea8ea0_8238, \9377 );
and \U$1674 ( \10738 , RIde85238_239, \9379 );
and \U$1675 ( \10739 , RIde813e0_220, \9381 );
and \U$1676 ( \10740 , RIfc938d8_6701, \9383 );
and \U$1677 ( \10741 , RIfce5e80_7638, \9385 );
and \U$1678 ( \10742 , RIfcbfd98_7205, \9387 );
and \U$1679 ( \10743 , RIfce8ce8_7671, \9389 );
and \U$1680 ( \10744 , RIe16b4e0_2598, \9391 );
and \U$1681 ( \10745 , RIfea8d38_8237, \9393 );
and \U$1682 ( \10746 , RIfea9f80_8250, \9395 );
and \U$1683 ( \10747 , RIe165108_2527, \9397 );
and \U$1684 ( \10748 , RIe162408_2495, \9399 );
and \U$1685 ( \10749 , RIfc779a8_6383, \9401 );
and \U$1686 ( \10750 , RIe15f708_2463, \9403 );
and \U$1687 ( \10751 , RIfe9dc08_8139, \9405 );
and \U$1688 ( \10752 , RIe15ca08_2431, \9407 );
and \U$1689 ( \10753 , RIe157008_2367, \9409 );
and \U$1690 ( \10754 , RIe154308_2335, \9411 );
and \U$1691 ( \10755 , RIfea7550_8220, \9413 );
and \U$1692 ( \10756 , RIe151608_2303, \9415 );
and \U$1693 ( \10757 , RIfcd6160_7458, \9417 );
and \U$1694 ( \10758 , RIe14e908_2271, \9419 );
and \U$1695 ( \10759 , RIfcd1408_7403, \9421 );
and \U$1696 ( \10760 , RIe14bc08_2239, \9423 );
and \U$1697 ( \10761 , RIe148f08_2207, \9425 );
and \U$1698 ( \10762 , RIe146208_2175, \9427 );
and \U$1699 ( \10763 , RIfceb718_7701, \9429 );
and \U$1700 ( \10764 , RIfcb19c8_7043, \9431 );
and \U$1701 ( \10765 , RIfc93e78_6705, \9433 );
and \U$1702 ( \10766 , RIfce7938_7657, \9435 );
and \U$1703 ( \10767 , RIe140da8_2115, \9437 );
and \U$1704 ( \10768 , RIdf3ecb0_2091, \9439 );
and \U$1705 ( \10769 , RIdf3c988_2066, \9441 );
and \U$1706 ( \10770 , RIfe9daa0_8138, \9443 );
and \U$1707 ( \10771 , RIfce8478_7665, \9445 );
and \U$1708 ( \10772 , RIfcdbf98_7525, \9447 );
and \U$1709 ( \10773 , RIfc776d8_6381, \9449 );
and \U$1710 ( \10774 , RIfc93fe0_6706, \9451 );
and \U$1711 ( \10775 , RIdf354d0_1983, \9453 );
and \U$1712 ( \10776 , RIdf33040_1957, \9455 );
and \U$1713 ( \10777 , RIdf30fe8_1934, \9457 );
and \U$1714 ( \10778 , RIdf2ee28_1910, \9459 );
or \U$1715 ( \10779 , \10715 , \10716 , \10717 , \10718 , \10719 , \10720 , \10721 , \10722 , \10723 , \10724 , \10725 , \10726 , \10727 , \10728 , \10729 , \10730 , \10731 , \10732 , \10733 , \10734 , \10735 , \10736 , \10737 , \10738 , \10739 , \10740 , \10741 , \10742 , \10743 , \10744 , \10745 , \10746 , \10747 , \10748 , \10749 , \10750 , \10751 , \10752 , \10753 , \10754 , \10755 , \10756 , \10757 , \10758 , \10759 , \10760 , \10761 , \10762 , \10763 , \10764 , \10765 , \10766 , \10767 , \10768 , \10769 , \10770 , \10771 , \10772 , \10773 , \10774 , \10775 , \10776 , \10777 , \10778 );
and \U$1716 ( \10780 , RIee2ba20_4955, \9462 );
and \U$1717 ( \10781 , RIfc93ba8_6703, \9464 );
and \U$1718 ( \10782 , RIfc77de0_6386, \9466 );
and \U$1719 ( \10783 , RIee27ad8_4910, \9468 );
and \U$1720 ( \10784 , RIfe9d668_8135, \9470 );
and \U$1721 ( \10785 , RIfea8bd0_8236, \9472 );
and \U$1722 ( \10786 , RIdf26458_1812, \9474 );
and \U$1723 ( \10787 , RIfe9d7d0_8136, \9476 );
and \U$1724 ( \10788 , RIfcb1c98_7045, \9478 );
and \U$1725 ( \10789 , RIee26cc8_4900, \9480 );
and \U$1726 ( \10790 , RIdf22ab0_1771, \9482 );
and \U$1727 ( \10791 , RIfcc0068_7207, \9484 );
and \U$1728 ( \10792 , RIdf21598_1756, \9486 );
and \U$1729 ( \10793 , RIdf1f6a8_1734, \9488 );
and \U$1730 ( \10794 , RIdf1aef0_1683, \9490 );
and \U$1731 ( \10795 , RIfe9d938_8137, \9492 );
and \U$1732 ( \10796 , RIdf16cd8_1636, \9494 );
and \U$1733 ( \10797 , RIdf13fd8_1604, \9496 );
and \U$1734 ( \10798 , RIdf112d8_1572, \9498 );
and \U$1735 ( \10799 , RIdf0e5d8_1540, \9500 );
and \U$1736 ( \10800 , RIdf0b8d8_1508, \9502 );
and \U$1737 ( \10801 , RIdf08bd8_1476, \9504 );
and \U$1738 ( \10802 , RIdf05ed8_1444, \9506 );
and \U$1739 ( \10803 , RIdf031d8_1412, \9508 );
and \U$1740 ( \10804 , RIdefd7d8_1348, \9510 );
and \U$1741 ( \10805 , RIdefaad8_1316, \9512 );
and \U$1742 ( \10806 , RIdef7dd8_1284, \9514 );
and \U$1743 ( \10807 , RIdef50d8_1252, \9516 );
and \U$1744 ( \10808 , RIdef23d8_1220, \9518 );
and \U$1745 ( \10809 , RIdeef6d8_1188, \9520 );
and \U$1746 ( \10810 , RIdeec9d8_1156, \9522 );
and \U$1747 ( \10811 , RIdee9cd8_1124, \9524 );
and \U$1748 ( \10812 , RIfc942b0_6708, \9526 );
and \U$1749 ( \10813 , RIfcde6f8_7553, \9528 );
and \U$1750 ( \10814 , RIfcd1138_7401, \9530 );
and \U$1751 ( \10815 , RIfcde860_7554, \9532 );
and \U$1752 ( \10816 , RIdee4878_1064, \9534 );
and \U$1753 ( \10817 , RIdee2af0_1043, \9536 );
and \U$1754 ( \10818 , RIdee0a98_1020, \9538 );
and \U$1755 ( \10819 , RIdede8d8_996, \9540 );
and \U$1756 ( \10820 , RIfc5c9f0_6076, \9542 );
and \U$1757 ( \10821 , RIee22240_4847, \9544 );
and \U$1758 ( \10822 , RIfcc8768_7303, \9546 );
and \U$1759 ( \10823 , RIee21160_4835, \9548 );
and \U$1760 ( \10824 , RIded95e0_937, \9550 );
and \U$1761 ( \10825 , RIded7150_911, \9552 );
and \U$1762 ( \10826 , RIded5260_889, \9554 );
and \U$1763 ( \10827 , RIfea76b8_8221, \9556 );
and \U$1764 ( \10828 , RIded0508_834, \9558 );
and \U$1765 ( \10829 , RIdecd808_802, \9560 );
and \U$1766 ( \10830 , RIdecab08_770, \9562 );
and \U$1767 ( \10831 , RIdec7e08_738, \9564 );
and \U$1768 ( \10832 , RIdeb4308_514, \9566 );
and \U$1769 ( \10833 , RIde96290_322, \9568 );
and \U$1770 ( \10834 , RIe16df10_2628, \9570 );
and \U$1771 ( \10835 , RIe159d08_2399, \9572 );
and \U$1772 ( \10836 , RIe143508_2143, \9574 );
and \U$1773 ( \10837 , RIdf37f00_2013, \9576 );
and \U$1774 ( \10838 , RIdf2c560_1881, \9578 );
and \U$1775 ( \10839 , RIdf1cde0_1705, \9580 );
and \U$1776 ( \10840 , RIdf004d8_1380, \9582 );
and \U$1777 ( \10841 , RIdee6fd8_1092, \9584 );
and \U$1778 ( \10842 , RIdedbd40_965, \9586 );
and \U$1779 ( \10843 , RIde7c1d8_195, \9588 );
or \U$1780 ( \10844 , \10780 , \10781 , \10782 , \10783 , \10784 , \10785 , \10786 , \10787 , \10788 , \10789 , \10790 , \10791 , \10792 , \10793 , \10794 , \10795 , \10796 , \10797 , \10798 , \10799 , \10800 , \10801 , \10802 , \10803 , \10804 , \10805 , \10806 , \10807 , \10808 , \10809 , \10810 , \10811 , \10812 , \10813 , \10814 , \10815 , \10816 , \10817 , \10818 , \10819 , \10820 , \10821 , \10822 , \10823 , \10824 , \10825 , \10826 , \10827 , \10828 , \10829 , \10830 , \10831 , \10832 , \10833 , \10834 , \10835 , \10836 , \10837 , \10838 , \10839 , \10840 , \10841 , \10842 , \10843 );
or \U$1781 ( \10845 , \10779 , \10844 );
_DC g45e3 ( \10846_nG45e3 , \10845 , \9597 );
and \U$1782 ( \10847 , RIe19d3a0_3166, \9059 );
and \U$1783 ( \10848 , RIe19a6a0_3134, \9061 );
and \U$1784 ( \10849 , RIfcb2c10_7056, \9063 );
and \U$1785 ( \10850 , RIe1979a0_3102, \9065 );
and \U$1786 ( \10851 , RIfc923c0_6686, \9067 );
and \U$1787 ( \10852 , RIe194ca0_3070, \9069 );
and \U$1788 ( \10853 , RIe191fa0_3038, \9071 );
and \U$1789 ( \10854 , RIe18f2a0_3006, \9073 );
and \U$1790 ( \10855 , RIe1898a0_2942, \9075 );
and \U$1791 ( \10856 , RIe186ba0_2910, \9077 );
and \U$1792 ( \10857 , RIfc422a8_5775, \9079 );
and \U$1793 ( \10858 , RIe183ea0_2878, \9081 );
and \U$1794 ( \10859 , RIfcbecb8_7193, \9083 );
and \U$1795 ( \10860 , RIe1811a0_2846, \9085 );
and \U$1796 ( \10861 , RIe17e4a0_2814, \9087 );
and \U$1797 ( \10862 , RIe17b7a0_2782, \9089 );
and \U$1798 ( \10863 , RIf142250_5212, \9091 );
and \U$1799 ( \10864 , RIf140bd0_5196, \9093 );
and \U$1800 ( \10865 , RIfec43f8_8353, \9095 );
and \U$1801 ( \10866 , RIe175968_2715, \9097 );
and \U$1802 ( \10867 , RIfc79b68_6407, \9099 );
and \U$1803 ( \10868 , RIf13efb0_5176, \9101 );
and \U$1804 ( \10869 , RIfc92528_6687, \9103 );
and \U$1805 ( \10870 , RIfcb2aa8_7055, \9105 );
and \U$1806 ( \10871 , RIfcd8320_7482, \9107 );
and \U$1807 ( \10872 , RIfcea200_7686, \9109 );
and \U$1808 ( \10873 , RIfc79898_6405, \9111 );
and \U$1809 ( \10874 , RIe1734d8_2689, \9113 );
and \U$1810 ( \10875 , RIfcd7948_7475, \9115 );
and \U$1811 ( \10876 , RIfcd7678_7473, \9117 );
and \U$1812 ( \10877 , RIf16e170_5712, \9119 );
and \U$1813 ( \10878 , RIfc927f8_6689, \9121 );
and \U$1814 ( \10879 , RIfc92960_6690, \9123 );
and \U$1815 ( \10880 , RIe2236f8_4693, \9125 );
and \U$1816 ( \10881 , RIfc795c8_6403, \9127 );
and \U$1817 ( \10882 , RIe2209f8_4661, \9129 );
and \U$1818 ( \10883 , RIf16ad68_5675, \9131 );
and \U$1819 ( \10884 , RIe21dcf8_4629, \9133 );
and \U$1820 ( \10885 , RIe2182f8_4565, \9135 );
and \U$1821 ( \10886 , RIe2155f8_4533, \9137 );
and \U$1822 ( \10887 , RIfe9d398_8133, \9139 );
and \U$1823 ( \10888 , RIe2128f8_4501, \9141 );
and \U$1824 ( \10889 , RIfcdb9f8_7521, \9143 );
and \U$1825 ( \10890 , RIe20fbf8_4469, \9145 );
and \U$1826 ( \10891 , RIfc41d08_5771, \9147 );
and \U$1827 ( \10892 , RIe20cef8_4437, \9149 );
and \U$1828 ( \10893 , RIe20a1f8_4405, \9151 );
and \U$1829 ( \10894 , RIe2074f8_4373, \9153 );
and \U$1830 ( \10895 , RIfcd7510_7472, \9155 );
and \U$1831 ( \10896 , RIf166010_5620, \9157 );
and \U$1832 ( \10897 , RIfe9d230_8132, \9159 );
and \U$1833 ( \10898 , RIe2008b0_4296, \9161 );
and \U$1834 ( \10899 , RIf165098_5609, \9163 );
and \U$1835 ( \10900 , RIfc41ba0_5770, \9165 );
and \U$1836 ( \10901 , RIfc41a38_5769, \9167 );
and \U$1837 ( \10902 , RIfc92c30_6692, \9169 );
and \U$1838 ( \10903 , RIfc418d0_5768, \9171 );
and \U$1839 ( \10904 , RIfc79190_6400, \9173 );
and \U$1840 ( \10905 , RIe1fcad0_4252, \9175 );
and \U$1841 ( \10906 , RIfec4560_8354, \9177 );
and \U$1842 ( \10907 , RIfc79028_6399, \9179 );
and \U$1843 ( \10908 , RIfcbf258_7197, \9181 );
and \U$1844 ( \10909 , RIfcc1df0_7228, \9183 );
and \U$1845 ( \10910 , RIfcd81b8_7481, \9185 );
or \U$1846 ( \10911 , \10847 , \10848 , \10849 , \10850 , \10851 , \10852 , \10853 , \10854 , \10855 , \10856 , \10857 , \10858 , \10859 , \10860 , \10861 , \10862 , \10863 , \10864 , \10865 , \10866 , \10867 , \10868 , \10869 , \10870 , \10871 , \10872 , \10873 , \10874 , \10875 , \10876 , \10877 , \10878 , \10879 , \10880 , \10881 , \10882 , \10883 , \10884 , \10885 , \10886 , \10887 , \10888 , \10889 , \10890 , \10891 , \10892 , \10893 , \10894 , \10895 , \10896 , \10897 , \10898 , \10899 , \10900 , \10901 , \10902 , \10903 , \10904 , \10905 , \10906 , \10907 , \10908 , \10909 , \10910 );
and \U$1847 ( \10912 , RIfc92d98_6693, \9188 );
and \U$1848 ( \10913 , RIfc5b4d8_6061, \9190 );
and \U$1849 ( \10914 , RIfcd77e0_7474, \9192 );
and \U$1850 ( \10915 , RIe1fa0a0_4222, \9194 );
and \U$1851 ( \10916 , RIf156188_5439, \9196 );
and \U$1852 ( \10917 , RIfe9d500_8134, \9198 );
and \U$1853 ( \10918 , RIf1546d0_5420, \9200 );
and \U$1854 ( \10919 , RIe1f5348_4167, \9202 );
and \U$1855 ( \10920 , RIfec4830_8356, \9204 );
and \U$1856 ( \10921 , RIfec46c8_8355, \9206 );
and \U$1857 ( \10922 , RIf1508f0_5376, \9208 );
and \U$1858 ( \10923 , RIe1f3020_4142, \9210 );
and \U$1859 ( \10924 , RIfce3180_7606, \9212 );
and \U$1860 ( \10925 , RIfce8fb8_7673, \9214 );
and \U$1861 ( \10926 , RIfcbf690_7200, \9216 );
and \U$1862 ( \10927 , RIe1edd28_4083, \9218 );
and \U$1863 ( \10928 , RIe1eb460_4054, \9220 );
and \U$1864 ( \10929 , RIe1e8760_4022, \9222 );
and \U$1865 ( \10930 , RIe1e5a60_3990, \9224 );
and \U$1866 ( \10931 , RIe1e2d60_3958, \9226 );
and \U$1867 ( \10932 , RIe1e0060_3926, \9228 );
and \U$1868 ( \10933 , RIe1dd360_3894, \9230 );
and \U$1869 ( \10934 , RIe1da660_3862, \9232 );
and \U$1870 ( \10935 , RIe1d7960_3830, \9234 );
and \U$1871 ( \10936 , RIe1d1f60_3766, \9236 );
and \U$1872 ( \10937 , RIe1cf260_3734, \9238 );
and \U$1873 ( \10938 , RIe1cc560_3702, \9240 );
and \U$1874 ( \10939 , RIe1c9860_3670, \9242 );
and \U$1875 ( \10940 , RIe1c6b60_3638, \9244 );
and \U$1876 ( \10941 , RIe1c3e60_3606, \9246 );
and \U$1877 ( \10942 , RIe1c1160_3574, \9248 );
and \U$1878 ( \10943 , RIe1be460_3542, \9250 );
and \U$1879 ( \10944 , RIfe9d0c8_8131, \9252 );
and \U$1880 ( \10945 , RIfe9cc90_8128, \9254 );
and \U$1881 ( \10946 , RIe1b9168_3483, \9256 );
and \U$1882 ( \10947 , RIe1b7110_3460, \9258 );
and \U$1883 ( \10948 , RIf14a3b0_5304, \9260 );
and \U$1884 ( \10949 , RIfe9cb28_8127, \9262 );
and \U$1885 ( \10950 , RIfe9cf60_8130, \9264 );
and \U$1886 ( \10951 , RIfe9c9c0_8126, \9266 );
and \U$1887 ( \10952 , RIfce2208_7595, \9268 );
and \U$1888 ( \10953 , RIfce9558_7677, \9270 );
and \U$1889 ( \10954 , RIfe9c858_8125, \9272 );
and \U$1890 ( \10955 , RIfe9cdf8_8129, \9274 );
and \U$1891 ( \10956 , RIf147110_5268, \9276 );
and \U$1892 ( \10957 , RIf146468_5259, \9278 );
and \U$1893 ( \10958 , RIe1ac2b0_3336, \9280 );
and \U$1894 ( \10959 , RIe1aaac8_3319, \9282 );
and \U$1895 ( \10960 , RIe1a87a0_3294, \9284 );
and \U$1896 ( \10961 , RIe1a5aa0_3262, \9286 );
and \U$1897 ( \10962 , RIe1a2da0_3230, \9288 );
and \U$1898 ( \10963 , RIe1a00a0_3198, \9290 );
and \U$1899 ( \10964 , RIe18c5a0_2974, \9292 );
and \U$1900 ( \10965 , RIe178aa0_2750, \9294 );
and \U$1901 ( \10966 , RIe2263f8_4725, \9296 );
and \U$1902 ( \10967 , RIe21aff8_4597, \9298 );
and \U$1903 ( \10968 , RIe2047f8_4341, \9300 );
and \U$1904 ( \10969 , RIe1fe858_4273, \9302 );
and \U$1905 ( \10970 , RIe1f7c10_4196, \9304 );
and \U$1906 ( \10971 , RIe1f0758_4113, \9306 );
and \U$1907 ( \10972 , RIe1d4c60_3798, \9308 );
and \U$1908 ( \10973 , RIe1bb760_3510, \9310 );
and \U$1909 ( \10974 , RIe1ae5d8_3361, \9312 );
and \U$1910 ( \10975 , RIe170c10_2660, \9314 );
or \U$1911 ( \10976 , \10912 , \10913 , \10914 , \10915 , \10916 , \10917 , \10918 , \10919 , \10920 , \10921 , \10922 , \10923 , \10924 , \10925 , \10926 , \10927 , \10928 , \10929 , \10930 , \10931 , \10932 , \10933 , \10934 , \10935 , \10936 , \10937 , \10938 , \10939 , \10940 , \10941 , \10942 , \10943 , \10944 , \10945 , \10946 , \10947 , \10948 , \10949 , \10950 , \10951 , \10952 , \10953 , \10954 , \10955 , \10956 , \10957 , \10958 , \10959 , \10960 , \10961 , \10962 , \10963 , \10964 , \10965 , \10966 , \10967 , \10968 , \10969 , \10970 , \10971 , \10972 , \10973 , \10974 , \10975 );
or \U$1912 ( \10977 , \10911 , \10976 );
_DC g4667 ( \10978_nG4667 , \10977 , \9323 );
xor g4668 ( \10979_nG4668 , \10846_nG45e3 , \10978_nG4667 );
buf \U$1913 ( \10980 , \10979_nG4668 );
xor \U$1914 ( \10981 , \10980 , \10691 );
not \U$1915 ( \10982 , \10691 );
and \U$1916 ( \10983 , \10981 , \10982 );
and \U$1917 ( \10984 , \10687 , \10983 );
_DC g657a ( \10985_nG657a , \10845 , \9597 );
_DC g657b ( \10986_nG657b , \10977 , \9323 );
and g657c ( \10987_nG657c , \10985_nG657a , \10986_nG657b );
buf \U$1918 ( \10988 , \10987_nG657c );
and \U$1919 ( \10989 , \10988 , \10691 );
nor \U$1920 ( \10990 , \10984 , \10989 );
xnor \U$1921 ( \10991 , \10990 , \10980 );
not \U$1922 ( \10992 , \10692 );
and \U$1923 ( \10993 , \10992 , \10980 );
xor \U$1924 ( \10994 , \10991 , \10993 );
buf g9c0b ( \10995_nG9c0b , \10994 );
and \U$1925 ( \10996 , \10704 , \10995_nG9c0b );
or \U$1926 ( \10997 , \10714 , \10996 );
xor \U$1927 ( \10998 , \10703 , \10997 );
buf \U$1928 ( \10999 , \10998 );
buf \U$1930 ( \11000 , \10999 );
and \U$1931 ( \11001 , \10713 , \11000 );
buf \U$1932 ( \11002 , \11001 );
and \U$1933 ( \11003 , \10707 , \10995_nG9c0b );
and \U$1934 ( \11004 , \10988 , \10983 );
and \U$1935 ( \11005 , RIdec6080_717, \9333 );
and \U$1936 ( \11006 , RIdec3380_685, \9335 );
and \U$1937 ( \11007 , RIee204b8_4826, \9337 );
and \U$1938 ( \11008 , RIdec0680_653, \9339 );
and \U$1939 ( \11009 , RIfcd70d8_7469, \9341 );
and \U$1940 ( \11010 , RIdebd980_621, \9343 );
and \U$1941 ( \11011 , RIdebac80_589, \9345 );
and \U$1942 ( \11012 , RIdeb7f80_557, \9347 );
and \U$1943 ( \11013 , RIfcbe448_7187, \9349 );
and \U$1944 ( \11014 , RIdeb2580_493, \9351 );
and \U$1945 ( \11015 , RIfcb3480_7062, \9353 );
and \U$1946 ( \11016 , RIdeaf880_461, \9355 );
and \U$1947 ( \11017 , RIfc43928_5791, \9357 );
and \U$1948 ( \11018 , RIdeac1a8_429, \9359 );
and \U$1949 ( \11019 , RIdea58a8_397, \9361 );
and \U$1950 ( \11020 , RIde9efa8_365, \9363 );
and \U$1951 ( \11021 , RIfcd88c0_7486, \9365 );
and \U$1952 ( \11022 , RIee1c408_4780, \9367 );
and \U$1953 ( \11023 , RIfcc77f0_7292, \9369 );
and \U$1954 ( \11024 , RIfea04d0_8168, \9371 );
and \U$1955 ( \11025 , RIde92438_303, \9373 );
and \U$1956 ( \11026 , RIde8ec70_286, \9375 );
and \U$1957 ( \11027 , RIde8aad0_266, \9377 );
and \U$1958 ( \11028 , RIde86930_246, \9379 );
and \U$1959 ( \11029 , RIfca31c0_6878, \9381 );
and \U$1960 ( \11030 , RIfc59a20_6042, \9383 );
and \U$1961 ( \11031 , RIfcd1de0_7410, \9385 );
and \U$1962 ( \11032 , RIfc91448_6675, \9387 );
and \U$1963 ( \11033 , RIfc97280_6742, \9389 );
and \U$1964 ( \11034 , RIe16c188_2607, \9391 );
and \U$1965 ( \11035 , RIfc97118_6741, \9393 );
and \U$1966 ( \11036 , RIe168948_2567, \9395 );
and \U$1967 ( \11037 , RIe166080_2538, \9397 );
and \U$1968 ( \11038 , RIe163380_2506, \9399 );
and \U$1969 ( \11039 , RIee37ac8_5092, \9401 );
and \U$1970 ( \11040 , RIe160680_2474, \9403 );
and \U$1971 ( \11041 , RIfcd1c78_7409, \9405 );
and \U$1972 ( \11042 , RIe15d980_2442, \9407 );
and \U$1973 ( \11043 , RIe157f80_2378, \9409 );
and \U$1974 ( \11044 , RIe155280_2346, \9411 );
and \U$1975 ( \11045 , RIfc3f530_5746, \9413 );
and \U$1976 ( \11046 , RIe152580_2314, \9415 );
and \U$1977 ( \11047 , RIee35368_5064, \9417 );
and \U$1978 ( \11048 , RIe14f880_2282, \9419 );
and \U$1979 ( \11049 , RIfc7a3d8_6413, \9421 );
and \U$1980 ( \11050 , RIe14cb80_2250, \9423 );
and \U$1981 ( \11051 , RIe149e80_2218, \9425 );
and \U$1982 ( \11052 , RIe147180_2186, \9427 );
and \U$1983 ( \11053 , RIfc42b18_5781, \9429 );
and \U$1984 ( \11054 , RIfc7a270_6412, \9431 );
and \U$1985 ( \11055 , RIfc5a560_6050, \9433 );
and \U$1986 ( \11056 , RIfc96b78_6737, \9435 );
and \U$1987 ( \11057 , RIfea6fb0_8216, \9437 );
and \U$1988 ( \11058 , RIe13f5c0_2098, \9439 );
and \U$1989 ( \11059 , RIdf3d4c8_2074, \9441 );
and \U$1990 ( \11060 , RIdf3b038_2048, \9443 );
and \U$1991 ( \11061 , RIfce5bb0_7636, \9445 );
and \U$1992 ( \11062 , RIee2fc38_5002, \9447 );
and \U$1993 ( \11063 , RIfc91cb8_6681, \9449 );
and \U$1994 ( \11064 , RIee2d910_4977, \9451 );
and \U$1995 ( \11065 , RIdf362e0_1993, \9453 );
and \U$1996 ( \11066 , RIdf33e50_1967, \9455 );
and \U$1997 ( \11067 , RIdf31c90_1943, \9457 );
and \U$1998 ( \11068 , RIdf2fda0_1921, \9459 );
or \U$1999 ( \11069 , \11005 , \11006 , \11007 , \11008 , \11009 , \11010 , \11011 , \11012 , \11013 , \11014 , \11015 , \11016 , \11017 , \11018 , \11019 , \11020 , \11021 , \11022 , \11023 , \11024 , \11025 , \11026 , \11027 , \11028 , \11029 , \11030 , \11031 , \11032 , \11033 , \11034 , \11035 , \11036 , \11037 , \11038 , \11039 , \11040 , \11041 , \11042 , \11043 , \11044 , \11045 , \11046 , \11047 , \11048 , \11049 , \11050 , \11051 , \11052 , \11053 , \11054 , \11055 , \11056 , \11057 , \11058 , \11059 , \11060 , \11061 , \11062 , \11063 , \11064 , \11065 , \11066 , \11067 , \11068 );
and \U$2000 ( \11070 , RIfc43658_5789, \9462 );
and \U$2001 ( \11071 , RIfc59e58_6045, \9464 );
and \U$2002 ( \11072 , RIfc96fb0_6740, \9466 );
and \U$2003 ( \11073 , RIfc7ac48_6419, \9468 );
and \U$2004 ( \11074 , RIfea0368_8167, \9470 );
and \U$2005 ( \11075 , RIdf28bb8_1840, \9472 );
and \U$2006 ( \11076 , RIdf26cc8_1818, \9474 );
and \U$2007 ( \11077 , RIdf25210_1799, \9476 );
and \U$2008 ( \11078 , RIfc91718_6677, \9478 );
and \U$2009 ( \11079 , RIfcb3318_7061, \9480 );
and \U$2010 ( \11080 , RIfc919e8_6679, \9482 );
and \U$2011 ( \11081 , RIfc91880_6678, \9484 );
and \U$2012 ( \11082 , RIfc430b8_5785, \9486 );
and \U$2013 ( \11083 , RIdf20350_1743, \9488 );
and \U$2014 ( \11084 , RIfc7a978_6417, \9490 );
and \U$2015 ( \11085 , RIdf19e10_1671, \9492 );
and \U$2016 ( \11086 , RIdf17c50_1647, \9494 );
and \U$2017 ( \11087 , RIdf14f50_1615, \9496 );
and \U$2018 ( \11088 , RIdf12250_1583, \9498 );
and \U$2019 ( \11089 , RIdf0f550_1551, \9500 );
and \U$2020 ( \11090 , RIdf0c850_1519, \9502 );
and \U$2021 ( \11091 , RIdf09b50_1487, \9504 );
and \U$2022 ( \11092 , RIdf06e50_1455, \9506 );
and \U$2023 ( \11093 , RIdf04150_1423, \9508 );
and \U$2024 ( \11094 , RIdefe750_1359, \9510 );
and \U$2025 ( \11095 , RIdefba50_1327, \9512 );
and \U$2026 ( \11096 , RIdef8d50_1295, \9514 );
and \U$2027 ( \11097 , RIdef6050_1263, \9516 );
and \U$2028 ( \11098 , RIdef3350_1231, \9518 );
and \U$2029 ( \11099 , RIdef0650_1199, \9520 );
and \U$2030 ( \11100 , RIdeed950_1167, \9522 );
and \U$2031 ( \11101 , RIdeeac50_1135, \9524 );
and \U$2032 ( \11102 , RIfcd1b10_7408, \9526 );
and \U$2033 ( \11103 , RIfc968a8_6735, \9528 );
and \U$2034 ( \11104 , RIfc91f88_6683, \9530 );
and \U$2035 ( \11105 , RIfcdfc10_7568, \9532 );
and \U$2036 ( \11106 , RIfea99e0_8246, \9534 );
and \U$2037 ( \11107 , RIdee3630_1051, \9536 );
and \U$2038 ( \11108 , RIdee1308_1026, \9538 );
and \U$2039 ( \11109 , RIdedf2b0_1003, \9540 );
and \U$2040 ( \11110 , RIfcc7d90_7296, \9542 );
and \U$2041 ( \11111 , RIfcd85f0_7484, \9544 );
and \U$2042 ( \11112 , RIfce3888_7611, \9546 );
and \U$2043 ( \11113 , RIfc5a830_6052, \9548 );
and \U$2044 ( \11114 , RIdeda3f0_947, \9550 );
and \U$2045 ( \11115 , RIfea9878_8245, \9552 );
and \U$2046 ( \11116 , RIded5f08_898, \9554 );
and \U$2047 ( \11117 , RIded37a8_870, \9556 );
and \U$2048 ( \11118 , RIded1480_845, \9558 );
and \U$2049 ( \11119 , RIdece780_813, \9560 );
and \U$2050 ( \11120 , RIdecba80_781, \9562 );
and \U$2051 ( \11121 , RIdec8d80_749, \9564 );
and \U$2052 ( \11122 , RIdeb5280_525, \9566 );
and \U$2053 ( \11123 , RIde986a8_333, \9568 );
and \U$2054 ( \11124 , RIe16ee88_2639, \9570 );
and \U$2055 ( \11125 , RIe15ac80_2410, \9572 );
and \U$2056 ( \11126 , RIe144480_2154, \9574 );
and \U$2057 ( \11127 , RIdf38e78_2024, \9576 );
and \U$2058 ( \11128 , RIdf2d4d8_1892, \9578 );
and \U$2059 ( \11129 , RIdf1dd58_1716, \9580 );
and \U$2060 ( \11130 , RIdf01450_1391, \9582 );
and \U$2061 ( \11131 , RIdee7f50_1103, \9584 );
and \U$2062 ( \11132 , RIdedccb8_976, \9586 );
and \U$2063 ( \11133 , RIde7e5f0_206, \9588 );
or \U$2064 ( \11134 , \11070 , \11071 , \11072 , \11073 , \11074 , \11075 , \11076 , \11077 , \11078 , \11079 , \11080 , \11081 , \11082 , \11083 , \11084 , \11085 , \11086 , \11087 , \11088 , \11089 , \11090 , \11091 , \11092 , \11093 , \11094 , \11095 , \11096 , \11097 , \11098 , \11099 , \11100 , \11101 , \11102 , \11103 , \11104 , \11105 , \11106 , \11107 , \11108 , \11109 , \11110 , \11111 , \11112 , \11113 , \11114 , \11115 , \11116 , \11117 , \11118 , \11119 , \11120 , \11121 , \11122 , \11123 , \11124 , \11125 , \11126 , \11127 , \11128 , \11129 , \11130 , \11131 , \11132 , \11133 );
or \U$2065 ( \11135 , \11069 , \11134 );
_DC g657d ( \11136_nG657d , \11135 , \9597 );
and \U$2066 ( \11137 , RIe19e318_3177, \9059 );
and \U$2067 ( \11138 , RIe19b618_3145, \9061 );
and \U$2068 ( \11139 , RIfc8f3f0_6652, \9063 );
and \U$2069 ( \11140 , RIe198918_3113, \9065 );
and \U$2070 ( \11141 , RIf144b18_5241, \9067 );
and \U$2071 ( \11142 , RIe195c18_3081, \9069 );
and \U$2072 ( \11143 , RIe192f18_3049, \9071 );
and \U$2073 ( \11144 , RIe190218_3017, \9073 );
and \U$2074 ( \11145 , RIe18a818_2953, \9075 );
and \U$2075 ( \11146 , RIe187b18_2921, \9077 );
and \U$2076 ( \11147 , RIf143d08_5231, \9079 );
and \U$2077 ( \11148 , RIe184e18_2889, \9081 );
and \U$2078 ( \11149 , RIfcb3cf0_7068, \9083 );
and \U$2079 ( \11150 , RIe182118_2857, \9085 );
and \U$2080 ( \11151 , RIe17f418_2825, \9087 );
and \U$2081 ( \11152 , RIe17c718_2793, \9089 );
and \U$2082 ( \11153 , RIfc448a0_5802, \9091 );
and \U$2083 ( \11154 , RIf141170_5200, \9093 );
and \U$2084 ( \11155 , RIfc7c9d0_6440, \9095 );
and \U$2085 ( \11156 , RIfea0098_8165, \9097 );
and \U$2086 ( \11157 , RIfc57e00_6022, \9099 );
and \U$2087 ( \11158 , RIf13f550_5180, \9101 );
and \U$2088 ( \11159 , RIfcd6e08_7467, \9103 );
and \U$2089 ( \11160 , RIee3d900_5159, \9105 );
and \U$2090 ( \11161 , RIfc8f6c0_6654, \9107 );
and \U$2091 ( \11162 , RIfce0048_7571, \9109 );
and \U$2092 ( \11163 , RIfca27e8_6871, \9111 );
and \U$2093 ( \11164 , RIe1742e8_2699, \9113 );
and \U$2094 ( \11165 , RIfc7c700_6438, \9115 );
and \U$2095 ( \11166 , RIfc8f990_6656, \9117 );
and \U$2096 ( \11167 , RIfce9828_7679, \9119 );
and \U$2097 ( \11168 , RIfc583a0_6026, \9121 );
and \U$2098 ( \11169 , RIf16cdc0_5698, \9123 );
and \U$2099 ( \11170 , RIe224670_4704, \9125 );
and \U$2100 ( \11171 , RIf16c118_5689, \9127 );
and \U$2101 ( \11172 , RIe221970_4672, \9129 );
and \U$2102 ( \11173 , RIfc58508_6027, \9131 );
and \U$2103 ( \11174 , RIe21ec70_4640, \9133 );
and \U$2104 ( \11175 , RIe219270_4576, \9135 );
and \U$2105 ( \11176 , RIe216570_4544, \9137 );
and \U$2106 ( \11177 , RIfc3ff08_5753, \9139 );
and \U$2107 ( \11178 , RIe213870_4512, \9141 );
and \U$2108 ( \11179 , RIf1696e8_5659, \9143 );
and \U$2109 ( \11180 , RIe210b70_4480, \9145 );
and \U$2110 ( \11181 , RIfc58940_6030, \9147 );
and \U$2111 ( \11182 , RIe20de70_4448, \9149 );
and \U$2112 ( \11183 , RIe20b170_4416, \9151 );
and \U$2113 ( \11184 , RIe208470_4384, \9153 );
and \U$2114 ( \11185 , RIfc8fc60_6658, \9155 );
and \U$2115 ( \11186 , RIfc97820_6746, \9157 );
and \U$2116 ( \11187 , RIe202ea8_4323, \9159 );
and \U$2117 ( \11188 , RIe201288_4303, \9161 );
and \U$2118 ( \11189 , RIfcc27c8_7235, \9163 );
and \U$2119 ( \11190 , RIfcdfee0_7570, \9165 );
and \U$2120 ( \11191 , RIfc44198_5797, \9167 );
and \U$2121 ( \11192 , RIfc58670_6028, \9169 );
and \U$2122 ( \11193 , RIf1608e0_5558, \9171 );
and \U$2123 ( \11194 , RIf15e9f0_5536, \9173 );
and \U$2124 ( \11195 , RIfe9ff30_8164, \9175 );
and \U$2125 ( \11196 , RIe1fc0f8_4245, \9177 );
and \U$2126 ( \11197 , RIfc7be90_6432, \9179 );
and \U$2127 ( \11198 , RIf15bb88_5503, \9181 );
and \U$2128 ( \11199 , RIfcd8cf8_7489, \9183 );
and \U$2129 ( \11200 , RIfcd8e60_7490, \9185 );
or \U$2130 ( \11201 , \11137 , \11138 , \11139 , \11140 , \11141 , \11142 , \11143 , \11144 , \11145 , \11146 , \11147 , \11148 , \11149 , \11150 , \11151 , \11152 , \11153 , \11154 , \11155 , \11156 , \11157 , \11158 , \11159 , \11160 , \11161 , \11162 , \11163 , \11164 , \11165 , \11166 , \11167 , \11168 , \11169 , \11170 , \11171 , \11172 , \11173 , \11174 , \11175 , \11176 , \11177 , \11178 , \11179 , \11180 , \11181 , \11182 , \11183 , \11184 , \11185 , \11186 , \11187 , \11188 , \11189 , \11190 , \11191 , \11192 , \11193 , \11194 , \11195 , \11196 , \11197 , \11198 , \11199 , \11200 );
and \U$2131 ( \11202 , RIfca2d88_6875, \9188 );
and \U$2132 ( \11203 , RIfcbdea8_7183, \9190 );
and \U$2133 ( \11204 , RIfcb3a20_7066, \9192 );
and \U$2134 ( \11205 , RIe1fabe0_4230, \9194 );
and \U$2135 ( \11206 , RIfc90098_6661, \9196 );
and \U$2136 ( \11207 , RIfc90200_6662, \9198 );
and \U$2137 ( \11208 , RIfcd20b0_7412, \9200 );
and \U$2138 ( \11209 , RIe1f6158_4177, \9202 );
and \U$2139 ( \11210 , RIfc904d0_6664, \9204 );
and \U$2140 ( \11211 , RIfca2ef0_6876, \9206 );
and \U$2141 ( \11212 , RIfc97550_6744, \9208 );
and \U$2142 ( \11213 , RIe1f3e30_4152, \9210 );
and \U$2143 ( \11214 , RIfc59048_6035, \9212 );
and \U$2144 ( \11215 , RIfc907a0_6666, \9214 );
and \U$2145 ( \11216 , RIfc90638_6665, \9216 );
and \U$2146 ( \11217 , RIe1eeb38_4093, \9218 );
and \U$2147 ( \11218 , RIe1ec3d8_4065, \9220 );
and \U$2148 ( \11219 , RIe1e96d8_4033, \9222 );
and \U$2149 ( \11220 , RIe1e69d8_4001, \9224 );
and \U$2150 ( \11221 , RIe1e3cd8_3969, \9226 );
and \U$2151 ( \11222 , RIe1e0fd8_3937, \9228 );
and \U$2152 ( \11223 , RIe1de2d8_3905, \9230 );
and \U$2153 ( \11224 , RIe1db5d8_3873, \9232 );
and \U$2154 ( \11225 , RIe1d88d8_3841, \9234 );
and \U$2155 ( \11226 , RIe1d2ed8_3777, \9236 );
and \U$2156 ( \11227 , RIe1d01d8_3745, \9238 );
and \U$2157 ( \11228 , RIe1cd4d8_3713, \9240 );
and \U$2158 ( \11229 , RIe1ca7d8_3681, \9242 );
and \U$2159 ( \11230 , RIe1c7ad8_3649, \9244 );
and \U$2160 ( \11231 , RIe1c4dd8_3617, \9246 );
and \U$2161 ( \11232 , RIe1c20d8_3585, \9248 );
and \U$2162 ( \11233 , RIe1bf3d8_3553, \9250 );
and \U$2163 ( \11234 , RIfcc73b8_7289, \9252 );
and \U$2164 ( \11235 , RIfce3cc0_7614, \9254 );
and \U$2165 ( \11236 , RIe1b9e10_3492, \9256 );
and \U$2166 ( \11237 , RIe1b7c50_3468, \9258 );
and \U$2167 ( \11238 , RIfcd6f70_7468, \9260 );
and \U$2168 ( \11239 , RIf149e10_5300, \9262 );
and \U$2169 ( \11240 , RIe1b5a90_3444, \9264 );
and \U$2170 ( \11241 , RIfea0200_8166, \9266 );
and \U$2171 ( \11242 , RIfc90bd8_6669, \9268 );
and \U$2172 ( \11243 , RIfcdfd78_7569, \9270 );
and \U$2173 ( \11244 , RIe1b2ef8_3413, \9272 );
and \U$2174 ( \11245 , RIe1b15a8_3395, \9274 );
and \U$2175 ( \11246 , RIfc973e8_6743, \9276 );
and \U$2176 ( \11247 , RIfcc7520_7290, \9278 );
and \U$2177 ( \11248 , RIe1acdf0_3344, \9280 );
and \U$2178 ( \11249 , RIe1ab608_3327, \9282 );
and \U$2179 ( \11250 , RIe1a9718_3305, \9284 );
and \U$2180 ( \11251 , RIe1a6a18_3273, \9286 );
and \U$2181 ( \11252 , RIe1a3d18_3241, \9288 );
and \U$2182 ( \11253 , RIe1a1018_3209, \9290 );
and \U$2183 ( \11254 , RIe18d518_2985, \9292 );
and \U$2184 ( \11255 , RIe179a18_2761, \9294 );
and \U$2185 ( \11256 , RIe227370_4736, \9296 );
and \U$2186 ( \11257 , RIe21bf70_4608, \9298 );
and \U$2187 ( \11258 , RIe205770_4352, \9300 );
and \U$2188 ( \11259 , RIe1ff7d0_4284, \9302 );
and \U$2189 ( \11260 , RIe1f8b88_4207, \9304 );
and \U$2190 ( \11261 , RIe1f16d0_4124, \9306 );
and \U$2191 ( \11262 , RIe1d5bd8_3809, \9308 );
and \U$2192 ( \11263 , RIe1bc6d8_3521, \9310 );
and \U$2193 ( \11264 , RIe1af550_3372, \9312 );
and \U$2194 ( \11265 , RIe171b88_2671, \9314 );
or \U$2195 ( \11266 , \11202 , \11203 , \11204 , \11205 , \11206 , \11207 , \11208 , \11209 , \11210 , \11211 , \11212 , \11213 , \11214 , \11215 , \11216 , \11217 , \11218 , \11219 , \11220 , \11221 , \11222 , \11223 , \11224 , \11225 , \11226 , \11227 , \11228 , \11229 , \11230 , \11231 , \11232 , \11233 , \11234 , \11235 , \11236 , \11237 , \11238 , \11239 , \11240 , \11241 , \11242 , \11243 , \11244 , \11245 , \11246 , \11247 , \11248 , \11249 , \11250 , \11251 , \11252 , \11253 , \11254 , \11255 , \11256 , \11257 , \11258 , \11259 , \11260 , \11261 , \11262 , \11263 , \11264 , \11265 );
or \U$2196 ( \11267 , \11201 , \11266 );
_DC g657e ( \11268_nG657e , \11267 , \9323 );
and g657f ( \11269_nG657f , \11136_nG657d , \11268_nG657e );
buf \U$2197 ( \11270 , \11269_nG657f );
and \U$2198 ( \11271 , \11270 , \10691 );
nor \U$2199 ( \11272 , \11004 , \11271 );
xnor \U$2200 ( \11273 , \11272 , \10980 );
_DC g46ec ( \11274_nG46ec , \11135 , \9597 );
_DC g4770 ( \11275_nG4770 , \11267 , \9323 );
xor g4771 ( \11276_nG4771 , \11274_nG46ec , \11275_nG4770 );
buf \U$2201 ( \11277 , \11276_nG4771 );
xor \U$2202 ( \11278 , \11277 , \10980 );
and \U$2203 ( \11279 , \10687 , \11278 );
xor \U$2204 ( \11280 , \11273 , \11279 );
and \U$2205 ( \11281 , \10991 , \10993 );
xor \U$2206 ( \11282 , \11280 , \11281 );
buf g9c08 ( \11283_nG9c08 , \11282 );
and \U$2207 ( \11284 , \10704 , \11283_nG9c08 );
or \U$2208 ( \11285 , \11003 , \11284 );
xor \U$2209 ( \11286 , \10703 , \11285 );
buf \U$2210 ( \11287 , \11286 );
buf \U$2212 ( \11288 , \11287 );
xor \U$2213 ( \11289 , \11002 , \11288 );
and \U$2214 ( \11290 , \10700 , \11289 );
and \U$2215 ( \11291 , \11002 , \11288 );
buf \U$2216 ( \11292 , \11291 );
and \U$2217 ( \11293 , \10417 , \10697 );
buf \U$2218 ( \11294 , \11293 );
buf \U$2220 ( \11295 , \11294 );
and \U$2221 ( \11296 , \10421 , \10694_nG9c0e );
and \U$2222 ( \11297 , \10418 , \10995_nG9c0b );
or \U$2223 ( \11298 , \11296 , \11297 );
xor \U$2224 ( \11299 , \10417 , \11298 );
buf \U$2225 ( \11300 , \11299 );
buf \U$2227 ( \11301 , \11300 );
xor \U$2228 ( \11302 , \11295 , \11301 );
buf \U$2229 ( \11303 , \11302 );
xor \U$2230 ( \11304 , \11292 , \11303 );
and \U$2231 ( \11305 , \10707 , \11283_nG9c08 );
and \U$2232 ( \11306 , RIdec64b8_720, \9333 );
and \U$2233 ( \11307 , RIdec37b8_688, \9335 );
and \U$2234 ( \11308 , RIfc8daa0_6634, \9337 );
and \U$2235 ( \11309 , RIdec0ab8_656, \9339 );
and \U$2236 ( \11310 , RIfc56348_6003, \9341 );
and \U$2237 ( \11311 , RIdebddb8_624, \9343 );
and \U$2238 ( \11312 , RIdebb0b8_592, \9345 );
and \U$2239 ( \11313 , RIdeb83b8_560, \9347 );
and \U$2240 ( \11314 , RIfc98798_6757, \9349 );
and \U$2241 ( \11315 , RIdeb29b8_496, \9351 );
and \U$2242 ( \11316 , RIfcbd098_7173, \9353 );
and \U$2243 ( \11317 , RIdeafcb8_464, \9355 );
and \U$2244 ( \11318 , RIfc8dc08_6635, \9357 );
and \U$2245 ( \11319 , RIdeacb80_432, \9359 );
and \U$2246 ( \11320 , RIdea6280_400, \9361 );
and \U$2247 ( \11321 , RIde9f980_368, \9363 );
and \U$2248 ( \11322 , RIfcd6868_7463, \9365 );
and \U$2249 ( \11323 , RIfc8ded8_6637, \9367 );
and \U$2250 ( \11324 , RIfc7dd80_6454, \9369 );
and \U$2251 ( \11325 , RIfc56618_6005, \9371 );
and \U$2252 ( \11326 , RIde92e10_306, \9373 );
and \U$2253 ( \11327 , RIde8f300_288, \9375 );
and \U$2254 ( \11328 , RIde8b160_268, \9377 );
and \U$2255 ( \11329 , RIde86fc0_248, \9379 );
and \U$2256 ( \11330 , RIde82ad8_227, \9381 );
and \U$2257 ( \11331 , RIfc8e040_6638, \9383 );
and \U$2258 ( \11332 , RIfcd96d0_7496, \9385 );
and \U$2259 ( \11333 , RIfca1e10_6864, \9387 );
and \U$2260 ( \11334 , RIfcbd200_7174, \9389 );
and \U$2261 ( \11335 , RIe16c5c0_2610, \9391 );
and \U$2262 ( \11336 , RIe16a298_2585, \9393 );
and \U$2263 ( \11337 , RIe168ab0_2568, \9395 );
and \U$2264 ( \11338 , RIe1664b8_2541, \9397 );
and \U$2265 ( \11339 , RIe1637b8_2509, \9399 );
and \U$2266 ( \11340 , RIee37f00_5095, \9401 );
and \U$2267 ( \11341 , RIe160ab8_2477, \9403 );
and \U$2268 ( \11342 , RIfc8ea18_6645, \9405 );
and \U$2269 ( \11343 , RIe15ddb8_2445, \9407 );
and \U$2270 ( \11344 , RIe1583b8_2381, \9409 );
and \U$2271 ( \11345 , RIe1556b8_2349, \9411 );
and \U$2272 ( \11346 , RIfe9f828_8159, \9413 );
and \U$2273 ( \11347 , RIe1529b8_2317, \9415 );
and \U$2274 ( \11348 , RIfe9f990_8160, \9417 );
and \U$2275 ( \11349 , RIe14fcb8_2285, \9419 );
and \U$2276 ( \11350 , RIfcbd368_7175, \9421 );
and \U$2277 ( \11351 , RIe14cfb8_2253, \9423 );
and \U$2278 ( \11352 , RIe14a2b8_2221, \9425 );
and \U$2279 ( \11353 , RIe1475b8_2189, \9427 );
and \U$2280 ( \11354 , RIfc8ee50_6648, \9429 );
and \U$2281 ( \11355 , RIfc45278_5809, \9431 );
and \U$2282 ( \11356 , RIfc98360_6754, \9433 );
and \U$2283 ( \11357 , RIfca2248_6867, \9435 );
and \U$2284 ( \11358 , RIe141d20_2126, \9437 );
and \U$2285 ( \11359 , RIe13f9f8_2101, \9439 );
and \U$2286 ( \11360 , RIdf3d900_2077, \9441 );
and \U$2287 ( \11361 , RIdf3b470_2051, \9443 );
and \U$2288 ( \11362 , RIfcd6ca0_7466, \9445 );
and \U$2289 ( \11363 , RIee2ff08_5004, \9447 );
and \U$2290 ( \11364 , RIfc8ece8_6647, \9449 );
and \U$2291 ( \11365 , RIee2dd48_4980, \9451 );
and \U$2292 ( \11366 , RIdf36718_1996, \9453 );
and \U$2293 ( \11367 , RIdf34120_1969, \9455 );
and \U$2294 ( \11368 , RIdf31f60_1945, \9457 );
and \U$2295 ( \11369 , RIfe9f6c0_8158, \9459 );
or \U$2296 ( \11370 , \11306 , \11307 , \11308 , \11309 , \11310 , \11311 , \11312 , \11313 , \11314 , \11315 , \11316 , \11317 , \11318 , \11319 , \11320 , \11321 , \11322 , \11323 , \11324 , \11325 , \11326 , \11327 , \11328 , \11329 , \11330 , \11331 , \11332 , \11333 , \11334 , \11335 , \11336 , \11337 , \11338 , \11339 , \11340 , \11341 , \11342 , \11343 , \11344 , \11345 , \11346 , \11347 , \11348 , \11349 , \11350 , \11351 , \11352 , \11353 , \11354 , \11355 , \11356 , \11357 , \11358 , \11359 , \11360 , \11361 , \11362 , \11363 , \11364 , \11365 , \11366 , \11367 , \11368 , \11369 );
and \U$2297 ( \11371 , RIfcb4560_7074, \9462 );
and \U$2298 ( \11372 , RIfc45db8_5817, \9464 );
and \U$2299 ( \11373 , RIfc8e1a8_6639, \9466 );
and \U$2300 ( \11374 , RIfc7d678_6449, \9468 );
and \U$2301 ( \11375 , RIdf2aee0_1865, \9470 );
and \U$2302 ( \11376 , RIdf28ff0_1843, \9472 );
and \U$2303 ( \11377 , RIdf26e30_1819, \9474 );
and \U$2304 ( \11378 , RIdf25378_1800, \9476 );
and \U$2305 ( \11379 , RIfcb43f8_7073, \9478 );
and \U$2306 ( \11380 , RIfc8e748_6643, \9480 );
and \U$2307 ( \11381 , RIdf23488_1778, \9482 );
and \U$2308 ( \11382 , RIfcc2c00_7238, \9484 );
and \U$2309 ( \11383 , RIdf21e08_1762, \9486 );
and \U$2310 ( \11384 , RIdf20788_1746, \9488 );
and \U$2311 ( \11385 , RIdf1b760_1689, \9490 );
and \U$2312 ( \11386 , RIdf1a248_1674, \9492 );
and \U$2313 ( \11387 , RIdf18088_1650, \9494 );
and \U$2314 ( \11388 , RIdf15388_1618, \9496 );
and \U$2315 ( \11389 , RIdf12688_1586, \9498 );
and \U$2316 ( \11390 , RIdf0f988_1554, \9500 );
and \U$2317 ( \11391 , RIdf0cc88_1522, \9502 );
and \U$2318 ( \11392 , RIdf09f88_1490, \9504 );
and \U$2319 ( \11393 , RIdf07288_1458, \9506 );
and \U$2320 ( \11394 , RIdf04588_1426, \9508 );
and \U$2321 ( \11395 , RIdefeb88_1362, \9510 );
and \U$2322 ( \11396 , RIdefbe88_1330, \9512 );
and \U$2323 ( \11397 , RIdef9188_1298, \9514 );
and \U$2324 ( \11398 , RIdef6488_1266, \9516 );
and \U$2325 ( \11399 , RIdef3788_1234, \9518 );
and \U$2326 ( \11400 , RIdef0a88_1202, \9520 );
and \U$2327 ( \11401 , RIdeedd88_1170, \9522 );
and \U$2328 ( \11402 , RIdeeb088_1138, \9524 );
and \U$2329 ( \11403 , RIfc8efb8_6649, \9526 );
and \U$2330 ( \11404 , RIfc44e40_5806, \9528 );
and \U$2331 ( \11405 , RIfc57860_6018, \9530 );
and \U$2332 ( \11406 , RIfca23b0_6868, \9532 );
and \U$2333 ( \11407 , RIfe9faf8_8161, \9534 );
and \U$2334 ( \11408 , RIdee3900_1053, \9536 );
and \U$2335 ( \11409 , RIdee1740_1029, \9538 );
and \U$2336 ( \11410 , RIdedf6e8_1006, \9540 );
and \U$2337 ( \11411 , RIfcbd4d0_7176, \9542 );
and \U$2338 ( \11412 , RIee22678_4850, \9544 );
and \U$2339 ( \11413 , RIfc98090_6752, \9546 );
and \U$2340 ( \11414 , RIee21598_4838, \9548 );
and \U$2341 ( \11415 , RIfe9fc60_8162, \9550 );
and \U$2342 ( \11416 , RIded80c8_922, \9552 );
and \U$2343 ( \11417 , RIfe9fdc8_8163, \9554 );
and \U$2344 ( \11418 , RIded3be0_873, \9556 );
and \U$2345 ( \11419 , RIded18b8_848, \9558 );
and \U$2346 ( \11420 , RIdecebb8_816, \9560 );
and \U$2347 ( \11421 , RIdecbeb8_784, \9562 );
and \U$2348 ( \11422 , RIdec91b8_752, \9564 );
and \U$2349 ( \11423 , RIdeb56b8_528, \9566 );
and \U$2350 ( \11424 , RIde99080_336, \9568 );
and \U$2351 ( \11425 , RIe16f2c0_2642, \9570 );
and \U$2352 ( \11426 , RIe15b0b8_2413, \9572 );
and \U$2353 ( \11427 , RIe1448b8_2157, \9574 );
and \U$2354 ( \11428 , RIdf392b0_2027, \9576 );
and \U$2355 ( \11429 , RIdf2d910_1895, \9578 );
and \U$2356 ( \11430 , RIdf1e190_1719, \9580 );
and \U$2357 ( \11431 , RIdf01888_1394, \9582 );
and \U$2358 ( \11432 , RIdee8388_1106, \9584 );
and \U$2359 ( \11433 , RIdedd0f0_979, \9586 );
and \U$2360 ( \11434 , RIde7efc8_209, \9588 );
or \U$2361 ( \11435 , \11371 , \11372 , \11373 , \11374 , \11375 , \11376 , \11377 , \11378 , \11379 , \11380 , \11381 , \11382 , \11383 , \11384 , \11385 , \11386 , \11387 , \11388 , \11389 , \11390 , \11391 , \11392 , \11393 , \11394 , \11395 , \11396 , \11397 , \11398 , \11399 , \11400 , \11401 , \11402 , \11403 , \11404 , \11405 , \11406 , \11407 , \11408 , \11409 , \11410 , \11411 , \11412 , \11413 , \11414 , \11415 , \11416 , \11417 , \11418 , \11419 , \11420 , \11421 , \11422 , \11423 , \11424 , \11425 , \11426 , \11427 , \11428 , \11429 , \11430 , \11431 , \11432 , \11433 , \11434 );
or \U$2362 ( \11436 , \11370 , \11435 );
_DC g47f5 ( \11437_nG47f5 , \11436 , \9597 );
and \U$2363 ( \11438 , RIe19e750_3180, \9059 );
and \U$2364 ( \11439 , RIe19ba50_3148, \9061 );
and \U$2365 ( \11440 , RIfc479d8_5837, \9063 );
and \U$2366 ( \11441 , RIe198d50_3116, \9065 );
and \U$2367 ( \11442 , RIfe9f558_8157, \9067 );
and \U$2368 ( \11443 , RIe196050_3084, \9069 );
and \U$2369 ( \11444 , RIe193350_3052, \9071 );
and \U$2370 ( \11445 , RIe190650_3020, \9073 );
and \U$2371 ( \11446 , RIe18ac50_2956, \9075 );
and \U$2372 ( \11447 , RIe187f50_2924, \9077 );
and \U$2373 ( \11448 , RIfc47870_5836, \9079 );
and \U$2374 ( \11449 , RIe185250_2892, \9081 );
and \U$2375 ( \11450 , RIf142ef8_5221, \9083 );
and \U$2376 ( \11451 , RIe182550_2860, \9085 );
and \U$2377 ( \11452 , RIe17f850_2828, \9087 );
and \U$2378 ( \11453 , RIe17cb50_2796, \9089 );
and \U$2379 ( \11454 , RIfcb5208_7083, \9091 );
and \U$2380 ( \11455 , RIfcbc6c0_7166, \9093 );
and \U$2381 ( \11456 , RIe177588_2735, \9095 );
and \U$2382 ( \11457 , RIe176610_2724, \9097 );
and \U$2383 ( \11458 , RIf13fdc0_5186, \9099 );
and \U$2384 ( \11459 , RIfe9f3f0_8156, \9101 );
and \U$2385 ( \11460 , RIfce40f8_7617, \9103 );
and \U$2386 ( \11461 , RIfc47708_5835, \9105 );
and \U$2387 ( \11462 , RIfc47438_5833, \9107 );
and \U$2388 ( \11463 , RIfca15a0_6858, \9109 );
and \U$2389 ( \11464 , RIfc99170_6764, \9111 );
and \U$2390 ( \11465 , RIe1745b8_2701, \9113 );
and \U$2391 ( \11466 , RIfc8cc90_6624, \9115 );
and \U$2392 ( \11467 , RIfc556a0_5994, \9117 );
and \U$2393 ( \11468 , RIfc7ee60_6466, \9119 );
and \U$2394 ( \11469 , RIfce8e50_7672, \9121 );
and \U$2395 ( \11470 , RIfe9f288_8155, \9123 );
and \U$2396 ( \11471 , RIe224aa8_4707, \9125 );
and \U$2397 ( \11472 , RIfc55808_5995, \9127 );
and \U$2398 ( \11473 , RIe221da8_4675, \9129 );
and \U$2399 ( \11474 , RIfcb50a0_7082, \9131 );
and \U$2400 ( \11475 , RIe21f0a8_4643, \9133 );
and \U$2401 ( \11476 , RIe2196a8_4579, \9135 );
and \U$2402 ( \11477 , RIe2169a8_4547, \9137 );
and \U$2403 ( \11478 , RIfcbc828_7167, \9139 );
and \U$2404 ( \11479 , RIe213ca8_4515, \9141 );
and \U$2405 ( \11480 , RIfc47000_5830, \9143 );
and \U$2406 ( \11481 , RIe210fa8_4483, \9145 );
and \U$2407 ( \11482 , RIfcbc990_7168, \9147 );
and \U$2408 ( \11483 , RIe20e2a8_4451, \9149 );
and \U$2409 ( \11484 , RIe20b5a8_4419, \9151 );
and \U$2410 ( \11485 , RIe2088a8_4387, \9153 );
and \U$2411 ( \11486 , RIfc46bc8_5827, \9155 );
and \U$2412 ( \11487 , RIfcd6598_7461, \9157 );
and \U$2413 ( \11488 , RIe2032e0_4326, \9159 );
and \U$2414 ( \11489 , RIe2016c0_4306, \9161 );
and \U$2415 ( \11490 , RIfc98ea0_6762, \9163 );
and \U$2416 ( \11491 , RIfc7eb90_6464, \9165 );
and \U$2417 ( \11492 , RIfce0318_7573, \9167 );
and \U$2418 ( \11493 , RIfcbcaf8_7169, \9169 );
and \U$2419 ( \11494 , RIfc8cf60_6626, \9171 );
and \U$2420 ( \11495 , RIfcb4dd0_7080, \9173 );
and \U$2421 ( \11496 , RIe1fd340_4258, \9175 );
and \U$2422 ( \11497 , RIe1fc260_4246, \9177 );
and \U$2423 ( \11498 , RIf15cf38_5517, \9179 );
and \U$2424 ( \11499 , RIfe9f120_8154, \9181 );
and \U$2425 ( \11500 , RIfc7ea28_6463, \9183 );
and \U$2426 ( \11501 , RIfc8d0c8_6627, \9185 );
or \U$2427 ( \11502 , \11438 , \11439 , \11440 , \11441 , \11442 , \11443 , \11444 , \11445 , \11446 , \11447 , \11448 , \11449 , \11450 , \11451 , \11452 , \11453 , \11454 , \11455 , \11456 , \11457 , \11458 , \11459 , \11460 , \11461 , \11462 , \11463 , \11464 , \11465 , \11466 , \11467 , \11468 , \11469 , \11470 , \11471 , \11472 , \11473 , \11474 , \11475 , \11476 , \11477 , \11478 , \11479 , \11480 , \11481 , \11482 , \11483 , \11484 , \11485 , \11486 , \11487 , \11488 , \11489 , \11490 , \11491 , \11492 , \11493 , \11494 , \11495 , \11496 , \11497 , \11498 , \11499 , \11500 , \11501 );
and \U$2428 ( \11503 , RIfcbcc60_7170, \9188 );
and \U$2429 ( \11504 , RIfc98bd0_6760, \9190 );
and \U$2430 ( \11505 , RIfce2d48_7603, \9192 );
and \U$2431 ( \11506 , RIe1fb018_4233, \9194 );
and \U$2432 ( \11507 , RIfc55f10_6000, \9196 );
and \U$2433 ( \11508 , RIfc7e8c0_6462, \9198 );
and \U$2434 ( \11509 , RIfc8d230_6628, \9200 );
and \U$2435 ( \11510 , RIe1f6590_4180, \9202 );
and \U$2436 ( \11511 , RIfce58e0_7634, \9204 );
and \U$2437 ( \11512 , RIfc468f8_5825, \9206 );
and \U$2438 ( \11513 , RIfcc2ed0_7240, \9208 );
and \U$2439 ( \11514 , RIe1f4100_4154, \9210 );
and \U$2440 ( \11515 , RIfceedf0_7740, \9212 );
and \U$2441 ( \11516 , RIfc8d398_6629, \9214 );
and \U$2442 ( \11517 , RIfc8d500_6630, \9216 );
and \U$2443 ( \11518 , RIe1eef70_4096, \9218 );
and \U$2444 ( \11519 , RIe1ec810_4068, \9220 );
and \U$2445 ( \11520 , RIe1e9b10_4036, \9222 );
and \U$2446 ( \11521 , RIe1e6e10_4004, \9224 );
and \U$2447 ( \11522 , RIe1e4110_3972, \9226 );
and \U$2448 ( \11523 , RIe1e1410_3940, \9228 );
and \U$2449 ( \11524 , RIe1de710_3908, \9230 );
and \U$2450 ( \11525 , RIe1dba10_3876, \9232 );
and \U$2451 ( \11526 , RIe1d8d10_3844, \9234 );
and \U$2452 ( \11527 , RIe1d3310_3780, \9236 );
and \U$2453 ( \11528 , RIe1d0610_3748, \9238 );
and \U$2454 ( \11529 , RIe1cd910_3716, \9240 );
and \U$2455 ( \11530 , RIe1cac10_3684, \9242 );
and \U$2456 ( \11531 , RIe1c7f10_3652, \9244 );
and \U$2457 ( \11532 , RIe1c5210_3620, \9246 );
and \U$2458 ( \11533 , RIe1c2510_3588, \9248 );
and \U$2459 ( \11534 , RIe1bf810_3556, \9250 );
and \U$2460 ( \11535 , RIf14d0b0_5336, \9252 );
and \U$2461 ( \11536 , RIfe9efb8_8153, \9254 );
and \U$2462 ( \11537 , RIe1ba248_3495, \9256 );
and \U$2463 ( \11538 , RIe1b8088_3471, \9258 );
and \U$2464 ( \11539 , RIfec4dd0_8360, \9260 );
and \U$2465 ( \11540 , RIfec50a0_8362, \9262 );
and \U$2466 ( \11541 , RIe1b5ec8_3447, \9264 );
and \U$2467 ( \11542 , RIe1b46e0_3430, \9266 );
and \U$2468 ( \11543 , RIfcb4998_7077, \9268 );
and \U$2469 ( \11544 , RIfcb4c68_7079, \9270 );
and \U$2470 ( \11545 , RIfec5370_8364, \9272 );
and \U$2471 ( \11546 , RIfe9ee50_8152, \9274 );
and \U$2472 ( \11547 , RIfcbcdc8_7171, \9276 );
and \U$2473 ( \11548 , RIfc46358_5821, \9278 );
and \U$2474 ( \11549 , RIfec5208_8363, \9280 );
and \U$2475 ( \11550 , RIfec4f38_8361, \9282 );
and \U$2476 ( \11551 , RIe1a9b50_3308, \9284 );
and \U$2477 ( \11552 , RIe1a6e50_3276, \9286 );
and \U$2478 ( \11553 , RIe1a4150_3244, \9288 );
and \U$2479 ( \11554 , RIe1a1450_3212, \9290 );
and \U$2480 ( \11555 , RIe18d950_2988, \9292 );
and \U$2481 ( \11556 , RIe179e50_2764, \9294 );
and \U$2482 ( \11557 , RIe2277a8_4739, \9296 );
and \U$2483 ( \11558 , RIe21c3a8_4611, \9298 );
and \U$2484 ( \11559 , RIe205ba8_4355, \9300 );
and \U$2485 ( \11560 , RIe1ffc08_4287, \9302 );
and \U$2486 ( \11561 , RIe1f8fc0_4210, \9304 );
and \U$2487 ( \11562 , RIe1f1b08_4127, \9306 );
and \U$2488 ( \11563 , RIe1d6010_3812, \9308 );
and \U$2489 ( \11564 , RIe1bcb10_3524, \9310 );
and \U$2490 ( \11565 , RIe1af988_3375, \9312 );
and \U$2491 ( \11566 , RIe171fc0_2674, \9314 );
or \U$2492 ( \11567 , \11503 , \11504 , \11505 , \11506 , \11507 , \11508 , \11509 , \11510 , \11511 , \11512 , \11513 , \11514 , \11515 , \11516 , \11517 , \11518 , \11519 , \11520 , \11521 , \11522 , \11523 , \11524 , \11525 , \11526 , \11527 , \11528 , \11529 , \11530 , \11531 , \11532 , \11533 , \11534 , \11535 , \11536 , \11537 , \11538 , \11539 , \11540 , \11541 , \11542 , \11543 , \11544 , \11545 , \11546 , \11547 , \11548 , \11549 , \11550 , \11551 , \11552 , \11553 , \11554 , \11555 , \11556 , \11557 , \11558 , \11559 , \11560 , \11561 , \11562 , \11563 , \11564 , \11565 , \11566 );
or \U$2493 ( \11568 , \11502 , \11567 );
_DC g4879 ( \11569_nG4879 , \11568 , \9323 );
xor g487a ( \11570_nG487a , \11437_nG47f5 , \11569_nG4879 );
buf \U$2494 ( \11571 , \11570_nG487a );
xor \U$2495 ( \11572 , \11571 , \11277 );
not \U$2496 ( \11573 , \11278 );
and \U$2497 ( \11574 , \11572 , \11573 );
and \U$2498 ( \11575 , \10687 , \11574 );
and \U$2499 ( \11576 , \10988 , \11278 );
nor \U$2500 ( \11577 , \11575 , \11576 );
and \U$2501 ( \11578 , \11277 , \10980 );
not \U$2502 ( \11579 , \11578 );
and \U$2503 ( \11580 , \11571 , \11579 );
xnor \U$2504 ( \11581 , \11577 , \11580 );
and \U$2505 ( \11582 , \11270 , \10983 );
_DC g6580 ( \11583_nG6580 , \11436 , \9597 );
_DC g6581 ( \11584_nG6581 , \11568 , \9323 );
and g6582 ( \11585_nG6582 , \11583_nG6580 , \11584_nG6581 );
buf \U$2506 ( \11586 , \11585_nG6582 );
and \U$2507 ( \11587 , \11586 , \10691 );
nor \U$2508 ( \11588 , \11582 , \11587 );
xnor \U$2509 ( \11589 , \11588 , \10980 );
not \U$2510 ( \11590 , \11279 );
and \U$2511 ( \11591 , \11590 , \11580 );
xor \U$2512 ( \11592 , \11589 , \11591 );
xor \U$2513 ( \11593 , \11581 , \11592 );
and \U$2514 ( \11594 , \11273 , \11279 );
and \U$2515 ( \11595 , \11280 , \11281 );
or \U$2516 ( \11596 , \11594 , \11595 );
xor \U$2517 ( \11597 , \11593 , \11596 );
buf g9c05 ( \11598_nG9c05 , \11597 );
and \U$2518 ( \11599 , \10704 , \11598_nG9c05 );
or \U$2519 ( \11600 , \11305 , \11599 );
xor \U$2520 ( \11601 , \10703 , \11600 );
buf \U$2521 ( \11602 , \11601 );
buf \U$2523 ( \11603 , \11602 );
xor \U$2524 ( \11604 , \11304 , \11603 );
and \U$2525 ( \11605 , \11290 , \11604 );
and \U$2526 ( \11606 , RIdec6788_722, \9059 );
and \U$2527 ( \11607 , RIdec3a88_690, \9061 );
and \U$2528 ( \11608 , RIee20788_4828, \9063 );
and \U$2529 ( \11609 , RIdec0d88_658, \9065 );
and \U$2530 ( \11610 , RIee1f810_4817, \9067 );
and \U$2531 ( \11611 , RIdebe088_626, \9069 );
and \U$2532 ( \11612 , RIdebb388_594, \9071 );
and \U$2533 ( \11613 , RIdeb8688_562, \9073 );
and \U$2534 ( \11614 , RIfc9b1c8_6787, \9075 );
and \U$2535 ( \11615 , RIdeb2c88_498, \9077 );
and \U$2536 ( \11616 , RIfce1f38_7593, \9079 );
and \U$2537 ( \11617 , RIdeaff88_466, \9081 );
and \U$2538 ( \11618 , RIfc892e8_6583, \9083 );
and \U$2539 ( \11619 , RIdead210_434, \9085 );
and \U$2540 ( \11620 , RIdea6910_402, \9087 );
and \U$2541 ( \11621 , RIdea0010_370, \9089 );
and \U$2542 ( \11622 , RIee1d650_4793, \9091 );
and \U$2543 ( \11623 , RIee1c570_4781, \9093 );
and \U$2544 ( \11624 , RIee1b5f8_4770, \9095 );
and \U$2545 ( \11625 , RIee1aef0_4765, \9097 );
and \U$2546 ( \11626 , RIfe99888_8091, \9099 );
and \U$2547 ( \11627 , RIfe99450_8088, \9101 );
and \U$2548 ( \11628 , RIfe99720_8090, \9103 );
and \U$2549 ( \11629 , RIfe995b8_8089, \9105 );
and \U$2550 ( \11630 , RIde83168_229, \9107 );
and \U$2551 ( \11631 , RIfcc43e8_7255, \9109 );
and \U$2552 ( \11632 , RIfcd5a58_7453, \9111 );
and \U$2553 ( \11633 , RIfc89450_6584, \9113 );
and \U$2554 ( \11634 , RIfcc5798_7269, \9115 );
and \U$2555 ( \11635 , RIe16c890_2612, \9117 );
and \U$2556 ( \11636 , RIe16a568_2587, \9119 );
and \U$2557 ( \11637 , RIe168d80_2570, \9121 );
and \U$2558 ( \11638 , RIe166788_2543, \9123 );
and \U$2559 ( \11639 , RIe163a88_2511, \9125 );
and \U$2560 ( \11640 , RIfc83618_6517, \9127 );
and \U$2561 ( \11641 , RIe160d88_2479, \9129 );
and \U$2562 ( \11642 , RIee36718_5078, \9131 );
and \U$2563 ( \11643 , RIe15e088_2447, \9133 );
and \U$2564 ( \11644 , RIe158688_2383, \9135 );
and \U$2565 ( \11645 , RIe155988_2351, \9137 );
and \U$2566 ( \11646 , RIfc3f800_5748, \9139 );
and \U$2567 ( \11647 , RIe152c88_2319, \9141 );
and \U$2568 ( \11648 , RIfc895b8_6585, \9143 );
and \U$2569 ( \11649 , RIe14ff88_2287, \9145 );
and \U$2570 ( \11650 , RIfc51cf8_5953, \9147 );
and \U$2571 ( \11651 , RIe14d288_2255, \9149 );
and \U$2572 ( \11652 , RIe14a588_2223, \9151 );
and \U$2573 ( \11653 , RIe147888_2191, \9153 );
and \U$2574 ( \11654 , RIee34990_5057, \9155 );
and \U$2575 ( \11655 , RIee338b0_5045, \9157 );
and \U$2576 ( \11656 , RIfc831e0_6514, \9159 );
and \U$2577 ( \11657 , RIfcd3b68_7431, \9161 );
and \U$2578 ( \11658 , RIe141ff0_2128, \9163 );
and \U$2579 ( \11659 , RIe13fcc8_2103, \9165 );
and \U$2580 ( \11660 , RIdf3dbd0_2079, \9167 );
and \U$2581 ( \11661 , RIdf3b740_2053, \9169 );
and \U$2582 ( \11662 , RIfcb6f90_7104, \9171 );
and \U$2583 ( \11663 , RIee301d8_5006, \9173 );
and \U$2584 ( \11664 , RIfcba938_7145, \9175 );
and \U$2585 ( \11665 , RIee2e018_4982, \9177 );
and \U$2586 ( \11666 , RIdf369e8_1998, \9179 );
and \U$2587 ( \11667 , RIdf343f0_1971, \9181 );
and \U$2588 ( \11668 , RIdf32230_1947, \9183 );
and \U$2589 ( \11669 , RIfe99e28_8095, \9185 );
or \U$2590 ( \11670 , \11606 , \11607 , \11608 , \11609 , \11610 , \11611 , \11612 , \11613 , \11614 , \11615 , \11616 , \11617 , \11618 , \11619 , \11620 , \11621 , \11622 , \11623 , \11624 , \11625 , \11626 , \11627 , \11628 , \11629 , \11630 , \11631 , \11632 , \11633 , \11634 , \11635 , \11636 , \11637 , \11638 , \11639 , \11640 , \11641 , \11642 , \11643 , \11644 , \11645 , \11646 , \11647 , \11648 , \11649 , \11650 , \11651 , \11652 , \11653 , \11654 , \11655 , \11656 , \11657 , \11658 , \11659 , \11660 , \11661 , \11662 , \11663 , \11664 , \11665 , \11666 , \11667 , \11668 , \11669 );
and \U$2591 ( \11671 , RIfc83078_6513, \9188 );
and \U$2592 ( \11672 , RIfcb6e28_7103, \9190 );
and \U$2593 ( \11673 , RIfc9ad90_6784, \9192 );
and \U$2594 ( \11674 , RIfcbad70_7148, \9194 );
and \U$2595 ( \11675 , RIdf2b1b0_1867, \9196 );
and \U$2596 ( \11676 , RIdf292c0_1845, \9198 );
and \U$2597 ( \11677 , RIfe99b58_8093, \9200 );
and \U$2598 ( \11678 , RIfe999f0_8092, \9202 );
and \U$2599 ( \11679 , RIfc9ac28_6783, \9204 );
and \U$2600 ( \11680 , RIfc4a9a8_5871, \9206 );
and \U$2601 ( \11681 , RIdf23758_1780, \9208 );
and \U$2602 ( \11682 , RIfc82da8_6511, \9210 );
and \U$2603 ( \11683 , RIdf220d8_1764, \9212 );
and \U$2604 ( \11684 , RIdf20a58_1748, \9214 );
and \U$2605 ( \11685 , RIdf1ba30_1691, \9216 );
and \U$2606 ( \11686 , RIfe99cc0_8094, \9218 );
and \U$2607 ( \11687 , RIdf18358_1652, \9220 );
and \U$2608 ( \11688 , RIdf15658_1620, \9222 );
and \U$2609 ( \11689 , RIdf12958_1588, \9224 );
and \U$2610 ( \11690 , RIdf0fc58_1556, \9226 );
and \U$2611 ( \11691 , RIdf0cf58_1524, \9228 );
and \U$2612 ( \11692 , RIdf0a258_1492, \9230 );
and \U$2613 ( \11693 , RIdf07558_1460, \9232 );
and \U$2614 ( \11694 , RIdf04858_1428, \9234 );
and \U$2615 ( \11695 , RIdefee58_1364, \9236 );
and \U$2616 ( \11696 , RIdefc158_1332, \9238 );
and \U$2617 ( \11697 , RIdef9458_1300, \9240 );
and \U$2618 ( \11698 , RIdef6758_1268, \9242 );
and \U$2619 ( \11699 , RIdef3a58_1236, \9244 );
and \U$2620 ( \11700 , RIdef0d58_1204, \9246 );
and \U$2621 ( \11701 , RIdeee058_1172, \9248 );
and \U$2622 ( \11702 , RIdeeb358_1140, \9250 );
and \U$2623 ( \11703 , RIee25918_4886, \9252 );
and \U$2624 ( \11704 , RIee24b08_4876, \9254 );
and \U$2625 ( \11705 , RIfc52568_5959, \9256 );
and \U$2626 ( \11706 , RIfc826a0_6506, \9258 );
and \U$2627 ( \11707 , RIdee5958_1076, \9260 );
and \U$2628 ( \11708 , RIdee3bd0_1055, \9262 );
and \U$2629 ( \11709 , RIfe99f90_8096, \9264 );
and \U$2630 ( \11710 , RIdedf9b8_1008, \9266 );
and \U$2631 ( \11711 , RIfce4800_7622, \9268 );
and \U$2632 ( \11712 , RIfc89b58_6589, \9270 );
and \U$2633 ( \11713 , RIfc9f3e0_6834, \9272 );
and \U$2634 ( \11714 , RIfc82538_6505, \9274 );
and \U$2635 ( \11715 , RIdeda828_950, \9276 );
and \U$2636 ( \11716 , RIded8398_924, \9278 );
and \U$2637 ( \11717 , RIfeabe70_8272, \9280 );
and \U$2638 ( \11718 , RIded3eb0_875, \9282 );
and \U$2639 ( \11719 , RIded1b88_850, \9284 );
and \U$2640 ( \11720 , RIdecee88_818, \9286 );
and \U$2641 ( \11721 , RIdecc188_786, \9288 );
and \U$2642 ( \11722 , RIdec9488_754, \9290 );
and \U$2643 ( \11723 , RIdeb5988_530, \9292 );
and \U$2644 ( \11724 , RIde99710_338, \9294 );
and \U$2645 ( \11725 , RIe16f590_2644, \9296 );
and \U$2646 ( \11726 , RIe15b388_2415, \9298 );
and \U$2647 ( \11727 , RIe144b88_2159, \9300 );
and \U$2648 ( \11728 , RIdf39580_2029, \9302 );
and \U$2649 ( \11729 , RIdf2dbe0_1897, \9304 );
and \U$2650 ( \11730 , RIdf1e460_1721, \9306 );
and \U$2651 ( \11731 , RIdf01b58_1396, \9308 );
and \U$2652 ( \11732 , RIdee8658_1108, \9310 );
and \U$2653 ( \11733 , RIdedd3c0_981, \9312 );
and \U$2654 ( \11734 , RIde7f658_211, \9314 );
or \U$2655 ( \11735 , \11671 , \11672 , \11673 , \11674 , \11675 , \11676 , \11677 , \11678 , \11679 , \11680 , \11681 , \11682 , \11683 , \11684 , \11685 , \11686 , \11687 , \11688 , \11689 , \11690 , \11691 , \11692 , \11693 , \11694 , \11695 , \11696 , \11697 , \11698 , \11699 , \11700 , \11701 , \11702 , \11703 , \11704 , \11705 , \11706 , \11707 , \11708 , \11709 , \11710 , \11711 , \11712 , \11713 , \11714 , \11715 , \11716 , \11717 , \11718 , \11719 , \11720 , \11721 , \11722 , \11723 , \11724 , \11725 , \11726 , \11727 , \11728 , \11729 , \11730 , \11731 , \11732 , \11733 , \11734 );
or \U$2656 ( \11736 , \11670 , \11735 );
_DC g2fb7 ( \11737_nG2fb7 , \11736 , \9323 );
buf \U$2657 ( \11738 , \11737_nG2fb7 );
and \U$2658 ( \11739 , RIe19ea20_3182, \9333 );
and \U$2659 ( \11740 , RIe19bd20_3150, \9335 );
and \U$2660 ( \11741 , RIf145928_5251, \9337 );
and \U$2661 ( \11742 , RIe199020_3118, \9339 );
and \U$2662 ( \11743 , RIfe98910_8080, \9341 );
and \U$2663 ( \11744 , RIe196320_3086, \9343 );
and \U$2664 ( \11745 , RIe193620_3054, \9345 );
and \U$2665 ( \11746 , RIe190920_3022, \9347 );
and \U$2666 ( \11747 , RIe18af20_2958, \9349 );
and \U$2667 ( \11748 , RIe188220_2926, \9351 );
and \U$2668 ( \11749 , RIf143e70_5232, \9353 );
and \U$2669 ( \11750 , RIe185520_2894, \9355 );
and \U$2670 ( \11751 , RIfc95c00_6726, \9357 );
and \U$2671 ( \11752 , RIe182820_2862, \9359 );
and \U$2672 ( \11753 , RIe17fb20_2830, \9361 );
and \U$2673 ( \11754 , RIe17ce20_2798, \9363 );
and \U$2674 ( \11755 , RIf142520_5214, \9365 );
and \U$2675 ( \11756 , RIf141440_5202, \9367 );
and \U$2676 ( \11757 , RIe1776f0_2736, \9369 );
and \U$2677 ( \11758 , RIfeab8d0_8268, \9371 );
and \U$2678 ( \11759 , RIfcc5bd0_7272, \9373 );
and \U$2679 ( \11760 , RIfc62dc8_6147, \9375 );
and \U$2680 ( \11761 , RIee3e710_5169, \9377 );
and \U$2681 ( \11762 , RIfc9cb18_6805, \9379 );
and \U$2682 ( \11763 , RIee3c820_5147, \9381 );
and \U$2683 ( \11764 , RIee3b470_5133, \9383 );
and \U$2684 ( \11765 , RIee3a390_5121, \9385 );
and \U$2685 ( \11766 , RIe174888_2703, \9387 );
and \U$2686 ( \11767 , RIf170498_5737, \9389 );
and \U$2687 ( \11768 , RIfc68660_6210, \9391 );
and \U$2688 ( \11769 , RIf16e878_5717, \9393 );
and \U$2689 ( \11770 , RIfc6ea38_6281, \9395 );
and \U$2690 ( \11771 , RIfe98d48_8083, \9397 );
and \U$2691 ( \11772 , RIe224d78_4709, \9399 );
and \U$2692 ( \11773 , RIf16c280_5690, \9401 );
and \U$2693 ( \11774 , RIe222078_4677, \9403 );
and \U$2694 ( \11775 , RIf16b308_5679, \9405 );
and \U$2695 ( \11776 , RIe21f378_4645, \9407 );
and \U$2696 ( \11777 , RIe219978_4581, \9409 );
and \U$2697 ( \11778 , RIe216c78_4549, \9411 );
and \U$2698 ( \11779 , RIf16a390_5668, \9413 );
and \U$2699 ( \11780 , RIe213f78_4517, \9415 );
and \U$2700 ( \11781 , RIf169b20_5662, \9417 );
and \U$2701 ( \11782 , RIe211278_4485, \9419 );
and \U$2702 ( \11783 , RIf1681d0_5644, \9421 );
and \U$2703 ( \11784 , RIe20e578_4453, \9423 );
and \U$2704 ( \11785 , RIe20b878_4421, \9425 );
and \U$2705 ( \11786 , RIe208b78_4389, \9427 );
and \U$2706 ( \11787 , RIfcd4ae0_7442, \9429 );
and \U$2707 ( \11788 , RIfc61478_6129, \9431 );
and \U$2708 ( \11789 , RIfeab060_8262, \9433 );
and \U$2709 ( \11790 , RIe201990_4308, \9435 );
and \U$2710 ( \11791 , RIfc70ec8_6307, \9437 );
and \U$2711 ( \11792 , RIfc70928_6303, \9439 );
and \U$2712 ( \11793 , RIfcec528_7711, \9441 );
and \U$2713 ( \11794 , RIfcbe880_7190, \9443 );
and \U$2714 ( \11795 , RIf160d18_5561, \9445 );
and \U$2715 ( \11796 , RIf15ee28_5539, \9447 );
and \U$2716 ( \11797 , RIfe98be0_8082, \9449 );
and \U$2717 ( \11798 , RIfe98eb0_8084, \9451 );
and \U$2718 ( \11799 , RIf15d0a0_5518, \9453 );
and \U$2719 ( \11800 , RIf15bcf0_5504, \9455 );
and \U$2720 ( \11801 , RIfcd4540_7438, \9457 );
and \U$2721 ( \11802 , RIf159e00_5482, \9459 );
or \U$2722 ( \11803 , \11739 , \11740 , \11741 , \11742 , \11743 , \11744 , \11745 , \11746 , \11747 , \11748 , \11749 , \11750 , \11751 , \11752 , \11753 , \11754 , \11755 , \11756 , \11757 , \11758 , \11759 , \11760 , \11761 , \11762 , \11763 , \11764 , \11765 , \11766 , \11767 , \11768 , \11769 , \11770 , \11771 , \11772 , \11773 , \11774 , \11775 , \11776 , \11777 , \11778 , \11779 , \11780 , \11781 , \11782 , \11783 , \11784 , \11785 , \11786 , \11787 , \11788 , \11789 , \11790 , \11791 , \11792 , \11793 , \11794 , \11795 , \11796 , \11797 , \11798 , \11799 , \11800 , \11801 , \11802 );
and \U$2723 ( \11804 , RIf1592c0_5474, \9462 );
and \U$2724 ( \11805 , RIf158078_5461, \9464 );
and \U$2725 ( \11806 , RIfca3a30_6884, \9466 );
and \U$2726 ( \11807 , RIfea7988_8223, \9468 );
and \U$2727 ( \11808 , RIf156728_5443, \9470 );
and \U$2728 ( \11809 , RIf155be8_5435, \9472 );
and \U$2729 ( \11810 , RIf154b08_5423, \9474 );
and \U$2730 ( \11811 , RIfe98a78_8081, \9476 );
and \U$2731 ( \11812 , RIf1538c0_5410, \9478 );
and \U$2732 ( \11813 , RIf1520d8_5393, \9480 );
and \U$2733 ( \11814 , RIf150e90_5380, \9482 );
and \U$2734 ( \11815 , RIe1f43d0_4156, \9484 );
and \U$2735 ( \11816 , RIf14fdb0_5368, \9486 );
and \U$2736 ( \11817 , RIfcd2380_7414, \9488 );
and \U$2737 ( \11818 , RIf14e2f8_5349, \9490 );
and \U$2738 ( \11819 , RIe1ef240_4098, \9492 );
and \U$2739 ( \11820 , RIe1ecae0_4070, \9494 );
and \U$2740 ( \11821 , RIe1e9de0_4038, \9496 );
and \U$2741 ( \11822 , RIe1e70e0_4006, \9498 );
and \U$2742 ( \11823 , RIe1e43e0_3974, \9500 );
and \U$2743 ( \11824 , RIe1e16e0_3942, \9502 );
and \U$2744 ( \11825 , RIe1de9e0_3910, \9504 );
and \U$2745 ( \11826 , RIe1dbce0_3878, \9506 );
and \U$2746 ( \11827 , RIe1d8fe0_3846, \9508 );
and \U$2747 ( \11828 , RIe1d35e0_3782, \9510 );
and \U$2748 ( \11829 , RIe1d08e0_3750, \9512 );
and \U$2749 ( \11830 , RIe1cdbe0_3718, \9514 );
and \U$2750 ( \11831 , RIe1caee0_3686, \9516 );
and \U$2751 ( \11832 , RIe1c81e0_3654, \9518 );
and \U$2752 ( \11833 , RIe1c54e0_3622, \9520 );
and \U$2753 ( \11834 , RIe1c27e0_3590, \9522 );
and \U$2754 ( \11835 , RIe1bfae0_3558, \9524 );
and \U$2755 ( \11836 , RIfc44b70_5804, \9526 );
and \U$2756 ( \11837 , RIf14bd00_5322, \9528 );
and \U$2757 ( \11838 , RIfe992e8_8087, \9530 );
and \U$2758 ( \11839 , RIfe987a8_8079, \9532 );
and \U$2759 ( \11840 , RIf14a950_5308, \9534 );
and \U$2760 ( \11841 , RIf149f78_5301, \9536 );
and \U$2761 ( \11842 , RIfe99180_8086, \9538 );
and \U$2762 ( \11843 , RIfe98640_8078, \9540 );
and \U$2763 ( \11844 , RIf149438_5293, \9542 );
and \U$2764 ( \11845 , RIfcec7f8_7713, \9544 );
and \U$2765 ( \11846 , RIfe984d8_8077, \9546 );
and \U$2766 ( \11847 , RIe1b1b48_3399, \9548 );
and \U$2767 ( \11848 , RIfc4b650_5880, \9550 );
and \U$2768 ( \11849 , RIfcda918_7509, \9552 );
and \U$2769 ( \11850 , RIfe98370_8076, \9554 );
and \U$2770 ( \11851 , RIfe99018_8085, \9556 );
and \U$2771 ( \11852 , RIe1a9e20_3310, \9558 );
and \U$2772 ( \11853 , RIe1a7120_3278, \9560 );
and \U$2773 ( \11854 , RIe1a4420_3246, \9562 );
and \U$2774 ( \11855 , RIe1a1720_3214, \9564 );
and \U$2775 ( \11856 , RIe18dc20_2990, \9566 );
and \U$2776 ( \11857 , RIe17a120_2766, \9568 );
and \U$2777 ( \11858 , RIe227a78_4741, \9570 );
and \U$2778 ( \11859 , RIe21c678_4613, \9572 );
and \U$2779 ( \11860 , RIe205e78_4357, \9574 );
and \U$2780 ( \11861 , RIe1ffed8_4289, \9576 );
and \U$2781 ( \11862 , RIe1f9290_4212, \9578 );
and \U$2782 ( \11863 , RIe1f1dd8_4129, \9580 );
and \U$2783 ( \11864 , RIe1d62e0_3814, \9582 );
and \U$2784 ( \11865 , RIe1bcde0_3526, \9584 );
and \U$2785 ( \11866 , RIe1afc58_3377, \9586 );
and \U$2786 ( \11867 , RIe172290_2676, \9588 );
or \U$2787 ( \11868 , \11804 , \11805 , \11806 , \11807 , \11808 , \11809 , \11810 , \11811 , \11812 , \11813 , \11814 , \11815 , \11816 , \11817 , \11818 , \11819 , \11820 , \11821 , \11822 , \11823 , \11824 , \11825 , \11826 , \11827 , \11828 , \11829 , \11830 , \11831 , \11832 , \11833 , \11834 , \11835 , \11836 , \11837 , \11838 , \11839 , \11840 , \11841 , \11842 , \11843 , \11844 , \11845 , \11846 , \11847 , \11848 , \11849 , \11850 , \11851 , \11852 , \11853 , \11854 , \11855 , \11856 , \11857 , \11858 , \11859 , \11860 , \11861 , \11862 , \11863 , \11864 , \11865 , \11866 , \11867 );
or \U$2788 ( \11869 , \11803 , \11868 );
_DC g40e4 ( \11870_nG40e4 , \11869 , \9597 );
buf \U$2789 ( \11871 , \11870_nG40e4 );
xor \U$2790 ( \11872 , \11738 , \11871 );
and \U$2791 ( \11873 , RIdec6620_721, \9059 );
and \U$2792 ( \11874 , RIdec3920_689, \9061 );
and \U$2793 ( \11875 , RIfc49328_5855, \9063 );
and \U$2794 ( \11876 , RIdec0c20_657, \9065 );
and \U$2795 ( \11877 , RIfc80eb8_6489, \9067 );
and \U$2796 ( \11878 , RIdebdf20_625, \9069 );
and \U$2797 ( \11879 , RIdebb220_593, \9071 );
and \U$2798 ( \11880 , RIdeb8520_561, \9073 );
and \U$2799 ( \11881 , RIfc80648_6483, \9075 );
and \U$2800 ( \11882 , RIdeb2b20_497, \9077 );
and \U$2801 ( \11883 , RIfc8b340_6606, \9079 );
and \U$2802 ( \11884 , RIdeafe20_465, \9081 );
and \U$2803 ( \11885 , RIfc491c0_5854, \9083 );
and \U$2804 ( \11886 , RIdeacec8_433, \9085 );
and \U$2805 ( \11887 , RIdea65c8_401, \9087 );
and \U$2806 ( \11888 , RIde9fcc8_369, \9089 );
and \U$2807 ( \11889 , RIfcd9c70_7500, \9091 );
and \U$2808 ( \11890 , RIfe98208_8075, \9093 );
and \U$2809 ( \11891 , RIfce4698_7621, \9095 );
and \U$2810 ( \11892 , RIfe980a0_8074, \9097 );
and \U$2811 ( \11893 , RIde93158_307, \9099 );
and \U$2812 ( \11894 , RIde8f648_289, \9101 );
and \U$2813 ( \11895 , RIde8b4a8_269, \9103 );
and \U$2814 ( \11896 , RIde87308_249, \9105 );
and \U$2815 ( \11897 , RIde82e20_228, \9107 );
and \U$2816 ( \11898 , RIfcbba18_7157, \9109 );
and \U$2817 ( \11899 , RIfc48d88_5851, \9111 );
and \U$2818 ( \11900 , RIfc99f80_6774, \9113 );
and \U$2819 ( \11901 , RIfc8b4a8_6607, \9115 );
and \U$2820 ( \11902 , RIe16c728_2611, \9117 );
and \U$2821 ( \11903 , RIe16a400_2586, \9119 );
and \U$2822 ( \11904 , RIe168c18_2569, \9121 );
and \U$2823 ( \11905 , RIe166620_2542, \9123 );
and \U$2824 ( \11906 , RIe163920_2510, \9125 );
and \U$2825 ( \11907 , RIee38068_5096, \9127 );
and \U$2826 ( \11908 , RIe160c20_2478, \9129 );
and \U$2827 ( \11909 , RIfc48248_5843, \9131 );
and \U$2828 ( \11910 , RIe15df20_2446, \9133 );
and \U$2829 ( \11911 , RIe158520_2382, \9135 );
and \U$2830 ( \11912 , RIe155820_2350, \9137 );
and \U$2831 ( \11913 , RIfcbbe50_7160, \9139 );
and \U$2832 ( \11914 , RIe152b20_2318, \9141 );
and \U$2833 ( \11915 , RIfc47e10_5840, \9143 );
and \U$2834 ( \11916 , RIe14fe20_2286, \9145 );
and \U$2835 ( \11917 , RIfca0e98_6853, \9147 );
and \U$2836 ( \11918 , RIe14d120_2254, \9149 );
and \U$2837 ( \11919 , RIe14a420_2222, \9151 );
and \U$2838 ( \11920 , RIe147720_2190, \9153 );
and \U$2839 ( \11921 , RIfc8be80_6614, \9155 );
and \U$2840 ( \11922 , RIfc7fb08_6475, \9157 );
and \U$2841 ( \11923 , RIfc480e0_5842, \9159 );
and \U$2842 ( \11924 , RIfc99878_6769, \9161 );
and \U$2843 ( \11925 , RIe141e88_2127, \9163 );
and \U$2844 ( \11926 , RIe13fb60_2102, \9165 );
and \U$2845 ( \11927 , RIdf3da68_2078, \9167 );
and \U$2846 ( \11928 , RIdf3b5d8_2052, \9169 );
and \U$2847 ( \11929 , RIfe97f38_8073, \9171 );
and \U$2848 ( \11930 , RIee30070_5005, \9173 );
and \U$2849 ( \11931 , RIee2eb58_4990, \9175 );
and \U$2850 ( \11932 , RIee2deb0_4981, \9177 );
and \U$2851 ( \11933 , RIdf36880_1997, \9179 );
and \U$2852 ( \11934 , RIdf34288_1970, \9181 );
and \U$2853 ( \11935 , RIdf320c8_1946, \9183 );
and \U$2854 ( \11936 , RIfe97dd0_8072, \9185 );
or \U$2855 ( \11937 , \11873 , \11874 , \11875 , \11876 , \11877 , \11878 , \11879 , \11880 , \11881 , \11882 , \11883 , \11884 , \11885 , \11886 , \11887 , \11888 , \11889 , \11890 , \11891 , \11892 , \11893 , \11894 , \11895 , \11896 , \11897 , \11898 , \11899 , \11900 , \11901 , \11902 , \11903 , \11904 , \11905 , \11906 , \11907 , \11908 , \11909 , \11910 , \11911 , \11912 , \11913 , \11914 , \11915 , \11916 , \11917 , \11918 , \11919 , \11920 , \11921 , \11922 , \11923 , \11924 , \11925 , \11926 , \11927 , \11928 , \11929 , \11930 , \11931 , \11932 , \11933 , \11934 , \11935 , \11936 );
and \U$2856 ( \11938 , RIfcc3740_7246, \9188 );
and \U$2857 ( \11939 , RIfc48ab8_5849, \9190 );
and \U$2858 ( \11940 , RIfce05e8_7575, \9192 );
and \U$2859 ( \11941 , RIfc80210_6480, \9194 );
and \U$2860 ( \11942 , RIdf2b048_1866, \9196 );
and \U$2861 ( \11943 , RIdf29158_1844, \9198 );
and \U$2862 ( \11944 , RIdf26f98_1820, \9200 );
and \U$2863 ( \11945 , RIdf254e0_1801, \9202 );
and \U$2864 ( \11946 , RIfc8bbb0_6612, \9204 );
and \U$2865 ( \11947 , RIfc48950_5848, \9206 );
and \U$2866 ( \11948 , RIdf235f0_1779, \9208 );
and \U$2867 ( \11949 , RIfc8bd18_6613, \9210 );
and \U$2868 ( \11950 , RIdf21f70_1763, \9212 );
and \U$2869 ( \11951 , RIdf208f0_1747, \9214 );
and \U$2870 ( \11952 , RIdf1b8c8_1690, \9216 );
and \U$2871 ( \11953 , RIdf1a3b0_1675, \9218 );
and \U$2872 ( \11954 , RIdf181f0_1651, \9220 );
and \U$2873 ( \11955 , RIdf154f0_1619, \9222 );
and \U$2874 ( \11956 , RIdf127f0_1587, \9224 );
and \U$2875 ( \11957 , RIdf0faf0_1555, \9226 );
and \U$2876 ( \11958 , RIdf0cdf0_1523, \9228 );
and \U$2877 ( \11959 , RIdf0a0f0_1491, \9230 );
and \U$2878 ( \11960 , RIdf073f0_1459, \9232 );
and \U$2879 ( \11961 , RIdf046f0_1427, \9234 );
and \U$2880 ( \11962 , RIdefecf0_1363, \9236 );
and \U$2881 ( \11963 , RIdefbff0_1331, \9238 );
and \U$2882 ( \11964 , RIdef92f0_1299, \9240 );
and \U$2883 ( \11965 , RIdef65f0_1267, \9242 );
and \U$2884 ( \11966 , RIdef38f0_1235, \9244 );
and \U$2885 ( \11967 , RIdef0bf0_1203, \9246 );
and \U$2886 ( \11968 , RIdeedef0_1171, \9248 );
and \U$2887 ( \11969 , RIdeeb1f0_1139, \9250 );
and \U$2888 ( \11970 , RIfcbc120_7162, \9252 );
and \U$2889 ( \11971 , RIfcd9838_7497, \9254 );
and \U$2890 ( \11972 , RIfc99710_6768, \9256 );
and \U$2891 ( \11973 , RIfca1168_6855, \9258 );
and \U$2892 ( \11974 , RIdee57f0_1075, \9260 );
and \U$2893 ( \11975 , RIdee3a68_1054, \9262 );
and \U$2894 ( \11976 , RIdee18a8_1030, \9264 );
and \U$2895 ( \11977 , RIdedf850_1007, \9266 );
and \U$2896 ( \11978 , RIfc549f8_5985, \9268 );
and \U$2897 ( \11979 , RIfcb5370_7084, \9270 );
and \U$2898 ( \11980 , RIfce43c8_7619, \9272 );
and \U$2899 ( \11981 , RIfce0480_7574, \9274 );
and \U$2900 ( \11982 , RIdeda6c0_949, \9276 );
and \U$2901 ( \11983 , RIded8230_923, \9278 );
and \U$2902 ( \11984 , RIded6070_899, \9280 );
and \U$2903 ( \11985 , RIded3d48_874, \9282 );
and \U$2904 ( \11986 , RIded1a20_849, \9284 );
and \U$2905 ( \11987 , RIdeced20_817, \9286 );
and \U$2906 ( \11988 , RIdecc020_785, \9288 );
and \U$2907 ( \11989 , RIdec9320_753, \9290 );
and \U$2908 ( \11990 , RIdeb5820_529, \9292 );
and \U$2909 ( \11991 , RIde993c8_337, \9294 );
and \U$2910 ( \11992 , RIe16f428_2643, \9296 );
and \U$2911 ( \11993 , RIe15b220_2414, \9298 );
and \U$2912 ( \11994 , RIe144a20_2158, \9300 );
and \U$2913 ( \11995 , RIdf39418_2028, \9302 );
and \U$2914 ( \11996 , RIdf2da78_1896, \9304 );
and \U$2915 ( \11997 , RIdf1e2f8_1720, \9306 );
and \U$2916 ( \11998 , RIdf019f0_1395, \9308 );
and \U$2917 ( \11999 , RIdee84f0_1107, \9310 );
and \U$2918 ( \12000 , RIdedd258_980, \9312 );
and \U$2919 ( \12001 , RIde7f310_210, \9314 );
or \U$2920 ( \12002 , \11938 , \11939 , \11940 , \11941 , \11942 , \11943 , \11944 , \11945 , \11946 , \11947 , \11948 , \11949 , \11950 , \11951 , \11952 , \11953 , \11954 , \11955 , \11956 , \11957 , \11958 , \11959 , \11960 , \11961 , \11962 , \11963 , \11964 , \11965 , \11966 , \11967 , \11968 , \11969 , \11970 , \11971 , \11972 , \11973 , \11974 , \11975 , \11976 , \11977 , \11978 , \11979 , \11980 , \11981 , \11982 , \11983 , \11984 , \11985 , \11986 , \11987 , \11988 , \11989 , \11990 , \11991 , \11992 , \11993 , \11994 , \11995 , \11996 , \11997 , \11998 , \11999 , \12000 , \12001 );
or \U$2921 ( \12003 , \11937 , \12002 );
_DC g303c ( \12004_nG303c , \12003 , \9323 );
buf \U$2922 ( \12005 , \12004_nG303c );
and \U$2923 ( \12006 , RIe19e8b8_3181, \9333 );
and \U$2924 ( \12007 , RIe19bbb8_3149, \9335 );
and \U$2925 ( \12008 , RIfe976c8_8067, \9337 );
and \U$2926 ( \12009 , RIe198eb8_3117, \9339 );
and \U$2927 ( \12010 , RIf144c80_5242, \9341 );
and \U$2928 ( \12011 , RIe1961b8_3085, \9343 );
and \U$2929 ( \12012 , RIe1934b8_3053, \9345 );
and \U$2930 ( \12013 , RIe1907b8_3021, \9347 );
and \U$2931 ( \12014 , RIe18adb8_2957, \9349 );
and \U$2932 ( \12015 , RIe1880b8_2925, \9351 );
and \U$2933 ( \12016 , RIfe97560_8066, \9353 );
and \U$2934 ( \12017 , RIe1853b8_2893, \9355 );
and \U$2935 ( \12018 , RIfcc3fb0_7252, \9357 );
and \U$2936 ( \12019 , RIe1826b8_2861, \9359 );
and \U$2937 ( \12020 , RIe17f9b8_2829, \9361 );
and \U$2938 ( \12021 , RIe17ccb8_2797, \9363 );
and \U$2939 ( \12022 , RIfcd3730_7428, \9365 );
and \U$2940 ( \12023 , RIf1412d8_5201, \9367 );
and \U$2941 ( \12024 , RIfcc4118_7253, \9369 );
and \U$2942 ( \12025 , RIfe97830_8068, \9371 );
and \U$2943 ( \12026 , RIfc4a6d8_5869, \9373 );
and \U$2944 ( \12027 , RIf13f6b8_5181, \9375 );
and \U$2945 ( \12028 , RIfc9f980_6838, \9377 );
and \U$2946 ( \12029 , RIfc9fae8_6839, \9379 );
and \U$2947 ( \12030 , RIfcc3e48_7251, \9381 );
and \U$2948 ( \12031 , RIfc89e28_6591, \9383 );
and \U$2949 ( \12032 , RIfc89cc0_6590, \9385 );
and \U$2950 ( \12033 , RIe174720_2702, \9387 );
and \U$2951 ( \12034 , RIfc4a408_5867, \9389 );
and \U$2952 ( \12035 , RIfce27a8_7599, \9391 );
and \U$2953 ( \12036 , RIfc530a8_5967, \9393 );
and \U$2954 ( \12037 , RIfcd5d28_7455, \9395 );
and \U$2955 ( \12038 , RIf16cf28_5699, \9397 );
and \U$2956 ( \12039 , RIe224c10_4708, \9399 );
and \U$2957 ( \12040 , RIfc53210_5968, \9401 );
and \U$2958 ( \12041 , RIe221f10_4676, \9403 );
and \U$2959 ( \12042 , RIf16b1a0_5678, \9405 );
and \U$2960 ( \12043 , RIe21f210_4644, \9407 );
and \U$2961 ( \12044 , RIe219810_4580, \9409 );
and \U$2962 ( \12045 , RIe216b10_4548, \9411 );
and \U$2963 ( \12046 , RIfc401d8_5755, \9413 );
and \U$2964 ( \12047 , RIe213e10_4516, \9415 );
and \U$2965 ( \12048 , RIf1699b8_5661, \9417 );
and \U$2966 ( \12049 , RIe211110_4484, \9419 );
and \U$2967 ( \12050 , RIfc81cc8_6499, \9421 );
and \U$2968 ( \12051 , RIe20e410_4452, \9423 );
and \U$2969 ( \12052 , RIe20b710_4420, \9425 );
and \U$2970 ( \12053 , RIe208a10_4388, \9427 );
and \U$2971 ( \12054 , RIfc8a0f8_6593, \9429 );
and \U$2972 ( \12055 , RIfcb6720_7098, \9431 );
and \U$2973 ( \12056 , RIe203448_4327, \9433 );
and \U$2974 ( \12057 , RIe201828_4307, \9435 );
and \U$2975 ( \12058 , RIfc53378_5969, \9437 );
and \U$2976 ( \12059 , RIfc8a3c8_6595, \9439 );
and \U$2977 ( \12060 , RIfcb65b8_7097, \9441 );
and \U$2978 ( \12061 , RIfc49fd0_5864, \9443 );
and \U$2979 ( \12062 , RIf160bb0_5560, \9445 );
and \U$2980 ( \12063 , RIf15ecc0_5538, \9447 );
and \U$2981 ( \12064 , RIe1fd4a8_4259, \9449 );
and \U$2982 ( \12065 , RIfe97b00_8070, \9451 );
and \U$2983 ( \12066 , RIfc8a530_6596, \9453 );
and \U$2984 ( \12067 , RIfe97c68_8071, \9455 );
and \U$2985 ( \12068 , RIfc8a800_6598, \9457 );
and \U$2986 ( \12069 , RIfc8a698_6597, \9459 );
or \U$2987 ( \12070 , \12006 , \12007 , \12008 , \12009 , \12010 , \12011 , \12012 , \12013 , \12014 , \12015 , \12016 , \12017 , \12018 , \12019 , \12020 , \12021 , \12022 , \12023 , \12024 , \12025 , \12026 , \12027 , \12028 , \12029 , \12030 , \12031 , \12032 , \12033 , \12034 , \12035 , \12036 , \12037 , \12038 , \12039 , \12040 , \12041 , \12042 , \12043 , \12044 , \12045 , \12046 , \12047 , \12048 , \12049 , \12050 , \12051 , \12052 , \12053 , \12054 , \12055 , \12056 , \12057 , \12058 , \12059 , \12060 , \12061 , \12062 , \12063 , \12064 , \12065 , \12066 , \12067 , \12068 , \12069 );
and \U$2988 ( \12071 , RIfc9a7f0_6780, \9462 );
and \U$2989 ( \12072 , RIfc81890_6496, \9464 );
and \U$2990 ( \12073 , RIfcd5e90_7456, \9466 );
and \U$2991 ( \12074 , RIe1fb180_4234, \9468 );
and \U$2992 ( \12075 , RIfc49e68_5863, \9470 );
and \U$2993 ( \12076 , RIfc81728_6495, \9472 );
and \U$2994 ( \12077 , RIfcbb1a8_7151, \9474 );
and \U$2995 ( \12078 , RIe1f66f8_4181, \9476 );
and \U$2996 ( \12079 , RIfcd3460_7426, \9478 );
and \U$2997 ( \12080 , RIfcb62e8_7095, \9480 );
and \U$2998 ( \12081 , RIfc9a520_6778, \9482 );
and \U$2999 ( \12082 , RIe1f4268_4155, \9484 );
and \U$3000 ( \12083 , RIfc49d00_5862, \9486 );
and \U$3001 ( \12084 , RIfcd9dd8_7501, \9488 );
and \U$3002 ( \12085 , RIfcbb310_7152, \9490 );
and \U$3003 ( \12086 , RIe1ef0d8_4097, \9492 );
and \U$3004 ( \12087 , RIe1ec978_4069, \9494 );
and \U$3005 ( \12088 , RIe1e9c78_4037, \9496 );
and \U$3006 ( \12089 , RIe1e6f78_4005, \9498 );
and \U$3007 ( \12090 , RIe1e4278_3973, \9500 );
and \U$3008 ( \12091 , RIe1e1578_3941, \9502 );
and \U$3009 ( \12092 , RIe1de878_3909, \9504 );
and \U$3010 ( \12093 , RIe1dbb78_3877, \9506 );
and \U$3011 ( \12094 , RIe1d8e78_3845, \9508 );
and \U$3012 ( \12095 , RIe1d3478_3781, \9510 );
and \U$3013 ( \12096 , RIe1d0778_3749, \9512 );
and \U$3014 ( \12097 , RIe1cda78_3717, \9514 );
and \U$3015 ( \12098 , RIe1cad78_3685, \9516 );
and \U$3016 ( \12099 , RIe1c8078_3653, \9518 );
and \U$3017 ( \12100 , RIe1c5378_3621, \9520 );
and \U$3018 ( \12101 , RIe1c2678_3589, \9522 );
and \U$3019 ( \12102 , RIe1bf978_3557, \9524 );
and \U$3020 ( \12103 , RIfc49a30_5860, \9526 );
and \U$3021 ( \12104 , RIfcb6018_7093, \9528 );
and \U$3022 ( \12105 , RIe1ba3b0_3496, \9530 );
and \U$3023 ( \12106 , RIe1b81f0_3472, \9532 );
and \U$3024 ( \12107 , RIfce0a20_7578, \9534 );
and \U$3025 ( \12108 , RIfcbb5e0_7154, \9536 );
and \U$3026 ( \12109 , RIe1b6030_3448, \9538 );
and \U$3027 ( \12110 , RIfe97998_8069, \9540 );
and \U$3028 ( \12111 , RIfce5610_7632, \9542 );
and \U$3029 ( \12112 , RIfcc3a10_7248, \9544 );
and \U$3030 ( \12113 , RIe1b3330_3416, \9546 );
and \U$3031 ( \12114 , RIe1b19e0_3398, \9548 );
and \U$3032 ( \12115 , RIfc495f8_5857, \9550 );
and \U$3033 ( \12116 , RIfc81188_6491, \9552 );
and \U$3034 ( \12117 , RIe1ad228_3347, \9554 );
and \U$3035 ( \12118 , RIe1aba40_3330, \9556 );
and \U$3036 ( \12119 , RIe1a9cb8_3309, \9558 );
and \U$3037 ( \12120 , RIe1a6fb8_3277, \9560 );
and \U$3038 ( \12121 , RIe1a42b8_3245, \9562 );
and \U$3039 ( \12122 , RIe1a15b8_3213, \9564 );
and \U$3040 ( \12123 , RIe18dab8_2989, \9566 );
and \U$3041 ( \12124 , RIe179fb8_2765, \9568 );
and \U$3042 ( \12125 , RIe227910_4740, \9570 );
and \U$3043 ( \12126 , RIe21c510_4612, \9572 );
and \U$3044 ( \12127 , RIe205d10_4356, \9574 );
and \U$3045 ( \12128 , RIe1ffd70_4288, \9576 );
and \U$3046 ( \12129 , RIe1f9128_4211, \9578 );
and \U$3047 ( \12130 , RIe1f1c70_4128, \9580 );
and \U$3048 ( \12131 , RIe1d6178_3813, \9582 );
and \U$3049 ( \12132 , RIe1bcc78_3525, \9584 );
and \U$3050 ( \12133 , RIe1afaf0_3376, \9586 );
and \U$3051 ( \12134 , RIe172128_2675, \9588 );
or \U$3052 ( \12135 , \12071 , \12072 , \12073 , \12074 , \12075 , \12076 , \12077 , \12078 , \12079 , \12080 , \12081 , \12082 , \12083 , \12084 , \12085 , \12086 , \12087 , \12088 , \12089 , \12090 , \12091 , \12092 , \12093 , \12094 , \12095 , \12096 , \12097 , \12098 , \12099 , \12100 , \12101 , \12102 , \12103 , \12104 , \12105 , \12106 , \12107 , \12108 , \12109 , \12110 , \12111 , \12112 , \12113 , \12114 , \12115 , \12116 , \12117 , \12118 , \12119 , \12120 , \12121 , \12122 , \12123 , \12124 , \12125 , \12126 , \12127 , \12128 , \12129 , \12130 , \12131 , \12132 , \12133 , \12134 );
or \U$3053 ( \12136 , \12070 , \12135 );
_DC g4169 ( \12137_nG4169 , \12136 , \9597 );
buf \U$3054 ( \12138 , \12137_nG4169 );
and \U$3055 ( \12139 , \12005 , \12138 );
and \U$3056 ( \12140 , \9325 , \9599 );
and \U$3057 ( \12141 , \9599 , \10407 );
and \U$3058 ( \12142 , \9325 , \10407 );
or \U$3059 ( \12143 , \12140 , \12141 , \12142 );
and \U$3060 ( \12144 , \12138 , \12143 );
and \U$3061 ( \12145 , \12005 , \12143 );
or \U$3062 ( \12146 , \12139 , \12144 , \12145 );
xor \U$3063 ( \12147 , \11872 , \12146 );
buf g4448 ( \12148_nG4448 , \12147 );
xor \U$3064 ( \12149 , \12005 , \12138 );
xor \U$3065 ( \12150 , \12149 , \12143 );
buf g444b ( \12151_nG444b , \12150 );
nand \U$3066 ( \12152 , \12151_nG444b , \10409_nG444e );
and \U$3067 ( \12153 , \12148_nG4448 , \12152 );
xor \U$3068 ( \12154 , \12151_nG444b , \10409_nG444e );
not \U$3069 ( \12155 , \12154 );
xor \U$3070 ( \12156 , \12148_nG4448 , \12151_nG444b );
and \U$3071 ( \12157 , \12155 , \12156 );
and \U$3073 ( \12158 , \12154 , \10694_nG9c0e );
or \U$3074 ( \12159 , 1'b0 , \12158 );
xor \U$3075 ( \12160 , \12153 , \12159 );
xor \U$3076 ( \12161 , \12153 , \12160 );
buf \U$3077 ( \12162 , \12161 );
buf \U$3078 ( \12163 , \12162 );
and \U$3079 ( \12164 , \11605 , \12163 );
and \U$3080 ( \12165 , \11295 , \11301 );
buf \U$3081 ( \12166 , \12165 );
and \U$3082 ( \12167 , \10421 , \10995_nG9c0b );
and \U$3083 ( \12168 , \10418 , \11283_nG9c08 );
or \U$3084 ( \12169 , \12167 , \12168 );
xor \U$3085 ( \12170 , \10417 , \12169 );
buf \U$3086 ( \12171 , \12170 );
buf \U$3088 ( \12172 , \12171 );
xor \U$3089 ( \12173 , \12166 , \12172 );
buf \U$3090 ( \12174 , \12173 );
and \U$3091 ( \12175 , \11292 , \11303 );
and \U$3092 ( \12176 , \11292 , \11603 );
and \U$3093 ( \12177 , \11303 , \11603 );
or \U$3094 ( \12178 , \12175 , \12176 , \12177 );
buf \U$3095 ( \12179 , \12178 );
xor \U$3096 ( \12180 , \12174 , \12179 );
and \U$3097 ( \12181 , \10707 , \11598_nG9c05 );
and \U$3098 ( \12182 , \11586 , \10983 );
and \U$3099 ( \12183 , RIdec6620_721, \9333 );
and \U$3100 ( \12184 , RIdec3920_689, \9335 );
and \U$3101 ( \12185 , RIfc49328_5855, \9337 );
and \U$3102 ( \12186 , RIdec0c20_657, \9339 );
and \U$3103 ( \12187 , RIfc80eb8_6489, \9341 );
and \U$3104 ( \12188 , RIdebdf20_625, \9343 );
and \U$3105 ( \12189 , RIdebb220_593, \9345 );
and \U$3106 ( \12190 , RIdeb8520_561, \9347 );
and \U$3107 ( \12191 , RIfc80648_6483, \9349 );
and \U$3108 ( \12192 , RIdeb2b20_497, \9351 );
and \U$3109 ( \12193 , RIfc8b340_6606, \9353 );
and \U$3110 ( \12194 , RIdeafe20_465, \9355 );
and \U$3111 ( \12195 , RIfc491c0_5854, \9357 );
and \U$3112 ( \12196 , RIdeacec8_433, \9359 );
and \U$3113 ( \12197 , RIdea65c8_401, \9361 );
and \U$3114 ( \12198 , RIde9fcc8_369, \9363 );
and \U$3115 ( \12199 , RIfcd9c70_7500, \9365 );
and \U$3116 ( \12200 , RIfe98208_8075, \9367 );
and \U$3117 ( \12201 , RIfce4698_7621, \9369 );
and \U$3118 ( \12202 , RIfe980a0_8074, \9371 );
and \U$3119 ( \12203 , RIde93158_307, \9373 );
and \U$3120 ( \12204 , RIde8f648_289, \9375 );
and \U$3121 ( \12205 , RIde8b4a8_269, \9377 );
and \U$3122 ( \12206 , RIde87308_249, \9379 );
and \U$3123 ( \12207 , RIde82e20_228, \9381 );
and \U$3124 ( \12208 , RIfcbba18_7157, \9383 );
and \U$3125 ( \12209 , RIfc48d88_5851, \9385 );
and \U$3126 ( \12210 , RIfc99f80_6774, \9387 );
and \U$3127 ( \12211 , RIfc8b4a8_6607, \9389 );
and \U$3128 ( \12212 , RIe16c728_2611, \9391 );
and \U$3129 ( \12213 , RIe16a400_2586, \9393 );
and \U$3130 ( \12214 , RIe168c18_2569, \9395 );
and \U$3131 ( \12215 , RIe166620_2542, \9397 );
and \U$3132 ( \12216 , RIe163920_2510, \9399 );
and \U$3133 ( \12217 , RIee38068_5096, \9401 );
and \U$3134 ( \12218 , RIe160c20_2478, \9403 );
and \U$3135 ( \12219 , RIfc48248_5843, \9405 );
and \U$3136 ( \12220 , RIe15df20_2446, \9407 );
and \U$3137 ( \12221 , RIe158520_2382, \9409 );
and \U$3138 ( \12222 , RIe155820_2350, \9411 );
and \U$3139 ( \12223 , RIfcbbe50_7160, \9413 );
and \U$3140 ( \12224 , RIe152b20_2318, \9415 );
and \U$3141 ( \12225 , RIfc47e10_5840, \9417 );
and \U$3142 ( \12226 , RIe14fe20_2286, \9419 );
and \U$3143 ( \12227 , RIfca0e98_6853, \9421 );
and \U$3144 ( \12228 , RIe14d120_2254, \9423 );
and \U$3145 ( \12229 , RIe14a420_2222, \9425 );
and \U$3146 ( \12230 , RIe147720_2190, \9427 );
and \U$3147 ( \12231 , RIfc8be80_6614, \9429 );
and \U$3148 ( \12232 , RIfc7fb08_6475, \9431 );
and \U$3149 ( \12233 , RIfc480e0_5842, \9433 );
and \U$3150 ( \12234 , RIfc99878_6769, \9435 );
and \U$3151 ( \12235 , RIe141e88_2127, \9437 );
and \U$3152 ( \12236 , RIe13fb60_2102, \9439 );
and \U$3153 ( \12237 , RIdf3da68_2078, \9441 );
and \U$3154 ( \12238 , RIdf3b5d8_2052, \9443 );
and \U$3155 ( \12239 , RIfe97f38_8073, \9445 );
and \U$3156 ( \12240 , RIee30070_5005, \9447 );
and \U$3157 ( \12241 , RIee2eb58_4990, \9449 );
and \U$3158 ( \12242 , RIee2deb0_4981, \9451 );
and \U$3159 ( \12243 , RIdf36880_1997, \9453 );
and \U$3160 ( \12244 , RIdf34288_1970, \9455 );
and \U$3161 ( \12245 , RIdf320c8_1946, \9457 );
and \U$3162 ( \12246 , RIfe97dd0_8072, \9459 );
or \U$3163 ( \12247 , \12183 , \12184 , \12185 , \12186 , \12187 , \12188 , \12189 , \12190 , \12191 , \12192 , \12193 , \12194 , \12195 , \12196 , \12197 , \12198 , \12199 , \12200 , \12201 , \12202 , \12203 , \12204 , \12205 , \12206 , \12207 , \12208 , \12209 , \12210 , \12211 , \12212 , \12213 , \12214 , \12215 , \12216 , \12217 , \12218 , \12219 , \12220 , \12221 , \12222 , \12223 , \12224 , \12225 , \12226 , \12227 , \12228 , \12229 , \12230 , \12231 , \12232 , \12233 , \12234 , \12235 , \12236 , \12237 , \12238 , \12239 , \12240 , \12241 , \12242 , \12243 , \12244 , \12245 , \12246 );
and \U$3164 ( \12248 , RIfcc3740_7246, \9462 );
and \U$3165 ( \12249 , RIfc48ab8_5849, \9464 );
and \U$3166 ( \12250 , RIfce05e8_7575, \9466 );
and \U$3167 ( \12251 , RIfc80210_6480, \9468 );
and \U$3168 ( \12252 , RIdf2b048_1866, \9470 );
and \U$3169 ( \12253 , RIdf29158_1844, \9472 );
and \U$3170 ( \12254 , RIdf26f98_1820, \9474 );
and \U$3171 ( \12255 , RIdf254e0_1801, \9476 );
and \U$3172 ( \12256 , RIfc8bbb0_6612, \9478 );
and \U$3173 ( \12257 , RIfc48950_5848, \9480 );
and \U$3174 ( \12258 , RIdf235f0_1779, \9482 );
and \U$3175 ( \12259 , RIfc8bd18_6613, \9484 );
and \U$3176 ( \12260 , RIdf21f70_1763, \9486 );
and \U$3177 ( \12261 , RIdf208f0_1747, \9488 );
and \U$3178 ( \12262 , RIdf1b8c8_1690, \9490 );
and \U$3179 ( \12263 , RIdf1a3b0_1675, \9492 );
and \U$3180 ( \12264 , RIdf181f0_1651, \9494 );
and \U$3181 ( \12265 , RIdf154f0_1619, \9496 );
and \U$3182 ( \12266 , RIdf127f0_1587, \9498 );
and \U$3183 ( \12267 , RIdf0faf0_1555, \9500 );
and \U$3184 ( \12268 , RIdf0cdf0_1523, \9502 );
and \U$3185 ( \12269 , RIdf0a0f0_1491, \9504 );
and \U$3186 ( \12270 , RIdf073f0_1459, \9506 );
and \U$3187 ( \12271 , RIdf046f0_1427, \9508 );
and \U$3188 ( \12272 , RIdefecf0_1363, \9510 );
and \U$3189 ( \12273 , RIdefbff0_1331, \9512 );
and \U$3190 ( \12274 , RIdef92f0_1299, \9514 );
and \U$3191 ( \12275 , RIdef65f0_1267, \9516 );
and \U$3192 ( \12276 , RIdef38f0_1235, \9518 );
and \U$3193 ( \12277 , RIdef0bf0_1203, \9520 );
and \U$3194 ( \12278 , RIdeedef0_1171, \9522 );
and \U$3195 ( \12279 , RIdeeb1f0_1139, \9524 );
and \U$3196 ( \12280 , RIfcbc120_7162, \9526 );
and \U$3197 ( \12281 , RIfcd9838_7497, \9528 );
and \U$3198 ( \12282 , RIfc99710_6768, \9530 );
and \U$3199 ( \12283 , RIfca1168_6855, \9532 );
and \U$3200 ( \12284 , RIdee57f0_1075, \9534 );
and \U$3201 ( \12285 , RIdee3a68_1054, \9536 );
and \U$3202 ( \12286 , RIdee18a8_1030, \9538 );
and \U$3203 ( \12287 , RIdedf850_1007, \9540 );
and \U$3204 ( \12288 , RIfc549f8_5985, \9542 );
and \U$3205 ( \12289 , RIfcb5370_7084, \9544 );
and \U$3206 ( \12290 , RIfce43c8_7619, \9546 );
and \U$3207 ( \12291 , RIfce0480_7574, \9548 );
and \U$3208 ( \12292 , RIdeda6c0_949, \9550 );
and \U$3209 ( \12293 , RIded8230_923, \9552 );
and \U$3210 ( \12294 , RIded6070_899, \9554 );
and \U$3211 ( \12295 , RIded3d48_874, \9556 );
and \U$3212 ( \12296 , RIded1a20_849, \9558 );
and \U$3213 ( \12297 , RIdeced20_817, \9560 );
and \U$3214 ( \12298 , RIdecc020_785, \9562 );
and \U$3215 ( \12299 , RIdec9320_753, \9564 );
and \U$3216 ( \12300 , RIdeb5820_529, \9566 );
and \U$3217 ( \12301 , RIde993c8_337, \9568 );
and \U$3218 ( \12302 , RIe16f428_2643, \9570 );
and \U$3219 ( \12303 , RIe15b220_2414, \9572 );
and \U$3220 ( \12304 , RIe144a20_2158, \9574 );
and \U$3221 ( \12305 , RIdf39418_2028, \9576 );
and \U$3222 ( \12306 , RIdf2da78_1896, \9578 );
and \U$3223 ( \12307 , RIdf1e2f8_1720, \9580 );
and \U$3224 ( \12308 , RIdf019f0_1395, \9582 );
and \U$3225 ( \12309 , RIdee84f0_1107, \9584 );
and \U$3226 ( \12310 , RIdedd258_980, \9586 );
and \U$3227 ( \12311 , RIde7f310_210, \9588 );
or \U$3228 ( \12312 , \12248 , \12249 , \12250 , \12251 , \12252 , \12253 , \12254 , \12255 , \12256 , \12257 , \12258 , \12259 , \12260 , \12261 , \12262 , \12263 , \12264 , \12265 , \12266 , \12267 , \12268 , \12269 , \12270 , \12271 , \12272 , \12273 , \12274 , \12275 , \12276 , \12277 , \12278 , \12279 , \12280 , \12281 , \12282 , \12283 , \12284 , \12285 , \12286 , \12287 , \12288 , \12289 , \12290 , \12291 , \12292 , \12293 , \12294 , \12295 , \12296 , \12297 , \12298 , \12299 , \12300 , \12301 , \12302 , \12303 , \12304 , \12305 , \12306 , \12307 , \12308 , \12309 , \12310 , \12311 );
or \U$3229 ( \12313 , \12247 , \12312 );
_DC g6583 ( \12314_nG6583 , \12313 , \9597 );
and \U$3230 ( \12315 , RIe19e8b8_3181, \9059 );
and \U$3231 ( \12316 , RIe19bbb8_3149, \9061 );
and \U$3232 ( \12317 , RIfe976c8_8067, \9063 );
and \U$3233 ( \12318 , RIe198eb8_3117, \9065 );
and \U$3234 ( \12319 , RIf144c80_5242, \9067 );
and \U$3235 ( \12320 , RIe1961b8_3085, \9069 );
and \U$3236 ( \12321 , RIe1934b8_3053, \9071 );
and \U$3237 ( \12322 , RIe1907b8_3021, \9073 );
and \U$3238 ( \12323 , RIe18adb8_2957, \9075 );
and \U$3239 ( \12324 , RIe1880b8_2925, \9077 );
and \U$3240 ( \12325 , RIfe97560_8066, \9079 );
and \U$3241 ( \12326 , RIe1853b8_2893, \9081 );
and \U$3242 ( \12327 , RIfcc3fb0_7252, \9083 );
and \U$3243 ( \12328 , RIe1826b8_2861, \9085 );
and \U$3244 ( \12329 , RIe17f9b8_2829, \9087 );
and \U$3245 ( \12330 , RIe17ccb8_2797, \9089 );
and \U$3246 ( \12331 , RIfcd3730_7428, \9091 );
and \U$3247 ( \12332 , RIf1412d8_5201, \9093 );
and \U$3248 ( \12333 , RIfcc4118_7253, \9095 );
and \U$3249 ( \12334 , RIfe97830_8068, \9097 );
and \U$3250 ( \12335 , RIfc4a6d8_5869, \9099 );
and \U$3251 ( \12336 , RIf13f6b8_5181, \9101 );
and \U$3252 ( \12337 , RIfc9f980_6838, \9103 );
and \U$3253 ( \12338 , RIfc9fae8_6839, \9105 );
and \U$3254 ( \12339 , RIfcc3e48_7251, \9107 );
and \U$3255 ( \12340 , RIfc89e28_6591, \9109 );
and \U$3256 ( \12341 , RIfc89cc0_6590, \9111 );
and \U$3257 ( \12342 , RIe174720_2702, \9113 );
and \U$3258 ( \12343 , RIfc4a408_5867, \9115 );
and \U$3259 ( \12344 , RIfce27a8_7599, \9117 );
and \U$3260 ( \12345 , RIfc530a8_5967, \9119 );
and \U$3261 ( \12346 , RIfcd5d28_7455, \9121 );
and \U$3262 ( \12347 , RIf16cf28_5699, \9123 );
and \U$3263 ( \12348 , RIe224c10_4708, \9125 );
and \U$3264 ( \12349 , RIfc53210_5968, \9127 );
and \U$3265 ( \12350 , RIe221f10_4676, \9129 );
and \U$3266 ( \12351 , RIf16b1a0_5678, \9131 );
and \U$3267 ( \12352 , RIe21f210_4644, \9133 );
and \U$3268 ( \12353 , RIe219810_4580, \9135 );
and \U$3269 ( \12354 , RIe216b10_4548, \9137 );
and \U$3270 ( \12355 , RIfc401d8_5755, \9139 );
and \U$3271 ( \12356 , RIe213e10_4516, \9141 );
and \U$3272 ( \12357 , RIf1699b8_5661, \9143 );
and \U$3273 ( \12358 , RIe211110_4484, \9145 );
and \U$3274 ( \12359 , RIfc81cc8_6499, \9147 );
and \U$3275 ( \12360 , RIe20e410_4452, \9149 );
and \U$3276 ( \12361 , RIe20b710_4420, \9151 );
and \U$3277 ( \12362 , RIe208a10_4388, \9153 );
and \U$3278 ( \12363 , RIfc8a0f8_6593, \9155 );
and \U$3279 ( \12364 , RIfcb6720_7098, \9157 );
and \U$3280 ( \12365 , RIe203448_4327, \9159 );
and \U$3281 ( \12366 , RIe201828_4307, \9161 );
and \U$3282 ( \12367 , RIfc53378_5969, \9163 );
and \U$3283 ( \12368 , RIfc8a3c8_6595, \9165 );
and \U$3284 ( \12369 , RIfcb65b8_7097, \9167 );
and \U$3285 ( \12370 , RIfc49fd0_5864, \9169 );
and \U$3286 ( \12371 , RIf160bb0_5560, \9171 );
and \U$3287 ( \12372 , RIf15ecc0_5538, \9173 );
and \U$3288 ( \12373 , RIe1fd4a8_4259, \9175 );
and \U$3289 ( \12374 , RIfe97b00_8070, \9177 );
and \U$3290 ( \12375 , RIfc8a530_6596, \9179 );
and \U$3291 ( \12376 , RIfe97c68_8071, \9181 );
and \U$3292 ( \12377 , RIfc8a800_6598, \9183 );
and \U$3293 ( \12378 , RIfc8a698_6597, \9185 );
or \U$3294 ( \12379 , \12315 , \12316 , \12317 , \12318 , \12319 , \12320 , \12321 , \12322 , \12323 , \12324 , \12325 , \12326 , \12327 , \12328 , \12329 , \12330 , \12331 , \12332 , \12333 , \12334 , \12335 , \12336 , \12337 , \12338 , \12339 , \12340 , \12341 , \12342 , \12343 , \12344 , \12345 , \12346 , \12347 , \12348 , \12349 , \12350 , \12351 , \12352 , \12353 , \12354 , \12355 , \12356 , \12357 , \12358 , \12359 , \12360 , \12361 , \12362 , \12363 , \12364 , \12365 , \12366 , \12367 , \12368 , \12369 , \12370 , \12371 , \12372 , \12373 , \12374 , \12375 , \12376 , \12377 , \12378 );
and \U$3295 ( \12380 , RIfc9a7f0_6780, \9188 );
and \U$3296 ( \12381 , RIfc81890_6496, \9190 );
and \U$3297 ( \12382 , RIfcd5e90_7456, \9192 );
and \U$3298 ( \12383 , RIe1fb180_4234, \9194 );
and \U$3299 ( \12384 , RIfc49e68_5863, \9196 );
and \U$3300 ( \12385 , RIfc81728_6495, \9198 );
and \U$3301 ( \12386 , RIfcbb1a8_7151, \9200 );
and \U$3302 ( \12387 , RIe1f66f8_4181, \9202 );
and \U$3303 ( \12388 , RIfcd3460_7426, \9204 );
and \U$3304 ( \12389 , RIfcb62e8_7095, \9206 );
and \U$3305 ( \12390 , RIfc9a520_6778, \9208 );
and \U$3306 ( \12391 , RIe1f4268_4155, \9210 );
and \U$3307 ( \12392 , RIfc49d00_5862, \9212 );
and \U$3308 ( \12393 , RIfcd9dd8_7501, \9214 );
and \U$3309 ( \12394 , RIfcbb310_7152, \9216 );
and \U$3310 ( \12395 , RIe1ef0d8_4097, \9218 );
and \U$3311 ( \12396 , RIe1ec978_4069, \9220 );
and \U$3312 ( \12397 , RIe1e9c78_4037, \9222 );
and \U$3313 ( \12398 , RIe1e6f78_4005, \9224 );
and \U$3314 ( \12399 , RIe1e4278_3973, \9226 );
and \U$3315 ( \12400 , RIe1e1578_3941, \9228 );
and \U$3316 ( \12401 , RIe1de878_3909, \9230 );
and \U$3317 ( \12402 , RIe1dbb78_3877, \9232 );
and \U$3318 ( \12403 , RIe1d8e78_3845, \9234 );
and \U$3319 ( \12404 , RIe1d3478_3781, \9236 );
and \U$3320 ( \12405 , RIe1d0778_3749, \9238 );
and \U$3321 ( \12406 , RIe1cda78_3717, \9240 );
and \U$3322 ( \12407 , RIe1cad78_3685, \9242 );
and \U$3323 ( \12408 , RIe1c8078_3653, \9244 );
and \U$3324 ( \12409 , RIe1c5378_3621, \9246 );
and \U$3325 ( \12410 , RIe1c2678_3589, \9248 );
and \U$3326 ( \12411 , RIe1bf978_3557, \9250 );
and \U$3327 ( \12412 , RIfc49a30_5860, \9252 );
and \U$3328 ( \12413 , RIfcb6018_7093, \9254 );
and \U$3329 ( \12414 , RIe1ba3b0_3496, \9256 );
and \U$3330 ( \12415 , RIe1b81f0_3472, \9258 );
and \U$3331 ( \12416 , RIfce0a20_7578, \9260 );
and \U$3332 ( \12417 , RIfcbb5e0_7154, \9262 );
and \U$3333 ( \12418 , RIe1b6030_3448, \9264 );
and \U$3334 ( \12419 , RIfe97998_8069, \9266 );
and \U$3335 ( \12420 , RIfce5610_7632, \9268 );
and \U$3336 ( \12421 , RIfcc3a10_7248, \9270 );
and \U$3337 ( \12422 , RIe1b3330_3416, \9272 );
and \U$3338 ( \12423 , RIe1b19e0_3398, \9274 );
and \U$3339 ( \12424 , RIfc495f8_5857, \9276 );
and \U$3340 ( \12425 , RIfc81188_6491, \9278 );
and \U$3341 ( \12426 , RIe1ad228_3347, \9280 );
and \U$3342 ( \12427 , RIe1aba40_3330, \9282 );
and \U$3343 ( \12428 , RIe1a9cb8_3309, \9284 );
and \U$3344 ( \12429 , RIe1a6fb8_3277, \9286 );
and \U$3345 ( \12430 , RIe1a42b8_3245, \9288 );
and \U$3346 ( \12431 , RIe1a15b8_3213, \9290 );
and \U$3347 ( \12432 , RIe18dab8_2989, \9292 );
and \U$3348 ( \12433 , RIe179fb8_2765, \9294 );
and \U$3349 ( \12434 , RIe227910_4740, \9296 );
and \U$3350 ( \12435 , RIe21c510_4612, \9298 );
and \U$3351 ( \12436 , RIe205d10_4356, \9300 );
and \U$3352 ( \12437 , RIe1ffd70_4288, \9302 );
and \U$3353 ( \12438 , RIe1f9128_4211, \9304 );
and \U$3354 ( \12439 , RIe1f1c70_4128, \9306 );
and \U$3355 ( \12440 , RIe1d6178_3813, \9308 );
and \U$3356 ( \12441 , RIe1bcc78_3525, \9310 );
and \U$3357 ( \12442 , RIe1afaf0_3376, \9312 );
and \U$3358 ( \12443 , RIe172128_2675, \9314 );
or \U$3359 ( \12444 , \12380 , \12381 , \12382 , \12383 , \12384 , \12385 , \12386 , \12387 , \12388 , \12389 , \12390 , \12391 , \12392 , \12393 , \12394 , \12395 , \12396 , \12397 , \12398 , \12399 , \12400 , \12401 , \12402 , \12403 , \12404 , \12405 , \12406 , \12407 , \12408 , \12409 , \12410 , \12411 , \12412 , \12413 , \12414 , \12415 , \12416 , \12417 , \12418 , \12419 , \12420 , \12421 , \12422 , \12423 , \12424 , \12425 , \12426 , \12427 , \12428 , \12429 , \12430 , \12431 , \12432 , \12433 , \12434 , \12435 , \12436 , \12437 , \12438 , \12439 , \12440 , \12441 , \12442 , \12443 );
or \U$3360 ( \12445 , \12379 , \12444 );
_DC g6584 ( \12446_nG6584 , \12445 , \9323 );
and g6585 ( \12447_nG6585 , \12314_nG6583 , \12446_nG6584 );
buf \U$3361 ( \12448 , \12447_nG6585 );
and \U$3362 ( \12449 , \12448 , \10691 );
nor \U$3363 ( \12450 , \12182 , \12449 );
xnor \U$3364 ( \12451 , \12450 , \10980 );
and \U$3365 ( \12452 , \10988 , \11574 );
and \U$3366 ( \12453 , \11270 , \11278 );
nor \U$3367 ( \12454 , \12452 , \12453 );
xnor \U$3368 ( \12455 , \12454 , \11580 );
xor \U$3369 ( \12456 , \12451 , \12455 );
_DC g48fe ( \12457_nG48fe , \12313 , \9597 );
_DC g4982 ( \12458_nG4982 , \12445 , \9323 );
xor g4983 ( \12459_nG4983 , \12457_nG48fe , \12458_nG4982 );
buf \U$3370 ( \12460 , \12459_nG4983 );
xor \U$3371 ( \12461 , \12460 , \11571 );
and \U$3372 ( \12462 , \10687 , \12461 );
xor \U$3373 ( \12463 , \12456 , \12462 );
and \U$3374 ( \12464 , \11589 , \11591 );
xor \U$3375 ( \12465 , \12463 , \12464 );
and \U$3376 ( \12466 , \11581 , \11592 );
and \U$3377 ( \12467 , \11593 , \11596 );
or \U$3378 ( \12468 , \12466 , \12467 );
xor \U$3379 ( \12469 , \12465 , \12468 );
buf g9c02 ( \12470_nG9c02 , \12469 );
and \U$3380 ( \12471 , \10704 , \12470_nG9c02 );
or \U$3381 ( \12472 , \12181 , \12471 );
xor \U$3382 ( \12473 , \10703 , \12472 );
buf \U$3383 ( \12474 , \12473 );
buf \U$3385 ( \12475 , \12474 );
xor \U$3386 ( \12476 , \12180 , \12475 );
and \U$3387 ( \12477 , \11605 , \12476 );
and \U$3388 ( \12478 , \12163 , \12476 );
or \U$3389 ( \12479 , \12164 , \12477 , \12478 );
and \U$3390 ( \12480 , \12153 , \12160 );
buf \U$3391 ( \12481 , \12480 );
buf \U$3393 ( \12482 , \12481 );
and \U$3394 ( \12483 , \12157 , \10694_nG9c0e );
and \U$3395 ( \12484 , \12154 , \10995_nG9c0b );
or \U$3396 ( \12485 , \12483 , \12484 );
xor \U$3397 ( \12486 , \12153 , \12485 );
buf \U$3398 ( \12487 , \12486 );
buf \U$3400 ( \12488 , \12487 );
xor \U$3401 ( \12489 , \12482 , \12488 );
buf \U$3402 ( \12490 , \12489 );
and \U$3403 ( \12491 , \10421 , \11283_nG9c08 );
and \U$3404 ( \12492 , \10418 , \11598_nG9c05 );
or \U$3405 ( \12493 , \12491 , \12492 );
xor \U$3406 ( \12494 , \10417 , \12493 );
buf \U$3407 ( \12495 , \12494 );
buf \U$3409 ( \12496 , \12495 );
xor \U$3410 ( \12497 , \12490 , \12496 );
and \U$3411 ( \12498 , \10707 , \12470_nG9c02 );
and \U$3412 ( \12499 , \12451 , \12455 );
and \U$3413 ( \12500 , \12455 , \12462 );
and \U$3414 ( \12501 , \12451 , \12462 );
or \U$3415 ( \12502 , \12499 , \12500 , \12501 );
and \U$3416 ( \12503 , \12448 , \10983 );
and \U$3417 ( \12504 , RIdec6788_722, \9333 );
and \U$3418 ( \12505 , RIdec3a88_690, \9335 );
and \U$3419 ( \12506 , RIee20788_4828, \9337 );
and \U$3420 ( \12507 , RIdec0d88_658, \9339 );
and \U$3421 ( \12508 , RIee1f810_4817, \9341 );
and \U$3422 ( \12509 , RIdebe088_626, \9343 );
and \U$3423 ( \12510 , RIdebb388_594, \9345 );
and \U$3424 ( \12511 , RIdeb8688_562, \9347 );
and \U$3425 ( \12512 , RIfc9b1c8_6787, \9349 );
and \U$3426 ( \12513 , RIdeb2c88_498, \9351 );
and \U$3427 ( \12514 , RIfce1f38_7593, \9353 );
and \U$3428 ( \12515 , RIdeaff88_466, \9355 );
and \U$3429 ( \12516 , RIfc892e8_6583, \9357 );
and \U$3430 ( \12517 , RIdead210_434, \9359 );
and \U$3431 ( \12518 , RIdea6910_402, \9361 );
and \U$3432 ( \12519 , RIdea0010_370, \9363 );
and \U$3433 ( \12520 , RIee1d650_4793, \9365 );
and \U$3434 ( \12521 , RIee1c570_4781, \9367 );
and \U$3435 ( \12522 , RIee1b5f8_4770, \9369 );
and \U$3436 ( \12523 , RIee1aef0_4765, \9371 );
and \U$3437 ( \12524 , RIfe99888_8091, \9373 );
and \U$3438 ( \12525 , RIfe99450_8088, \9375 );
and \U$3439 ( \12526 , RIfe99720_8090, \9377 );
and \U$3440 ( \12527 , RIfe995b8_8089, \9379 );
and \U$3441 ( \12528 , RIde83168_229, \9381 );
and \U$3442 ( \12529 , RIfcc43e8_7255, \9383 );
and \U$3443 ( \12530 , RIfcd5a58_7453, \9385 );
and \U$3444 ( \12531 , RIfc89450_6584, \9387 );
and \U$3445 ( \12532 , RIfcc5798_7269, \9389 );
and \U$3446 ( \12533 , RIe16c890_2612, \9391 );
and \U$3447 ( \12534 , RIe16a568_2587, \9393 );
and \U$3448 ( \12535 , RIe168d80_2570, \9395 );
and \U$3449 ( \12536 , RIe166788_2543, \9397 );
and \U$3450 ( \12537 , RIe163a88_2511, \9399 );
and \U$3451 ( \12538 , RIfc83618_6517, \9401 );
and \U$3452 ( \12539 , RIe160d88_2479, \9403 );
and \U$3453 ( \12540 , RIee36718_5078, \9405 );
and \U$3454 ( \12541 , RIe15e088_2447, \9407 );
and \U$3455 ( \12542 , RIe158688_2383, \9409 );
and \U$3456 ( \12543 , RIe155988_2351, \9411 );
and \U$3457 ( \12544 , RIfc3f800_5748, \9413 );
and \U$3458 ( \12545 , RIe152c88_2319, \9415 );
and \U$3459 ( \12546 , RIfc895b8_6585, \9417 );
and \U$3460 ( \12547 , RIe14ff88_2287, \9419 );
and \U$3461 ( \12548 , RIfc51cf8_5953, \9421 );
and \U$3462 ( \12549 , RIe14d288_2255, \9423 );
and \U$3463 ( \12550 , RIe14a588_2223, \9425 );
and \U$3464 ( \12551 , RIe147888_2191, \9427 );
and \U$3465 ( \12552 , RIee34990_5057, \9429 );
and \U$3466 ( \12553 , RIee338b0_5045, \9431 );
and \U$3467 ( \12554 , RIfc831e0_6514, \9433 );
and \U$3468 ( \12555 , RIfcd3b68_7431, \9435 );
and \U$3469 ( \12556 , RIe141ff0_2128, \9437 );
and \U$3470 ( \12557 , RIe13fcc8_2103, \9439 );
and \U$3471 ( \12558 , RIdf3dbd0_2079, \9441 );
and \U$3472 ( \12559 , RIdf3b740_2053, \9443 );
and \U$3473 ( \12560 , RIfcb6f90_7104, \9445 );
and \U$3474 ( \12561 , RIee301d8_5006, \9447 );
and \U$3475 ( \12562 , RIfcba938_7145, \9449 );
and \U$3476 ( \12563 , RIee2e018_4982, \9451 );
and \U$3477 ( \12564 , RIdf369e8_1998, \9453 );
and \U$3478 ( \12565 , RIdf343f0_1971, \9455 );
and \U$3479 ( \12566 , RIdf32230_1947, \9457 );
and \U$3480 ( \12567 , RIfe99e28_8095, \9459 );
or \U$3481 ( \12568 , \12504 , \12505 , \12506 , \12507 , \12508 , \12509 , \12510 , \12511 , \12512 , \12513 , \12514 , \12515 , \12516 , \12517 , \12518 , \12519 , \12520 , \12521 , \12522 , \12523 , \12524 , \12525 , \12526 , \12527 , \12528 , \12529 , \12530 , \12531 , \12532 , \12533 , \12534 , \12535 , \12536 , \12537 , \12538 , \12539 , \12540 , \12541 , \12542 , \12543 , \12544 , \12545 , \12546 , \12547 , \12548 , \12549 , \12550 , \12551 , \12552 , \12553 , \12554 , \12555 , \12556 , \12557 , \12558 , \12559 , \12560 , \12561 , \12562 , \12563 , \12564 , \12565 , \12566 , \12567 );
and \U$3482 ( \12569 , RIfc83078_6513, \9462 );
and \U$3483 ( \12570 , RIfcb6e28_7103, \9464 );
and \U$3484 ( \12571 , RIfc9ad90_6784, \9466 );
and \U$3485 ( \12572 , RIfcbad70_7148, \9468 );
and \U$3486 ( \12573 , RIdf2b1b0_1867, \9470 );
and \U$3487 ( \12574 , RIdf292c0_1845, \9472 );
and \U$3488 ( \12575 , RIfe99b58_8093, \9474 );
and \U$3489 ( \12576 , RIfe999f0_8092, \9476 );
and \U$3490 ( \12577 , RIfc9ac28_6783, \9478 );
and \U$3491 ( \12578 , RIfc4a9a8_5871, \9480 );
and \U$3492 ( \12579 , RIdf23758_1780, \9482 );
and \U$3493 ( \12580 , RIfc82da8_6511, \9484 );
and \U$3494 ( \12581 , RIdf220d8_1764, \9486 );
and \U$3495 ( \12582 , RIdf20a58_1748, \9488 );
and \U$3496 ( \12583 , RIdf1ba30_1691, \9490 );
and \U$3497 ( \12584 , RIfe99cc0_8094, \9492 );
and \U$3498 ( \12585 , RIdf18358_1652, \9494 );
and \U$3499 ( \12586 , RIdf15658_1620, \9496 );
and \U$3500 ( \12587 , RIdf12958_1588, \9498 );
and \U$3501 ( \12588 , RIdf0fc58_1556, \9500 );
and \U$3502 ( \12589 , RIdf0cf58_1524, \9502 );
and \U$3503 ( \12590 , RIdf0a258_1492, \9504 );
and \U$3504 ( \12591 , RIdf07558_1460, \9506 );
and \U$3505 ( \12592 , RIdf04858_1428, \9508 );
and \U$3506 ( \12593 , RIdefee58_1364, \9510 );
and \U$3507 ( \12594 , RIdefc158_1332, \9512 );
and \U$3508 ( \12595 , RIdef9458_1300, \9514 );
and \U$3509 ( \12596 , RIdef6758_1268, \9516 );
and \U$3510 ( \12597 , RIdef3a58_1236, \9518 );
and \U$3511 ( \12598 , RIdef0d58_1204, \9520 );
and \U$3512 ( \12599 , RIdeee058_1172, \9522 );
and \U$3513 ( \12600 , RIdeeb358_1140, \9524 );
and \U$3514 ( \12601 , RIee25918_4886, \9526 );
and \U$3515 ( \12602 , RIee24b08_4876, \9528 );
and \U$3516 ( \12603 , RIfc52568_5959, \9530 );
and \U$3517 ( \12604 , RIfc826a0_6506, \9532 );
and \U$3518 ( \12605 , RIdee5958_1076, \9534 );
and \U$3519 ( \12606 , RIdee3bd0_1055, \9536 );
and \U$3520 ( \12607 , RIfe99f90_8096, \9538 );
and \U$3521 ( \12608 , RIdedf9b8_1008, \9540 );
and \U$3522 ( \12609 , RIfce4800_7622, \9542 );
and \U$3523 ( \12610 , RIfc89b58_6589, \9544 );
and \U$3524 ( \12611 , RIfc9f3e0_6834, \9546 );
and \U$3525 ( \12612 , RIfc82538_6505, \9548 );
and \U$3526 ( \12613 , RIdeda828_950, \9550 );
and \U$3527 ( \12614 , RIded8398_924, \9552 );
and \U$3528 ( \12615 , RIfeabe70_8272, \9554 );
and \U$3529 ( \12616 , RIded3eb0_875, \9556 );
and \U$3530 ( \12617 , RIded1b88_850, \9558 );
and \U$3531 ( \12618 , RIdecee88_818, \9560 );
and \U$3532 ( \12619 , RIdecc188_786, \9562 );
and \U$3533 ( \12620 , RIdec9488_754, \9564 );
and \U$3534 ( \12621 , RIdeb5988_530, \9566 );
and \U$3535 ( \12622 , RIde99710_338, \9568 );
and \U$3536 ( \12623 , RIe16f590_2644, \9570 );
and \U$3537 ( \12624 , RIe15b388_2415, \9572 );
and \U$3538 ( \12625 , RIe144b88_2159, \9574 );
and \U$3539 ( \12626 , RIdf39580_2029, \9576 );
and \U$3540 ( \12627 , RIdf2dbe0_1897, \9578 );
and \U$3541 ( \12628 , RIdf1e460_1721, \9580 );
and \U$3542 ( \12629 , RIdf01b58_1396, \9582 );
and \U$3543 ( \12630 , RIdee8658_1108, \9584 );
and \U$3544 ( \12631 , RIdedd3c0_981, \9586 );
and \U$3545 ( \12632 , RIde7f658_211, \9588 );
or \U$3546 ( \12633 , \12569 , \12570 , \12571 , \12572 , \12573 , \12574 , \12575 , \12576 , \12577 , \12578 , \12579 , \12580 , \12581 , \12582 , \12583 , \12584 , \12585 , \12586 , \12587 , \12588 , \12589 , \12590 , \12591 , \12592 , \12593 , \12594 , \12595 , \12596 , \12597 , \12598 , \12599 , \12600 , \12601 , \12602 , \12603 , \12604 , \12605 , \12606 , \12607 , \12608 , \12609 , \12610 , \12611 , \12612 , \12613 , \12614 , \12615 , \12616 , \12617 , \12618 , \12619 , \12620 , \12621 , \12622 , \12623 , \12624 , \12625 , \12626 , \12627 , \12628 , \12629 , \12630 , \12631 , \12632 );
or \U$3547 ( \12634 , \12568 , \12633 );
_DC g6586 ( \12635_nG6586 , \12634 , \9597 );
and \U$3548 ( \12636 , RIe19ea20_3182, \9059 );
and \U$3549 ( \12637 , RIe19bd20_3150, \9061 );
and \U$3550 ( \12638 , RIf145928_5251, \9063 );
and \U$3551 ( \12639 , RIe199020_3118, \9065 );
and \U$3552 ( \12640 , RIfe98910_8080, \9067 );
and \U$3553 ( \12641 , RIe196320_3086, \9069 );
and \U$3554 ( \12642 , RIe193620_3054, \9071 );
and \U$3555 ( \12643 , RIe190920_3022, \9073 );
and \U$3556 ( \12644 , RIe18af20_2958, \9075 );
and \U$3557 ( \12645 , RIe188220_2926, \9077 );
and \U$3558 ( \12646 , RIf143e70_5232, \9079 );
and \U$3559 ( \12647 , RIe185520_2894, \9081 );
and \U$3560 ( \12648 , RIfc95c00_6726, \9083 );
and \U$3561 ( \12649 , RIe182820_2862, \9085 );
and \U$3562 ( \12650 , RIe17fb20_2830, \9087 );
and \U$3563 ( \12651 , RIe17ce20_2798, \9089 );
and \U$3564 ( \12652 , RIf142520_5214, \9091 );
and \U$3565 ( \12653 , RIf141440_5202, \9093 );
and \U$3566 ( \12654 , RIe1776f0_2736, \9095 );
and \U$3567 ( \12655 , RIfeab8d0_8268, \9097 );
and \U$3568 ( \12656 , RIfcc5bd0_7272, \9099 );
and \U$3569 ( \12657 , RIfc62dc8_6147, \9101 );
and \U$3570 ( \12658 , RIee3e710_5169, \9103 );
and \U$3571 ( \12659 , RIfc9cb18_6805, \9105 );
and \U$3572 ( \12660 , RIee3c820_5147, \9107 );
and \U$3573 ( \12661 , RIee3b470_5133, \9109 );
and \U$3574 ( \12662 , RIee3a390_5121, \9111 );
and \U$3575 ( \12663 , RIe174888_2703, \9113 );
and \U$3576 ( \12664 , RIf170498_5737, \9115 );
and \U$3577 ( \12665 , RIfc68660_6210, \9117 );
and \U$3578 ( \12666 , RIf16e878_5717, \9119 );
and \U$3579 ( \12667 , RIfc6ea38_6281, \9121 );
and \U$3580 ( \12668 , RIfe98d48_8083, \9123 );
and \U$3581 ( \12669 , RIe224d78_4709, \9125 );
and \U$3582 ( \12670 , RIf16c280_5690, \9127 );
and \U$3583 ( \12671 , RIe222078_4677, \9129 );
and \U$3584 ( \12672 , RIf16b308_5679, \9131 );
and \U$3585 ( \12673 , RIe21f378_4645, \9133 );
and \U$3586 ( \12674 , RIe219978_4581, \9135 );
and \U$3587 ( \12675 , RIe216c78_4549, \9137 );
and \U$3588 ( \12676 , RIf16a390_5668, \9139 );
and \U$3589 ( \12677 , RIe213f78_4517, \9141 );
and \U$3590 ( \12678 , RIf169b20_5662, \9143 );
and \U$3591 ( \12679 , RIe211278_4485, \9145 );
and \U$3592 ( \12680 , RIf1681d0_5644, \9147 );
and \U$3593 ( \12681 , RIe20e578_4453, \9149 );
and \U$3594 ( \12682 , RIe20b878_4421, \9151 );
and \U$3595 ( \12683 , RIe208b78_4389, \9153 );
and \U$3596 ( \12684 , RIfcd4ae0_7442, \9155 );
and \U$3597 ( \12685 , RIfc61478_6129, \9157 );
and \U$3598 ( \12686 , RIfeab060_8262, \9159 );
and \U$3599 ( \12687 , RIe201990_4308, \9161 );
and \U$3600 ( \12688 , RIfc70ec8_6307, \9163 );
and \U$3601 ( \12689 , RIfc70928_6303, \9165 );
and \U$3602 ( \12690 , RIfcec528_7711, \9167 );
and \U$3603 ( \12691 , RIfcbe880_7190, \9169 );
and \U$3604 ( \12692 , RIf160d18_5561, \9171 );
and \U$3605 ( \12693 , RIf15ee28_5539, \9173 );
and \U$3606 ( \12694 , RIfe98be0_8082, \9175 );
and \U$3607 ( \12695 , RIfe98eb0_8084, \9177 );
and \U$3608 ( \12696 , RIf15d0a0_5518, \9179 );
and \U$3609 ( \12697 , RIf15bcf0_5504, \9181 );
and \U$3610 ( \12698 , RIfcd4540_7438, \9183 );
and \U$3611 ( \12699 , RIf159e00_5482, \9185 );
or \U$3612 ( \12700 , \12636 , \12637 , \12638 , \12639 , \12640 , \12641 , \12642 , \12643 , \12644 , \12645 , \12646 , \12647 , \12648 , \12649 , \12650 , \12651 , \12652 , \12653 , \12654 , \12655 , \12656 , \12657 , \12658 , \12659 , \12660 , \12661 , \12662 , \12663 , \12664 , \12665 , \12666 , \12667 , \12668 , \12669 , \12670 , \12671 , \12672 , \12673 , \12674 , \12675 , \12676 , \12677 , \12678 , \12679 , \12680 , \12681 , \12682 , \12683 , \12684 , \12685 , \12686 , \12687 , \12688 , \12689 , \12690 , \12691 , \12692 , \12693 , \12694 , \12695 , \12696 , \12697 , \12698 , \12699 );
and \U$3613 ( \12701 , RIf1592c0_5474, \9188 );
and \U$3614 ( \12702 , RIf158078_5461, \9190 );
and \U$3615 ( \12703 , RIfca3a30_6884, \9192 );
and \U$3616 ( \12704 , RIfea7988_8223, \9194 );
and \U$3617 ( \12705 , RIf156728_5443, \9196 );
and \U$3618 ( \12706 , RIf155be8_5435, \9198 );
and \U$3619 ( \12707 , RIf154b08_5423, \9200 );
and \U$3620 ( \12708 , RIfe98a78_8081, \9202 );
and \U$3621 ( \12709 , RIf1538c0_5410, \9204 );
and \U$3622 ( \12710 , RIf1520d8_5393, \9206 );
and \U$3623 ( \12711 , RIf150e90_5380, \9208 );
and \U$3624 ( \12712 , RIe1f43d0_4156, \9210 );
and \U$3625 ( \12713 , RIf14fdb0_5368, \9212 );
and \U$3626 ( \12714 , RIfcd2380_7414, \9214 );
and \U$3627 ( \12715 , RIf14e2f8_5349, \9216 );
and \U$3628 ( \12716 , RIe1ef240_4098, \9218 );
and \U$3629 ( \12717 , RIe1ecae0_4070, \9220 );
and \U$3630 ( \12718 , RIe1e9de0_4038, \9222 );
and \U$3631 ( \12719 , RIe1e70e0_4006, \9224 );
and \U$3632 ( \12720 , RIe1e43e0_3974, \9226 );
and \U$3633 ( \12721 , RIe1e16e0_3942, \9228 );
and \U$3634 ( \12722 , RIe1de9e0_3910, \9230 );
and \U$3635 ( \12723 , RIe1dbce0_3878, \9232 );
and \U$3636 ( \12724 , RIe1d8fe0_3846, \9234 );
and \U$3637 ( \12725 , RIe1d35e0_3782, \9236 );
and \U$3638 ( \12726 , RIe1d08e0_3750, \9238 );
and \U$3639 ( \12727 , RIe1cdbe0_3718, \9240 );
and \U$3640 ( \12728 , RIe1caee0_3686, \9242 );
and \U$3641 ( \12729 , RIe1c81e0_3654, \9244 );
and \U$3642 ( \12730 , RIe1c54e0_3622, \9246 );
and \U$3643 ( \12731 , RIe1c27e0_3590, \9248 );
and \U$3644 ( \12732 , RIe1bfae0_3558, \9250 );
and \U$3645 ( \12733 , RIfc44b70_5804, \9252 );
and \U$3646 ( \12734 , RIf14bd00_5322, \9254 );
and \U$3647 ( \12735 , RIfe992e8_8087, \9256 );
and \U$3648 ( \12736 , RIfe987a8_8079, \9258 );
and \U$3649 ( \12737 , RIf14a950_5308, \9260 );
and \U$3650 ( \12738 , RIf149f78_5301, \9262 );
and \U$3651 ( \12739 , RIfe99180_8086, \9264 );
and \U$3652 ( \12740 , RIfe98640_8078, \9266 );
and \U$3653 ( \12741 , RIf149438_5293, \9268 );
and \U$3654 ( \12742 , RIfcec7f8_7713, \9270 );
and \U$3655 ( \12743 , RIfe984d8_8077, \9272 );
and \U$3656 ( \12744 , RIe1b1b48_3399, \9274 );
and \U$3657 ( \12745 , RIfc4b650_5880, \9276 );
and \U$3658 ( \12746 , RIfcda918_7509, \9278 );
and \U$3659 ( \12747 , RIfe98370_8076, \9280 );
and \U$3660 ( \12748 , RIfe99018_8085, \9282 );
and \U$3661 ( \12749 , RIe1a9e20_3310, \9284 );
and \U$3662 ( \12750 , RIe1a7120_3278, \9286 );
and \U$3663 ( \12751 , RIe1a4420_3246, \9288 );
and \U$3664 ( \12752 , RIe1a1720_3214, \9290 );
and \U$3665 ( \12753 , RIe18dc20_2990, \9292 );
and \U$3666 ( \12754 , RIe17a120_2766, \9294 );
and \U$3667 ( \12755 , RIe227a78_4741, \9296 );
and \U$3668 ( \12756 , RIe21c678_4613, \9298 );
and \U$3669 ( \12757 , RIe205e78_4357, \9300 );
and \U$3670 ( \12758 , RIe1ffed8_4289, \9302 );
and \U$3671 ( \12759 , RIe1f9290_4212, \9304 );
and \U$3672 ( \12760 , RIe1f1dd8_4129, \9306 );
and \U$3673 ( \12761 , RIe1d62e0_3814, \9308 );
and \U$3674 ( \12762 , RIe1bcde0_3526, \9310 );
and \U$3675 ( \12763 , RIe1afc58_3377, \9312 );
and \U$3676 ( \12764 , RIe172290_2676, \9314 );
or \U$3677 ( \12765 , \12701 , \12702 , \12703 , \12704 , \12705 , \12706 , \12707 , \12708 , \12709 , \12710 , \12711 , \12712 , \12713 , \12714 , \12715 , \12716 , \12717 , \12718 , \12719 , \12720 , \12721 , \12722 , \12723 , \12724 , \12725 , \12726 , \12727 , \12728 , \12729 , \12730 , \12731 , \12732 , \12733 , \12734 , \12735 , \12736 , \12737 , \12738 , \12739 , \12740 , \12741 , \12742 , \12743 , \12744 , \12745 , \12746 , \12747 , \12748 , \12749 , \12750 , \12751 , \12752 , \12753 , \12754 , \12755 , \12756 , \12757 , \12758 , \12759 , \12760 , \12761 , \12762 , \12763 , \12764 );
or \U$3678 ( \12766 , \12700 , \12765 );
_DC g6587 ( \12767_nG6587 , \12766 , \9323 );
and g6588 ( \12768_nG6588 , \12635_nG6586 , \12767_nG6587 );
buf \U$3679 ( \12769 , \12768_nG6588 );
and \U$3680 ( \12770 , \12769 , \10691 );
nor \U$3681 ( \12771 , \12503 , \12770 );
xnor \U$3682 ( \12772 , \12771 , \10980 );
not \U$3683 ( \12773 , \12462 );
_DC g4a07 ( \12774_nG4a07 , \12634 , \9597 );
_DC g4a8b ( \12775_nG4a8b , \12766 , \9323 );
xor g4a8c ( \12776_nG4a8c , \12774_nG4a07 , \12775_nG4a8b );
buf \U$3684 ( \12777 , \12776_nG4a8c );
and \U$3685 ( \12778 , \12460 , \11571 );
not \U$3686 ( \12779 , \12778 );
and \U$3687 ( \12780 , \12777 , \12779 );
and \U$3688 ( \12781 , \12773 , \12780 );
xor \U$3689 ( \12782 , \12772 , \12781 );
and \U$3690 ( \12783 , \11270 , \11574 );
and \U$3691 ( \12784 , \11586 , \11278 );
nor \U$3692 ( \12785 , \12783 , \12784 );
xnor \U$3693 ( \12786 , \12785 , \11580 );
xor \U$3694 ( \12787 , \12782 , \12786 );
xor \U$3695 ( \12788 , \12777 , \12460 );
not \U$3696 ( \12789 , \12461 );
and \U$3697 ( \12790 , \12788 , \12789 );
and \U$3698 ( \12791 , \10687 , \12790 );
and \U$3699 ( \12792 , \10988 , \12461 );
nor \U$3700 ( \12793 , \12791 , \12792 );
xnor \U$3701 ( \12794 , \12793 , \12780 );
xor \U$3702 ( \12795 , \12787 , \12794 );
xor \U$3703 ( \12796 , \12502 , \12795 );
and \U$3704 ( \12797 , \12463 , \12464 );
and \U$3705 ( \12798 , \12465 , \12468 );
or \U$3706 ( \12799 , \12797 , \12798 );
xor \U$3707 ( \12800 , \12796 , \12799 );
buf g9bff ( \12801_nG9bff , \12800 );
and \U$3708 ( \12802 , \10704 , \12801_nG9bff );
or \U$3709 ( \12803 , \12498 , \12802 );
xor \U$3710 ( \12804 , \10703 , \12803 );
buf \U$3711 ( \12805 , \12804 );
buf \U$3713 ( \12806 , \12805 );
xor \U$3714 ( \12807 , \12497 , \12806 );
buf \U$3715 ( \12808 , \12807 );
and \U$3716 ( \12809 , \12174 , \12179 );
and \U$3717 ( \12810 , \12174 , \12475 );
and \U$3718 ( \12811 , \12179 , \12475 );
or \U$3719 ( \12812 , \12809 , \12810 , \12811 );
buf \U$3720 ( \12813 , \12812 );
xor \U$3721 ( \12814 , \12808 , \12813 );
and \U$3722 ( \12815 , \12166 , \12172 );
buf \U$3723 ( \12816 , \12815 );
xor \U$3724 ( \12817 , \12814 , \12816 );
and \U$3725 ( \12818 , \12479 , \12817 );
and \U$3726 ( \12819 , RIdec6a58_724, \9059 );
and \U$3727 ( \12820 , RIdec3d58_692, \9061 );
and \U$3728 ( \12821 , RIfc723e0_6322, \9063 );
and \U$3729 ( \12822 , RIdec1058_660, \9065 );
and \U$3730 ( \12823 , RIfc59fc0_6046, \9067 );
and \U$3731 ( \12824 , RIdebe358_628, \9069 );
and \U$3732 ( \12825 , RIdebb658_596, \9071 );
and \U$3733 ( \12826 , RIdeb8958_564, \9073 );
and \U$3734 ( \12827 , RIfcb96f0_7132, \9075 );
and \U$3735 ( \12828 , RIdeb2f58_500, \9077 );
and \U$3736 ( \12829 , RIfce1c68_7591, \9079 );
and \U$3737 ( \12830 , RIdeb0258_468, \9081 );
and \U$3738 ( \12831 , RIfc9b498_6789, \9083 );
and \U$3739 ( \12832 , RIdead558_436, \9085 );
and \U$3740 ( \12833 , RIdea6fa0_404, \9087 );
and \U$3741 ( \12834 , RIdea06a0_372, \9089 );
and \U$3742 ( \12835 , RIfc81458_6493, \9091 );
and \U$3743 ( \12836 , RIfc83780_6518, \9093 );
and \U$3744 ( \12837 , RIfc4e620_5914, \9095 );
and \U$3745 ( \12838 , RIfcd3e38_7433, \9097 );
and \U$3746 ( \12839 , RIde937e8_309, \9099 );
and \U$3747 ( \12840 , RIde8f990_290, \9101 );
and \U$3748 ( \12841 , RIde8bb38_271, \9103 );
and \U$3749 ( \12842 , RIde87650_250, \9105 );
and \U$3750 ( \12843 , RIde834b0_230, \9107 );
and \U$3751 ( \12844 , RIfc42c80_5782, \9109 );
and \U$3752 ( \12845 , RIfc65960_6178, \9111 );
and \U$3753 ( \12846 , RIfc6c710_6256, \9113 );
and \U$3754 ( \12847 , RIee392b0_5109, \9115 );
and \U$3755 ( \12848 , RIe16cb60_2614, \9117 );
and \U$3756 ( \12849 , RIe16a6d0_2588, \9119 );
and \U$3757 ( \12850 , RIe169050_2572, \9121 );
and \U$3758 ( \12851 , RIe166a58_2545, \9123 );
and \U$3759 ( \12852 , RIe163d58_2513, \9125 );
and \U$3760 ( \12853 , RIfec3cf0_8348, \9127 );
and \U$3761 ( \12854 , RIe161058_2481, \9129 );
and \U$3762 ( \12855 , RIfcd54b8_7449, \9131 );
and \U$3763 ( \12856 , RIe15e358_2449, \9133 );
and \U$3764 ( \12857 , RIe158958_2385, \9135 );
and \U$3765 ( \12858 , RIe155c58_2353, \9137 );
and \U$3766 ( \12859 , RIfe9ba48_8115, \9139 );
and \U$3767 ( \12860 , RIe152f58_2321, \9141 );
and \U$3768 ( \12861 , RIfec4128_8351, \9143 );
and \U$3769 ( \12862 , RIe150258_2289, \9145 );
and \U$3770 ( \12863 , RIfcb9b28_7135, \9147 );
and \U$3771 ( \12864 , RIe14d558_2257, \9149 );
and \U$3772 ( \12865 , RIe14a858_2225, \9151 );
and \U$3773 ( \12866 , RIe147b58_2193, \9153 );
and \U$3774 ( \12867 , RIfcdb2f0_7516, \9155 );
and \U$3775 ( \12868 , RIfc553d0_5992, \9157 );
and \U$3776 ( \12869 , RIfc9a0e8_6775, \9159 );
and \U$3777 ( \12870 , RIfcbd908_7179, \9161 );
and \U$3778 ( \12871 , RIe1422c0_2130, \9163 );
and \U$3779 ( \12872 , RIe13ff98_2105, \9165 );
and \U$3780 ( \12873 , RIdf3dea0_2081, \9167 );
and \U$3781 ( \12874 , RIdf3ba10_2055, \9169 );
and \U$3782 ( \12875 , RIfc87128_6559, \9171 );
and \U$3783 ( \12876 , RIee304a8_5008, \9173 );
and \U$3784 ( \12877 , RIfcc51f8_7265, \9175 );
and \U$3785 ( \12878 , RIee2e2e8_4984, \9177 );
and \U$3786 ( \12879 , RIdf36cb8_2000, \9179 );
and \U$3787 ( \12880 , RIfec3fc0_8350, \9181 );
and \U$3788 ( \12881 , RIdf32500_1949, \9183 );
and \U$3789 ( \12882 , RIfec3e58_8349, \9185 );
or \U$3790 ( \12883 , \12819 , \12820 , \12821 , \12822 , \12823 , \12824 , \12825 , \12826 , \12827 , \12828 , \12829 , \12830 , \12831 , \12832 , \12833 , \12834 , \12835 , \12836 , \12837 , \12838 , \12839 , \12840 , \12841 , \12842 , \12843 , \12844 , \12845 , \12846 , \12847 , \12848 , \12849 , \12850 , \12851 , \12852 , \12853 , \12854 , \12855 , \12856 , \12857 , \12858 , \12859 , \12860 , \12861 , \12862 , \12863 , \12864 , \12865 , \12866 , \12867 , \12868 , \12869 , \12870 , \12871 , \12872 , \12873 , \12874 , \12875 , \12876 , \12877 , \12878 , \12879 , \12880 , \12881 , \12882 );
and \U$3791 ( \12884 , RIee2c830_4965, \9188 );
and \U$3792 ( \12885 , RIee2ad78_4946, \9190 );
and \U$3793 ( \12886 , RIee296f8_4930, \9192 );
and \U$3794 ( \12887 , RIee284b0_4917, \9194 );
and \U$3795 ( \12888 , RIfe9b8e0_8114, \9196 );
and \U$3796 ( \12889 , RIfe9b610_8112, \9198 );
and \U$3797 ( \12890 , RIfe9b778_8113, \9200 );
and \U$3798 ( \12891 , RIfe9b4a8_8111, \9202 );
and \U$3799 ( \12892 , RIfcb7c38_7113, \9204 );
and \U$3800 ( \12893 , RIfc86b88_6555, \9206 );
and \U$3801 ( \12894 , RIdf238c0_1781, \9208 );
and \U$3802 ( \12895 , RIfc75ab8_6361, \9210 );
and \U$3803 ( \12896 , RIdf22240_1765, \9212 );
and \U$3804 ( \12897 , RIfeaa3b8_8253, \9214 );
and \U$3805 ( \12898 , RIdf1bb98_1692, \9216 );
and \U$3806 ( \12899 , RIdf1a680_1677, \9218 );
and \U$3807 ( \12900 , RIdf18628_1654, \9220 );
and \U$3808 ( \12901 , RIdf15928_1622, \9222 );
and \U$3809 ( \12902 , RIdf12c28_1590, \9224 );
and \U$3810 ( \12903 , RIdf0ff28_1558, \9226 );
and \U$3811 ( \12904 , RIdf0d228_1526, \9228 );
and \U$3812 ( \12905 , RIdf0a528_1494, \9230 );
and \U$3813 ( \12906 , RIdf07828_1462, \9232 );
and \U$3814 ( \12907 , RIdf04b28_1430, \9234 );
and \U$3815 ( \12908 , RIdeff128_1366, \9236 );
and \U$3816 ( \12909 , RIdefc428_1334, \9238 );
and \U$3817 ( \12910 , RIdef9728_1302, \9240 );
and \U$3818 ( \12911 , RIdef6a28_1270, \9242 );
and \U$3819 ( \12912 , RIdef3d28_1238, \9244 );
and \U$3820 ( \12913 , RIdef1028_1206, \9246 );
and \U$3821 ( \12914 , RIdeee328_1174, \9248 );
and \U$3822 ( \12915 , RIdeeb628_1142, \9250 );
and \U$3823 ( \12916 , RIee25a80_4887, \9252 );
and \U$3824 ( \12917 , RIee24c70_4877, \9254 );
and \U$3825 ( \12918 , RIfcddd20_7546, \9256 );
and \U$3826 ( \12919 , RIfccc110_7344, \9258 );
and \U$3827 ( \12920 , RIdee5c28_1078, \9260 );
and \U$3828 ( \12921 , RIdee3ea0_1057, \9262 );
and \U$3829 ( \12922 , RIdee1b78_1032, \9264 );
and \U$3830 ( \12923 , RIdedfc88_1010, \9266 );
and \U$3831 ( \12924 , RIfc6a6b8_6233, \9268 );
and \U$3832 ( \12925 , RIee227e0_4851, \9270 );
and \U$3833 ( \12926 , RIfc88be0_6578, \9272 );
and \U$3834 ( \12927 , RIee21868_4840, \9274 );
and \U$3835 ( \12928 , RIdedaaf8_952, \9276 );
and \U$3836 ( \12929 , RIded8668_926, \9278 );
and \U$3837 ( \12930 , RIded6340_901, \9280 );
and \U$3838 ( \12931 , RIded4180_877, \9282 );
and \U$3839 ( \12932 , RIded1e58_852, \9284 );
and \U$3840 ( \12933 , RIdecf158_820, \9286 );
and \U$3841 ( \12934 , RIdecc458_788, \9288 );
and \U$3842 ( \12935 , RIdec9758_756, \9290 );
and \U$3843 ( \12936 , RIdeb5c58_532, \9292 );
and \U$3844 ( \12937 , RIde99da0_340, \9294 );
and \U$3845 ( \12938 , RIe16f860_2646, \9296 );
and \U$3846 ( \12939 , RIe15b658_2417, \9298 );
and \U$3847 ( \12940 , RIe144e58_2161, \9300 );
and \U$3848 ( \12941 , RIdf39850_2031, \9302 );
and \U$3849 ( \12942 , RIdf2deb0_1899, \9304 );
and \U$3850 ( \12943 , RIdf1e730_1723, \9306 );
and \U$3851 ( \12944 , RIdf01e28_1398, \9308 );
and \U$3852 ( \12945 , RIdee8928_1110, \9310 );
and \U$3853 ( \12946 , RIdedd690_983, \9312 );
and \U$3854 ( \12947 , RIde7fce8_213, \9314 );
or \U$3855 ( \12948 , \12884 , \12885 , \12886 , \12887 , \12888 , \12889 , \12890 , \12891 , \12892 , \12893 , \12894 , \12895 , \12896 , \12897 , \12898 , \12899 , \12900 , \12901 , \12902 , \12903 , \12904 , \12905 , \12906 , \12907 , \12908 , \12909 , \12910 , \12911 , \12912 , \12913 , \12914 , \12915 , \12916 , \12917 , \12918 , \12919 , \12920 , \12921 , \12922 , \12923 , \12924 , \12925 , \12926 , \12927 , \12928 , \12929 , \12930 , \12931 , \12932 , \12933 , \12934 , \12935 , \12936 , \12937 , \12938 , \12939 , \12940 , \12941 , \12942 , \12943 , \12944 , \12945 , \12946 , \12947 );
or \U$3856 ( \12949 , \12883 , \12948 );
_DC g2ead ( \12950_nG2ead , \12949 , \9323 );
buf \U$3857 ( \12951 , \12950_nG2ead );
and \U$3858 ( \12952 , RIe19ecf0_3184, \9333 );
and \U$3859 ( \12953 , RIe19bff0_3152, \9335 );
and \U$3860 ( \12954 , RIf145a90_5252, \9337 );
and \U$3861 ( \12955 , RIe1992f0_3120, \9339 );
and \U$3862 ( \12956 , RIf144de8_5243, \9341 );
and \U$3863 ( \12957 , RIe1965f0_3088, \9343 );
and \U$3864 ( \12958 , RIe1938f0_3056, \9345 );
and \U$3865 ( \12959 , RIe190bf0_3024, \9347 );
and \U$3866 ( \12960 , RIe18b1f0_2960, \9349 );
and \U$3867 ( \12961 , RIe1884f0_2928, \9351 );
and \U$3868 ( \12962 , RIfc72980_6326, \9353 );
and \U$3869 ( \12963 , RIe1857f0_2896, \9355 );
and \U$3870 ( \12964 , RIf143060_5222, \9357 );
and \U$3871 ( \12965 , RIe182af0_2864, \9359 );
and \U$3872 ( \12966 , RIe17fdf0_2832, \9361 );
and \U$3873 ( \12967 , RIe17d0f0_2800, \9363 );
and \U$3874 ( \12968 , RIf142688_5215, \9365 );
and \U$3875 ( \12969 , RIf141710_5204, \9367 );
and \U$3876 ( \12970 , RIe177858_2737, \9369 );
and \U$3877 ( \12971 , RIe176778_2725, \9371 );
and \U$3878 ( \12972 , RIfcea638_7689, \9373 );
and \U$3879 ( \12973 , RIfca54e8_6903, \9375 );
and \U$3880 ( \12974 , RIee3e878_5170, \9377 );
and \U$3881 ( \12975 , RIee3dbd0_5161, \9379 );
and \U$3882 ( \12976 , RIee3c988_5148, \9381 );
and \U$3883 ( \12977 , RIee3b5d8_5134, \9383 );
and \U$3884 ( \12978 , RIee3a4f8_5122, \9385 );
and \U$3885 ( \12979 , RIe174b58_2705, \9387 );
and \U$3886 ( \12980 , RIf170600_5738, \9389 );
and \U$3887 ( \12981 , RIfc76fd0_6376, \9391 );
and \U$3888 ( \12982 , RIf16e9e0_5718, \9393 );
and \U$3889 ( \12983 , RIfced608_7723, \9395 );
and \U$3890 ( \12984 , RIf16d090_5700, \9397 );
and \U$3891 ( \12985 , RIe225048_4711, \9399 );
and \U$3892 ( \12986 , RIf16c550_5692, \9401 );
and \U$3893 ( \12987 , RIe222348_4679, \9403 );
and \U$3894 ( \12988 , RIf16b470_5680, \9405 );
and \U$3895 ( \12989 , RIe21f648_4647, \9407 );
and \U$3896 ( \12990 , RIe219c48_4583, \9409 );
and \U$3897 ( \12991 , RIe216f48_4551, \9411 );
and \U$3898 ( \12992 , RIf16a4f8_5669, \9413 );
and \U$3899 ( \12993 , RIe214248_4519, \9415 );
and \U$3900 ( \12994 , RIf169df0_5664, \9417 );
and \U$3901 ( \12995 , RIe211548_4487, \9419 );
and \U$3902 ( \12996 , RIf1684a0_5646, \9421 );
and \U$3903 ( \12997 , RIe20e848_4455, \9423 );
and \U$3904 ( \12998 , RIe20bb48_4423, \9425 );
and \U$3905 ( \12999 , RIe208e48_4391, \9427 );
and \U$3906 ( \13000 , RIf1673c0_5634, \9429 );
and \U$3907 ( \13001 , RIf166448_5623, \9431 );
and \U$3908 ( \13002 , RIfe9c6f0_8124, \9433 );
and \U$3909 ( \13003 , RIfe9c150_8120, \9435 );
and \U$3910 ( \13004 , RIf1654d0_5612, \9437 );
and \U$3911 ( \13005 , RIfcc4550_7256, \9439 );
and \U$3912 ( \13006 , RIf1635e0_5590, \9441 );
and \U$3913 ( \13007 , RIf162500_5578, \9443 );
and \U$3914 ( \13008 , RIf160fe8_5563, \9445 );
and \U$3915 ( \13009 , RIf15f0f8_5541, \9447 );
and \U$3916 ( \13010 , RIfe9bfe8_8119, \9449 );
and \U$3917 ( \13011 , RIfe9c588_8123, \9451 );
and \U$3918 ( \13012 , RIf15d208_5519, \9453 );
and \U$3919 ( \13013 , RIf15bfc0_5506, \9455 );
and \U$3920 ( \13014 , RIfc4d540_5902, \9457 );
and \U$3921 ( \13015 , RIfc9c848_6803, \9459 );
or \U$3922 ( \13016 , \12952 , \12953 , \12954 , \12955 , \12956 , \12957 , \12958 , \12959 , \12960 , \12961 , \12962 , \12963 , \12964 , \12965 , \12966 , \12967 , \12968 , \12969 , \12970 , \12971 , \12972 , \12973 , \12974 , \12975 , \12976 , \12977 , \12978 , \12979 , \12980 , \12981 , \12982 , \12983 , \12984 , \12985 , \12986 , \12987 , \12988 , \12989 , \12990 , \12991 , \12992 , \12993 , \12994 , \12995 , \12996 , \12997 , \12998 , \12999 , \13000 , \13001 , \13002 , \13003 , \13004 , \13005 , \13006 , \13007 , \13008 , \13009 , \13010 , \13011 , \13012 , \13013 , \13014 , \13015 );
and \U$3923 ( \13017 , RIfec4290_8352, \9462 );
and \U$3924 ( \13018 , RIfe9c2b8_8121, \9464 );
and \U$3925 ( \13019 , RIfcc01d0_7208, \9466 );
and \U$3926 ( \13020 , RIe1fb2e8_4235, \9468 );
and \U$3927 ( \13021 , RIfe9c420_8122, \9470 );
and \U$3928 ( \13022 , RIfca3e68_6887, \9472 );
and \U$3929 ( \13023 , RIf154c70_5424, \9474 );
and \U$3930 ( \13024 , RIe1f69c8_4183, \9476 );
and \U$3931 ( \13025 , RIf153a28_5411, \9478 );
and \U$3932 ( \13026 , RIf152240_5394, \9480 );
and \U$3933 ( \13027 , RIf150ff8_5381, \9482 );
and \U$3934 ( \13028 , RIe1f46a0_4158, \9484 );
and \U$3935 ( \13029 , RIfca6028_6911, \9486 );
and \U$3936 ( \13030 , RIfc43bf8_5793, \9488 );
and \U$3937 ( \13031 , RIf14e460_5350, \9490 );
and \U$3938 ( \13032 , RIe1ef3a8_4099, \9492 );
and \U$3939 ( \13033 , RIe1ecdb0_4072, \9494 );
and \U$3940 ( \13034 , RIe1ea0b0_4040, \9496 );
and \U$3941 ( \13035 , RIe1e73b0_4008, \9498 );
and \U$3942 ( \13036 , RIe1e46b0_3976, \9500 );
and \U$3943 ( \13037 , RIe1e19b0_3944, \9502 );
and \U$3944 ( \13038 , RIe1decb0_3912, \9504 );
and \U$3945 ( \13039 , RIe1dbfb0_3880, \9506 );
and \U$3946 ( \13040 , RIe1d92b0_3848, \9508 );
and \U$3947 ( \13041 , RIe1d38b0_3784, \9510 );
and \U$3948 ( \13042 , RIe1d0bb0_3752, \9512 );
and \U$3949 ( \13043 , RIe1cdeb0_3720, \9514 );
and \U$3950 ( \13044 , RIe1cb1b0_3688, \9516 );
and \U$3951 ( \13045 , RIe1c84b0_3656, \9518 );
and \U$3952 ( \13046 , RIe1c57b0_3624, \9520 );
and \U$3953 ( \13047 , RIe1c2ab0_3592, \9522 );
and \U$3954 ( \13048 , RIe1bfdb0_3560, \9524 );
and \U$3955 ( \13049 , RIfc4d6a8_5903, \9526 );
and \U$3956 ( \13050 , RIf14be68_5323, \9528 );
and \U$3957 ( \13051 , RIe1ba680_3498, \9530 );
and \U$3958 ( \13052 , RIfe9be80_8118, \9532 );
and \U$3959 ( \13053 , RIfc86e58_6557, \9534 );
and \U$3960 ( \13054 , RIfcd46a8_7439, \9536 );
and \U$3961 ( \13055 , RIe1b6300_3450, \9538 );
and \U$3962 ( \13056 , RIfe9bd18_8117, \9540 );
and \U$3963 ( \13057 , RIf1495a0_5294, \9542 );
and \U$3964 ( \13058 , RIf1481f0_5280, \9544 );
and \U$3965 ( \13059 , RIe1b3600_3418, \9546 );
and \U$3966 ( \13060 , RIe1b1e18_3401, \9548 );
and \U$3967 ( \13061 , RIfc69470_6220, \9550 );
and \U$3968 ( \13062 , RIfcbfac8_7203, \9552 );
and \U$3969 ( \13063 , RIfe9bbb0_8116, \9554 );
and \U$3970 ( \13064 , RIe1abd10_3332, \9556 );
and \U$3971 ( \13065 , RIe1aa0f0_3312, \9558 );
and \U$3972 ( \13066 , RIe1a73f0_3280, \9560 );
and \U$3973 ( \13067 , RIe1a46f0_3248, \9562 );
and \U$3974 ( \13068 , RIe1a19f0_3216, \9564 );
and \U$3975 ( \13069 , RIe18def0_2992, \9566 );
and \U$3976 ( \13070 , RIe17a3f0_2768, \9568 );
and \U$3977 ( \13071 , RIe227d48_4743, \9570 );
and \U$3978 ( \13072 , RIe21c948_4615, \9572 );
and \U$3979 ( \13073 , RIe206148_4359, \9574 );
and \U$3980 ( \13074 , RIe2001a8_4291, \9576 );
and \U$3981 ( \13075 , RIe1f9560_4214, \9578 );
and \U$3982 ( \13076 , RIe1f20a8_4131, \9580 );
and \U$3983 ( \13077 , RIe1d65b0_3816, \9582 );
and \U$3984 ( \13078 , RIe1bd0b0_3528, \9584 );
and \U$3985 ( \13079 , RIe1aff28_3379, \9586 );
and \U$3986 ( \13080 , RIe172560_2678, \9588 );
or \U$3987 ( \13081 , \13017 , \13018 , \13019 , \13020 , \13021 , \13022 , \13023 , \13024 , \13025 , \13026 , \13027 , \13028 , \13029 , \13030 , \13031 , \13032 , \13033 , \13034 , \13035 , \13036 , \13037 , \13038 , \13039 , \13040 , \13041 , \13042 , \13043 , \13044 , \13045 , \13046 , \13047 , \13048 , \13049 , \13050 , \13051 , \13052 , \13053 , \13054 , \13055 , \13056 , \13057 , \13058 , \13059 , \13060 , \13061 , \13062 , \13063 , \13064 , \13065 , \13066 , \13067 , \13068 , \13069 , \13070 , \13071 , \13072 , \13073 , \13074 , \13075 , \13076 , \13077 , \13078 , \13079 , \13080 );
or \U$3988 ( \13082 , \13016 , \13081 );
_DC g3fda ( \13083_nG3fda , \13082 , \9597 );
buf \U$3989 ( \13084 , \13083_nG3fda );
xor \U$3990 ( \13085 , \12951 , \13084 );
and \U$3991 ( \13086 , RIdec68f0_723, \9059 );
and \U$3992 ( \13087 , RIdec3bf0_691, \9061 );
and \U$3993 ( \13088 , RIee208f0_4829, \9063 );
and \U$3994 ( \13089 , RIdec0ef0_659, \9065 );
and \U$3995 ( \13090 , RIfc7ce08_6443, \9067 );
and \U$3996 ( \13091 , RIdebe1f0_627, \9069 );
and \U$3997 ( \13092 , RIdebb4f0_595, \9071 );
and \U$3998 ( \13093 , RIdeb87f0_563, \9073 );
and \U$3999 ( \13094 , RIfc9b8d0_6792, \9075 );
and \U$4000 ( \13095 , RIdeb2df0_499, \9077 );
and \U$4001 ( \13096 , RIfcc6710_7280, \9079 );
and \U$4002 ( \13097 , RIdeb00f0_467, \9081 );
and \U$4003 ( \13098 , RIfc5ff60_6114, \9083 );
and \U$4004 ( \13099 , RIdead3f0_435, \9085 );
and \U$4005 ( \13100 , RIdea6c58_403, \9087 );
and \U$4006 ( \13101 , RIdea0358_371, \9089 );
and \U$4007 ( \13102 , RIfce5070_7628, \9091 );
and \U$4008 ( \13103 , RIee1c6d8_4782, \9093 );
and \U$4009 ( \13104 , RIfce70c8_7651, \9095 );
and \U$4010 ( \13105 , RIee1b058_4766, \9097 );
and \U$4011 ( \13106 , RIde934a0_308, \9099 );
and \U$4012 ( \13107 , RIfe9b1d8_8109, \9101 );
and \U$4013 ( \13108 , RIde8b7f0_270, \9103 );
and \U$4014 ( \13109 , RIfe9b340_8110, \9105 );
and \U$4015 ( \13110 , RIfc6b798_6245, \9107 );
and \U$4016 ( \13111 , RIfcb2238_7049, \9109 );
and \U$4017 ( \13112 , RIfcd3a00_7430, \9111 );
and \U$4018 ( \13113 , RIfcdb020_7514, \9113 );
and \U$4019 ( \13114 , RIfc511b8_5945, \9115 );
and \U$4020 ( \13115 , RIe16c9f8_2613, \9117 );
and \U$4021 ( \13116 , RIfcb27d8_7053, \9119 );
and \U$4022 ( \13117 , RIe168ee8_2571, \9121 );
and \U$4023 ( \13118 , RIe1668f0_2544, \9123 );
and \U$4024 ( \13119 , RIe163bf0_2512, \9125 );
and \U$4025 ( \13120 , RIee381d0_5097, \9127 );
and \U$4026 ( \13121 , RIe160ef0_2480, \9129 );
and \U$4027 ( \13122 , RIfcdfaa8_7567, \9131 );
and \U$4028 ( \13123 , RIe15e1f0_2448, \9133 );
and \U$4029 ( \13124 , RIe1587f0_2384, \9135 );
and \U$4030 ( \13125 , RIe155af0_2352, \9137 );
and \U$4031 ( \13126 , RIfc3f968_5749, \9139 );
and \U$4032 ( \13127 , RIe152df0_2320, \9141 );
and \U$4033 ( \13128 , RIfcd5080_7446, \9143 );
and \U$4034 ( \13129 , RIe1500f0_2288, \9145 );
and \U$4035 ( \13130 , RIfc84b30_6532, \9147 );
and \U$4036 ( \13131 , RIe14d3f0_2256, \9149 );
and \U$4037 ( \13132 , RIe14a6f0_2224, \9151 );
and \U$4038 ( \13133 , RIe1479f0_2192, \9153 );
and \U$4039 ( \13134 , RIfcea098_7685, \9155 );
and \U$4040 ( \13135 , RIfc92f00_6694, \9157 );
and \U$4041 ( \13136 , RIfc54890_5984, \9159 );
and \U$4042 ( \13137 , RIfcdcc40_7534, \9161 );
and \U$4043 ( \13138 , RIe142158_2129, \9163 );
and \U$4044 ( \13139 , RIe13fe30_2104, \9165 );
and \U$4045 ( \13140 , RIdf3dd38_2080, \9167 );
and \U$4046 ( \13141 , RIdf3b8a8_2054, \9169 );
and \U$4047 ( \13142 , RIfc57590_6016, \9171 );
and \U$4048 ( \13143 , RIee30340_5007, \9173 );
and \U$4049 ( \13144 , RIfcd0490_7392, \9175 );
and \U$4050 ( \13145 , RIee2e180_4983, \9177 );
and \U$4051 ( \13146 , RIdf36b50_1999, \9179 );
and \U$4052 ( \13147 , RIdf34558_1972, \9181 );
and \U$4053 ( \13148 , RIdf32398_1948, \9183 );
and \U$4054 ( \13149 , RIfe9b070_8108, \9185 );
or \U$4055 ( \13150 , \13086 , \13087 , \13088 , \13089 , \13090 , \13091 , \13092 , \13093 , \13094 , \13095 , \13096 , \13097 , \13098 , \13099 , \13100 , \13101 , \13102 , \13103 , \13104 , \13105 , \13106 , \13107 , \13108 , \13109 , \13110 , \13111 , \13112 , \13113 , \13114 , \13115 , \13116 , \13117 , \13118 , \13119 , \13120 , \13121 , \13122 , \13123 , \13124 , \13125 , \13126 , \13127 , \13128 , \13129 , \13130 , \13131 , \13132 , \13133 , \13134 , \13135 , \13136 , \13137 , \13138 , \13139 , \13140 , \13141 , \13142 , \13143 , \13144 , \13145 , \13146 , \13147 , \13148 , \13149 );
and \U$4056 ( \13151 , RIfcb1860_7042, \9188 );
and \U$4057 ( \13152 , RIfca1b40_6862, \9190 );
and \U$4058 ( \13153 , RIfc5c018_6069, \9192 );
and \U$4059 ( \13154 , RIfe9ada0_8106, \9194 );
and \U$4060 ( \13155 , RIdf2b318_1868, \9196 );
and \U$4061 ( \13156 , RIdf29428_1846, \9198 );
and \U$4062 ( \13157 , RIdf27100_1821, \9200 );
and \U$4063 ( \13158 , RIfe9af08_8107, \9202 );
and \U$4064 ( \13159 , RIfc5e1d8_6093, \9204 );
and \U$4065 ( \13160 , RIfcdcda8_7535, \9206 );
and \U$4066 ( \13161 , RIfcac400_6982, \9208 );
and \U$4067 ( \13162 , RIfc691a0_6218, \9210 );
and \U$4068 ( \13163 , RIfcaad80_6966, \9212 );
and \U$4069 ( \13164 , RIdf20bc0_1749, \9214 );
and \U$4070 ( \13165 , RIfc61b80_6134, \9216 );
and \U$4071 ( \13166 , RIdf1a518_1676, \9218 );
and \U$4072 ( \13167 , RIdf184c0_1653, \9220 );
and \U$4073 ( \13168 , RIdf157c0_1621, \9222 );
and \U$4074 ( \13169 , RIdf12ac0_1589, \9224 );
and \U$4075 ( \13170 , RIdf0fdc0_1557, \9226 );
and \U$4076 ( \13171 , RIdf0d0c0_1525, \9228 );
and \U$4077 ( \13172 , RIdf0a3c0_1493, \9230 );
and \U$4078 ( \13173 , RIdf076c0_1461, \9232 );
and \U$4079 ( \13174 , RIdf049c0_1429, \9234 );
and \U$4080 ( \13175 , RIdefefc0_1365, \9236 );
and \U$4081 ( \13176 , RIdefc2c0_1333, \9238 );
and \U$4082 ( \13177 , RIdef95c0_1301, \9240 );
and \U$4083 ( \13178 , RIdef68c0_1269, \9242 );
and \U$4084 ( \13179 , RIdef3bc0_1237, \9244 );
and \U$4085 ( \13180 , RIdef0ec0_1205, \9246 );
and \U$4086 ( \13181 , RIdeee1c0_1173, \9248 );
and \U$4087 ( \13182 , RIdeeb4c0_1141, \9250 );
and \U$4088 ( \13183 , RIfc69b78_6225, \9252 );
and \U$4089 ( \13184 , RIfc6b900_6246, \9254 );
and \U$4090 ( \13185 , RIfc4d270_5900, \9256 );
and \U$4091 ( \13186 , RIfced770_7724, \9258 );
and \U$4092 ( \13187 , RIdee5ac0_1077, \9260 );
and \U$4093 ( \13188 , RIdee3d38_1056, \9262 );
and \U$4094 ( \13189 , RIdee1a10_1031, \9264 );
and \U$4095 ( \13190 , RIdedfb20_1009, \9266 );
and \U$4096 ( \13191 , RIfc7ff40_6478, \9268 );
and \U$4097 ( \13192 , RIfca4408_6891, \9270 );
and \U$4098 ( \13193 , RIfcb5640_7086, \9272 );
and \U$4099 ( \13194 , RIee21700_4839, \9274 );
and \U$4100 ( \13195 , RIdeda990_951, \9276 );
and \U$4101 ( \13196 , RIded8500_925, \9278 );
and \U$4102 ( \13197 , RIded61d8_900, \9280 );
and \U$4103 ( \13198 , RIded4018_876, \9282 );
and \U$4104 ( \13199 , RIded1cf0_851, \9284 );
and \U$4105 ( \13200 , RIdeceff0_819, \9286 );
and \U$4106 ( \13201 , RIdecc2f0_787, \9288 );
and \U$4107 ( \13202 , RIdec95f0_755, \9290 );
and \U$4108 ( \13203 , RIdeb5af0_531, \9292 );
and \U$4109 ( \13204 , RIde99a58_339, \9294 );
and \U$4110 ( \13205 , RIe16f6f8_2645, \9296 );
and \U$4111 ( \13206 , RIe15b4f0_2416, \9298 );
and \U$4112 ( \13207 , RIe144cf0_2160, \9300 );
and \U$4113 ( \13208 , RIdf396e8_2030, \9302 );
and \U$4114 ( \13209 , RIdf2dd48_1898, \9304 );
and \U$4115 ( \13210 , RIdf1e5c8_1722, \9306 );
and \U$4116 ( \13211 , RIdf01cc0_1397, \9308 );
and \U$4117 ( \13212 , RIdee87c0_1109, \9310 );
and \U$4118 ( \13213 , RIdedd528_982, \9312 );
and \U$4119 ( \13214 , RIde7f9a0_212, \9314 );
or \U$4120 ( \13215 , \13151 , \13152 , \13153 , \13154 , \13155 , \13156 , \13157 , \13158 , \13159 , \13160 , \13161 , \13162 , \13163 , \13164 , \13165 , \13166 , \13167 , \13168 , \13169 , \13170 , \13171 , \13172 , \13173 , \13174 , \13175 , \13176 , \13177 , \13178 , \13179 , \13180 , \13181 , \13182 , \13183 , \13184 , \13185 , \13186 , \13187 , \13188 , \13189 , \13190 , \13191 , \13192 , \13193 , \13194 , \13195 , \13196 , \13197 , \13198 , \13199 , \13200 , \13201 , \13202 , \13203 , \13204 , \13205 , \13206 , \13207 , \13208 , \13209 , \13210 , \13211 , \13212 , \13213 , \13214 );
or \U$4121 ( \13216 , \13150 , \13215 );
_DC g2f32 ( \13217_nG2f32 , \13216 , \9323 );
buf \U$4122 ( \13218 , \13217_nG2f32 );
and \U$4123 ( \13219 , RIe19eb88_3183, \9333 );
and \U$4124 ( \13220 , RIe19be88_3151, \9335 );
and \U$4125 ( \13221 , RIfe9a698_8101, \9337 );
and \U$4126 ( \13222 , RIe199188_3119, \9339 );
and \U$4127 ( \13223 , RIfe9a530_8100, \9341 );
and \U$4128 ( \13224 , RIe196488_3087, \9343 );
and \U$4129 ( \13225 , RIe193788_3055, \9345 );
and \U$4130 ( \13226 , RIe190a88_3023, \9347 );
and \U$4131 ( \13227 , RIe18b088_2959, \9349 );
and \U$4132 ( \13228 , RIe188388_2927, \9351 );
and \U$4133 ( \13229 , RIfe9a800_8102, \9353 );
and \U$4134 ( \13230 , RIe185688_2895, \9355 );
and \U$4135 ( \13231 , RIfc8d938_6633, \9357 );
and \U$4136 ( \13232 , RIe182988_2863, \9359 );
and \U$4137 ( \13233 , RIe17fc88_2831, \9361 );
and \U$4138 ( \13234 , RIe17cf88_2799, \9363 );
and \U$4139 ( \13235 , RIfe9a3c8_8099, \9365 );
and \U$4140 ( \13236 , RIf1415a8_5203, \9367 );
and \U$4141 ( \13237 , RIfe9a260_8098, \9369 );
and \U$4142 ( \13238 , RIfe9a0f8_8097, \9371 );
and \U$4143 ( \13239 , RIfcb9150_7128, \9373 );
and \U$4144 ( \13240 , RIf13f820_5182, \9375 );
and \U$4145 ( \13241 , RIfc9fc50_6840, \9377 );
and \U$4146 ( \13242 , RIfce5340_7630, \9379 );
and \U$4147 ( \13243 , RIfc5cb58_6077, \9381 );
and \U$4148 ( \13244 , RIfc576f8_6017, \9383 );
and \U$4149 ( \13245 , RIfc780b0_6388, \9385 );
and \U$4150 ( \13246 , RIe1749f0_2704, \9387 );
and \U$4151 ( \13247 , RIfc7adb0_6420, \9389 );
and \U$4152 ( \13248 , RIfc7c2c8_6435, \9391 );
and \U$4153 ( \13249 , RIfcb2d78_7057, \9393 );
and \U$4154 ( \13250 , RIfc7e758_6461, \9395 );
and \U$4155 ( \13251 , RIfe9aad0_8104, \9397 );
and \U$4156 ( \13252 , RIe224ee0_4710, \9399 );
and \U$4157 ( \13253 , RIf16c3e8_5691, \9401 );
and \U$4158 ( \13254 , RIe2221e0_4678, \9403 );
and \U$4159 ( \13255 , RIfcd3898_7429, \9405 );
and \U$4160 ( \13256 , RIe21f4e0_4646, \9407 );
and \U$4161 ( \13257 , RIe219ae0_4582, \9409 );
and \U$4162 ( \13258 , RIe216de0_4550, \9411 );
and \U$4163 ( \13259 , RIfc880a0_6570, \9413 );
and \U$4164 ( \13260 , RIe2140e0_4518, \9415 );
and \U$4165 ( \13261 , RIf169c88_5663, \9417 );
and \U$4166 ( \13262 , RIe2113e0_4486, \9419 );
and \U$4167 ( \13263 , RIf168338_5645, \9421 );
and \U$4168 ( \13264 , RIe20e6e0_4454, \9423 );
and \U$4169 ( \13265 , RIe20b9e0_4422, \9425 );
and \U$4170 ( \13266 , RIe208ce0_4390, \9427 );
and \U$4171 ( \13267 , RIfce4c38_7625, \9429 );
and \U$4172 ( \13268 , RIfc9c6e0_6802, \9431 );
and \U$4173 ( \13269 , RIe2035b0_4328, \9433 );
and \U$4174 ( \13270 , RIe201af8_4309, \9435 );
and \U$4175 ( \13271 , RIfc500d8_5933, \9437 );
and \U$4176 ( \13272 , RIfc85c10_6544, \9439 );
and \U$4177 ( \13273 , RIfce81a8_7663, \9441 );
and \U$4178 ( \13274 , RIfce9c60_7682, \9443 );
and \U$4179 ( \13275 , RIf160e80_5562, \9445 );
and \U$4180 ( \13276 , RIf15ef90_5540, \9447 );
and \U$4181 ( \13277 , RIfe9a968_8103, \9449 );
and \U$4182 ( \13278 , RIfe9ac38_8105, \9451 );
and \U$4183 ( \13279 , RIfca8d28_6943, \9453 );
and \U$4184 ( \13280 , RIf15be58_5505, \9455 );
and \U$4185 ( \13281 , RIfcedba8_7727, \9457 );
and \U$4186 ( \13282 , RIfc6a988_6235, \9459 );
or \U$4187 ( \13283 , \13219 , \13220 , \13221 , \13222 , \13223 , \13224 , \13225 , \13226 , \13227 , \13228 , \13229 , \13230 , \13231 , \13232 , \13233 , \13234 , \13235 , \13236 , \13237 , \13238 , \13239 , \13240 , \13241 , \13242 , \13243 , \13244 , \13245 , \13246 , \13247 , \13248 , \13249 , \13250 , \13251 , \13252 , \13253 , \13254 , \13255 , \13256 , \13257 , \13258 , \13259 , \13260 , \13261 , \13262 , \13263 , \13264 , \13265 , \13266 , \13267 , \13268 , \13269 , \13270 , \13271 , \13272 , \13273 , \13274 , \13275 , \13276 , \13277 , \13278 , \13279 , \13280 , \13281 , \13282 );
and \U$4188 ( \13284 , RIfc71cd8_6317, \9462 );
and \U$4189 ( \13285 , RIfccb198_7333, \9464 );
and \U$4190 ( \13286 , RIfcaa3a8_6959, \9466 );
and \U$4191 ( \13287 , RIfec3b88_8347, \9468 );
and \U$4192 ( \13288 , RIfc4c730_5892, \9470 );
and \U$4193 ( \13289 , RIfc6d688_6267, \9472 );
and \U$4194 ( \13290 , RIfca8e90_6944, \9474 );
and \U$4195 ( \13291 , RIe1f6860_4182, \9476 );
and \U$4196 ( \13292 , RIfc64e20_6170, \9478 );
and \U$4197 ( \13293 , RIfcaee30_7012, \9480 );
and \U$4198 ( \13294 , RIfccee10_7376, \9482 );
and \U$4199 ( \13295 , RIe1f4538_4157, \9484 );
and \U$4200 ( \13296 , RIfc63ea8_6159, \9486 );
and \U$4201 ( \13297 , RIfcaecc8_7011, \9488 );
and \U$4202 ( \13298 , RIfcae458_7005, \9490 );
and \U$4203 ( \13299 , RIfeab1c8_8263, \9492 );
and \U$4204 ( \13300 , RIe1ecc48_4071, \9494 );
and \U$4205 ( \13301 , RIe1e9f48_4039, \9496 );
and \U$4206 ( \13302 , RIe1e7248_4007, \9498 );
and \U$4207 ( \13303 , RIe1e4548_3975, \9500 );
and \U$4208 ( \13304 , RIe1e1848_3943, \9502 );
and \U$4209 ( \13305 , RIe1deb48_3911, \9504 );
and \U$4210 ( \13306 , RIe1dbe48_3879, \9506 );
and \U$4211 ( \13307 , RIe1d9148_3847, \9508 );
and \U$4212 ( \13308 , RIe1d3748_3783, \9510 );
and \U$4213 ( \13309 , RIe1d0a48_3751, \9512 );
and \U$4214 ( \13310 , RIe1cdd48_3719, \9514 );
and \U$4215 ( \13311 , RIe1cb048_3687, \9516 );
and \U$4216 ( \13312 , RIe1c8348_3655, \9518 );
and \U$4217 ( \13313 , RIe1c5648_3623, \9520 );
and \U$4218 ( \13314 , RIe1c2948_3591, \9522 );
and \U$4219 ( \13315 , RIe1bfc48_3559, \9524 );
and \U$4220 ( \13316 , RIfcc70e8_7287, \9526 );
and \U$4221 ( \13317 , RIfca7ae0_6930, \9528 );
and \U$4222 ( \13318 , RIe1ba518_3497, \9530 );
and \U$4223 ( \13319 , RIe1b8358_3473, \9532 );
and \U$4224 ( \13320 , RIfc598b8_6041, \9534 );
and \U$4225 ( \13321 , RIfcc2228_7231, \9536 );
and \U$4226 ( \13322 , RIe1b6198_3449, \9538 );
and \U$4227 ( \13323 , RIe1b4848_3431, \9540 );
and \U$4228 ( \13324 , RIfc82f10_6512, \9542 );
and \U$4229 ( \13325 , RIfc55970_5996, \9544 );
and \U$4230 ( \13326 , RIe1b3498_3417, \9546 );
and \U$4231 ( \13327 , RIe1b1cb0_3400, \9548 );
and \U$4232 ( \13328 , RIfcb7698_7109, \9550 );
and \U$4233 ( \13329 , RIfc4b4e8_5879, \9552 );
and \U$4234 ( \13330 , RIe1ad390_3348, \9554 );
and \U$4235 ( \13331 , RIe1abba8_3331, \9556 );
and \U$4236 ( \13332 , RIe1a9f88_3311, \9558 );
and \U$4237 ( \13333 , RIe1a7288_3279, \9560 );
and \U$4238 ( \13334 , RIe1a4588_3247, \9562 );
and \U$4239 ( \13335 , RIe1a1888_3215, \9564 );
and \U$4240 ( \13336 , RIe18dd88_2991, \9566 );
and \U$4241 ( \13337 , RIe17a288_2767, \9568 );
and \U$4242 ( \13338 , RIe227be0_4742, \9570 );
and \U$4243 ( \13339 , RIe21c7e0_4614, \9572 );
and \U$4244 ( \13340 , RIe205fe0_4358, \9574 );
and \U$4245 ( \13341 , RIe200040_4290, \9576 );
and \U$4246 ( \13342 , RIe1f93f8_4213, \9578 );
and \U$4247 ( \13343 , RIe1f1f40_4130, \9580 );
and \U$4248 ( \13344 , RIe1d6448_3815, \9582 );
and \U$4249 ( \13345 , RIe1bcf48_3527, \9584 );
and \U$4250 ( \13346 , RIe1afdc0_3378, \9586 );
and \U$4251 ( \13347 , RIe1723f8_2677, \9588 );
or \U$4252 ( \13348 , \13284 , \13285 , \13286 , \13287 , \13288 , \13289 , \13290 , \13291 , \13292 , \13293 , \13294 , \13295 , \13296 , \13297 , \13298 , \13299 , \13300 , \13301 , \13302 , \13303 , \13304 , \13305 , \13306 , \13307 , \13308 , \13309 , \13310 , \13311 , \13312 , \13313 , \13314 , \13315 , \13316 , \13317 , \13318 , \13319 , \13320 , \13321 , \13322 , \13323 , \13324 , \13325 , \13326 , \13327 , \13328 , \13329 , \13330 , \13331 , \13332 , \13333 , \13334 , \13335 , \13336 , \13337 , \13338 , \13339 , \13340 , \13341 , \13342 , \13343 , \13344 , \13345 , \13346 , \13347 );
or \U$4253 ( \13349 , \13283 , \13348 );
_DC g405f ( \13350_nG405f , \13349 , \9597 );
buf \U$4254 ( \13351 , \13350_nG405f );
and \U$4255 ( \13352 , \13218 , \13351 );
and \U$4256 ( \13353 , \11738 , \11871 );
and \U$4257 ( \13354 , \11871 , \12146 );
and \U$4258 ( \13355 , \11738 , \12146 );
or \U$4259 ( \13356 , \13353 , \13354 , \13355 );
and \U$4260 ( \13357 , \13351 , \13356 );
and \U$4261 ( \13358 , \13218 , \13356 );
or \U$4262 ( \13359 , \13352 , \13357 , \13358 );
xor \U$4263 ( \13360 , \13085 , \13359 );
buf g4442 ( \13361_nG4442 , \13360 );
xor \U$4264 ( \13362 , \13218 , \13351 );
xor \U$4265 ( \13363 , \13362 , \13356 );
buf g4445 ( \13364_nG4445 , \13363 );
nand \U$4266 ( \13365 , \13364_nG4445 , \12148_nG4448 );
and \U$4267 ( \13366 , \13361_nG4442 , \13365 );
xor \U$4268 ( \13367 , \13364_nG4445 , \12148_nG4448 );
not \U$4269 ( \13368 , \13367 );
xor \U$4270 ( \13369 , \13361_nG4442 , \13364_nG4445 );
and \U$4271 ( \13370 , \13368 , \13369 );
and \U$4273 ( \13371 , \13367 , \10694_nG9c0e );
or \U$4274 ( \13372 , 1'b0 , \13371 );
xor \U$4275 ( \13373 , \13366 , \13372 );
xor \U$4276 ( \13374 , \13366 , \13373 );
buf \U$4277 ( \13375 , \13374 );
buf \U$4278 ( \13376 , \13375 );
and \U$4279 ( \13377 , \12818 , \13376 );
and \U$4280 ( \13378 , \12808 , \12813 );
and \U$4281 ( \13379 , \12808 , \12816 );
and \U$4282 ( \13380 , \12813 , \12816 );
or \U$4283 ( \13381 , \13378 , \13379 , \13380 );
buf \U$4284 ( \13382 , \13381 );
and \U$4285 ( \13383 , \12490 , \12496 );
and \U$4286 ( \13384 , \12490 , \12806 );
and \U$4287 ( \13385 , \12496 , \12806 );
or \U$4288 ( \13386 , \13383 , \13384 , \13385 );
buf \U$4289 ( \13387 , \13386 );
xor \U$4290 ( \13388 , \13382 , \13387 );
and \U$4291 ( \13389 , \12482 , \12488 );
buf \U$4292 ( \13390 , \13389 );
and \U$4293 ( \13391 , \12157 , \10995_nG9c0b );
and \U$4294 ( \13392 , \12154 , \11283_nG9c08 );
or \U$4295 ( \13393 , \13391 , \13392 );
xor \U$4296 ( \13394 , \12153 , \13393 );
buf \U$4297 ( \13395 , \13394 );
buf \U$4299 ( \13396 , \13395 );
xor \U$4300 ( \13397 , \13390 , \13396 );
buf \U$4301 ( \13398 , \13397 );
and \U$4302 ( \13399 , \10421 , \11598_nG9c05 );
and \U$4303 ( \13400 , \10418 , \12470_nG9c02 );
or \U$4304 ( \13401 , \13399 , \13400 );
xor \U$4305 ( \13402 , \10417 , \13401 );
buf \U$4306 ( \13403 , \13402 );
buf \U$4308 ( \13404 , \13403 );
xor \U$4309 ( \13405 , \13398 , \13404 );
and \U$4310 ( \13406 , \10707 , \12801_nG9bff );
and \U$4311 ( \13407 , \12772 , \12781 );
and \U$4312 ( \13408 , \10988 , \12790 );
and \U$4313 ( \13409 , \11270 , \12461 );
nor \U$4314 ( \13410 , \13408 , \13409 );
xnor \U$4315 ( \13411 , \13410 , \12780 );
xor \U$4316 ( \13412 , \13407 , \13411 );
and \U$4317 ( \13413 , \12769 , \10983 );
and \U$4318 ( \13414 , RIdec68f0_723, \9333 );
and \U$4319 ( \13415 , RIdec3bf0_691, \9335 );
and \U$4320 ( \13416 , RIee208f0_4829, \9337 );
and \U$4321 ( \13417 , RIdec0ef0_659, \9339 );
and \U$4322 ( \13418 , RIfc7ce08_6443, \9341 );
and \U$4323 ( \13419 , RIdebe1f0_627, \9343 );
and \U$4324 ( \13420 , RIdebb4f0_595, \9345 );
and \U$4325 ( \13421 , RIdeb87f0_563, \9347 );
and \U$4326 ( \13422 , RIfc9b8d0_6792, \9349 );
and \U$4327 ( \13423 , RIdeb2df0_499, \9351 );
and \U$4328 ( \13424 , RIfcc6710_7280, \9353 );
and \U$4329 ( \13425 , RIdeb00f0_467, \9355 );
and \U$4330 ( \13426 , RIfc5ff60_6114, \9357 );
and \U$4331 ( \13427 , RIdead3f0_435, \9359 );
and \U$4332 ( \13428 , RIdea6c58_403, \9361 );
and \U$4333 ( \13429 , RIdea0358_371, \9363 );
and \U$4334 ( \13430 , RIfce5070_7628, \9365 );
and \U$4335 ( \13431 , RIee1c6d8_4782, \9367 );
and \U$4336 ( \13432 , RIfce70c8_7651, \9369 );
and \U$4337 ( \13433 , RIee1b058_4766, \9371 );
and \U$4338 ( \13434 , RIde934a0_308, \9373 );
and \U$4339 ( \13435 , RIfe9b1d8_8109, \9375 );
and \U$4340 ( \13436 , RIde8b7f0_270, \9377 );
and \U$4341 ( \13437 , RIfe9b340_8110, \9379 );
and \U$4342 ( \13438 , RIfc6b798_6245, \9381 );
and \U$4343 ( \13439 , RIfcb2238_7049, \9383 );
and \U$4344 ( \13440 , RIfcd3a00_7430, \9385 );
and \U$4345 ( \13441 , RIfcdb020_7514, \9387 );
and \U$4346 ( \13442 , RIfc511b8_5945, \9389 );
and \U$4347 ( \13443 , RIe16c9f8_2613, \9391 );
and \U$4348 ( \13444 , RIfcb27d8_7053, \9393 );
and \U$4349 ( \13445 , RIe168ee8_2571, \9395 );
and \U$4350 ( \13446 , RIe1668f0_2544, \9397 );
and \U$4351 ( \13447 , RIe163bf0_2512, \9399 );
and \U$4352 ( \13448 , RIee381d0_5097, \9401 );
and \U$4353 ( \13449 , RIe160ef0_2480, \9403 );
and \U$4354 ( \13450 , RIfcdfaa8_7567, \9405 );
and \U$4355 ( \13451 , RIe15e1f0_2448, \9407 );
and \U$4356 ( \13452 , RIe1587f0_2384, \9409 );
and \U$4357 ( \13453 , RIe155af0_2352, \9411 );
and \U$4358 ( \13454 , RIfc3f968_5749, \9413 );
and \U$4359 ( \13455 , RIe152df0_2320, \9415 );
and \U$4360 ( \13456 , RIfcd5080_7446, \9417 );
and \U$4361 ( \13457 , RIe1500f0_2288, \9419 );
and \U$4362 ( \13458 , RIfc84b30_6532, \9421 );
and \U$4363 ( \13459 , RIe14d3f0_2256, \9423 );
and \U$4364 ( \13460 , RIe14a6f0_2224, \9425 );
and \U$4365 ( \13461 , RIe1479f0_2192, \9427 );
and \U$4366 ( \13462 , RIfcea098_7685, \9429 );
and \U$4367 ( \13463 , RIfc92f00_6694, \9431 );
and \U$4368 ( \13464 , RIfc54890_5984, \9433 );
and \U$4369 ( \13465 , RIfcdcc40_7534, \9435 );
and \U$4370 ( \13466 , RIe142158_2129, \9437 );
and \U$4371 ( \13467 , RIe13fe30_2104, \9439 );
and \U$4372 ( \13468 , RIdf3dd38_2080, \9441 );
and \U$4373 ( \13469 , RIdf3b8a8_2054, \9443 );
and \U$4374 ( \13470 , RIfc57590_6016, \9445 );
and \U$4375 ( \13471 , RIee30340_5007, \9447 );
and \U$4376 ( \13472 , RIfcd0490_7392, \9449 );
and \U$4377 ( \13473 , RIee2e180_4983, \9451 );
and \U$4378 ( \13474 , RIdf36b50_1999, \9453 );
and \U$4379 ( \13475 , RIdf34558_1972, \9455 );
and \U$4380 ( \13476 , RIdf32398_1948, \9457 );
and \U$4381 ( \13477 , RIfe9b070_8108, \9459 );
or \U$4382 ( \13478 , \13414 , \13415 , \13416 , \13417 , \13418 , \13419 , \13420 , \13421 , \13422 , \13423 , \13424 , \13425 , \13426 , \13427 , \13428 , \13429 , \13430 , \13431 , \13432 , \13433 , \13434 , \13435 , \13436 , \13437 , \13438 , \13439 , \13440 , \13441 , \13442 , \13443 , \13444 , \13445 , \13446 , \13447 , \13448 , \13449 , \13450 , \13451 , \13452 , \13453 , \13454 , \13455 , \13456 , \13457 , \13458 , \13459 , \13460 , \13461 , \13462 , \13463 , \13464 , \13465 , \13466 , \13467 , \13468 , \13469 , \13470 , \13471 , \13472 , \13473 , \13474 , \13475 , \13476 , \13477 );
and \U$4383 ( \13479 , RIfcb1860_7042, \9462 );
and \U$4384 ( \13480 , RIfca1b40_6862, \9464 );
and \U$4385 ( \13481 , RIfc5c018_6069, \9466 );
and \U$4386 ( \13482 , RIfe9ada0_8106, \9468 );
and \U$4387 ( \13483 , RIdf2b318_1868, \9470 );
and \U$4388 ( \13484 , RIdf29428_1846, \9472 );
and \U$4389 ( \13485 , RIdf27100_1821, \9474 );
and \U$4390 ( \13486 , RIfe9af08_8107, \9476 );
and \U$4391 ( \13487 , RIfc5e1d8_6093, \9478 );
and \U$4392 ( \13488 , RIfcdcda8_7535, \9480 );
and \U$4393 ( \13489 , RIfcac400_6982, \9482 );
and \U$4394 ( \13490 , RIfc691a0_6218, \9484 );
and \U$4395 ( \13491 , RIfcaad80_6966, \9486 );
and \U$4396 ( \13492 , RIdf20bc0_1749, \9488 );
and \U$4397 ( \13493 , RIfc61b80_6134, \9490 );
and \U$4398 ( \13494 , RIdf1a518_1676, \9492 );
and \U$4399 ( \13495 , RIdf184c0_1653, \9494 );
and \U$4400 ( \13496 , RIdf157c0_1621, \9496 );
and \U$4401 ( \13497 , RIdf12ac0_1589, \9498 );
and \U$4402 ( \13498 , RIdf0fdc0_1557, \9500 );
and \U$4403 ( \13499 , RIdf0d0c0_1525, \9502 );
and \U$4404 ( \13500 , RIdf0a3c0_1493, \9504 );
and \U$4405 ( \13501 , RIdf076c0_1461, \9506 );
and \U$4406 ( \13502 , RIdf049c0_1429, \9508 );
and \U$4407 ( \13503 , RIdefefc0_1365, \9510 );
and \U$4408 ( \13504 , RIdefc2c0_1333, \9512 );
and \U$4409 ( \13505 , RIdef95c0_1301, \9514 );
and \U$4410 ( \13506 , RIdef68c0_1269, \9516 );
and \U$4411 ( \13507 , RIdef3bc0_1237, \9518 );
and \U$4412 ( \13508 , RIdef0ec0_1205, \9520 );
and \U$4413 ( \13509 , RIdeee1c0_1173, \9522 );
and \U$4414 ( \13510 , RIdeeb4c0_1141, \9524 );
and \U$4415 ( \13511 , RIfc69b78_6225, \9526 );
and \U$4416 ( \13512 , RIfc6b900_6246, \9528 );
and \U$4417 ( \13513 , RIfc4d270_5900, \9530 );
and \U$4418 ( \13514 , RIfced770_7724, \9532 );
and \U$4419 ( \13515 , RIdee5ac0_1077, \9534 );
and \U$4420 ( \13516 , RIdee3d38_1056, \9536 );
and \U$4421 ( \13517 , RIdee1a10_1031, \9538 );
and \U$4422 ( \13518 , RIdedfb20_1009, \9540 );
and \U$4423 ( \13519 , RIfc7ff40_6478, \9542 );
and \U$4424 ( \13520 , RIfca4408_6891, \9544 );
and \U$4425 ( \13521 , RIfcb5640_7086, \9546 );
and \U$4426 ( \13522 , RIee21700_4839, \9548 );
and \U$4427 ( \13523 , RIdeda990_951, \9550 );
and \U$4428 ( \13524 , RIded8500_925, \9552 );
and \U$4429 ( \13525 , RIded61d8_900, \9554 );
and \U$4430 ( \13526 , RIded4018_876, \9556 );
and \U$4431 ( \13527 , RIded1cf0_851, \9558 );
and \U$4432 ( \13528 , RIdeceff0_819, \9560 );
and \U$4433 ( \13529 , RIdecc2f0_787, \9562 );
and \U$4434 ( \13530 , RIdec95f0_755, \9564 );
and \U$4435 ( \13531 , RIdeb5af0_531, \9566 );
and \U$4436 ( \13532 , RIde99a58_339, \9568 );
and \U$4437 ( \13533 , RIe16f6f8_2645, \9570 );
and \U$4438 ( \13534 , RIe15b4f0_2416, \9572 );
and \U$4439 ( \13535 , RIe144cf0_2160, \9574 );
and \U$4440 ( \13536 , RIdf396e8_2030, \9576 );
and \U$4441 ( \13537 , RIdf2dd48_1898, \9578 );
and \U$4442 ( \13538 , RIdf1e5c8_1722, \9580 );
and \U$4443 ( \13539 , RIdf01cc0_1397, \9582 );
and \U$4444 ( \13540 , RIdee87c0_1109, \9584 );
and \U$4445 ( \13541 , RIdedd528_982, \9586 );
and \U$4446 ( \13542 , RIde7f9a0_212, \9588 );
or \U$4447 ( \13543 , \13479 , \13480 , \13481 , \13482 , \13483 , \13484 , \13485 , \13486 , \13487 , \13488 , \13489 , \13490 , \13491 , \13492 , \13493 , \13494 , \13495 , \13496 , \13497 , \13498 , \13499 , \13500 , \13501 , \13502 , \13503 , \13504 , \13505 , \13506 , \13507 , \13508 , \13509 , \13510 , \13511 , \13512 , \13513 , \13514 , \13515 , \13516 , \13517 , \13518 , \13519 , \13520 , \13521 , \13522 , \13523 , \13524 , \13525 , \13526 , \13527 , \13528 , \13529 , \13530 , \13531 , \13532 , \13533 , \13534 , \13535 , \13536 , \13537 , \13538 , \13539 , \13540 , \13541 , \13542 );
or \U$4448 ( \13544 , \13478 , \13543 );
_DC g6589 ( \13545_nG6589 , \13544 , \9597 );
and \U$4449 ( \13546 , RIe19eb88_3183, \9059 );
and \U$4450 ( \13547 , RIe19be88_3151, \9061 );
and \U$4451 ( \13548 , RIfe9a698_8101, \9063 );
and \U$4452 ( \13549 , RIe199188_3119, \9065 );
and \U$4453 ( \13550 , RIfe9a530_8100, \9067 );
and \U$4454 ( \13551 , RIe196488_3087, \9069 );
and \U$4455 ( \13552 , RIe193788_3055, \9071 );
and \U$4456 ( \13553 , RIe190a88_3023, \9073 );
and \U$4457 ( \13554 , RIe18b088_2959, \9075 );
and \U$4458 ( \13555 , RIe188388_2927, \9077 );
and \U$4459 ( \13556 , RIfe9a800_8102, \9079 );
and \U$4460 ( \13557 , RIe185688_2895, \9081 );
and \U$4461 ( \13558 , RIfc8d938_6633, \9083 );
and \U$4462 ( \13559 , RIe182988_2863, \9085 );
and \U$4463 ( \13560 , RIe17fc88_2831, \9087 );
and \U$4464 ( \13561 , RIe17cf88_2799, \9089 );
and \U$4465 ( \13562 , RIfe9a3c8_8099, \9091 );
and \U$4466 ( \13563 , RIf1415a8_5203, \9093 );
and \U$4467 ( \13564 , RIfe9a260_8098, \9095 );
and \U$4468 ( \13565 , RIfe9a0f8_8097, \9097 );
and \U$4469 ( \13566 , RIfcb9150_7128, \9099 );
and \U$4470 ( \13567 , RIf13f820_5182, \9101 );
and \U$4471 ( \13568 , RIfc9fc50_6840, \9103 );
and \U$4472 ( \13569 , RIfce5340_7630, \9105 );
and \U$4473 ( \13570 , RIfc5cb58_6077, \9107 );
and \U$4474 ( \13571 , RIfc576f8_6017, \9109 );
and \U$4475 ( \13572 , RIfc780b0_6388, \9111 );
and \U$4476 ( \13573 , RIe1749f0_2704, \9113 );
and \U$4477 ( \13574 , RIfc7adb0_6420, \9115 );
and \U$4478 ( \13575 , RIfc7c2c8_6435, \9117 );
and \U$4479 ( \13576 , RIfcb2d78_7057, \9119 );
and \U$4480 ( \13577 , RIfc7e758_6461, \9121 );
and \U$4481 ( \13578 , RIfe9aad0_8104, \9123 );
and \U$4482 ( \13579 , RIe224ee0_4710, \9125 );
and \U$4483 ( \13580 , RIf16c3e8_5691, \9127 );
and \U$4484 ( \13581 , RIe2221e0_4678, \9129 );
and \U$4485 ( \13582 , RIfcd3898_7429, \9131 );
and \U$4486 ( \13583 , RIe21f4e0_4646, \9133 );
and \U$4487 ( \13584 , RIe219ae0_4582, \9135 );
and \U$4488 ( \13585 , RIe216de0_4550, \9137 );
and \U$4489 ( \13586 , RIfc880a0_6570, \9139 );
and \U$4490 ( \13587 , RIe2140e0_4518, \9141 );
and \U$4491 ( \13588 , RIf169c88_5663, \9143 );
and \U$4492 ( \13589 , RIe2113e0_4486, \9145 );
and \U$4493 ( \13590 , RIf168338_5645, \9147 );
and \U$4494 ( \13591 , RIe20e6e0_4454, \9149 );
and \U$4495 ( \13592 , RIe20b9e0_4422, \9151 );
and \U$4496 ( \13593 , RIe208ce0_4390, \9153 );
and \U$4497 ( \13594 , RIfce4c38_7625, \9155 );
and \U$4498 ( \13595 , RIfc9c6e0_6802, \9157 );
and \U$4499 ( \13596 , RIe2035b0_4328, \9159 );
and \U$4500 ( \13597 , RIe201af8_4309, \9161 );
and \U$4501 ( \13598 , RIfc500d8_5933, \9163 );
and \U$4502 ( \13599 , RIfc85c10_6544, \9165 );
and \U$4503 ( \13600 , RIfce81a8_7663, \9167 );
and \U$4504 ( \13601 , RIfce9c60_7682, \9169 );
and \U$4505 ( \13602 , RIf160e80_5562, \9171 );
and \U$4506 ( \13603 , RIf15ef90_5540, \9173 );
and \U$4507 ( \13604 , RIfe9a968_8103, \9175 );
and \U$4508 ( \13605 , RIfe9ac38_8105, \9177 );
and \U$4509 ( \13606 , RIfca8d28_6943, \9179 );
and \U$4510 ( \13607 , RIf15be58_5505, \9181 );
and \U$4511 ( \13608 , RIfcedba8_7727, \9183 );
and \U$4512 ( \13609 , RIfc6a988_6235, \9185 );
or \U$4513 ( \13610 , \13546 , \13547 , \13548 , \13549 , \13550 , \13551 , \13552 , \13553 , \13554 , \13555 , \13556 , \13557 , \13558 , \13559 , \13560 , \13561 , \13562 , \13563 , \13564 , \13565 , \13566 , \13567 , \13568 , \13569 , \13570 , \13571 , \13572 , \13573 , \13574 , \13575 , \13576 , \13577 , \13578 , \13579 , \13580 , \13581 , \13582 , \13583 , \13584 , \13585 , \13586 , \13587 , \13588 , \13589 , \13590 , \13591 , \13592 , \13593 , \13594 , \13595 , \13596 , \13597 , \13598 , \13599 , \13600 , \13601 , \13602 , \13603 , \13604 , \13605 , \13606 , \13607 , \13608 , \13609 );
and \U$4514 ( \13611 , RIfc71cd8_6317, \9188 );
and \U$4515 ( \13612 , RIfccb198_7333, \9190 );
and \U$4516 ( \13613 , RIfcaa3a8_6959, \9192 );
and \U$4517 ( \13614 , RIfec3b88_8347, \9194 );
and \U$4518 ( \13615 , RIfc4c730_5892, \9196 );
and \U$4519 ( \13616 , RIfc6d688_6267, \9198 );
and \U$4520 ( \13617 , RIfca8e90_6944, \9200 );
and \U$4521 ( \13618 , RIe1f6860_4182, \9202 );
and \U$4522 ( \13619 , RIfc64e20_6170, \9204 );
and \U$4523 ( \13620 , RIfcaee30_7012, \9206 );
and \U$4524 ( \13621 , RIfccee10_7376, \9208 );
and \U$4525 ( \13622 , RIe1f4538_4157, \9210 );
and \U$4526 ( \13623 , RIfc63ea8_6159, \9212 );
and \U$4527 ( \13624 , RIfcaecc8_7011, \9214 );
and \U$4528 ( \13625 , RIfcae458_7005, \9216 );
and \U$4529 ( \13626 , RIfeab1c8_8263, \9218 );
and \U$4530 ( \13627 , RIe1ecc48_4071, \9220 );
and \U$4531 ( \13628 , RIe1e9f48_4039, \9222 );
and \U$4532 ( \13629 , RIe1e7248_4007, \9224 );
and \U$4533 ( \13630 , RIe1e4548_3975, \9226 );
and \U$4534 ( \13631 , RIe1e1848_3943, \9228 );
and \U$4535 ( \13632 , RIe1deb48_3911, \9230 );
and \U$4536 ( \13633 , RIe1dbe48_3879, \9232 );
and \U$4537 ( \13634 , RIe1d9148_3847, \9234 );
and \U$4538 ( \13635 , RIe1d3748_3783, \9236 );
and \U$4539 ( \13636 , RIe1d0a48_3751, \9238 );
and \U$4540 ( \13637 , RIe1cdd48_3719, \9240 );
and \U$4541 ( \13638 , RIe1cb048_3687, \9242 );
and \U$4542 ( \13639 , RIe1c8348_3655, \9244 );
and \U$4543 ( \13640 , RIe1c5648_3623, \9246 );
and \U$4544 ( \13641 , RIe1c2948_3591, \9248 );
and \U$4545 ( \13642 , RIe1bfc48_3559, \9250 );
and \U$4546 ( \13643 , RIfcc70e8_7287, \9252 );
and \U$4547 ( \13644 , RIfca7ae0_6930, \9254 );
and \U$4548 ( \13645 , RIe1ba518_3497, \9256 );
and \U$4549 ( \13646 , RIe1b8358_3473, \9258 );
and \U$4550 ( \13647 , RIfc598b8_6041, \9260 );
and \U$4551 ( \13648 , RIfcc2228_7231, \9262 );
and \U$4552 ( \13649 , RIe1b6198_3449, \9264 );
and \U$4553 ( \13650 , RIe1b4848_3431, \9266 );
and \U$4554 ( \13651 , RIfc82f10_6512, \9268 );
and \U$4555 ( \13652 , RIfc55970_5996, \9270 );
and \U$4556 ( \13653 , RIe1b3498_3417, \9272 );
and \U$4557 ( \13654 , RIe1b1cb0_3400, \9274 );
and \U$4558 ( \13655 , RIfcb7698_7109, \9276 );
and \U$4559 ( \13656 , RIfc4b4e8_5879, \9278 );
and \U$4560 ( \13657 , RIe1ad390_3348, \9280 );
and \U$4561 ( \13658 , RIe1abba8_3331, \9282 );
and \U$4562 ( \13659 , RIe1a9f88_3311, \9284 );
and \U$4563 ( \13660 , RIe1a7288_3279, \9286 );
and \U$4564 ( \13661 , RIe1a4588_3247, \9288 );
and \U$4565 ( \13662 , RIe1a1888_3215, \9290 );
and \U$4566 ( \13663 , RIe18dd88_2991, \9292 );
and \U$4567 ( \13664 , RIe17a288_2767, \9294 );
and \U$4568 ( \13665 , RIe227be0_4742, \9296 );
and \U$4569 ( \13666 , RIe21c7e0_4614, \9298 );
and \U$4570 ( \13667 , RIe205fe0_4358, \9300 );
and \U$4571 ( \13668 , RIe200040_4290, \9302 );
and \U$4572 ( \13669 , RIe1f93f8_4213, \9304 );
and \U$4573 ( \13670 , RIe1f1f40_4130, \9306 );
and \U$4574 ( \13671 , RIe1d6448_3815, \9308 );
and \U$4575 ( \13672 , RIe1bcf48_3527, \9310 );
and \U$4576 ( \13673 , RIe1afdc0_3378, \9312 );
and \U$4577 ( \13674 , RIe1723f8_2677, \9314 );
or \U$4578 ( \13675 , \13611 , \13612 , \13613 , \13614 , \13615 , \13616 , \13617 , \13618 , \13619 , \13620 , \13621 , \13622 , \13623 , \13624 , \13625 , \13626 , \13627 , \13628 , \13629 , \13630 , \13631 , \13632 , \13633 , \13634 , \13635 , \13636 , \13637 , \13638 , \13639 , \13640 , \13641 , \13642 , \13643 , \13644 , \13645 , \13646 , \13647 , \13648 , \13649 , \13650 , \13651 , \13652 , \13653 , \13654 , \13655 , \13656 , \13657 , \13658 , \13659 , \13660 , \13661 , \13662 , \13663 , \13664 , \13665 , \13666 , \13667 , \13668 , \13669 , \13670 , \13671 , \13672 , \13673 , \13674 );
or \U$4579 ( \13676 , \13610 , \13675 );
_DC g658a ( \13677_nG658a , \13676 , \9323 );
and g658b ( \13678_nG658b , \13545_nG6589 , \13677_nG658a );
buf \U$4580 ( \13679 , \13678_nG658b );
and \U$4581 ( \13680 , \13679 , \10691 );
nor \U$4582 ( \13681 , \13413 , \13680 );
xnor \U$4583 ( \13682 , \13681 , \10980 );
and \U$4584 ( \13683 , \11586 , \11574 );
and \U$4585 ( \13684 , \12448 , \11278 );
nor \U$4586 ( \13685 , \13683 , \13684 );
xnor \U$4587 ( \13686 , \13685 , \11580 );
xor \U$4588 ( \13687 , \13682 , \13686 );
_DC g4b10 ( \13688_nG4b10 , \13544 , \9597 );
_DC g4b94 ( \13689_nG4b94 , \13676 , \9323 );
xor g4b95 ( \13690_nG4b95 , \13688_nG4b10 , \13689_nG4b94 );
buf \U$4589 ( \13691 , \13690_nG4b95 );
xor \U$4590 ( \13692 , \13691 , \12777 );
and \U$4591 ( \13693 , \10687 , \13692 );
xor \U$4592 ( \13694 , \13687 , \13693 );
xor \U$4593 ( \13695 , \13412 , \13694 );
and \U$4594 ( \13696 , \12782 , \12786 );
and \U$4595 ( \13697 , \12786 , \12794 );
and \U$4596 ( \13698 , \12782 , \12794 );
or \U$4597 ( \13699 , \13696 , \13697 , \13698 );
xor \U$4598 ( \13700 , \13695 , \13699 );
and \U$4599 ( \13701 , \12502 , \12795 );
and \U$4600 ( \13702 , \12796 , \12799 );
or \U$4601 ( \13703 , \13701 , \13702 );
xor \U$4602 ( \13704 , \13700 , \13703 );
buf g9bfc ( \13705_nG9bfc , \13704 );
and \U$4603 ( \13706 , \10704 , \13705_nG9bfc );
or \U$4604 ( \13707 , \13406 , \13706 );
xor \U$4605 ( \13708 , \10703 , \13707 );
buf \U$4606 ( \13709 , \13708 );
buf \U$4608 ( \13710 , \13709 );
xor \U$4609 ( \13711 , \13405 , \13710 );
buf \U$4610 ( \13712 , \13711 );
xor \U$4611 ( \13713 , \13388 , \13712 );
and \U$4612 ( \13714 , \12818 , \13713 );
and \U$4613 ( \13715 , \13376 , \13713 );
or \U$4614 ( \13716 , \13377 , \13714 , \13715 );
and \U$4615 ( \13717 , \13382 , \13387 );
and \U$4616 ( \13718 , \13382 , \13712 );
and \U$4617 ( \13719 , \13387 , \13712 );
or \U$4618 ( \13720 , \13717 , \13718 , \13719 );
buf \U$4619 ( \13721 , \13720 );
and \U$4620 ( \13722 , \13398 , \13404 );
and \U$4621 ( \13723 , \13398 , \13710 );
and \U$4622 ( \13724 , \13404 , \13710 );
or \U$4623 ( \13725 , \13722 , \13723 , \13724 );
buf \U$4624 ( \13726 , \13725 );
xor \U$4625 ( \13727 , \13721 , \13726 );
and \U$4626 ( \13728 , \13366 , \13373 );
buf \U$4627 ( \13729 , \13728 );
buf \U$4629 ( \13730 , \13729 );
and \U$4630 ( \13731 , \13370 , \10694_nG9c0e );
and \U$4631 ( \13732 , \13367 , \10995_nG9c0b );
or \U$4632 ( \13733 , \13731 , \13732 );
xor \U$4633 ( \13734 , \13366 , \13733 );
buf \U$4634 ( \13735 , \13734 );
buf \U$4636 ( \13736 , \13735 );
xor \U$4637 ( \13737 , \13730 , \13736 );
buf \U$4638 ( \13738 , \13737 );
and \U$4639 ( \13739 , \12157 , \11283_nG9c08 );
and \U$4640 ( \13740 , \12154 , \11598_nG9c05 );
or \U$4641 ( \13741 , \13739 , \13740 );
xor \U$4642 ( \13742 , \12153 , \13741 );
buf \U$4643 ( \13743 , \13742 );
buf \U$4645 ( \13744 , \13743 );
xor \U$4646 ( \13745 , \13738 , \13744 );
and \U$4647 ( \13746 , \10421 , \12470_nG9c02 );
and \U$4648 ( \13747 , \10418 , \12801_nG9bff );
or \U$4649 ( \13748 , \13746 , \13747 );
xor \U$4650 ( \13749 , \10417 , \13748 );
buf \U$4651 ( \13750 , \13749 );
buf \U$4653 ( \13751 , \13750 );
xor \U$4654 ( \13752 , \13745 , \13751 );
buf \U$4655 ( \13753 , \13752 );
and \U$4656 ( \13754 , \13390 , \13396 );
buf \U$4657 ( \13755 , \13754 );
xor \U$4658 ( \13756 , \13753 , \13755 );
and \U$4659 ( \13757 , \10707 , \13705_nG9bfc );
and \U$4660 ( \13758 , \13679 , \10983 );
and \U$4661 ( \13759 , RIdec6a58_724, \9333 );
and \U$4662 ( \13760 , RIdec3d58_692, \9335 );
and \U$4663 ( \13761 , RIfc723e0_6322, \9337 );
and \U$4664 ( \13762 , RIdec1058_660, \9339 );
and \U$4665 ( \13763 , RIfc59fc0_6046, \9341 );
and \U$4666 ( \13764 , RIdebe358_628, \9343 );
and \U$4667 ( \13765 , RIdebb658_596, \9345 );
and \U$4668 ( \13766 , RIdeb8958_564, \9347 );
and \U$4669 ( \13767 , RIfcb96f0_7132, \9349 );
and \U$4670 ( \13768 , RIdeb2f58_500, \9351 );
and \U$4671 ( \13769 , RIfce1c68_7591, \9353 );
and \U$4672 ( \13770 , RIdeb0258_468, \9355 );
and \U$4673 ( \13771 , RIfc9b498_6789, \9357 );
and \U$4674 ( \13772 , RIdead558_436, \9359 );
and \U$4675 ( \13773 , RIdea6fa0_404, \9361 );
and \U$4676 ( \13774 , RIdea06a0_372, \9363 );
and \U$4677 ( \13775 , RIfc81458_6493, \9365 );
and \U$4678 ( \13776 , RIfc83780_6518, \9367 );
and \U$4679 ( \13777 , RIfc4e620_5914, \9369 );
and \U$4680 ( \13778 , RIfcd3e38_7433, \9371 );
and \U$4681 ( \13779 , RIde937e8_309, \9373 );
and \U$4682 ( \13780 , RIde8f990_290, \9375 );
and \U$4683 ( \13781 , RIde8bb38_271, \9377 );
and \U$4684 ( \13782 , RIde87650_250, \9379 );
and \U$4685 ( \13783 , RIde834b0_230, \9381 );
and \U$4686 ( \13784 , RIfc42c80_5782, \9383 );
and \U$4687 ( \13785 , RIfc65960_6178, \9385 );
and \U$4688 ( \13786 , RIfc6c710_6256, \9387 );
and \U$4689 ( \13787 , RIee392b0_5109, \9389 );
and \U$4690 ( \13788 , RIe16cb60_2614, \9391 );
and \U$4691 ( \13789 , RIe16a6d0_2588, \9393 );
and \U$4692 ( \13790 , RIe169050_2572, \9395 );
and \U$4693 ( \13791 , RIe166a58_2545, \9397 );
and \U$4694 ( \13792 , RIe163d58_2513, \9399 );
and \U$4695 ( \13793 , RIfec3cf0_8348, \9401 );
and \U$4696 ( \13794 , RIe161058_2481, \9403 );
and \U$4697 ( \13795 , RIfcd54b8_7449, \9405 );
and \U$4698 ( \13796 , RIe15e358_2449, \9407 );
and \U$4699 ( \13797 , RIe158958_2385, \9409 );
and \U$4700 ( \13798 , RIe155c58_2353, \9411 );
and \U$4701 ( \13799 , RIfe9ba48_8115, \9413 );
and \U$4702 ( \13800 , RIe152f58_2321, \9415 );
and \U$4703 ( \13801 , RIfec4128_8351, \9417 );
and \U$4704 ( \13802 , RIe150258_2289, \9419 );
and \U$4705 ( \13803 , RIfcb9b28_7135, \9421 );
and \U$4706 ( \13804 , RIe14d558_2257, \9423 );
and \U$4707 ( \13805 , RIe14a858_2225, \9425 );
and \U$4708 ( \13806 , RIe147b58_2193, \9427 );
and \U$4709 ( \13807 , RIfcdb2f0_7516, \9429 );
and \U$4710 ( \13808 , RIfc553d0_5992, \9431 );
and \U$4711 ( \13809 , RIfc9a0e8_6775, \9433 );
and \U$4712 ( \13810 , RIfcbd908_7179, \9435 );
and \U$4713 ( \13811 , RIe1422c0_2130, \9437 );
and \U$4714 ( \13812 , RIe13ff98_2105, \9439 );
and \U$4715 ( \13813 , RIdf3dea0_2081, \9441 );
and \U$4716 ( \13814 , RIdf3ba10_2055, \9443 );
and \U$4717 ( \13815 , RIfc87128_6559, \9445 );
and \U$4718 ( \13816 , RIee304a8_5008, \9447 );
and \U$4719 ( \13817 , RIfcc51f8_7265, \9449 );
and \U$4720 ( \13818 , RIee2e2e8_4984, \9451 );
and \U$4721 ( \13819 , RIdf36cb8_2000, \9453 );
and \U$4722 ( \13820 , RIfec3fc0_8350, \9455 );
and \U$4723 ( \13821 , RIdf32500_1949, \9457 );
and \U$4724 ( \13822 , RIfec3e58_8349, \9459 );
or \U$4725 ( \13823 , \13759 , \13760 , \13761 , \13762 , \13763 , \13764 , \13765 , \13766 , \13767 , \13768 , \13769 , \13770 , \13771 , \13772 , \13773 , \13774 , \13775 , \13776 , \13777 , \13778 , \13779 , \13780 , \13781 , \13782 , \13783 , \13784 , \13785 , \13786 , \13787 , \13788 , \13789 , \13790 , \13791 , \13792 , \13793 , \13794 , \13795 , \13796 , \13797 , \13798 , \13799 , \13800 , \13801 , \13802 , \13803 , \13804 , \13805 , \13806 , \13807 , \13808 , \13809 , \13810 , \13811 , \13812 , \13813 , \13814 , \13815 , \13816 , \13817 , \13818 , \13819 , \13820 , \13821 , \13822 );
and \U$4726 ( \13824 , RIee2c830_4965, \9462 );
and \U$4727 ( \13825 , RIee2ad78_4946, \9464 );
and \U$4728 ( \13826 , RIee296f8_4930, \9466 );
and \U$4729 ( \13827 , RIee284b0_4917, \9468 );
and \U$4730 ( \13828 , RIfe9b8e0_8114, \9470 );
and \U$4731 ( \13829 , RIfe9b610_8112, \9472 );
and \U$4732 ( \13830 , RIfe9b778_8113, \9474 );
and \U$4733 ( \13831 , RIfe9b4a8_8111, \9476 );
and \U$4734 ( \13832 , RIfcb7c38_7113, \9478 );
and \U$4735 ( \13833 , RIfc86b88_6555, \9480 );
and \U$4736 ( \13834 , RIdf238c0_1781, \9482 );
and \U$4737 ( \13835 , RIfc75ab8_6361, \9484 );
and \U$4738 ( \13836 , RIdf22240_1765, \9486 );
and \U$4739 ( \13837 , RIfeaa3b8_8253, \9488 );
and \U$4740 ( \13838 , RIdf1bb98_1692, \9490 );
and \U$4741 ( \13839 , RIdf1a680_1677, \9492 );
and \U$4742 ( \13840 , RIdf18628_1654, \9494 );
and \U$4743 ( \13841 , RIdf15928_1622, \9496 );
and \U$4744 ( \13842 , RIdf12c28_1590, \9498 );
and \U$4745 ( \13843 , RIdf0ff28_1558, \9500 );
and \U$4746 ( \13844 , RIdf0d228_1526, \9502 );
and \U$4747 ( \13845 , RIdf0a528_1494, \9504 );
and \U$4748 ( \13846 , RIdf07828_1462, \9506 );
and \U$4749 ( \13847 , RIdf04b28_1430, \9508 );
and \U$4750 ( \13848 , RIdeff128_1366, \9510 );
and \U$4751 ( \13849 , RIdefc428_1334, \9512 );
and \U$4752 ( \13850 , RIdef9728_1302, \9514 );
and \U$4753 ( \13851 , RIdef6a28_1270, \9516 );
and \U$4754 ( \13852 , RIdef3d28_1238, \9518 );
and \U$4755 ( \13853 , RIdef1028_1206, \9520 );
and \U$4756 ( \13854 , RIdeee328_1174, \9522 );
and \U$4757 ( \13855 , RIdeeb628_1142, \9524 );
and \U$4758 ( \13856 , RIee25a80_4887, \9526 );
and \U$4759 ( \13857 , RIee24c70_4877, \9528 );
and \U$4760 ( \13858 , RIfcddd20_7546, \9530 );
and \U$4761 ( \13859 , RIfccc110_7344, \9532 );
and \U$4762 ( \13860 , RIdee5c28_1078, \9534 );
and \U$4763 ( \13861 , RIdee3ea0_1057, \9536 );
and \U$4764 ( \13862 , RIdee1b78_1032, \9538 );
and \U$4765 ( \13863 , RIdedfc88_1010, \9540 );
and \U$4766 ( \13864 , RIfc6a6b8_6233, \9542 );
and \U$4767 ( \13865 , RIee227e0_4851, \9544 );
and \U$4768 ( \13866 , RIfc88be0_6578, \9546 );
and \U$4769 ( \13867 , RIee21868_4840, \9548 );
and \U$4770 ( \13868 , RIdedaaf8_952, \9550 );
and \U$4771 ( \13869 , RIded8668_926, \9552 );
and \U$4772 ( \13870 , RIded6340_901, \9554 );
and \U$4773 ( \13871 , RIded4180_877, \9556 );
and \U$4774 ( \13872 , RIded1e58_852, \9558 );
and \U$4775 ( \13873 , RIdecf158_820, \9560 );
and \U$4776 ( \13874 , RIdecc458_788, \9562 );
and \U$4777 ( \13875 , RIdec9758_756, \9564 );
and \U$4778 ( \13876 , RIdeb5c58_532, \9566 );
and \U$4779 ( \13877 , RIde99da0_340, \9568 );
and \U$4780 ( \13878 , RIe16f860_2646, \9570 );
and \U$4781 ( \13879 , RIe15b658_2417, \9572 );
and \U$4782 ( \13880 , RIe144e58_2161, \9574 );
and \U$4783 ( \13881 , RIdf39850_2031, \9576 );
and \U$4784 ( \13882 , RIdf2deb0_1899, \9578 );
and \U$4785 ( \13883 , RIdf1e730_1723, \9580 );
and \U$4786 ( \13884 , RIdf01e28_1398, \9582 );
and \U$4787 ( \13885 , RIdee8928_1110, \9584 );
and \U$4788 ( \13886 , RIdedd690_983, \9586 );
and \U$4789 ( \13887 , RIde7fce8_213, \9588 );
or \U$4790 ( \13888 , \13824 , \13825 , \13826 , \13827 , \13828 , \13829 , \13830 , \13831 , \13832 , \13833 , \13834 , \13835 , \13836 , \13837 , \13838 , \13839 , \13840 , \13841 , \13842 , \13843 , \13844 , \13845 , \13846 , \13847 , \13848 , \13849 , \13850 , \13851 , \13852 , \13853 , \13854 , \13855 , \13856 , \13857 , \13858 , \13859 , \13860 , \13861 , \13862 , \13863 , \13864 , \13865 , \13866 , \13867 , \13868 , \13869 , \13870 , \13871 , \13872 , \13873 , \13874 , \13875 , \13876 , \13877 , \13878 , \13879 , \13880 , \13881 , \13882 , \13883 , \13884 , \13885 , \13886 , \13887 );
or \U$4791 ( \13889 , \13823 , \13888 );
_DC g658c ( \13890_nG658c , \13889 , \9597 );
and \U$4792 ( \13891 , RIe19ecf0_3184, \9059 );
and \U$4793 ( \13892 , RIe19bff0_3152, \9061 );
and \U$4794 ( \13893 , RIf145a90_5252, \9063 );
and \U$4795 ( \13894 , RIe1992f0_3120, \9065 );
and \U$4796 ( \13895 , RIf144de8_5243, \9067 );
and \U$4797 ( \13896 , RIe1965f0_3088, \9069 );
and \U$4798 ( \13897 , RIe1938f0_3056, \9071 );
and \U$4799 ( \13898 , RIe190bf0_3024, \9073 );
and \U$4800 ( \13899 , RIe18b1f0_2960, \9075 );
and \U$4801 ( \13900 , RIe1884f0_2928, \9077 );
and \U$4802 ( \13901 , RIfc72980_6326, \9079 );
and \U$4803 ( \13902 , RIe1857f0_2896, \9081 );
and \U$4804 ( \13903 , RIf143060_5222, \9083 );
and \U$4805 ( \13904 , RIe182af0_2864, \9085 );
and \U$4806 ( \13905 , RIe17fdf0_2832, \9087 );
and \U$4807 ( \13906 , RIe17d0f0_2800, \9089 );
and \U$4808 ( \13907 , RIf142688_5215, \9091 );
and \U$4809 ( \13908 , RIf141710_5204, \9093 );
and \U$4810 ( \13909 , RIe177858_2737, \9095 );
and \U$4811 ( \13910 , RIe176778_2725, \9097 );
and \U$4812 ( \13911 , RIfcea638_7689, \9099 );
and \U$4813 ( \13912 , RIfca54e8_6903, \9101 );
and \U$4814 ( \13913 , RIee3e878_5170, \9103 );
and \U$4815 ( \13914 , RIee3dbd0_5161, \9105 );
and \U$4816 ( \13915 , RIee3c988_5148, \9107 );
and \U$4817 ( \13916 , RIee3b5d8_5134, \9109 );
and \U$4818 ( \13917 , RIee3a4f8_5122, \9111 );
and \U$4819 ( \13918 , RIe174b58_2705, \9113 );
and \U$4820 ( \13919 , RIf170600_5738, \9115 );
and \U$4821 ( \13920 , RIfc76fd0_6376, \9117 );
and \U$4822 ( \13921 , RIf16e9e0_5718, \9119 );
and \U$4823 ( \13922 , RIfced608_7723, \9121 );
and \U$4824 ( \13923 , RIf16d090_5700, \9123 );
and \U$4825 ( \13924 , RIe225048_4711, \9125 );
and \U$4826 ( \13925 , RIf16c550_5692, \9127 );
and \U$4827 ( \13926 , RIe222348_4679, \9129 );
and \U$4828 ( \13927 , RIf16b470_5680, \9131 );
and \U$4829 ( \13928 , RIe21f648_4647, \9133 );
and \U$4830 ( \13929 , RIe219c48_4583, \9135 );
and \U$4831 ( \13930 , RIe216f48_4551, \9137 );
and \U$4832 ( \13931 , RIf16a4f8_5669, \9139 );
and \U$4833 ( \13932 , RIe214248_4519, \9141 );
and \U$4834 ( \13933 , RIf169df0_5664, \9143 );
and \U$4835 ( \13934 , RIe211548_4487, \9145 );
and \U$4836 ( \13935 , RIf1684a0_5646, \9147 );
and \U$4837 ( \13936 , RIe20e848_4455, \9149 );
and \U$4838 ( \13937 , RIe20bb48_4423, \9151 );
and \U$4839 ( \13938 , RIe208e48_4391, \9153 );
and \U$4840 ( \13939 , RIf1673c0_5634, \9155 );
and \U$4841 ( \13940 , RIf166448_5623, \9157 );
and \U$4842 ( \13941 , RIfe9c6f0_8124, \9159 );
and \U$4843 ( \13942 , RIfe9c150_8120, \9161 );
and \U$4844 ( \13943 , RIf1654d0_5612, \9163 );
and \U$4845 ( \13944 , RIfcc4550_7256, \9165 );
and \U$4846 ( \13945 , RIf1635e0_5590, \9167 );
and \U$4847 ( \13946 , RIf162500_5578, \9169 );
and \U$4848 ( \13947 , RIf160fe8_5563, \9171 );
and \U$4849 ( \13948 , RIf15f0f8_5541, \9173 );
and \U$4850 ( \13949 , RIfe9bfe8_8119, \9175 );
and \U$4851 ( \13950 , RIfe9c588_8123, \9177 );
and \U$4852 ( \13951 , RIf15d208_5519, \9179 );
and \U$4853 ( \13952 , RIf15bfc0_5506, \9181 );
and \U$4854 ( \13953 , RIfc4d540_5902, \9183 );
and \U$4855 ( \13954 , RIfc9c848_6803, \9185 );
or \U$4856 ( \13955 , \13891 , \13892 , \13893 , \13894 , \13895 , \13896 , \13897 , \13898 , \13899 , \13900 , \13901 , \13902 , \13903 , \13904 , \13905 , \13906 , \13907 , \13908 , \13909 , \13910 , \13911 , \13912 , \13913 , \13914 , \13915 , \13916 , \13917 , \13918 , \13919 , \13920 , \13921 , \13922 , \13923 , \13924 , \13925 , \13926 , \13927 , \13928 , \13929 , \13930 , \13931 , \13932 , \13933 , \13934 , \13935 , \13936 , \13937 , \13938 , \13939 , \13940 , \13941 , \13942 , \13943 , \13944 , \13945 , \13946 , \13947 , \13948 , \13949 , \13950 , \13951 , \13952 , \13953 , \13954 );
and \U$4857 ( \13956 , RIfec4290_8352, \9188 );
and \U$4858 ( \13957 , RIfe9c2b8_8121, \9190 );
and \U$4859 ( \13958 , RIfcc01d0_7208, \9192 );
and \U$4860 ( \13959 , RIe1fb2e8_4235, \9194 );
and \U$4861 ( \13960 , RIfe9c420_8122, \9196 );
and \U$4862 ( \13961 , RIfca3e68_6887, \9198 );
and \U$4863 ( \13962 , RIf154c70_5424, \9200 );
and \U$4864 ( \13963 , RIe1f69c8_4183, \9202 );
and \U$4865 ( \13964 , RIf153a28_5411, \9204 );
and \U$4866 ( \13965 , RIf152240_5394, \9206 );
and \U$4867 ( \13966 , RIf150ff8_5381, \9208 );
and \U$4868 ( \13967 , RIe1f46a0_4158, \9210 );
and \U$4869 ( \13968 , RIfca6028_6911, \9212 );
and \U$4870 ( \13969 , RIfc43bf8_5793, \9214 );
and \U$4871 ( \13970 , RIf14e460_5350, \9216 );
and \U$4872 ( \13971 , RIe1ef3a8_4099, \9218 );
and \U$4873 ( \13972 , RIe1ecdb0_4072, \9220 );
and \U$4874 ( \13973 , RIe1ea0b0_4040, \9222 );
and \U$4875 ( \13974 , RIe1e73b0_4008, \9224 );
and \U$4876 ( \13975 , RIe1e46b0_3976, \9226 );
and \U$4877 ( \13976 , RIe1e19b0_3944, \9228 );
and \U$4878 ( \13977 , RIe1decb0_3912, \9230 );
and \U$4879 ( \13978 , RIe1dbfb0_3880, \9232 );
and \U$4880 ( \13979 , RIe1d92b0_3848, \9234 );
and \U$4881 ( \13980 , RIe1d38b0_3784, \9236 );
and \U$4882 ( \13981 , RIe1d0bb0_3752, \9238 );
and \U$4883 ( \13982 , RIe1cdeb0_3720, \9240 );
and \U$4884 ( \13983 , RIe1cb1b0_3688, \9242 );
and \U$4885 ( \13984 , RIe1c84b0_3656, \9244 );
and \U$4886 ( \13985 , RIe1c57b0_3624, \9246 );
and \U$4887 ( \13986 , RIe1c2ab0_3592, \9248 );
and \U$4888 ( \13987 , RIe1bfdb0_3560, \9250 );
and \U$4889 ( \13988 , RIfc4d6a8_5903, \9252 );
and \U$4890 ( \13989 , RIf14be68_5323, \9254 );
and \U$4891 ( \13990 , RIe1ba680_3498, \9256 );
and \U$4892 ( \13991 , RIfe9be80_8118, \9258 );
and \U$4893 ( \13992 , RIfc86e58_6557, \9260 );
and \U$4894 ( \13993 , RIfcd46a8_7439, \9262 );
and \U$4895 ( \13994 , RIe1b6300_3450, \9264 );
and \U$4896 ( \13995 , RIfe9bd18_8117, \9266 );
and \U$4897 ( \13996 , RIf1495a0_5294, \9268 );
and \U$4898 ( \13997 , RIf1481f0_5280, \9270 );
and \U$4899 ( \13998 , RIe1b3600_3418, \9272 );
and \U$4900 ( \13999 , RIe1b1e18_3401, \9274 );
and \U$4901 ( \14000 , RIfc69470_6220, \9276 );
and \U$4902 ( \14001 , RIfcbfac8_7203, \9278 );
and \U$4903 ( \14002 , RIfe9bbb0_8116, \9280 );
and \U$4904 ( \14003 , RIe1abd10_3332, \9282 );
and \U$4905 ( \14004 , RIe1aa0f0_3312, \9284 );
and \U$4906 ( \14005 , RIe1a73f0_3280, \9286 );
and \U$4907 ( \14006 , RIe1a46f0_3248, \9288 );
and \U$4908 ( \14007 , RIe1a19f0_3216, \9290 );
and \U$4909 ( \14008 , RIe18def0_2992, \9292 );
and \U$4910 ( \14009 , RIe17a3f0_2768, \9294 );
and \U$4911 ( \14010 , RIe227d48_4743, \9296 );
and \U$4912 ( \14011 , RIe21c948_4615, \9298 );
and \U$4913 ( \14012 , RIe206148_4359, \9300 );
and \U$4914 ( \14013 , RIe2001a8_4291, \9302 );
and \U$4915 ( \14014 , RIe1f9560_4214, \9304 );
and \U$4916 ( \14015 , RIe1f20a8_4131, \9306 );
and \U$4917 ( \14016 , RIe1d65b0_3816, \9308 );
and \U$4918 ( \14017 , RIe1bd0b0_3528, \9310 );
and \U$4919 ( \14018 , RIe1aff28_3379, \9312 );
and \U$4920 ( \14019 , RIe172560_2678, \9314 );
or \U$4921 ( \14020 , \13956 , \13957 , \13958 , \13959 , \13960 , \13961 , \13962 , \13963 , \13964 , \13965 , \13966 , \13967 , \13968 , \13969 , \13970 , \13971 , \13972 , \13973 , \13974 , \13975 , \13976 , \13977 , \13978 , \13979 , \13980 , \13981 , \13982 , \13983 , \13984 , \13985 , \13986 , \13987 , \13988 , \13989 , \13990 , \13991 , \13992 , \13993 , \13994 , \13995 , \13996 , \13997 , \13998 , \13999 , \14000 , \14001 , \14002 , \14003 , \14004 , \14005 , \14006 , \14007 , \14008 , \14009 , \14010 , \14011 , \14012 , \14013 , \14014 , \14015 , \14016 , \14017 , \14018 , \14019 );
or \U$4922 ( \14021 , \13955 , \14020 );
_DC g658d ( \14022_nG658d , \14021 , \9323 );
and g658e ( \14023_nG658e , \13890_nG658c , \14022_nG658d );
buf \U$4923 ( \14024 , \14023_nG658e );
and \U$4924 ( \14025 , \14024 , \10691 );
nor \U$4925 ( \14026 , \13758 , \14025 );
xnor \U$4926 ( \14027 , \14026 , \10980 );
not \U$4927 ( \14028 , \13693 );
_DC g4c19 ( \14029_nG4c19 , \13889 , \9597 );
_DC g4c9d ( \14030_nG4c9d , \14021 , \9323 );
xor g4c9e ( \14031_nG4c9e , \14029_nG4c19 , \14030_nG4c9d );
buf \U$4928 ( \14032 , \14031_nG4c9e );
and \U$4929 ( \14033 , \13691 , \12777 );
not \U$4930 ( \14034 , \14033 );
and \U$4931 ( \14035 , \14032 , \14034 );
and \U$4932 ( \14036 , \14028 , \14035 );
xor \U$4933 ( \14037 , \14027 , \14036 );
and \U$4934 ( \14038 , \13682 , \13686 );
and \U$4935 ( \14039 , \13686 , \13693 );
and \U$4936 ( \14040 , \13682 , \13693 );
or \U$4937 ( \14041 , \14038 , \14039 , \14040 );
xor \U$4938 ( \14042 , \14037 , \14041 );
and \U$4939 ( \14043 , \12448 , \11574 );
and \U$4940 ( \14044 , \12769 , \11278 );
nor \U$4941 ( \14045 , \14043 , \14044 );
xnor \U$4942 ( \14046 , \14045 , \11580 );
and \U$4943 ( \14047 , \11270 , \12790 );
and \U$4944 ( \14048 , \11586 , \12461 );
nor \U$4945 ( \14049 , \14047 , \14048 );
xnor \U$4946 ( \14050 , \14049 , \12780 );
xor \U$4947 ( \14051 , \14046 , \14050 );
xor \U$4948 ( \14052 , \14032 , \13691 );
not \U$4949 ( \14053 , \13692 );
and \U$4950 ( \14054 , \14052 , \14053 );
and \U$4951 ( \14055 , \10687 , \14054 );
and \U$4952 ( \14056 , \10988 , \13692 );
nor \U$4953 ( \14057 , \14055 , \14056 );
xnor \U$4954 ( \14058 , \14057 , \14035 );
xor \U$4955 ( \14059 , \14051 , \14058 );
xor \U$4956 ( \14060 , \14042 , \14059 );
and \U$4957 ( \14061 , \13407 , \13411 );
and \U$4958 ( \14062 , \13411 , \13694 );
and \U$4959 ( \14063 , \13407 , \13694 );
or \U$4960 ( \14064 , \14061 , \14062 , \14063 );
xor \U$4961 ( \14065 , \14060 , \14064 );
and \U$4962 ( \14066 , \13695 , \13699 );
and \U$4963 ( \14067 , \13700 , \13703 );
or \U$4964 ( \14068 , \14066 , \14067 );
xor \U$4965 ( \14069 , \14065 , \14068 );
buf g9bf9 ( \14070_nG9bf9 , \14069 );
and \U$4966 ( \14071 , \10704 , \14070_nG9bf9 );
or \U$4967 ( \14072 , \13757 , \14071 );
xor \U$4968 ( \14073 , \10703 , \14072 );
buf \U$4969 ( \14074 , \14073 );
buf \U$4971 ( \14075 , \14074 );
xor \U$4972 ( \14076 , \13756 , \14075 );
buf \U$4973 ( \14077 , \14076 );
xor \U$4974 ( \14078 , \13727 , \14077 );
and \U$4975 ( \14079 , \13716 , \14078 );
and \U$4976 ( \14080 , RIdec6d28_726, \9059 );
and \U$4977 ( \14081 , RIdec4028_694, \9061 );
and \U$4978 ( \14082 , RIee20bc0_4831, \9063 );
and \U$4979 ( \14083 , RIdec1328_662, \9065 );
and \U$4980 ( \14084 , RIfcbaed8_7149, \9067 );
and \U$4981 ( \14085 , RIdebe628_630, \9069 );
and \U$4982 ( \14086 , RIdebb928_598, \9071 );
and \U$4983 ( \14087 , RIdeb8c28_566, \9073 );
and \U$4984 ( \14088 , RIfc412b8_5767, \9075 );
and \U$4985 ( \14089 , RIdeb3228_502, \9077 );
and \U$4986 ( \14090 , RIfc9ea08_6827, \9079 );
and \U$4987 ( \14091 , RIdeb0528_470, \9081 );
and \U$4988 ( \14092 , RIee1e028_4800, \9083 );
and \U$4989 ( \14093 , RIdead828_438, \9085 );
and \U$4990 ( \14094 , RIdea7630_406, \9087 );
and \U$4991 ( \14095 , RIdea0d30_374, \9089 );
and \U$4992 ( \14096 , RIfcbac08_7147, \9091 );
and \U$4993 ( \14097 , RIfc55538_5993, \9093 );
and \U$4994 ( \14098 , RIfcba668_7143, \9095 );
and \U$4995 ( \14099 , RIfc4af48_5875, \9097 );
and \U$4996 ( \14100 , RIfe912f0_7996, \9099 );
and \U$4997 ( \14101 , RIfe91458_7997, \9101 );
and \U$4998 ( \14102 , RIde8be80_272, \9103 );
and \U$4999 ( \14103 , RIde87ce0_252, \9105 );
and \U$5000 ( \14104 , RIfc85238_6537, \9107 );
and \U$5001 ( \14105 , RIfc88640_6574, \9109 );
and \U$5002 ( \14106 , RIfcda210_7504, \9111 );
and \U$5003 ( \14107 , RIfcd5788_7451, \9113 );
and \U$5004 ( \14108 , RIee39418_5110, \9115 );
and \U$5005 ( \14109 , RIe16ce30_2616, \9117 );
and \U$5006 ( \14110 , RIfc884d8_6573, \9119 );
and \U$5007 ( \14111 , RIe169320_2574, \9121 );
and \U$5008 ( \14112 , RIe166d28_2547, \9123 );
and \U$5009 ( \14113 , RIe164028_2515, \9125 );
and \U$5010 ( \14114 , RIfe90918_7989, \9127 );
and \U$5011 ( \14115 , RIe161328_2483, \9129 );
and \U$5012 ( \14116 , RIee36880_5079, \9131 );
and \U$5013 ( \14117 , RIe15e628_2451, \9133 );
and \U$5014 ( \14118 , RIe158c28_2387, \9135 );
and \U$5015 ( \14119 , RIe155f28_2355, \9137 );
and \U$5016 ( \14120 , RIfe91188_7995, \9139 );
and \U$5017 ( \14121 , RIe153228_2323, \9141 );
and \U$5018 ( \14122 , RIfe91020_7994, \9143 );
and \U$5019 ( \14123 , RIe150528_2291, \9145 );
and \U$5020 ( \14124 , RIfcda378_7505, \9147 );
and \U$5021 ( \14125 , RIe14d828_2259, \9149 );
and \U$5022 ( \14126 , RIe14ab28_2227, \9151 );
and \U$5023 ( \14127 , RIe147e28_2195, \9153 );
and \U$5024 ( \14128 , RIfe90eb8_7993, \9155 );
and \U$5025 ( \14129 , RIfe90d50_7992, \9157 );
and \U$5026 ( \14130 , RIfcb99c0_7134, \9159 );
and \U$5027 ( \14131 , RIfc9c2a8_6799, \9161 );
and \U$5028 ( \14132 , RIfe90be8_7991, \9163 );
and \U$5029 ( \14133 , RIfe90a80_7990, \9165 );
and \U$5030 ( \14134 , RIdf3e008_2082, \9167 );
and \U$5031 ( \14135 , RIdf3bce0_2057, \9169 );
and \U$5032 ( \14136 , RIfcec690_7712, \9171 );
and \U$5033 ( \14137 , RIee30778_5010, \9173 );
and \U$5034 ( \14138 , RIfc87dd0_6568, \9175 );
and \U$5035 ( \14139 , RIee2e5b8_4986, \9177 );
and \U$5036 ( \14140 , RIdf36e20_2001, \9179 );
and \U$5037 ( \14141 , RIdf346c0_1973, \9181 );
and \U$5038 ( \14142 , RIdf32668_1950, \9183 );
and \U$5039 ( \14143 , RIdf30070_1923, \9185 );
or \U$5040 ( \14144 , \14080 , \14081 , \14082 , \14083 , \14084 , \14085 , \14086 , \14087 , \14088 , \14089 , \14090 , \14091 , \14092 , \14093 , \14094 , \14095 , \14096 , \14097 , \14098 , \14099 , \14100 , \14101 , \14102 , \14103 , \14104 , \14105 , \14106 , \14107 , \14108 , \14109 , \14110 , \14111 , \14112 , \14113 , \14114 , \14115 , \14116 , \14117 , \14118 , \14119 , \14120 , \14121 , \14122 , \14123 , \14124 , \14125 , \14126 , \14127 , \14128 , \14129 , \14130 , \14131 , \14132 , \14133 , \14134 , \14135 , \14136 , \14137 , \14138 , \14139 , \14140 , \14141 , \14142 , \14143 );
and \U$5041 ( \14145 , RIee2c998_4966, \9188 );
and \U$5042 ( \14146 , RIee2aee0_4947, \9190 );
and \U$5043 ( \14147 , RIee299c8_4932, \9192 );
and \U$5044 ( \14148 , RIee28618_4918, \9194 );
and \U$5045 ( \14149 , RIfe90378_7985, \9196 );
and \U$5046 ( \14150 , RIfe907b0_7988, \9198 );
and \U$5047 ( \14151 , RIfe904e0_7986, \9200 );
and \U$5048 ( \14152 , RIfe90648_7987, \9202 );
and \U$5049 ( \14153 , RIfc9d928_6815, \9204 );
and \U$5050 ( \14154 , RIfc86048_6547, \9206 );
and \U$5051 ( \14155 , RIfcb92b8_7129, \9208 );
and \U$5052 ( \14156 , RIfc4ee90_5920, \9210 );
and \U$5053 ( \14157 , RIfc86a20_6554, \9212 );
and \U$5054 ( \14158 , RIdf20e90_1751, \9214 );
and \U$5055 ( \14159 , RIfcb8fe8_7127, \9216 );
and \U$5056 ( \14160 , RIdf1a950_1679, \9218 );
and \U$5057 ( \14161 , RIdf188f8_1656, \9220 );
and \U$5058 ( \14162 , RIdf15bf8_1624, \9222 );
and \U$5059 ( \14163 , RIdf12ef8_1592, \9224 );
and \U$5060 ( \14164 , RIdf101f8_1560, \9226 );
and \U$5061 ( \14165 , RIdf0d4f8_1528, \9228 );
and \U$5062 ( \14166 , RIdf0a7f8_1496, \9230 );
and \U$5063 ( \14167 , RIdf07af8_1464, \9232 );
and \U$5064 ( \14168 , RIdf04df8_1432, \9234 );
and \U$5065 ( \14169 , RIdeff3f8_1368, \9236 );
and \U$5066 ( \14170 , RIdefc6f8_1336, \9238 );
and \U$5067 ( \14171 , RIdef99f8_1304, \9240 );
and \U$5068 ( \14172 , RIdef6cf8_1272, \9242 );
and \U$5069 ( \14173 , RIdef3ff8_1240, \9244 );
and \U$5070 ( \14174 , RIdef12f8_1208, \9246 );
and \U$5071 ( \14175 , RIdeee5f8_1176, \9248 );
and \U$5072 ( \14176 , RIdeeb8f8_1144, \9250 );
and \U$5073 ( \14177 , RIfc857d8_6541, \9252 );
and \U$5074 ( \14178 , RIee24dd8_4878, \9254 );
and \U$5075 ( \14179 , RIfc4ff70_5932, \9256 );
and \U$5076 ( \14180 , RIfc50240_5934, \9258 );
and \U$5077 ( \14181 , RIdee5ef8_1080, \9260 );
and \U$5078 ( \14182 , RIdee4170_1059, \9262 );
and \U$5079 ( \14183 , RIfe915c0_7998, \9264 );
and \U$5080 ( \14184 , RIdedff58_1012, \9266 );
and \U$5081 ( \14185 , RIfcd4810_7440, \9268 );
and \U$5082 ( \14186 , RIee22948_4852, \9270 );
and \U$5083 ( \14187 , RIfce1560_7586, \9272 );
and \U$5084 ( \14188 , RIee219d0_4841, \9274 );
and \U$5085 ( \14189 , RIdedac60_953, \9276 );
and \U$5086 ( \14190 , RIfe91728_7999, \9278 );
and \U$5087 ( \14191 , RIded64a8_902, \9280 );
and \U$5088 ( \14192 , RIfe91890_8000, \9282 );
and \U$5089 ( \14193 , RIded2128_854, \9284 );
and \U$5090 ( \14194 , RIdecf428_822, \9286 );
and \U$5091 ( \14195 , RIdecc728_790, \9288 );
and \U$5092 ( \14196 , RIdec9a28_758, \9290 );
and \U$5093 ( \14197 , RIdeb5f28_534, \9292 );
and \U$5094 ( \14198 , RIde9a430_342, \9294 );
and \U$5095 ( \14199 , RIe16fb30_2648, \9296 );
and \U$5096 ( \14200 , RIe15b928_2419, \9298 );
and \U$5097 ( \14201 , RIe145128_2163, \9300 );
and \U$5098 ( \14202 , RIdf39b20_2033, \9302 );
and \U$5099 ( \14203 , RIdf2e180_1901, \9304 );
and \U$5100 ( \14204 , RIdf1ea00_1725, \9306 );
and \U$5101 ( \14205 , RIdf020f8_1400, \9308 );
and \U$5102 ( \14206 , RIdee8bf8_1112, \9310 );
and \U$5103 ( \14207 , RIdedd960_985, \9312 );
and \U$5104 ( \14208 , RIde80378_215, \9314 );
or \U$5105 ( \14209 , \14145 , \14146 , \14147 , \14148 , \14149 , \14150 , \14151 , \14152 , \14153 , \14154 , \14155 , \14156 , \14157 , \14158 , \14159 , \14160 , \14161 , \14162 , \14163 , \14164 , \14165 , \14166 , \14167 , \14168 , \14169 , \14170 , \14171 , \14172 , \14173 , \14174 , \14175 , \14176 , \14177 , \14178 , \14179 , \14180 , \14181 , \14182 , \14183 , \14184 , \14185 , \14186 , \14187 , \14188 , \14189 , \14190 , \14191 , \14192 , \14193 , \14194 , \14195 , \14196 , \14197 , \14198 , \14199 , \14200 , \14201 , \14202 , \14203 , \14204 , \14205 , \14206 , \14207 , \14208 );
or \U$5106 ( \14210 , \14144 , \14209 );
_DC g2da3 ( \14211_nG2da3 , \14210 , \9323 );
buf \U$5107 ( \14212 , \14211_nG2da3 );
and \U$5108 ( \14213 , RIe19efc0_3186, \9333 );
and \U$5109 ( \14214 , RIe19c2c0_3154, \9335 );
and \U$5110 ( \14215 , RIf145d60_5254, \9337 );
and \U$5111 ( \14216 , RIe1995c0_3122, \9339 );
and \U$5112 ( \14217 , RIfc637a0_6154, \9341 );
and \U$5113 ( \14218 , RIe1968c0_3090, \9343 );
and \U$5114 ( \14219 , RIe193bc0_3058, \9345 );
and \U$5115 ( \14220 , RIe190ec0_3026, \9347 );
and \U$5116 ( \14221 , RIe18b4c0_2962, \9349 );
and \U$5117 ( \14222 , RIe1887c0_2930, \9351 );
and \U$5118 ( \14223 , RIfc62af8_6145, \9353 );
and \U$5119 ( \14224 , RIe185ac0_2898, \9355 );
and \U$5120 ( \14225 , RIfe8fc70_7980, \9357 );
and \U$5121 ( \14226 , RIe182dc0_2866, \9359 );
and \U$5122 ( \14227 , RIe1800c0_2834, \9361 );
and \U$5123 ( \14228 , RIe17d3c0_2802, \9363 );
and \U$5124 ( \14229 , RIfe90210_7984, \9365 );
and \U$5125 ( \14230 , RIfe8ff40_7982, \9367 );
and \U$5126 ( \14231 , RIfc72f20_6330, \9369 );
and \U$5127 ( \14232 , RIe176a48_2727, \9371 );
and \U$5128 ( \14233 , RIfcaf6a0_7018, \9373 );
and \U$5129 ( \14234 , RIfc61040_6126, \9375 );
and \U$5130 ( \14235 , RIf13e8a8_5171, \9377 );
and \U$5131 ( \14236 , RIfe900a8_7983, \9379 );
and \U$5132 ( \14237 , RIee3caf0_5149, \9381 );
and \U$5133 ( \14238 , RIee3b740_5135, \9383 );
and \U$5134 ( \14239 , RIee3a660_5123, \9385 );
and \U$5135 ( \14240 , RIe174e28_2707, \9387 );
and \U$5136 ( \14241 , RIf170768_5739, \9389 );
and \U$5137 ( \14242 , RIfc5fdf8_6113, \9391 );
and \U$5138 ( \14243 , RIf16eb48_5719, \9393 );
and \U$5139 ( \14244 , RIfcaaab0_6964, \9395 );
and \U$5140 ( \14245 , RIf16d1f8_5701, \9397 );
and \U$5141 ( \14246 , RIe225318_4713, \9399 );
and \U$5142 ( \14247 , RIf16c6b8_5693, \9401 );
and \U$5143 ( \14248 , RIe222618_4681, \9403 );
and \U$5144 ( \14249 , RIf16b5d8_5681, \9405 );
and \U$5145 ( \14250 , RIe21f918_4649, \9407 );
and \U$5146 ( \14251 , RIe219f18_4585, \9409 );
and \U$5147 ( \14252 , RIe217218_4553, \9411 );
and \U$5148 ( \14253 , RIfca62f8_6913, \9413 );
and \U$5149 ( \14254 , RIe214518_4521, \9415 );
and \U$5150 ( \14255 , RIfcc9578_7313, \9417 );
and \U$5151 ( \14256 , RIe211818_4489, \9419 );
and \U$5152 ( \14257 , RIfca5a88_6907, \9421 );
and \U$5153 ( \14258 , RIe20eb18_4457, \9423 );
and \U$5154 ( \14259 , RIe20be18_4425, \9425 );
and \U$5155 ( \14260 , RIe209118_4393, \9427 );
and \U$5156 ( \14261 , RIf167690_5636, \9429 );
and \U$5157 ( \14262 , RIf166718_5625, \9431 );
and \U$5158 ( \14263 , RIfe8f9a0_7978, \9433 );
and \U$5159 ( \14264 , RIfe8f838_7977, \9435 );
and \U$5160 ( \14265 , RIf165638_5613, \9437 );
and \U$5161 ( \14266 , RIf164990_5604, \9439 );
and \U$5162 ( \14267 , RIf1638b0_5592, \9441 );
and \U$5163 ( \14268 , RIf1627d0_5580, \9443 );
and \U$5164 ( \14269 , RIf161150_5564, \9445 );
and \U$5165 ( \14270 , RIf15f260_5542, \9447 );
and \U$5166 ( \14271 , RIe1fd778_4261, \9449 );
and \U$5167 ( \14272 , RIe1fc530_4248, \9451 );
and \U$5168 ( \14273 , RIf15d4d8_5521, \9453 );
and \U$5169 ( \14274 , RIf15c290_5508, \9455 );
and \U$5170 ( \14275 , RIfca20e0_6866, \9457 );
and \U$5171 ( \14276 , RIf159f68_5483, \9459 );
or \U$5172 ( \14277 , \14213 , \14214 , \14215 , \14216 , \14217 , \14218 , \14219 , \14220 , \14221 , \14222 , \14223 , \14224 , \14225 , \14226 , \14227 , \14228 , \14229 , \14230 , \14231 , \14232 , \14233 , \14234 , \14235 , \14236 , \14237 , \14238 , \14239 , \14240 , \14241 , \14242 , \14243 , \14244 , \14245 , \14246 , \14247 , \14248 , \14249 , \14250 , \14251 , \14252 , \14253 , \14254 , \14255 , \14256 , \14257 , \14258 , \14259 , \14260 , \14261 , \14262 , \14263 , \14264 , \14265 , \14266 , \14267 , \14268 , \14269 , \14270 , \14271 , \14272 , \14273 , \14274 , \14275 , \14276 );
and \U$5173 ( \14278 , RIf159428_5475, \9462 );
and \U$5174 ( \14279 , RIf1581e0_5462, \9464 );
and \U$5175 ( \14280 , RIfc5ebb0_6100, \9466 );
and \U$5176 ( \14281 , RIfe8fdd8_7981, \9468 );
and \U$5177 ( \14282 , RIfc69e48_6227, \9470 );
and \U$5178 ( \14283 , RIfc5e8e0_6098, \9472 );
and \U$5179 ( \14284 , RIf154f40_5426, \9474 );
and \U$5180 ( \14285 , RIe1f6b30_4184, \9476 );
and \U$5181 ( \14286 , RIf153b90_5412, \9478 );
and \U$5182 ( \14287 , RIf1523a8_5395, \9480 );
and \U$5183 ( \14288 , RIfce88b0_7668, \9482 );
and \U$5184 ( \14289 , RIfe8fb08_7979, \9484 );
and \U$5185 ( \14290 , RIfcebe20_7706, \9486 );
and \U$5186 ( \14291 , RIfcb1158_7037, \9488 );
and \U$5187 ( \14292 , RIf14e730_5352, \9490 );
and \U$5188 ( \14293 , RIe1ef678_4101, \9492 );
and \U$5189 ( \14294 , RIe1ed080_4074, \9494 );
and \U$5190 ( \14295 , RIe1ea380_4042, \9496 );
and \U$5191 ( \14296 , RIe1e7680_4010, \9498 );
and \U$5192 ( \14297 , RIe1e4980_3978, \9500 );
and \U$5193 ( \14298 , RIe1e1c80_3946, \9502 );
and \U$5194 ( \14299 , RIe1def80_3914, \9504 );
and \U$5195 ( \14300 , RIe1dc280_3882, \9506 );
and \U$5196 ( \14301 , RIe1d9580_3850, \9508 );
and \U$5197 ( \14302 , RIe1d3b80_3786, \9510 );
and \U$5198 ( \14303 , RIe1d0e80_3754, \9512 );
and \U$5199 ( \14304 , RIe1ce180_3722, \9514 );
and \U$5200 ( \14305 , RIe1cb480_3690, \9516 );
and \U$5201 ( \14306 , RIe1c8780_3658, \9518 );
and \U$5202 ( \14307 , RIe1c5a80_3626, \9520 );
and \U$5203 ( \14308 , RIe1c2d80_3594, \9522 );
and \U$5204 ( \14309 , RIe1c0080_3562, \9524 );
and \U$5205 ( \14310 , RIfcc8ba0_7306, \9526 );
and \U$5206 ( \14311 , RIfc5d698_6085, \9528 );
and \U$5207 ( \14312 , RIfec35e8_8343, \9530 );
and \U$5208 ( \14313 , RIfeabd08_8271, \9532 );
and \U$5209 ( \14314 , RIfc5cf90_6080, \9534 );
and \U$5210 ( \14315 , RIfc5ce28_6079, \9536 );
and \U$5211 ( \14316 , RIfec31b0_8340, \9538 );
and \U$5212 ( \14317 , RIe1b4b18_3433, \9540 );
and \U$5213 ( \14318 , RIf149708_5295, \9542 );
and \U$5214 ( \14319 , RIf148358_5281, \9544 );
and \U$5215 ( \14320 , RIe1b3768_3419, \9546 );
and \U$5216 ( \14321 , RIfec3480_8342, \9548 );
and \U$5217 ( \14322 , RIfc483b0_5844, \9550 );
and \U$5218 ( \14323 , RIfc80be8_6487, \9552 );
and \U$5219 ( \14324 , RIe1ad4f8_3349, \9554 );
and \U$5220 ( \14325 , RIfec3318_8341, \9556 );
and \U$5221 ( \14326 , RIe1aa3c0_3314, \9558 );
and \U$5222 ( \14327 , RIe1a76c0_3282, \9560 );
and \U$5223 ( \14328 , RIe1a49c0_3250, \9562 );
and \U$5224 ( \14329 , RIe1a1cc0_3218, \9564 );
and \U$5225 ( \14330 , RIe18e1c0_2994, \9566 );
and \U$5226 ( \14331 , RIe17a6c0_2770, \9568 );
and \U$5227 ( \14332 , RIe228018_4745, \9570 );
and \U$5228 ( \14333 , RIe21cc18_4617, \9572 );
and \U$5229 ( \14334 , RIe206418_4361, \9574 );
and \U$5230 ( \14335 , RIe200478_4293, \9576 );
and \U$5231 ( \14336 , RIe1f9830_4216, \9578 );
and \U$5232 ( \14337 , RIe1f2378_4133, \9580 );
and \U$5233 ( \14338 , RIe1d6880_3818, \9582 );
and \U$5234 ( \14339 , RIe1bd380_3530, \9584 );
and \U$5235 ( \14340 , RIe1b01f8_3381, \9586 );
and \U$5236 ( \14341 , RIe172830_2680, \9588 );
or \U$5237 ( \14342 , \14278 , \14279 , \14280 , \14281 , \14282 , \14283 , \14284 , \14285 , \14286 , \14287 , \14288 , \14289 , \14290 , \14291 , \14292 , \14293 , \14294 , \14295 , \14296 , \14297 , \14298 , \14299 , \14300 , \14301 , \14302 , \14303 , \14304 , \14305 , \14306 , \14307 , \14308 , \14309 , \14310 , \14311 , \14312 , \14313 , \14314 , \14315 , \14316 , \14317 , \14318 , \14319 , \14320 , \14321 , \14322 , \14323 , \14324 , \14325 , \14326 , \14327 , \14328 , \14329 , \14330 , \14331 , \14332 , \14333 , \14334 , \14335 , \14336 , \14337 , \14338 , \14339 , \14340 , \14341 );
or \U$5238 ( \14343 , \14277 , \14342 );
_DC g3ed0 ( \14344_nG3ed0 , \14343 , \9597 );
buf \U$5239 ( \14345 , \14344_nG3ed0 );
xor \U$5240 ( \14346 , \14212 , \14345 );
and \U$5241 ( \14347 , RIdec6bc0_725, \9059 );
and \U$5242 ( \14348 , RIdec3ec0_693, \9061 );
and \U$5243 ( \14349 , RIee20a58_4830, \9063 );
and \U$5244 ( \14350 , RIdec11c0_661, \9065 );
and \U$5245 ( \14351 , RIee1f978_4818, \9067 );
and \U$5246 ( \14352 , RIdebe4c0_629, \9069 );
and \U$5247 ( \14353 , RIdebb7c0_597, \9071 );
and \U$5248 ( \14354 , RIdeb8ac0_565, \9073 );
and \U$5249 ( \14355 , RIee1efa0_4811, \9075 );
and \U$5250 ( \14356 , RIdeb30c0_501, \9077 );
and \U$5251 ( \14357 , RIfcb04b0_7028, \9079 );
and \U$5252 ( \14358 , RIdeb03c0_469, \9081 );
and \U$5253 ( \14359 , RIfc5e4a8_6095, \9083 );
and \U$5254 ( \14360 , RIdead6c0_437, \9085 );
and \U$5255 ( \14361 , RIdea72e8_405, \9087 );
and \U$5256 ( \14362 , RIdea09e8_373, \9089 );
and \U$5257 ( \14363 , RIfcb2508_7051, \9091 );
and \U$5258 ( \14364 , RIfcd16d8_7405, \9093 );
and \U$5259 ( \14365 , RIfc5d800_6086, \9095 );
and \U$5260 ( \14366 , RIfc63d40_6158, \9097 );
and \U$5261 ( \14367 , RIde93b30_310, \9099 );
and \U$5262 ( \14368 , RIfea7820_8222, \9101 );
and \U$5263 ( \14369 , RIfea73e8_8219, \9103 );
and \U$5264 ( \14370 , RIde87998_251, \9105 );
and \U$5265 ( \14371 , RIde837f8_231, \9107 );
and \U$5266 ( \14372 , RIfc7bd28_6431, \9109 );
and \U$5267 ( \14373 , RIfcc7ef8_7297, \9111 );
and \U$5268 ( \14374 , RIfc7a108_6411, \9113 );
and \U$5269 ( \14375 , RIfc7a6a8_6415, \9115 );
and \U$5270 ( \14376 , RIe16ccc8_2615, \9117 );
and \U$5271 ( \14377 , RIe16a838_2589, \9119 );
and \U$5272 ( \14378 , RIe1691b8_2573, \9121 );
and \U$5273 ( \14379 , RIe166bc0_2546, \9123 );
and \U$5274 ( \14380 , RIe163ec0_2514, \9125 );
and \U$5275 ( \14381 , RIee38338_5098, \9127 );
and \U$5276 ( \14382 , RIe1611c0_2482, \9129 );
and \U$5277 ( \14383 , RIfc54b60_5986, \9131 );
and \U$5278 ( \14384 , RIe15e4c0_2450, \9133 );
and \U$5279 ( \14385 , RIe158ac0_2386, \9135 );
and \U$5280 ( \14386 , RIe155dc0_2354, \9137 );
and \U$5281 ( \14387 , RIee35a70_5069, \9139 );
and \U$5282 ( \14388 , RIe1530c0_2322, \9141 );
and \U$5283 ( \14389 , RIee357a0_5067, \9143 );
and \U$5284 ( \14390 , RIe1503c0_2290, \9145 );
and \U$5285 ( \14391 , RIfc9fdb8_6841, \9147 );
and \U$5286 ( \14392 , RIe14d6c0_2258, \9149 );
and \U$5287 ( \14393 , RIe14a9c0_2226, \9151 );
and \U$5288 ( \14394 , RIe147cc0_2194, \9153 );
and \U$5289 ( \14395 , RIee34af8_5058, \9155 );
and \U$5290 ( \14396 , RIee33a18_5046, \9157 );
and \U$5291 ( \14397 , RIee327d0_5033, \9159 );
and \U$5292 ( \14398 , RIfcbcf30_7172, \9161 );
and \U$5293 ( \14399 , RIe142428_2131, \9163 );
and \U$5294 ( \14400 , RIe140100_2106, \9165 );
and \U$5295 ( \14401 , RIfea7280_8218, \9167 );
and \U$5296 ( \14402 , RIdf3bb78_2056, \9169 );
and \U$5297 ( \14403 , RIfc731f0_6332, \9171 );
and \U$5298 ( \14404 , RIee30610_5009, \9173 );
and \U$5299 ( \14405 , RIfcbe010_7184, \9175 );
and \U$5300 ( \14406 , RIee2e450_4985, \9177 );
and \U$5301 ( \14407 , RIfec2ee0_8338, \9179 );
and \U$5302 ( \14408 , RIfec3048_8339, \9181 );
and \U$5303 ( \14409 , RIfec2c10_8336, \9183 );
and \U$5304 ( \14410 , RIfec2d78_8337, \9185 );
or \U$5305 ( \14411 , \14347 , \14348 , \14349 , \14350 , \14351 , \14352 , \14353 , \14354 , \14355 , \14356 , \14357 , \14358 , \14359 , \14360 , \14361 , \14362 , \14363 , \14364 , \14365 , \14366 , \14367 , \14368 , \14369 , \14370 , \14371 , \14372 , \14373 , \14374 , \14375 , \14376 , \14377 , \14378 , \14379 , \14380 , \14381 , \14382 , \14383 , \14384 , \14385 , \14386 , \14387 , \14388 , \14389 , \14390 , \14391 , \14392 , \14393 , \14394 , \14395 , \14396 , \14397 , \14398 , \14399 , \14400 , \14401 , \14402 , \14403 , \14404 , \14405 , \14406 , \14407 , \14408 , \14409 , \14410 );
and \U$5306 ( \14412 , RIfcb46c8_7075, \9188 );
and \U$5307 ( \14413 , RIfcb4830_7076, \9190 );
and \U$5308 ( \14414 , RIee29860_4931, \9192 );
and \U$5309 ( \14415 , RIfcb88e0_7122, \9194 );
and \U$5310 ( \14416 , RIdf2b480_1869, \9196 );
and \U$5311 ( \14417 , RIdf29590_1847, \9198 );
and \U$5312 ( \14418 , RIdf27268_1822, \9200 );
and \U$5313 ( \14419 , RIdf25648_1802, \9202 );
and \U$5314 ( \14420 , RIfcc9de8_7319, \9204 );
and \U$5315 ( \14421 , RIfc53648_5971, \9206 );
and \U$5316 ( \14422 , RIdf23a28_1782, \9208 );
and \U$5317 ( \14423 , RIfc823d0_6504, \9210 );
and \U$5318 ( \14424 , RIdf223a8_1766, \9212 );
and \U$5319 ( \14425 , RIdf20d28_1750, \9214 );
and \U$5320 ( \14426 , RIdf1bd00_1693, \9216 );
and \U$5321 ( \14427 , RIdf1a7e8_1678, \9218 );
and \U$5322 ( \14428 , RIdf18790_1655, \9220 );
and \U$5323 ( \14429 , RIdf15a90_1623, \9222 );
and \U$5324 ( \14430 , RIdf12d90_1591, \9224 );
and \U$5325 ( \14431 , RIdf10090_1559, \9226 );
and \U$5326 ( \14432 , RIdf0d390_1527, \9228 );
and \U$5327 ( \14433 , RIdf0a690_1495, \9230 );
and \U$5328 ( \14434 , RIdf07990_1463, \9232 );
and \U$5329 ( \14435 , RIdf04c90_1431, \9234 );
and \U$5330 ( \14436 , RIdeff290_1367, \9236 );
and \U$5331 ( \14437 , RIdefc590_1335, \9238 );
and \U$5332 ( \14438 , RIdef9890_1303, \9240 );
and \U$5333 ( \14439 , RIdef6b90_1271, \9242 );
and \U$5334 ( \14440 , RIdef3e90_1239, \9244 );
and \U$5335 ( \14441 , RIdef1190_1207, \9246 );
and \U$5336 ( \14442 , RIdeee490_1175, \9248 );
and \U$5337 ( \14443 , RIdeeb790_1143, \9250 );
and \U$5338 ( \14444 , RIee25be8_4888, \9252 );
and \U$5339 ( \14445 , RIfc6af28_6239, \9254 );
and \U$5340 ( \14446 , RIee23fc8_4868, \9256 );
and \U$5341 ( \14447 , RIfccf680_7382, \9258 );
and \U$5342 ( \14448 , RIdee5d90_1079, \9260 );
and \U$5343 ( \14449 , RIdee4008_1058, \9262 );
and \U$5344 ( \14450 , RIdee1ce0_1033, \9264 );
and \U$5345 ( \14451 , RIdedfdf0_1011, \9266 );
and \U$5346 ( \14452 , RIfc6b090_6240, \9268 );
and \U$5347 ( \14453 , RIfc534e0_5970, \9270 );
and \U$5348 ( \14454 , RIfca5920_6906, \9272 );
and \U$5349 ( \14455 , RIfc66770_6188, \9274 );
and \U$5350 ( \14456 , RIfe8f6d0_7976, \9276 );
and \U$5351 ( \14457 , RIded87d0_927, \9278 );
and \U$5352 ( \14458 , RIfe8f568_7975, \9280 );
and \U$5353 ( \14459 , RIded42e8_878, \9282 );
and \U$5354 ( \14460 , RIded1fc0_853, \9284 );
and \U$5355 ( \14461 , RIdecf2c0_821, \9286 );
and \U$5356 ( \14462 , RIdecc5c0_789, \9288 );
and \U$5357 ( \14463 , RIdec98c0_757, \9290 );
and \U$5358 ( \14464 , RIdeb5dc0_533, \9292 );
and \U$5359 ( \14465 , RIde9a0e8_341, \9294 );
and \U$5360 ( \14466 , RIe16f9c8_2647, \9296 );
and \U$5361 ( \14467 , RIe15b7c0_2418, \9298 );
and \U$5362 ( \14468 , RIe144fc0_2162, \9300 );
and \U$5363 ( \14469 , RIdf399b8_2032, \9302 );
and \U$5364 ( \14470 , RIdf2e018_1900, \9304 );
and \U$5365 ( \14471 , RIdf1e898_1724, \9306 );
and \U$5366 ( \14472 , RIdf01f90_1399, \9308 );
and \U$5367 ( \14473 , RIdee8a90_1111, \9310 );
and \U$5368 ( \14474 , RIdedd7f8_984, \9312 );
and \U$5369 ( \14475 , RIde80030_214, \9314 );
or \U$5370 ( \14476 , \14412 , \14413 , \14414 , \14415 , \14416 , \14417 , \14418 , \14419 , \14420 , \14421 , \14422 , \14423 , \14424 , \14425 , \14426 , \14427 , \14428 , \14429 , \14430 , \14431 , \14432 , \14433 , \14434 , \14435 , \14436 , \14437 , \14438 , \14439 , \14440 , \14441 , \14442 , \14443 , \14444 , \14445 , \14446 , \14447 , \14448 , \14449 , \14450 , \14451 , \14452 , \14453 , \14454 , \14455 , \14456 , \14457 , \14458 , \14459 , \14460 , \14461 , \14462 , \14463 , \14464 , \14465 , \14466 , \14467 , \14468 , \14469 , \14470 , \14471 , \14472 , \14473 , \14474 , \14475 );
or \U$5371 ( \14477 , \14411 , \14476 );
_DC g2e28 ( \14478_nG2e28 , \14477 , \9323 );
buf \U$5372 ( \14479 , \14478_nG2e28 );
and \U$5373 ( \14480 , RIe19ee58_3185, \9333 );
and \U$5374 ( \14481 , RIe19c158_3153, \9335 );
and \U$5375 ( \14482 , RIf145bf8_5253, \9337 );
and \U$5376 ( \14483 , RIe199458_3121, \9339 );
and \U$5377 ( \14484 , RIfe8f298_7973, \9341 );
and \U$5378 ( \14485 , RIe196758_3089, \9343 );
and \U$5379 ( \14486 , RIe193a58_3057, \9345 );
and \U$5380 ( \14487 , RIe190d58_3025, \9347 );
and \U$5381 ( \14488 , RIe18b358_2961, \9349 );
and \U$5382 ( \14489 , RIe188658_2929, \9351 );
and \U$5383 ( \14490 , RIfe8f130_7972, \9353 );
and \U$5384 ( \14491 , RIe185958_2897, \9355 );
and \U$5385 ( \14492 , RIfc9f278_6833, \9357 );
and \U$5386 ( \14493 , RIe182c58_2865, \9359 );
and \U$5387 ( \14494 , RIe17ff58_2833, \9361 );
and \U$5388 ( \14495 , RIe17d258_2801, \9363 );
and \U$5389 ( \14496 , RIf1427f0_5216, \9365 );
and \U$5390 ( \14497 , RIfe8efc8_7971, \9367 );
and \U$5391 ( \14498 , RIe1779c0_2738, \9369 );
and \U$5392 ( \14499 , RIe1768e0_2726, \9371 );
and \U$5393 ( \14500 , RIfc81e30_6500, \9373 );
and \U$5394 ( \14501 , RIfc9ff20_6842, \9375 );
and \U$5395 ( \14502 , RIfca0088_6843, \9377 );
and \U$5396 ( \14503 , RIfc81b60_6498, \9379 );
and \U$5397 ( \14504 , RIfce5778_7633, \9381 );
and \U$5398 ( \14505 , RIfce08b8_7577, \9383 );
and \U$5399 ( \14506 , RIfc815c0_6494, \9385 );
and \U$5400 ( \14507 , RIe174cc0_2706, \9387 );
and \U$5401 ( \14508 , RIfca04c0_6846, \9389 );
and \U$5402 ( \14509 , RIfc53eb8_5977, \9391 );
and \U$5403 ( \14510 , RIfcc65a8_7279, \9393 );
and \U$5404 ( \14511 , RIfc80d50_6488, \9395 );
and \U$5405 ( \14512 , RIfc804e0_6482, \9397 );
and \U$5406 ( \14513 , RIe2251b0_4712, \9399 );
and \U$5407 ( \14514 , RIfc80378_6481, \9401 );
and \U$5408 ( \14515 , RIe2224b0_4680, \9403 );
and \U$5409 ( \14516 , RIfcb5910_7088, \9405 );
and \U$5410 ( \14517 , RIe21f7b0_4648, \9407 );
and \U$5411 ( \14518 , RIe219db0_4584, \9409 );
and \U$5412 ( \14519 , RIe2170b0_4552, \9411 );
and \U$5413 ( \14520 , RIfca01f0_6844, \9413 );
and \U$5414 ( \14521 , RIe2143b0_4520, \9415 );
and \U$5415 ( \14522 , RIfc82c40_6510, \9417 );
and \U$5416 ( \14523 , RIe2116b0_4488, \9419 );
and \U$5417 ( \14524 , RIfc7f6d0_6472, \9421 );
and \U$5418 ( \14525 , RIe20e9b0_4456, \9423 );
and \U$5419 ( \14526 , RIe20bcb0_4424, \9425 );
and \U$5420 ( \14527 , RIe208fb0_4392, \9427 );
and \U$5421 ( \14528 , RIf167528_5635, \9429 );
and \U$5422 ( \14529 , RIf1665b0_5624, \9431 );
and \U$5423 ( \14530 , RIe203718_4329, \9433 );
and \U$5424 ( \14531 , RIe201c60_4310, \9435 );
and \U$5425 ( \14532 , RIfc9da90_6816, \9437 );
and \U$5426 ( \14533 , RIfcc5360_7266, \9439 );
and \U$5427 ( \14534 , RIf163748_5591, \9441 );
and \U$5428 ( \14535 , RIf162668_5579, \9443 );
and \U$5429 ( \14536 , RIfc7e320_6458, \9445 );
and \U$5430 ( \14537 , RIfc87998_6565, \9447 );
and \U$5431 ( \14538 , RIe1fd610_4260, \9449 );
and \U$5432 ( \14539 , RIe1fc3c8_4247, \9451 );
and \U$5433 ( \14540 , RIf15d370_5520, \9453 );
and \U$5434 ( \14541 , RIf15c128_5507, \9455 );
and \U$5435 ( \14542 , RIfcc5d38_7273, \9457 );
and \U$5436 ( \14543 , RIfce7d70_7660, \9459 );
or \U$5437 ( \14544 , \14480 , \14481 , \14482 , \14483 , \14484 , \14485 , \14486 , \14487 , \14488 , \14489 , \14490 , \14491 , \14492 , \14493 , \14494 , \14495 , \14496 , \14497 , \14498 , \14499 , \14500 , \14501 , \14502 , \14503 , \14504 , \14505 , \14506 , \14507 , \14508 , \14509 , \14510 , \14511 , \14512 , \14513 , \14514 , \14515 , \14516 , \14517 , \14518 , \14519 , \14520 , \14521 , \14522 , \14523 , \14524 , \14525 , \14526 , \14527 , \14528 , \14529 , \14530 , \14531 , \14532 , \14533 , \14534 , \14535 , \14536 , \14537 , \14538 , \14539 , \14540 , \14541 , \14542 , \14543 );
and \U$5438 ( \14545 , RIfc4bd58_5885, \9462 );
and \U$5439 ( \14546 , RIfc55c40_5998, \9464 );
and \U$5440 ( \14547 , RIfca2ab8_6873, \9466 );
and \U$5441 ( \14548 , RIe1fb450_4236, \9468 );
and \U$5442 ( \14549 , RIf156890_5444, \9470 );
and \U$5443 ( \14550 , RIfcd5ff8_7457, \9472 );
and \U$5444 ( \14551 , RIf154dd8_5425, \9474 );
and \U$5445 ( \14552 , RIfec2aa8_8335, \9476 );
and \U$5446 ( \14553 , RIfcb4b00_7078, \9478 );
and \U$5447 ( \14554 , RIfcd9400_7494, \9480 );
and \U$5448 ( \14555 , RIf151160_5382, \9482 );
and \U$5449 ( \14556 , RIe1f4808_4159, \9484 );
and \U$5450 ( \14557 , RIfc44738_5801, \9486 );
and \U$5451 ( \14558 , RIfc90908_6667, \9488 );
and \U$5452 ( \14559 , RIf14e5c8_5351, \9490 );
and \U$5453 ( \14560 , RIe1ef510_4100, \9492 );
and \U$5454 ( \14561 , RIe1ecf18_4073, \9494 );
and \U$5455 ( \14562 , RIe1ea218_4041, \9496 );
and \U$5456 ( \14563 , RIe1e7518_4009, \9498 );
and \U$5457 ( \14564 , RIe1e4818_3977, \9500 );
and \U$5458 ( \14565 , RIe1e1b18_3945, \9502 );
and \U$5459 ( \14566 , RIe1dee18_3913, \9504 );
and \U$5460 ( \14567 , RIe1dc118_3881, \9506 );
and \U$5461 ( \14568 , RIe1d9418_3849, \9508 );
and \U$5462 ( \14569 , RIe1d3a18_3785, \9510 );
and \U$5463 ( \14570 , RIe1d0d18_3753, \9512 );
and \U$5464 ( \14571 , RIe1ce018_3721, \9514 );
and \U$5465 ( \14572 , RIe1cb318_3689, \9516 );
and \U$5466 ( \14573 , RIe1c8618_3657, \9518 );
and \U$5467 ( \14574 , RIe1c5918_3625, \9520 );
and \U$5468 ( \14575 , RIe1c2c18_3593, \9522 );
and \U$5469 ( \14576 , RIe1bff18_3561, \9524 );
and \U$5470 ( \14577 , RIf14d218_5337, \9526 );
and \U$5471 ( \14578 , RIfe8ee60_7970, \9528 );
and \U$5472 ( \14579 , RIfea8090_8228, \9530 );
and \U$5473 ( \14580 , RIe1b84c0_3474, \9532 );
and \U$5474 ( \14581 , RIf14aab8_5309, \9534 );
and \U$5475 ( \14582 , RIfc6c170_6252, \9536 );
and \U$5476 ( \14583 , RIe1b6468_3451, \9538 );
and \U$5477 ( \14584 , RIe1b49b0_3432, \9540 );
and \U$5478 ( \14585 , RIfcafad8_7021, \9542 );
and \U$5479 ( \14586 , RIfcaa948_6963, \9544 );
and \U$5480 ( \14587 , RIfe8ecf8_7969, \9546 );
and \U$5481 ( \14588 , RIfe8f400_7974, \9548 );
and \U$5482 ( \14589 , RIfc67f58_6205, \9550 );
and \U$5483 ( \14590 , RIfca8ff8_6945, \9552 );
and \U$5484 ( \14591 , RIfe8eb90_7968, \9554 );
and \U$5485 ( \14592 , RIe1abe78_3333, \9556 );
and \U$5486 ( \14593 , RIe1aa258_3313, \9558 );
and \U$5487 ( \14594 , RIe1a7558_3281, \9560 );
and \U$5488 ( \14595 , RIe1a4858_3249, \9562 );
and \U$5489 ( \14596 , RIe1a1b58_3217, \9564 );
and \U$5490 ( \14597 , RIe18e058_2993, \9566 );
and \U$5491 ( \14598 , RIe17a558_2769, \9568 );
and \U$5492 ( \14599 , RIe227eb0_4744, \9570 );
and \U$5493 ( \14600 , RIe21cab0_4616, \9572 );
and \U$5494 ( \14601 , RIe2062b0_4360, \9574 );
and \U$5495 ( \14602 , RIe200310_4292, \9576 );
and \U$5496 ( \14603 , RIe1f96c8_4215, \9578 );
and \U$5497 ( \14604 , RIe1f2210_4132, \9580 );
and \U$5498 ( \14605 , RIe1d6718_3817, \9582 );
and \U$5499 ( \14606 , RIe1bd218_3529, \9584 );
and \U$5500 ( \14607 , RIe1b0090_3380, \9586 );
and \U$5501 ( \14608 , RIe1726c8_2679, \9588 );
or \U$5502 ( \14609 , \14545 , \14546 , \14547 , \14548 , \14549 , \14550 , \14551 , \14552 , \14553 , \14554 , \14555 , \14556 , \14557 , \14558 , \14559 , \14560 , \14561 , \14562 , \14563 , \14564 , \14565 , \14566 , \14567 , \14568 , \14569 , \14570 , \14571 , \14572 , \14573 , \14574 , \14575 , \14576 , \14577 , \14578 , \14579 , \14580 , \14581 , \14582 , \14583 , \14584 , \14585 , \14586 , \14587 , \14588 , \14589 , \14590 , \14591 , \14592 , \14593 , \14594 , \14595 , \14596 , \14597 , \14598 , \14599 , \14600 , \14601 , \14602 , \14603 , \14604 , \14605 , \14606 , \14607 , \14608 );
or \U$5503 ( \14610 , \14544 , \14609 );
_DC g3f55 ( \14611_nG3f55 , \14610 , \9597 );
buf \U$5504 ( \14612 , \14611_nG3f55 );
and \U$5505 ( \14613 , \14479 , \14612 );
and \U$5506 ( \14614 , \12951 , \13084 );
and \U$5507 ( \14615 , \13084 , \13359 );
and \U$5508 ( \14616 , \12951 , \13359 );
or \U$5509 ( \14617 , \14614 , \14615 , \14616 );
and \U$5510 ( \14618 , \14612 , \14617 );
and \U$5511 ( \14619 , \14479 , \14617 );
or \U$5512 ( \14620 , \14613 , \14618 , \14619 );
xor \U$5513 ( \14621 , \14346 , \14620 );
buf g443c ( \14622_nG443c , \14621 );
xor \U$5514 ( \14623 , \14479 , \14612 );
xor \U$5515 ( \14624 , \14623 , \14617 );
buf g443f ( \14625_nG443f , \14624 );
nand \U$5516 ( \14626 , \14625_nG443f , \13361_nG4442 );
and \U$5517 ( \14627 , \14622_nG443c , \14626 );
xor \U$5518 ( \14628 , \14625_nG443f , \13361_nG4442 );
not \U$5519 ( \14629 , \14628 );
xor \U$5520 ( \14630 , \14622_nG443c , \14625_nG443f );
and \U$5521 ( \14631 , \14629 , \14630 );
and \U$5523 ( \14632 , \14628 , \10694_nG9c0e );
or \U$5524 ( \14633 , 1'b0 , \14632 );
xor \U$5525 ( \14634 , \14627 , \14633 );
xor \U$5526 ( \14635 , \14627 , \14634 );
buf \U$5527 ( \14636 , \14635 );
buf \U$5528 ( \14637 , \14636 );
and \U$5529 ( \14638 , \14079 , \14637 );
and \U$5530 ( \14639 , \13721 , \13726 );
and \U$5531 ( \14640 , \13721 , \14077 );
and \U$5532 ( \14641 , \13726 , \14077 );
or \U$5533 ( \14642 , \14639 , \14640 , \14641 );
buf \U$5534 ( \14643 , \14642 );
and \U$5535 ( \14644 , \13730 , \13736 );
buf \U$5536 ( \14645 , \14644 );
and \U$5537 ( \14646 , \13370 , \10995_nG9c0b );
and \U$5538 ( \14647 , \13367 , \11283_nG9c08 );
or \U$5539 ( \14648 , \14646 , \14647 );
xor \U$5540 ( \14649 , \13366 , \14648 );
buf \U$5541 ( \14650 , \14649 );
buf \U$5543 ( \14651 , \14650 );
xor \U$5544 ( \14652 , \14645 , \14651 );
buf \U$5545 ( \14653 , \14652 );
and \U$5546 ( \14654 , \12157 , \11598_nG9c05 );
and \U$5547 ( \14655 , \12154 , \12470_nG9c02 );
or \U$5548 ( \14656 , \14654 , \14655 );
xor \U$5549 ( \14657 , \12153 , \14656 );
buf \U$5550 ( \14658 , \14657 );
buf \U$5552 ( \14659 , \14658 );
xor \U$5553 ( \14660 , \14653 , \14659 );
and \U$5554 ( \14661 , \10421 , \12801_nG9bff );
and \U$5555 ( \14662 , \10418 , \13705_nG9bfc );
or \U$5556 ( \14663 , \14661 , \14662 );
xor \U$5557 ( \14664 , \10417 , \14663 );
buf \U$5558 ( \14665 , \14664 );
buf \U$5560 ( \14666 , \14665 );
xor \U$5561 ( \14667 , \14660 , \14666 );
buf \U$5562 ( \14668 , \14667 );
and \U$5563 ( \14669 , \13738 , \13744 );
and \U$5564 ( \14670 , \13738 , \13751 );
and \U$5565 ( \14671 , \13744 , \13751 );
or \U$5566 ( \14672 , \14669 , \14670 , \14671 );
buf \U$5567 ( \14673 , \14672 );
xor \U$5568 ( \14674 , \14668 , \14673 );
and \U$5569 ( \14675 , \10707 , \14070_nG9bf9 );
and \U$5570 ( \14676 , \14037 , \14041 );
and \U$5571 ( \14677 , \14041 , \14059 );
and \U$5572 ( \14678 , \14037 , \14059 );
or \U$5573 ( \14679 , \14676 , \14677 , \14678 );
and \U$5574 ( \14680 , \14046 , \14050 );
and \U$5575 ( \14681 , \14050 , \14058 );
and \U$5576 ( \14682 , \14046 , \14058 );
or \U$5577 ( \14683 , \14680 , \14681 , \14682 );
and \U$5578 ( \14684 , \14024 , \10983 );
and \U$5579 ( \14685 , RIdec6bc0_725, \9333 );
and \U$5580 ( \14686 , RIdec3ec0_693, \9335 );
and \U$5581 ( \14687 , RIee20a58_4830, \9337 );
and \U$5582 ( \14688 , RIdec11c0_661, \9339 );
and \U$5583 ( \14689 , RIee1f978_4818, \9341 );
and \U$5584 ( \14690 , RIdebe4c0_629, \9343 );
and \U$5585 ( \14691 , RIdebb7c0_597, \9345 );
and \U$5586 ( \14692 , RIdeb8ac0_565, \9347 );
and \U$5587 ( \14693 , RIee1efa0_4811, \9349 );
and \U$5588 ( \14694 , RIdeb30c0_501, \9351 );
and \U$5589 ( \14695 , RIfcb04b0_7028, \9353 );
and \U$5590 ( \14696 , RIdeb03c0_469, \9355 );
and \U$5591 ( \14697 , RIfc5e4a8_6095, \9357 );
and \U$5592 ( \14698 , RIdead6c0_437, \9359 );
and \U$5593 ( \14699 , RIdea72e8_405, \9361 );
and \U$5594 ( \14700 , RIdea09e8_373, \9363 );
and \U$5595 ( \14701 , RIfcb2508_7051, \9365 );
and \U$5596 ( \14702 , RIfcd16d8_7405, \9367 );
and \U$5597 ( \14703 , RIfc5d800_6086, \9369 );
and \U$5598 ( \14704 , RIfc63d40_6158, \9371 );
and \U$5599 ( \14705 , RIde93b30_310, \9373 );
and \U$5600 ( \14706 , RIfea7820_8222, \9375 );
and \U$5601 ( \14707 , RIfea73e8_8219, \9377 );
and \U$5602 ( \14708 , RIde87998_251, \9379 );
and \U$5603 ( \14709 , RIde837f8_231, \9381 );
and \U$5604 ( \14710 , RIfc7bd28_6431, \9383 );
and \U$5605 ( \14711 , RIfcc7ef8_7297, \9385 );
and \U$5606 ( \14712 , RIfc7a108_6411, \9387 );
and \U$5607 ( \14713 , RIfc7a6a8_6415, \9389 );
and \U$5608 ( \14714 , RIe16ccc8_2615, \9391 );
and \U$5609 ( \14715 , RIe16a838_2589, \9393 );
and \U$5610 ( \14716 , RIe1691b8_2573, \9395 );
and \U$5611 ( \14717 , RIe166bc0_2546, \9397 );
and \U$5612 ( \14718 , RIe163ec0_2514, \9399 );
and \U$5613 ( \14719 , RIee38338_5098, \9401 );
and \U$5614 ( \14720 , RIe1611c0_2482, \9403 );
and \U$5615 ( \14721 , RIfc54b60_5986, \9405 );
and \U$5616 ( \14722 , RIe15e4c0_2450, \9407 );
and \U$5617 ( \14723 , RIe158ac0_2386, \9409 );
and \U$5618 ( \14724 , RIe155dc0_2354, \9411 );
and \U$5619 ( \14725 , RIee35a70_5069, \9413 );
and \U$5620 ( \14726 , RIe1530c0_2322, \9415 );
and \U$5621 ( \14727 , RIee357a0_5067, \9417 );
and \U$5622 ( \14728 , RIe1503c0_2290, \9419 );
and \U$5623 ( \14729 , RIfc9fdb8_6841, \9421 );
and \U$5624 ( \14730 , RIe14d6c0_2258, \9423 );
and \U$5625 ( \14731 , RIe14a9c0_2226, \9425 );
and \U$5626 ( \14732 , RIe147cc0_2194, \9427 );
and \U$5627 ( \14733 , RIee34af8_5058, \9429 );
and \U$5628 ( \14734 , RIee33a18_5046, \9431 );
and \U$5629 ( \14735 , RIee327d0_5033, \9433 );
and \U$5630 ( \14736 , RIfcbcf30_7172, \9435 );
and \U$5631 ( \14737 , RIe142428_2131, \9437 );
and \U$5632 ( \14738 , RIe140100_2106, \9439 );
and \U$5633 ( \14739 , RIfea7280_8218, \9441 );
and \U$5634 ( \14740 , RIdf3bb78_2056, \9443 );
and \U$5635 ( \14741 , RIfc731f0_6332, \9445 );
and \U$5636 ( \14742 , RIee30610_5009, \9447 );
and \U$5637 ( \14743 , RIfcbe010_7184, \9449 );
and \U$5638 ( \14744 , RIee2e450_4985, \9451 );
and \U$5639 ( \14745 , RIfec2ee0_8338, \9453 );
and \U$5640 ( \14746 , RIfec3048_8339, \9455 );
and \U$5641 ( \14747 , RIfec2c10_8336, \9457 );
and \U$5642 ( \14748 , RIfec2d78_8337, \9459 );
or \U$5643 ( \14749 , \14685 , \14686 , \14687 , \14688 , \14689 , \14690 , \14691 , \14692 , \14693 , \14694 , \14695 , \14696 , \14697 , \14698 , \14699 , \14700 , \14701 , \14702 , \14703 , \14704 , \14705 , \14706 , \14707 , \14708 , \14709 , \14710 , \14711 , \14712 , \14713 , \14714 , \14715 , \14716 , \14717 , \14718 , \14719 , \14720 , \14721 , \14722 , \14723 , \14724 , \14725 , \14726 , \14727 , \14728 , \14729 , \14730 , \14731 , \14732 , \14733 , \14734 , \14735 , \14736 , \14737 , \14738 , \14739 , \14740 , \14741 , \14742 , \14743 , \14744 , \14745 , \14746 , \14747 , \14748 );
and \U$5644 ( \14750 , RIfcb46c8_7075, \9462 );
and \U$5645 ( \14751 , RIfcb4830_7076, \9464 );
and \U$5646 ( \14752 , RIee29860_4931, \9466 );
and \U$5647 ( \14753 , RIfcb88e0_7122, \9468 );
and \U$5648 ( \14754 , RIdf2b480_1869, \9470 );
and \U$5649 ( \14755 , RIdf29590_1847, \9472 );
and \U$5650 ( \14756 , RIdf27268_1822, \9474 );
and \U$5651 ( \14757 , RIdf25648_1802, \9476 );
and \U$5652 ( \14758 , RIfcc9de8_7319, \9478 );
and \U$5653 ( \14759 , RIfc53648_5971, \9480 );
and \U$5654 ( \14760 , RIdf23a28_1782, \9482 );
and \U$5655 ( \14761 , RIfc823d0_6504, \9484 );
and \U$5656 ( \14762 , RIdf223a8_1766, \9486 );
and \U$5657 ( \14763 , RIdf20d28_1750, \9488 );
and \U$5658 ( \14764 , RIdf1bd00_1693, \9490 );
and \U$5659 ( \14765 , RIdf1a7e8_1678, \9492 );
and \U$5660 ( \14766 , RIdf18790_1655, \9494 );
and \U$5661 ( \14767 , RIdf15a90_1623, \9496 );
and \U$5662 ( \14768 , RIdf12d90_1591, \9498 );
and \U$5663 ( \14769 , RIdf10090_1559, \9500 );
and \U$5664 ( \14770 , RIdf0d390_1527, \9502 );
and \U$5665 ( \14771 , RIdf0a690_1495, \9504 );
and \U$5666 ( \14772 , RIdf07990_1463, \9506 );
and \U$5667 ( \14773 , RIdf04c90_1431, \9508 );
and \U$5668 ( \14774 , RIdeff290_1367, \9510 );
and \U$5669 ( \14775 , RIdefc590_1335, \9512 );
and \U$5670 ( \14776 , RIdef9890_1303, \9514 );
and \U$5671 ( \14777 , RIdef6b90_1271, \9516 );
and \U$5672 ( \14778 , RIdef3e90_1239, \9518 );
and \U$5673 ( \14779 , RIdef1190_1207, \9520 );
and \U$5674 ( \14780 , RIdeee490_1175, \9522 );
and \U$5675 ( \14781 , RIdeeb790_1143, \9524 );
and \U$5676 ( \14782 , RIee25be8_4888, \9526 );
and \U$5677 ( \14783 , RIfc6af28_6239, \9528 );
and \U$5678 ( \14784 , RIee23fc8_4868, \9530 );
and \U$5679 ( \14785 , RIfccf680_7382, \9532 );
and \U$5680 ( \14786 , RIdee5d90_1079, \9534 );
and \U$5681 ( \14787 , RIdee4008_1058, \9536 );
and \U$5682 ( \14788 , RIdee1ce0_1033, \9538 );
and \U$5683 ( \14789 , RIdedfdf0_1011, \9540 );
and \U$5684 ( \14790 , RIfc6b090_6240, \9542 );
and \U$5685 ( \14791 , RIfc534e0_5970, \9544 );
and \U$5686 ( \14792 , RIfca5920_6906, \9546 );
and \U$5687 ( \14793 , RIfc66770_6188, \9548 );
and \U$5688 ( \14794 , RIfe8f6d0_7976, \9550 );
and \U$5689 ( \14795 , RIded87d0_927, \9552 );
and \U$5690 ( \14796 , RIfe8f568_7975, \9554 );
and \U$5691 ( \14797 , RIded42e8_878, \9556 );
and \U$5692 ( \14798 , RIded1fc0_853, \9558 );
and \U$5693 ( \14799 , RIdecf2c0_821, \9560 );
and \U$5694 ( \14800 , RIdecc5c0_789, \9562 );
and \U$5695 ( \14801 , RIdec98c0_757, \9564 );
and \U$5696 ( \14802 , RIdeb5dc0_533, \9566 );
and \U$5697 ( \14803 , RIde9a0e8_341, \9568 );
and \U$5698 ( \14804 , RIe16f9c8_2647, \9570 );
and \U$5699 ( \14805 , RIe15b7c0_2418, \9572 );
and \U$5700 ( \14806 , RIe144fc0_2162, \9574 );
and \U$5701 ( \14807 , RIdf399b8_2032, \9576 );
and \U$5702 ( \14808 , RIdf2e018_1900, \9578 );
and \U$5703 ( \14809 , RIdf1e898_1724, \9580 );
and \U$5704 ( \14810 , RIdf01f90_1399, \9582 );
and \U$5705 ( \14811 , RIdee8a90_1111, \9584 );
and \U$5706 ( \14812 , RIdedd7f8_984, \9586 );
and \U$5707 ( \14813 , RIde80030_214, \9588 );
or \U$5708 ( \14814 , \14750 , \14751 , \14752 , \14753 , \14754 , \14755 , \14756 , \14757 , \14758 , \14759 , \14760 , \14761 , \14762 , \14763 , \14764 , \14765 , \14766 , \14767 , \14768 , \14769 , \14770 , \14771 , \14772 , \14773 , \14774 , \14775 , \14776 , \14777 , \14778 , \14779 , \14780 , \14781 , \14782 , \14783 , \14784 , \14785 , \14786 , \14787 , \14788 , \14789 , \14790 , \14791 , \14792 , \14793 , \14794 , \14795 , \14796 , \14797 , \14798 , \14799 , \14800 , \14801 , \14802 , \14803 , \14804 , \14805 , \14806 , \14807 , \14808 , \14809 , \14810 , \14811 , \14812 , \14813 );
or \U$5709 ( \14815 , \14749 , \14814 );
_DC g658f ( \14816_nG658f , \14815 , \9597 );
and \U$5710 ( \14817 , RIe19ee58_3185, \9059 );
and \U$5711 ( \14818 , RIe19c158_3153, \9061 );
and \U$5712 ( \14819 , RIf145bf8_5253, \9063 );
and \U$5713 ( \14820 , RIe199458_3121, \9065 );
and \U$5714 ( \14821 , RIfe8f298_7973, \9067 );
and \U$5715 ( \14822 , RIe196758_3089, \9069 );
and \U$5716 ( \14823 , RIe193a58_3057, \9071 );
and \U$5717 ( \14824 , RIe190d58_3025, \9073 );
and \U$5718 ( \14825 , RIe18b358_2961, \9075 );
and \U$5719 ( \14826 , RIe188658_2929, \9077 );
and \U$5720 ( \14827 , RIfe8f130_7972, \9079 );
and \U$5721 ( \14828 , RIe185958_2897, \9081 );
and \U$5722 ( \14829 , RIfc9f278_6833, \9083 );
and \U$5723 ( \14830 , RIe182c58_2865, \9085 );
and \U$5724 ( \14831 , RIe17ff58_2833, \9087 );
and \U$5725 ( \14832 , RIe17d258_2801, \9089 );
and \U$5726 ( \14833 , RIf1427f0_5216, \9091 );
and \U$5727 ( \14834 , RIfe8efc8_7971, \9093 );
and \U$5728 ( \14835 , RIe1779c0_2738, \9095 );
and \U$5729 ( \14836 , RIe1768e0_2726, \9097 );
and \U$5730 ( \14837 , RIfc81e30_6500, \9099 );
and \U$5731 ( \14838 , RIfc9ff20_6842, \9101 );
and \U$5732 ( \14839 , RIfca0088_6843, \9103 );
and \U$5733 ( \14840 , RIfc81b60_6498, \9105 );
and \U$5734 ( \14841 , RIfce5778_7633, \9107 );
and \U$5735 ( \14842 , RIfce08b8_7577, \9109 );
and \U$5736 ( \14843 , RIfc815c0_6494, \9111 );
and \U$5737 ( \14844 , RIe174cc0_2706, \9113 );
and \U$5738 ( \14845 , RIfca04c0_6846, \9115 );
and \U$5739 ( \14846 , RIfc53eb8_5977, \9117 );
and \U$5740 ( \14847 , RIfcc65a8_7279, \9119 );
and \U$5741 ( \14848 , RIfc80d50_6488, \9121 );
and \U$5742 ( \14849 , RIfc804e0_6482, \9123 );
and \U$5743 ( \14850 , RIe2251b0_4712, \9125 );
and \U$5744 ( \14851 , RIfc80378_6481, \9127 );
and \U$5745 ( \14852 , RIe2224b0_4680, \9129 );
and \U$5746 ( \14853 , RIfcb5910_7088, \9131 );
and \U$5747 ( \14854 , RIe21f7b0_4648, \9133 );
and \U$5748 ( \14855 , RIe219db0_4584, \9135 );
and \U$5749 ( \14856 , RIe2170b0_4552, \9137 );
and \U$5750 ( \14857 , RIfca01f0_6844, \9139 );
and \U$5751 ( \14858 , RIe2143b0_4520, \9141 );
and \U$5752 ( \14859 , RIfc82c40_6510, \9143 );
and \U$5753 ( \14860 , RIe2116b0_4488, \9145 );
and \U$5754 ( \14861 , RIfc7f6d0_6472, \9147 );
and \U$5755 ( \14862 , RIe20e9b0_4456, \9149 );
and \U$5756 ( \14863 , RIe20bcb0_4424, \9151 );
and \U$5757 ( \14864 , RIe208fb0_4392, \9153 );
and \U$5758 ( \14865 , RIf167528_5635, \9155 );
and \U$5759 ( \14866 , RIf1665b0_5624, \9157 );
and \U$5760 ( \14867 , RIe203718_4329, \9159 );
and \U$5761 ( \14868 , RIe201c60_4310, \9161 );
and \U$5762 ( \14869 , RIfc9da90_6816, \9163 );
and \U$5763 ( \14870 , RIfcc5360_7266, \9165 );
and \U$5764 ( \14871 , RIf163748_5591, \9167 );
and \U$5765 ( \14872 , RIf162668_5579, \9169 );
and \U$5766 ( \14873 , RIfc7e320_6458, \9171 );
and \U$5767 ( \14874 , RIfc87998_6565, \9173 );
and \U$5768 ( \14875 , RIe1fd610_4260, \9175 );
and \U$5769 ( \14876 , RIe1fc3c8_4247, \9177 );
and \U$5770 ( \14877 , RIf15d370_5520, \9179 );
and \U$5771 ( \14878 , RIf15c128_5507, \9181 );
and \U$5772 ( \14879 , RIfcc5d38_7273, \9183 );
and \U$5773 ( \14880 , RIfce7d70_7660, \9185 );
or \U$5774 ( \14881 , \14817 , \14818 , \14819 , \14820 , \14821 , \14822 , \14823 , \14824 , \14825 , \14826 , \14827 , \14828 , \14829 , \14830 , \14831 , \14832 , \14833 , \14834 , \14835 , \14836 , \14837 , \14838 , \14839 , \14840 , \14841 , \14842 , \14843 , \14844 , \14845 , \14846 , \14847 , \14848 , \14849 , \14850 , \14851 , \14852 , \14853 , \14854 , \14855 , \14856 , \14857 , \14858 , \14859 , \14860 , \14861 , \14862 , \14863 , \14864 , \14865 , \14866 , \14867 , \14868 , \14869 , \14870 , \14871 , \14872 , \14873 , \14874 , \14875 , \14876 , \14877 , \14878 , \14879 , \14880 );
and \U$5775 ( \14882 , RIfc4bd58_5885, \9188 );
and \U$5776 ( \14883 , RIfc55c40_5998, \9190 );
and \U$5777 ( \14884 , RIfca2ab8_6873, \9192 );
and \U$5778 ( \14885 , RIe1fb450_4236, \9194 );
and \U$5779 ( \14886 , RIf156890_5444, \9196 );
and \U$5780 ( \14887 , RIfcd5ff8_7457, \9198 );
and \U$5781 ( \14888 , RIf154dd8_5425, \9200 );
and \U$5782 ( \14889 , RIfec2aa8_8335, \9202 );
and \U$5783 ( \14890 , RIfcb4b00_7078, \9204 );
and \U$5784 ( \14891 , RIfcd9400_7494, \9206 );
and \U$5785 ( \14892 , RIf151160_5382, \9208 );
and \U$5786 ( \14893 , RIe1f4808_4159, \9210 );
and \U$5787 ( \14894 , RIfc44738_5801, \9212 );
and \U$5788 ( \14895 , RIfc90908_6667, \9214 );
and \U$5789 ( \14896 , RIf14e5c8_5351, \9216 );
and \U$5790 ( \14897 , RIe1ef510_4100, \9218 );
and \U$5791 ( \14898 , RIe1ecf18_4073, \9220 );
and \U$5792 ( \14899 , RIe1ea218_4041, \9222 );
and \U$5793 ( \14900 , RIe1e7518_4009, \9224 );
and \U$5794 ( \14901 , RIe1e4818_3977, \9226 );
and \U$5795 ( \14902 , RIe1e1b18_3945, \9228 );
and \U$5796 ( \14903 , RIe1dee18_3913, \9230 );
and \U$5797 ( \14904 , RIe1dc118_3881, \9232 );
and \U$5798 ( \14905 , RIe1d9418_3849, \9234 );
and \U$5799 ( \14906 , RIe1d3a18_3785, \9236 );
and \U$5800 ( \14907 , RIe1d0d18_3753, \9238 );
and \U$5801 ( \14908 , RIe1ce018_3721, \9240 );
and \U$5802 ( \14909 , RIe1cb318_3689, \9242 );
and \U$5803 ( \14910 , RIe1c8618_3657, \9244 );
and \U$5804 ( \14911 , RIe1c5918_3625, \9246 );
and \U$5805 ( \14912 , RIe1c2c18_3593, \9248 );
and \U$5806 ( \14913 , RIe1bff18_3561, \9250 );
and \U$5807 ( \14914 , RIf14d218_5337, \9252 );
and \U$5808 ( \14915 , RIfe8ee60_7970, \9254 );
and \U$5809 ( \14916 , RIfea8090_8228, \9256 );
and \U$5810 ( \14917 , RIe1b84c0_3474, \9258 );
and \U$5811 ( \14918 , RIf14aab8_5309, \9260 );
and \U$5812 ( \14919 , RIfc6c170_6252, \9262 );
and \U$5813 ( \14920 , RIe1b6468_3451, \9264 );
and \U$5814 ( \14921 , RIe1b49b0_3432, \9266 );
and \U$5815 ( \14922 , RIfcafad8_7021, \9268 );
and \U$5816 ( \14923 , RIfcaa948_6963, \9270 );
and \U$5817 ( \14924 , RIfe8ecf8_7969, \9272 );
and \U$5818 ( \14925 , RIfe8f400_7974, \9274 );
and \U$5819 ( \14926 , RIfc67f58_6205, \9276 );
and \U$5820 ( \14927 , RIfca8ff8_6945, \9278 );
and \U$5821 ( \14928 , RIfe8eb90_7968, \9280 );
and \U$5822 ( \14929 , RIe1abe78_3333, \9282 );
and \U$5823 ( \14930 , RIe1aa258_3313, \9284 );
and \U$5824 ( \14931 , RIe1a7558_3281, \9286 );
and \U$5825 ( \14932 , RIe1a4858_3249, \9288 );
and \U$5826 ( \14933 , RIe1a1b58_3217, \9290 );
and \U$5827 ( \14934 , RIe18e058_2993, \9292 );
and \U$5828 ( \14935 , RIe17a558_2769, \9294 );
and \U$5829 ( \14936 , RIe227eb0_4744, \9296 );
and \U$5830 ( \14937 , RIe21cab0_4616, \9298 );
and \U$5831 ( \14938 , RIe2062b0_4360, \9300 );
and \U$5832 ( \14939 , RIe200310_4292, \9302 );
and \U$5833 ( \14940 , RIe1f96c8_4215, \9304 );
and \U$5834 ( \14941 , RIe1f2210_4132, \9306 );
and \U$5835 ( \14942 , RIe1d6718_3817, \9308 );
and \U$5836 ( \14943 , RIe1bd218_3529, \9310 );
and \U$5837 ( \14944 , RIe1b0090_3380, \9312 );
and \U$5838 ( \14945 , RIe1726c8_2679, \9314 );
or \U$5839 ( \14946 , \14882 , \14883 , \14884 , \14885 , \14886 , \14887 , \14888 , \14889 , \14890 , \14891 , \14892 , \14893 , \14894 , \14895 , \14896 , \14897 , \14898 , \14899 , \14900 , \14901 , \14902 , \14903 , \14904 , \14905 , \14906 , \14907 , \14908 , \14909 , \14910 , \14911 , \14912 , \14913 , \14914 , \14915 , \14916 , \14917 , \14918 , \14919 , \14920 , \14921 , \14922 , \14923 , \14924 , \14925 , \14926 , \14927 , \14928 , \14929 , \14930 , \14931 , \14932 , \14933 , \14934 , \14935 , \14936 , \14937 , \14938 , \14939 , \14940 , \14941 , \14942 , \14943 , \14944 , \14945 );
or \U$5840 ( \14947 , \14881 , \14946 );
_DC g6590 ( \14948_nG6590 , \14947 , \9323 );
and g6591 ( \14949_nG6591 , \14816_nG658f , \14948_nG6590 );
buf \U$5841 ( \14950 , \14949_nG6591 );
and \U$5842 ( \14951 , \14950 , \10691 );
nor \U$5843 ( \14952 , \14684 , \14951 );
xnor \U$5844 ( \14953 , \14952 , \10980 );
and \U$5845 ( \14954 , \10988 , \14054 );
and \U$5846 ( \14955 , \11270 , \13692 );
nor \U$5847 ( \14956 , \14954 , \14955 );
xnor \U$5848 ( \14957 , \14956 , \14035 );
xor \U$5849 ( \14958 , \14953 , \14957 );
_DC g4d22 ( \14959_nG4d22 , \14815 , \9597 );
_DC g4da6 ( \14960_nG4da6 , \14947 , \9323 );
xor g4da7 ( \14961_nG4da7 , \14959_nG4d22 , \14960_nG4da6 );
buf \U$5850 ( \14962 , \14961_nG4da7 );
xor \U$5851 ( \14963 , \14962 , \14032 );
and \U$5852 ( \14964 , \10687 , \14963 );
xor \U$5853 ( \14965 , \14958 , \14964 );
xor \U$5854 ( \14966 , \14683 , \14965 );
and \U$5855 ( \14967 , \14027 , \14036 );
and \U$5856 ( \14968 , \12769 , \11574 );
and \U$5857 ( \14969 , \13679 , \11278 );
nor \U$5858 ( \14970 , \14968 , \14969 );
xnor \U$5859 ( \14971 , \14970 , \11580 );
xor \U$5860 ( \14972 , \14967 , \14971 );
and \U$5861 ( \14973 , \11586 , \12790 );
and \U$5862 ( \14974 , \12448 , \12461 );
nor \U$5863 ( \14975 , \14973 , \14974 );
xnor \U$5864 ( \14976 , \14975 , \12780 );
xor \U$5865 ( \14977 , \14972 , \14976 );
xor \U$5866 ( \14978 , \14966 , \14977 );
xor \U$5867 ( \14979 , \14679 , \14978 );
and \U$5868 ( \14980 , \14060 , \14064 );
and \U$5869 ( \14981 , \14065 , \14068 );
or \U$5870 ( \14982 , \14980 , \14981 );
xor \U$5871 ( \14983 , \14979 , \14982 );
buf g9bf6 ( \14984_nG9bf6 , \14983 );
and \U$5872 ( \14985 , \10704 , \14984_nG9bf6 );
or \U$5873 ( \14986 , \14675 , \14985 );
xor \U$5874 ( \14987 , \10703 , \14986 );
buf \U$5875 ( \14988 , \14987 );
buf \U$5877 ( \14989 , \14988 );
xor \U$5878 ( \14990 , \14674 , \14989 );
buf \U$5879 ( \14991 , \14990 );
xor \U$5880 ( \14992 , \14643 , \14991 );
and \U$5881 ( \14993 , \13753 , \13755 );
and \U$5882 ( \14994 , \13753 , \14075 );
and \U$5883 ( \14995 , \13755 , \14075 );
or \U$5884 ( \14996 , \14993 , \14994 , \14995 );
buf \U$5885 ( \14997 , \14996 );
xor \U$5886 ( \14998 , \14992 , \14997 );
and \U$5887 ( \14999 , \14079 , \14998 );
and \U$5888 ( \15000 , \14637 , \14998 );
or \U$5889 ( \15001 , \14638 , \14999 , \15000 );
and \U$5890 ( \15002 , \14668 , \14673 );
and \U$5891 ( \15003 , \14668 , \14989 );
and \U$5892 ( \15004 , \14673 , \14989 );
or \U$5893 ( \15005 , \15002 , \15003 , \15004 );
buf \U$5894 ( \15006 , \15005 );
and \U$5895 ( \15007 , \14627 , \14634 );
buf \U$5896 ( \15008 , \15007 );
buf \U$5898 ( \15009 , \15008 );
and \U$5899 ( \15010 , \14631 , \10694_nG9c0e );
and \U$5900 ( \15011 , \14628 , \10995_nG9c0b );
or \U$5901 ( \15012 , \15010 , \15011 );
xor \U$5902 ( \15013 , \14627 , \15012 );
buf \U$5903 ( \15014 , \15013 );
buf \U$5905 ( \15015 , \15014 );
xor \U$5906 ( \15016 , \15009 , \15015 );
buf \U$5907 ( \15017 , \15016 );
and \U$5908 ( \15018 , \13370 , \11283_nG9c08 );
and \U$5909 ( \15019 , \13367 , \11598_nG9c05 );
or \U$5910 ( \15020 , \15018 , \15019 );
xor \U$5911 ( \15021 , \13366 , \15020 );
buf \U$5912 ( \15022 , \15021 );
buf \U$5914 ( \15023 , \15022 );
xor \U$5915 ( \15024 , \15017 , \15023 );
and \U$5916 ( \15025 , \12157 , \12470_nG9c02 );
and \U$5917 ( \15026 , \12154 , \12801_nG9bff );
or \U$5918 ( \15027 , \15025 , \15026 );
xor \U$5919 ( \15028 , \12153 , \15027 );
buf \U$5920 ( \15029 , \15028 );
buf \U$5922 ( \15030 , \15029 );
xor \U$5923 ( \15031 , \15024 , \15030 );
buf \U$5924 ( \15032 , \15031 );
and \U$5925 ( \15033 , \14653 , \14659 );
and \U$5926 ( \15034 , \14653 , \14666 );
and \U$5927 ( \15035 , \14659 , \14666 );
or \U$5928 ( \15036 , \15033 , \15034 , \15035 );
buf \U$5929 ( \15037 , \15036 );
and \U$5930 ( \15038 , \14645 , \14651 );
buf \U$5931 ( \15039 , \15038 );
xor \U$5932 ( \15040 , \15037 , \15039 );
and \U$5933 ( \15041 , \10421 , \13705_nG9bfc );
and \U$5934 ( \15042 , \10418 , \14070_nG9bf9 );
or \U$5935 ( \15043 , \15041 , \15042 );
xor \U$5936 ( \15044 , \10417 , \15043 );
buf \U$5937 ( \15045 , \15044 );
buf \U$5939 ( \15046 , \15045 );
xor \U$5940 ( \15047 , \15040 , \15046 );
buf \U$5941 ( \15048 , \15047 );
xor \U$5942 ( \15049 , \15032 , \15048 );
and \U$5943 ( \15050 , \10707 , \14984_nG9bf6 );
and \U$5944 ( \15051 , \14967 , \14971 );
and \U$5945 ( \15052 , \14971 , \14976 );
and \U$5946 ( \15053 , \14967 , \14976 );
or \U$5947 ( \15054 , \15051 , \15052 , \15053 );
and \U$5948 ( \15055 , \14950 , \10983 );
and \U$5949 ( \15056 , RIdec6d28_726, \9333 );
and \U$5950 ( \15057 , RIdec4028_694, \9335 );
and \U$5951 ( \15058 , RIee20bc0_4831, \9337 );
and \U$5952 ( \15059 , RIdec1328_662, \9339 );
and \U$5953 ( \15060 , RIfcbaed8_7149, \9341 );
and \U$5954 ( \15061 , RIdebe628_630, \9343 );
and \U$5955 ( \15062 , RIdebb928_598, \9345 );
and \U$5956 ( \15063 , RIdeb8c28_566, \9347 );
and \U$5957 ( \15064 , RIfc412b8_5767, \9349 );
and \U$5958 ( \15065 , RIdeb3228_502, \9351 );
and \U$5959 ( \15066 , RIfc9ea08_6827, \9353 );
and \U$5960 ( \15067 , RIdeb0528_470, \9355 );
and \U$5961 ( \15068 , RIee1e028_4800, \9357 );
and \U$5962 ( \15069 , RIdead828_438, \9359 );
and \U$5963 ( \15070 , RIdea7630_406, \9361 );
and \U$5964 ( \15071 , RIdea0d30_374, \9363 );
and \U$5965 ( \15072 , RIfcbac08_7147, \9365 );
and \U$5966 ( \15073 , RIfc55538_5993, \9367 );
and \U$5967 ( \15074 , RIfcba668_7143, \9369 );
and \U$5968 ( \15075 , RIfc4af48_5875, \9371 );
and \U$5969 ( \15076 , RIfe912f0_7996, \9373 );
and \U$5970 ( \15077 , RIfe91458_7997, \9375 );
and \U$5971 ( \15078 , RIde8be80_272, \9377 );
and \U$5972 ( \15079 , RIde87ce0_252, \9379 );
and \U$5973 ( \15080 , RIfc85238_6537, \9381 );
and \U$5974 ( \15081 , RIfc88640_6574, \9383 );
and \U$5975 ( \15082 , RIfcda210_7504, \9385 );
and \U$5976 ( \15083 , RIfcd5788_7451, \9387 );
and \U$5977 ( \15084 , RIee39418_5110, \9389 );
and \U$5978 ( \15085 , RIe16ce30_2616, \9391 );
and \U$5979 ( \15086 , RIfc884d8_6573, \9393 );
and \U$5980 ( \15087 , RIe169320_2574, \9395 );
and \U$5981 ( \15088 , RIe166d28_2547, \9397 );
and \U$5982 ( \15089 , RIe164028_2515, \9399 );
and \U$5983 ( \15090 , RIfe90918_7989, \9401 );
and \U$5984 ( \15091 , RIe161328_2483, \9403 );
and \U$5985 ( \15092 , RIee36880_5079, \9405 );
and \U$5986 ( \15093 , RIe15e628_2451, \9407 );
and \U$5987 ( \15094 , RIe158c28_2387, \9409 );
and \U$5988 ( \15095 , RIe155f28_2355, \9411 );
and \U$5989 ( \15096 , RIfe91188_7995, \9413 );
and \U$5990 ( \15097 , RIe153228_2323, \9415 );
and \U$5991 ( \15098 , RIfe91020_7994, \9417 );
and \U$5992 ( \15099 , RIe150528_2291, \9419 );
and \U$5993 ( \15100 , RIfcda378_7505, \9421 );
and \U$5994 ( \15101 , RIe14d828_2259, \9423 );
and \U$5995 ( \15102 , RIe14ab28_2227, \9425 );
and \U$5996 ( \15103 , RIe147e28_2195, \9427 );
and \U$5997 ( \15104 , RIfe90eb8_7993, \9429 );
and \U$5998 ( \15105 , RIfe90d50_7992, \9431 );
and \U$5999 ( \15106 , RIfcb99c0_7134, \9433 );
and \U$6000 ( \15107 , RIfc9c2a8_6799, \9435 );
and \U$6001 ( \15108 , RIfe90be8_7991, \9437 );
and \U$6002 ( \15109 , RIfe90a80_7990, \9439 );
and \U$6003 ( \15110 , RIdf3e008_2082, \9441 );
and \U$6004 ( \15111 , RIdf3bce0_2057, \9443 );
and \U$6005 ( \15112 , RIfcec690_7712, \9445 );
and \U$6006 ( \15113 , RIee30778_5010, \9447 );
and \U$6007 ( \15114 , RIfc87dd0_6568, \9449 );
and \U$6008 ( \15115 , RIee2e5b8_4986, \9451 );
and \U$6009 ( \15116 , RIdf36e20_2001, \9453 );
and \U$6010 ( \15117 , RIdf346c0_1973, \9455 );
and \U$6011 ( \15118 , RIdf32668_1950, \9457 );
and \U$6012 ( \15119 , RIdf30070_1923, \9459 );
or \U$6013 ( \15120 , \15056 , \15057 , \15058 , \15059 , \15060 , \15061 , \15062 , \15063 , \15064 , \15065 , \15066 , \15067 , \15068 , \15069 , \15070 , \15071 , \15072 , \15073 , \15074 , \15075 , \15076 , \15077 , \15078 , \15079 , \15080 , \15081 , \15082 , \15083 , \15084 , \15085 , \15086 , \15087 , \15088 , \15089 , \15090 , \15091 , \15092 , \15093 , \15094 , \15095 , \15096 , \15097 , \15098 , \15099 , \15100 , \15101 , \15102 , \15103 , \15104 , \15105 , \15106 , \15107 , \15108 , \15109 , \15110 , \15111 , \15112 , \15113 , \15114 , \15115 , \15116 , \15117 , \15118 , \15119 );
and \U$6014 ( \15121 , RIee2c998_4966, \9462 );
and \U$6015 ( \15122 , RIee2aee0_4947, \9464 );
and \U$6016 ( \15123 , RIee299c8_4932, \9466 );
and \U$6017 ( \15124 , RIee28618_4918, \9468 );
and \U$6018 ( \15125 , RIfe90378_7985, \9470 );
and \U$6019 ( \15126 , RIfe907b0_7988, \9472 );
and \U$6020 ( \15127 , RIfe904e0_7986, \9474 );
and \U$6021 ( \15128 , RIfe90648_7987, \9476 );
and \U$6022 ( \15129 , RIfc9d928_6815, \9478 );
and \U$6023 ( \15130 , RIfc86048_6547, \9480 );
and \U$6024 ( \15131 , RIfcb92b8_7129, \9482 );
and \U$6025 ( \15132 , RIfc4ee90_5920, \9484 );
and \U$6026 ( \15133 , RIfc86a20_6554, \9486 );
and \U$6027 ( \15134 , RIdf20e90_1751, \9488 );
and \U$6028 ( \15135 , RIfcb8fe8_7127, \9490 );
and \U$6029 ( \15136 , RIdf1a950_1679, \9492 );
and \U$6030 ( \15137 , RIdf188f8_1656, \9494 );
and \U$6031 ( \15138 , RIdf15bf8_1624, \9496 );
and \U$6032 ( \15139 , RIdf12ef8_1592, \9498 );
and \U$6033 ( \15140 , RIdf101f8_1560, \9500 );
and \U$6034 ( \15141 , RIdf0d4f8_1528, \9502 );
and \U$6035 ( \15142 , RIdf0a7f8_1496, \9504 );
and \U$6036 ( \15143 , RIdf07af8_1464, \9506 );
and \U$6037 ( \15144 , RIdf04df8_1432, \9508 );
and \U$6038 ( \15145 , RIdeff3f8_1368, \9510 );
and \U$6039 ( \15146 , RIdefc6f8_1336, \9512 );
and \U$6040 ( \15147 , RIdef99f8_1304, \9514 );
and \U$6041 ( \15148 , RIdef6cf8_1272, \9516 );
and \U$6042 ( \15149 , RIdef3ff8_1240, \9518 );
and \U$6043 ( \15150 , RIdef12f8_1208, \9520 );
and \U$6044 ( \15151 , RIdeee5f8_1176, \9522 );
and \U$6045 ( \15152 , RIdeeb8f8_1144, \9524 );
and \U$6046 ( \15153 , RIfc857d8_6541, \9526 );
and \U$6047 ( \15154 , RIee24dd8_4878, \9528 );
and \U$6048 ( \15155 , RIfc4ff70_5932, \9530 );
and \U$6049 ( \15156 , RIfc50240_5934, \9532 );
and \U$6050 ( \15157 , RIdee5ef8_1080, \9534 );
and \U$6051 ( \15158 , RIdee4170_1059, \9536 );
and \U$6052 ( \15159 , RIfe915c0_7998, \9538 );
and \U$6053 ( \15160 , RIdedff58_1012, \9540 );
and \U$6054 ( \15161 , RIfcd4810_7440, \9542 );
and \U$6055 ( \15162 , RIee22948_4852, \9544 );
and \U$6056 ( \15163 , RIfce1560_7586, \9546 );
and \U$6057 ( \15164 , RIee219d0_4841, \9548 );
and \U$6058 ( \15165 , RIdedac60_953, \9550 );
and \U$6059 ( \15166 , RIfe91728_7999, \9552 );
and \U$6060 ( \15167 , RIded64a8_902, \9554 );
and \U$6061 ( \15168 , RIfe91890_8000, \9556 );
and \U$6062 ( \15169 , RIded2128_854, \9558 );
and \U$6063 ( \15170 , RIdecf428_822, \9560 );
and \U$6064 ( \15171 , RIdecc728_790, \9562 );
and \U$6065 ( \15172 , RIdec9a28_758, \9564 );
and \U$6066 ( \15173 , RIdeb5f28_534, \9566 );
and \U$6067 ( \15174 , RIde9a430_342, \9568 );
and \U$6068 ( \15175 , RIe16fb30_2648, \9570 );
and \U$6069 ( \15176 , RIe15b928_2419, \9572 );
and \U$6070 ( \15177 , RIe145128_2163, \9574 );
and \U$6071 ( \15178 , RIdf39b20_2033, \9576 );
and \U$6072 ( \15179 , RIdf2e180_1901, \9578 );
and \U$6073 ( \15180 , RIdf1ea00_1725, \9580 );
and \U$6074 ( \15181 , RIdf020f8_1400, \9582 );
and \U$6075 ( \15182 , RIdee8bf8_1112, \9584 );
and \U$6076 ( \15183 , RIdedd960_985, \9586 );
and \U$6077 ( \15184 , RIde80378_215, \9588 );
or \U$6078 ( \15185 , \15121 , \15122 , \15123 , \15124 , \15125 , \15126 , \15127 , \15128 , \15129 , \15130 , \15131 , \15132 , \15133 , \15134 , \15135 , \15136 , \15137 , \15138 , \15139 , \15140 , \15141 , \15142 , \15143 , \15144 , \15145 , \15146 , \15147 , \15148 , \15149 , \15150 , \15151 , \15152 , \15153 , \15154 , \15155 , \15156 , \15157 , \15158 , \15159 , \15160 , \15161 , \15162 , \15163 , \15164 , \15165 , \15166 , \15167 , \15168 , \15169 , \15170 , \15171 , \15172 , \15173 , \15174 , \15175 , \15176 , \15177 , \15178 , \15179 , \15180 , \15181 , \15182 , \15183 , \15184 );
or \U$6079 ( \15186 , \15120 , \15185 );
_DC g6592 ( \15187_nG6592 , \15186 , \9597 );
and \U$6080 ( \15188 , RIe19efc0_3186, \9059 );
and \U$6081 ( \15189 , RIe19c2c0_3154, \9061 );
and \U$6082 ( \15190 , RIf145d60_5254, \9063 );
and \U$6083 ( \15191 , RIe1995c0_3122, \9065 );
and \U$6084 ( \15192 , RIfc637a0_6154, \9067 );
and \U$6085 ( \15193 , RIe1968c0_3090, \9069 );
and \U$6086 ( \15194 , RIe193bc0_3058, \9071 );
and \U$6087 ( \15195 , RIe190ec0_3026, \9073 );
and \U$6088 ( \15196 , RIe18b4c0_2962, \9075 );
and \U$6089 ( \15197 , RIe1887c0_2930, \9077 );
and \U$6090 ( \15198 , RIfc62af8_6145, \9079 );
and \U$6091 ( \15199 , RIe185ac0_2898, \9081 );
and \U$6092 ( \15200 , RIfe8fc70_7980, \9083 );
and \U$6093 ( \15201 , RIe182dc0_2866, \9085 );
and \U$6094 ( \15202 , RIe1800c0_2834, \9087 );
and \U$6095 ( \15203 , RIe17d3c0_2802, \9089 );
and \U$6096 ( \15204 , RIfe90210_7984, \9091 );
and \U$6097 ( \15205 , RIfe8ff40_7982, \9093 );
and \U$6098 ( \15206 , RIfc72f20_6330, \9095 );
and \U$6099 ( \15207 , RIe176a48_2727, \9097 );
and \U$6100 ( \15208 , RIfcaf6a0_7018, \9099 );
and \U$6101 ( \15209 , RIfc61040_6126, \9101 );
and \U$6102 ( \15210 , RIf13e8a8_5171, \9103 );
and \U$6103 ( \15211 , RIfe900a8_7983, \9105 );
and \U$6104 ( \15212 , RIee3caf0_5149, \9107 );
and \U$6105 ( \15213 , RIee3b740_5135, \9109 );
and \U$6106 ( \15214 , RIee3a660_5123, \9111 );
and \U$6107 ( \15215 , RIe174e28_2707, \9113 );
and \U$6108 ( \15216 , RIf170768_5739, \9115 );
and \U$6109 ( \15217 , RIfc5fdf8_6113, \9117 );
and \U$6110 ( \15218 , RIf16eb48_5719, \9119 );
and \U$6111 ( \15219 , RIfcaaab0_6964, \9121 );
and \U$6112 ( \15220 , RIf16d1f8_5701, \9123 );
and \U$6113 ( \15221 , RIe225318_4713, \9125 );
and \U$6114 ( \15222 , RIf16c6b8_5693, \9127 );
and \U$6115 ( \15223 , RIe222618_4681, \9129 );
and \U$6116 ( \15224 , RIf16b5d8_5681, \9131 );
and \U$6117 ( \15225 , RIe21f918_4649, \9133 );
and \U$6118 ( \15226 , RIe219f18_4585, \9135 );
and \U$6119 ( \15227 , RIe217218_4553, \9137 );
and \U$6120 ( \15228 , RIfca62f8_6913, \9139 );
and \U$6121 ( \15229 , RIe214518_4521, \9141 );
and \U$6122 ( \15230 , RIfcc9578_7313, \9143 );
and \U$6123 ( \15231 , RIe211818_4489, \9145 );
and \U$6124 ( \15232 , RIfca5a88_6907, \9147 );
and \U$6125 ( \15233 , RIe20eb18_4457, \9149 );
and \U$6126 ( \15234 , RIe20be18_4425, \9151 );
and \U$6127 ( \15235 , RIe209118_4393, \9153 );
and \U$6128 ( \15236 , RIf167690_5636, \9155 );
and \U$6129 ( \15237 , RIf166718_5625, \9157 );
and \U$6130 ( \15238 , RIfe8f9a0_7978, \9159 );
and \U$6131 ( \15239 , RIfe8f838_7977, \9161 );
and \U$6132 ( \15240 , RIf165638_5613, \9163 );
and \U$6133 ( \15241 , RIf164990_5604, \9165 );
and \U$6134 ( \15242 , RIf1638b0_5592, \9167 );
and \U$6135 ( \15243 , RIf1627d0_5580, \9169 );
and \U$6136 ( \15244 , RIf161150_5564, \9171 );
and \U$6137 ( \15245 , RIf15f260_5542, \9173 );
and \U$6138 ( \15246 , RIe1fd778_4261, \9175 );
and \U$6139 ( \15247 , RIe1fc530_4248, \9177 );
and \U$6140 ( \15248 , RIf15d4d8_5521, \9179 );
and \U$6141 ( \15249 , RIf15c290_5508, \9181 );
and \U$6142 ( \15250 , RIfca20e0_6866, \9183 );
and \U$6143 ( \15251 , RIf159f68_5483, \9185 );
or \U$6144 ( \15252 , \15188 , \15189 , \15190 , \15191 , \15192 , \15193 , \15194 , \15195 , \15196 , \15197 , \15198 , \15199 , \15200 , \15201 , \15202 , \15203 , \15204 , \15205 , \15206 , \15207 , \15208 , \15209 , \15210 , \15211 , \15212 , \15213 , \15214 , \15215 , \15216 , \15217 , \15218 , \15219 , \15220 , \15221 , \15222 , \15223 , \15224 , \15225 , \15226 , \15227 , \15228 , \15229 , \15230 , \15231 , \15232 , \15233 , \15234 , \15235 , \15236 , \15237 , \15238 , \15239 , \15240 , \15241 , \15242 , \15243 , \15244 , \15245 , \15246 , \15247 , \15248 , \15249 , \15250 , \15251 );
and \U$6145 ( \15253 , RIf159428_5475, \9188 );
and \U$6146 ( \15254 , RIf1581e0_5462, \9190 );
and \U$6147 ( \15255 , RIfc5ebb0_6100, \9192 );
and \U$6148 ( \15256 , RIfe8fdd8_7981, \9194 );
and \U$6149 ( \15257 , RIfc69e48_6227, \9196 );
and \U$6150 ( \15258 , RIfc5e8e0_6098, \9198 );
and \U$6151 ( \15259 , RIf154f40_5426, \9200 );
and \U$6152 ( \15260 , RIe1f6b30_4184, \9202 );
and \U$6153 ( \15261 , RIf153b90_5412, \9204 );
and \U$6154 ( \15262 , RIf1523a8_5395, \9206 );
and \U$6155 ( \15263 , RIfce88b0_7668, \9208 );
and \U$6156 ( \15264 , RIfe8fb08_7979, \9210 );
and \U$6157 ( \15265 , RIfcebe20_7706, \9212 );
and \U$6158 ( \15266 , RIfcb1158_7037, \9214 );
and \U$6159 ( \15267 , RIf14e730_5352, \9216 );
and \U$6160 ( \15268 , RIe1ef678_4101, \9218 );
and \U$6161 ( \15269 , RIe1ed080_4074, \9220 );
and \U$6162 ( \15270 , RIe1ea380_4042, \9222 );
and \U$6163 ( \15271 , RIe1e7680_4010, \9224 );
and \U$6164 ( \15272 , RIe1e4980_3978, \9226 );
and \U$6165 ( \15273 , RIe1e1c80_3946, \9228 );
and \U$6166 ( \15274 , RIe1def80_3914, \9230 );
and \U$6167 ( \15275 , RIe1dc280_3882, \9232 );
and \U$6168 ( \15276 , RIe1d9580_3850, \9234 );
and \U$6169 ( \15277 , RIe1d3b80_3786, \9236 );
and \U$6170 ( \15278 , RIe1d0e80_3754, \9238 );
and \U$6171 ( \15279 , RIe1ce180_3722, \9240 );
and \U$6172 ( \15280 , RIe1cb480_3690, \9242 );
and \U$6173 ( \15281 , RIe1c8780_3658, \9244 );
and \U$6174 ( \15282 , RIe1c5a80_3626, \9246 );
and \U$6175 ( \15283 , RIe1c2d80_3594, \9248 );
and \U$6176 ( \15284 , RIe1c0080_3562, \9250 );
and \U$6177 ( \15285 , RIfcc8ba0_7306, \9252 );
and \U$6178 ( \15286 , RIfc5d698_6085, \9254 );
and \U$6179 ( \15287 , RIfec35e8_8343, \9256 );
and \U$6180 ( \15288 , RIfeabd08_8271, \9258 );
and \U$6181 ( \15289 , RIfc5cf90_6080, \9260 );
and \U$6182 ( \15290 , RIfc5ce28_6079, \9262 );
and \U$6183 ( \15291 , RIfec31b0_8340, \9264 );
and \U$6184 ( \15292 , RIe1b4b18_3433, \9266 );
and \U$6185 ( \15293 , RIf149708_5295, \9268 );
and \U$6186 ( \15294 , RIf148358_5281, \9270 );
and \U$6187 ( \15295 , RIe1b3768_3419, \9272 );
and \U$6188 ( \15296 , RIfec3480_8342, \9274 );
and \U$6189 ( \15297 , RIfc483b0_5844, \9276 );
and \U$6190 ( \15298 , RIfc80be8_6487, \9278 );
and \U$6191 ( \15299 , RIe1ad4f8_3349, \9280 );
and \U$6192 ( \15300 , RIfec3318_8341, \9282 );
and \U$6193 ( \15301 , RIe1aa3c0_3314, \9284 );
and \U$6194 ( \15302 , RIe1a76c0_3282, \9286 );
and \U$6195 ( \15303 , RIe1a49c0_3250, \9288 );
and \U$6196 ( \15304 , RIe1a1cc0_3218, \9290 );
and \U$6197 ( \15305 , RIe18e1c0_2994, \9292 );
and \U$6198 ( \15306 , RIe17a6c0_2770, \9294 );
and \U$6199 ( \15307 , RIe228018_4745, \9296 );
and \U$6200 ( \15308 , RIe21cc18_4617, \9298 );
and \U$6201 ( \15309 , RIe206418_4361, \9300 );
and \U$6202 ( \15310 , RIe200478_4293, \9302 );
and \U$6203 ( \15311 , RIe1f9830_4216, \9304 );
and \U$6204 ( \15312 , RIe1f2378_4133, \9306 );
and \U$6205 ( \15313 , RIe1d6880_3818, \9308 );
and \U$6206 ( \15314 , RIe1bd380_3530, \9310 );
and \U$6207 ( \15315 , RIe1b01f8_3381, \9312 );
and \U$6208 ( \15316 , RIe172830_2680, \9314 );
or \U$6209 ( \15317 , \15253 , \15254 , \15255 , \15256 , \15257 , \15258 , \15259 , \15260 , \15261 , \15262 , \15263 , \15264 , \15265 , \15266 , \15267 , \15268 , \15269 , \15270 , \15271 , \15272 , \15273 , \15274 , \15275 , \15276 , \15277 , \15278 , \15279 , \15280 , \15281 , \15282 , \15283 , \15284 , \15285 , \15286 , \15287 , \15288 , \15289 , \15290 , \15291 , \15292 , \15293 , \15294 , \15295 , \15296 , \15297 , \15298 , \15299 , \15300 , \15301 , \15302 , \15303 , \15304 , \15305 , \15306 , \15307 , \15308 , \15309 , \15310 , \15311 , \15312 , \15313 , \15314 , \15315 , \15316 );
or \U$6210 ( \15318 , \15252 , \15317 );
_DC g6593 ( \15319_nG6593 , \15318 , \9323 );
and g6594 ( \15320_nG6594 , \15187_nG6592 , \15319_nG6593 );
buf \U$6211 ( \15321 , \15320_nG6594 );
and \U$6212 ( \15322 , \15321 , \10691 );
nor \U$6213 ( \15323 , \15055 , \15322 );
xnor \U$6214 ( \15324 , \15323 , \10980 );
and \U$6215 ( \15325 , \11270 , \14054 );
and \U$6216 ( \15326 , \11586 , \13692 );
nor \U$6217 ( \15327 , \15325 , \15326 );
xnor \U$6218 ( \15328 , \15327 , \14035 );
xor \U$6219 ( \15329 , \15324 , \15328 );
_DC g4e2b ( \15330_nG4e2b , \15186 , \9597 );
_DC g4eaf ( \15331_nG4eaf , \15318 , \9323 );
xor g4eb0 ( \15332_nG4eb0 , \15330_nG4e2b , \15331_nG4eaf );
buf \U$6220 ( \15333 , \15332_nG4eb0 );
xor \U$6221 ( \15334 , \15333 , \14962 );
not \U$6222 ( \15335 , \14963 );
and \U$6223 ( \15336 , \15334 , \15335 );
and \U$6224 ( \15337 , \10687 , \15336 );
and \U$6225 ( \15338 , \10988 , \14963 );
nor \U$6226 ( \15339 , \15337 , \15338 );
and \U$6227 ( \15340 , \14962 , \14032 );
not \U$6228 ( \15341 , \15340 );
and \U$6229 ( \15342 , \15333 , \15341 );
xnor \U$6230 ( \15343 , \15339 , \15342 );
xor \U$6231 ( \15344 , \15329 , \15343 );
xor \U$6232 ( \15345 , \15054 , \15344 );
and \U$6233 ( \15346 , \13679 , \11574 );
and \U$6234 ( \15347 , \14024 , \11278 );
nor \U$6235 ( \15348 , \15346 , \15347 );
xnor \U$6236 ( \15349 , \15348 , \11580 );
not \U$6237 ( \15350 , \14964 );
and \U$6238 ( \15351 , \15350 , \15342 );
xor \U$6239 ( \15352 , \15349 , \15351 );
and \U$6240 ( \15353 , \14953 , \14957 );
and \U$6241 ( \15354 , \14957 , \14964 );
and \U$6242 ( \15355 , \14953 , \14964 );
or \U$6243 ( \15356 , \15353 , \15354 , \15355 );
xor \U$6244 ( \15357 , \15352 , \15356 );
and \U$6245 ( \15358 , \12448 , \12790 );
and \U$6246 ( \15359 , \12769 , \12461 );
nor \U$6247 ( \15360 , \15358 , \15359 );
xnor \U$6248 ( \15361 , \15360 , \12780 );
xor \U$6249 ( \15362 , \15357 , \15361 );
xor \U$6250 ( \15363 , \15345 , \15362 );
and \U$6251 ( \15364 , \14683 , \14965 );
and \U$6252 ( \15365 , \14965 , \14977 );
and \U$6253 ( \15366 , \14683 , \14977 );
or \U$6254 ( \15367 , \15364 , \15365 , \15366 );
xor \U$6255 ( \15368 , \15363 , \15367 );
and \U$6256 ( \15369 , \14679 , \14978 );
and \U$6257 ( \15370 , \14979 , \14982 );
or \U$6258 ( \15371 , \15369 , \15370 );
xor \U$6259 ( \15372 , \15368 , \15371 );
buf g9bf3 ( \15373_nG9bf3 , \15372 );
and \U$6260 ( \15374 , \10704 , \15373_nG9bf3 );
or \U$6261 ( \15375 , \15050 , \15374 );
xor \U$6262 ( \15376 , \10703 , \15375 );
buf \U$6263 ( \15377 , \15376 );
buf \U$6265 ( \15378 , \15377 );
xor \U$6266 ( \15379 , \15049 , \15378 );
buf \U$6267 ( \15380 , \15379 );
xor \U$6268 ( \15381 , \15006 , \15380 );
and \U$6269 ( \15382 , \14643 , \14991 );
and \U$6270 ( \15383 , \14643 , \14997 );
and \U$6271 ( \15384 , \14991 , \14997 );
or \U$6272 ( \15385 , \15382 , \15383 , \15384 );
buf \U$6273 ( \15386 , \15385 );
xor \U$6274 ( \15387 , \15381 , \15386 );
and \U$6275 ( \15388 , \15001 , \15387 );
and \U$6276 ( \15389 , RIdec4460_697, \9059 );
and \U$6277 ( \15390 , RIdec1760_665, \9061 );
and \U$6278 ( \15391 , RIee1fae0_4819, \9063 );
and \U$6279 ( \15392 , RIdebea60_633, \9065 );
and \U$6280 ( \15393 , RIee1f108_4812, \9067 );
and \U$6281 ( \15394 , RIdebbd60_601, \9069 );
and \U$6282 ( \15395 , RIdeb9060_569, \9071 );
and \U$6283 ( \15396 , RIdeb6360_537, \9073 );
and \U$6284 ( \15397 , RIee1eb68_4808, \9075 );
and \U$6285 ( \15398 , RIdeb0960_473, \9077 );
and \U$6286 ( \15399 , RIee1e460_4803, \9079 );
and \U$6287 ( \15400 , RIdeadc60_441, \9081 );
and \U$6288 ( \15401 , RIee1d7b8_4794, \9083 );
and \U$6289 ( \15402 , RIdea8008_409, \9085 );
and \U$6290 ( \15403 , RIdea1708_377, \9087 );
and \U$6291 ( \15404 , RIde9ae08_345, \9089 );
and \U$6292 ( \15405 , RIfe957d8_8045, \9091 );
and \U$6293 ( \15406 , RIfe95508_8043, \9093 );
and \U$6294 ( \15407 , RIfe95670_8044, \9095 );
and \U$6295 ( \15408 , RIee1a7e8_4760, \9097 );
and \U$6296 ( \15409 , RIfe95aa8_8047, \9099 );
and \U$6297 ( \15410 , RIfe95238_8041, \9101 );
and \U$6298 ( \15411 , RIfe95940_8046, \9103 );
and \U$6299 ( \15412 , RIfe953a0_8042, \9105 );
and \U$6300 ( \15413 , RIee1a0e0_4755, \9107 );
and \U$6301 ( \15414 , RIee19ca8_4752, \9109 );
and \U$6302 ( \15415 , RIee19870_4749, \9111 );
and \U$6303 ( \15416 , RIee19438_4746, \9113 );
and \U$6304 ( \15417 , RIee38ba8_5104, \9115 );
and \U$6305 ( \15418 , RIfe95c10_8048, \9117 );
and \U$6306 ( \15419 , RIee384a0_5099, \9119 );
and \U$6307 ( \15420 , RIfea9440_8242, \9121 );
and \U$6308 ( \15421 , RIe164460_2518, \9123 );
and \U$6309 ( \15422 , RIe161760_2486, \9125 );
and \U$6310 ( \15423 , RIfe942c0_8030, \9127 );
and \U$6311 ( \15424 , RIe15ea60_2454, \9129 );
and \U$6312 ( \15425 , RIfe94158_8029, \9131 );
and \U$6313 ( \15426 , RIe15bd60_2422, \9133 );
and \U$6314 ( \15427 , RIe156360_2358, \9135 );
and \U$6315 ( \15428 , RIe153660_2326, \9137 );
and \U$6316 ( \15429 , RIfe94428_8031, \9139 );
and \U$6317 ( \15430 , RIe150960_2294, \9141 );
and \U$6318 ( \15431 , RIfe94590_8032, \9143 );
and \U$6319 ( \15432 , RIe14dc60_2262, \9145 );
and \U$6320 ( \15433 , RIfc5c2e8_6071, \9147 );
and \U$6321 ( \15434 , RIe14af60_2230, \9149 );
and \U$6322 ( \15435 , RIe148260_2198, \9151 );
and \U$6323 ( \15436 , RIe145560_2166, \9153 );
and \U$6324 ( \15437 , RIee33ce8_5048, \9155 );
and \U$6325 ( \15438 , RIee32aa0_5035, \9157 );
and \U$6326 ( \15439 , RIee31858_5022, \9159 );
and \U$6327 ( \15440 , RIfc5d530_6084, \9161 );
and \U$6328 ( \15441 , RIe140538_2109, \9163 );
and \U$6329 ( \15442 , RIdf3e2d8_2084, \9165 );
and \U$6330 ( \15443 , RIdf3c118_2060, \9167 );
and \U$6331 ( \15444 , RIdf39df0_2035, \9169 );
and \U$6332 ( \15445 , RIfcdd780_7542, \9171 );
and \U$6333 ( \15446 , RIee2ee28_4992, \9173 );
and \U$6334 ( \15447 , RIfcc88d0_7304, \9175 );
and \U$6335 ( \15448 , RIee2cc68_4968, \9177 );
and \U$6336 ( \15449 , RIdf34990_1975, \9179 );
and \U$6337 ( \15450 , RIdf32aa0_1953, \9181 );
and \U$6338 ( \15451 , RIdf304a8_1926, \9183 );
and \U$6339 ( \15452 , RIdf2e5b8_1904, \9185 );
or \U$6340 ( \15453 , \15389 , \15390 , \15391 , \15392 , \15393 , \15394 , \15395 , \15396 , \15397 , \15398 , \15399 , \15400 , \15401 , \15402 , \15403 , \15404 , \15405 , \15406 , \15407 , \15408 , \15409 , \15410 , \15411 , \15412 , \15413 , \15414 , \15415 , \15416 , \15417 , \15418 , \15419 , \15420 , \15421 , \15422 , \15423 , \15424 , \15425 , \15426 , \15427 , \15428 , \15429 , \15430 , \15431 , \15432 , \15433 , \15434 , \15435 , \15436 , \15437 , \15438 , \15439 , \15440 , \15441 , \15442 , \15443 , \15444 , \15445 , \15446 , \15447 , \15448 , \15449 , \15450 , \15451 , \15452 );
and \U$6341 ( \15454 , RIee2b1b0_4949, \9188 );
and \U$6342 ( \15455 , RIfe946f8_8033, \9190 );
and \U$6343 ( \15456 , RIfcb2940_7054, \9192 );
and \U$6344 ( \15457 , RIee273d0_4905, \9194 );
and \U$6345 ( \15458 , RIfe949c8_8035, \9196 );
and \U$6346 ( \15459 , RIdf27538_1824, \9198 );
and \U$6347 ( \15460 , RIfe94b30_8036, \9200 );
and \U$6348 ( \15461 , RIfe94860_8034, \9202 );
and \U$6349 ( \15462 , RIee26f98_4902, \9204 );
and \U$6350 ( \15463 , RIee269f8_4898, \9206 );
and \U$6351 ( \15464 , RIee26728_4896, \9208 );
and \U$6352 ( \15465 , RIee26458_4894, \9210 );
and \U$6353 ( \15466 , RIee26188_4892, \9212 );
and \U$6354 ( \15467 , RIfe94c98_8037, \9214 );
and \U$6355 ( \15468 , RIee25d50_4889, \9216 );
and \U$6356 ( \15469 , RIfea9170_8240, \9218 );
and \U$6357 ( \15470 , RIdf16030_1627, \9220 );
and \U$6358 ( \15471 , RIdf13330_1595, \9222 );
and \U$6359 ( \15472 , RIdf10630_1563, \9224 );
and \U$6360 ( \15473 , RIdf0d930_1531, \9226 );
and \U$6361 ( \15474 , RIdf0ac30_1499, \9228 );
and \U$6362 ( \15475 , RIdf07f30_1467, \9230 );
and \U$6363 ( \15476 , RIdf05230_1435, \9232 );
and \U$6364 ( \15477 , RIdf02530_1403, \9234 );
and \U$6365 ( \15478 , RIdefcb30_1339, \9236 );
and \U$6366 ( \15479 , RIdef9e30_1307, \9238 );
and \U$6367 ( \15480 , RIdef7130_1275, \9240 );
and \U$6368 ( \15481 , RIdef4430_1243, \9242 );
and \U$6369 ( \15482 , RIdef1730_1211, \9244 );
and \U$6370 ( \15483 , RIdeeea30_1179, \9246 );
and \U$6371 ( \15484 , RIdeebd30_1147, \9248 );
and \U$6372 ( \15485 , RIdee9030_1115, \9250 );
and \U$6373 ( \15486 , RIee250a8_4880, \9252 );
and \U$6374 ( \15487 , RIee24298_4870, \9254 );
and \U$6375 ( \15488 , RIee23758_4862, \9256 );
and \U$6376 ( \15489 , RIee22d80_4855, \9258 );
and \U$6377 ( \15490 , RIfe950d0_8040, \9260 );
and \U$6378 ( \15491 , RIfe94f68_8039, \9262 );
and \U$6379 ( \15492 , RIfe94e00_8038, \9264 );
and \U$6380 ( \15493 , RIdeddd98_988, \9266 );
and \U$6381 ( \15494 , RIee22ab0_4853, \9268 );
and \U$6382 ( \15495 , RIee21e08_4844, \9270 );
and \U$6383 ( \15496 , RIfca46d8_6893, \9272 );
and \U$6384 ( \15497 , RIfc5dad0_6088, \9274 );
and \U$6385 ( \15498 , RIfeaa250_8252, \9276 );
and \U$6386 ( \15499 , RIfe96048_8051, \9278 );
and \U$6387 ( \15500 , RIfe95d78_8049, \9280 );
and \U$6388 ( \15501 , RIfe95ee0_8050, \9282 );
and \U$6389 ( \15502 , RIdecf860_825, \9284 );
and \U$6390 ( \15503 , RIdeccb60_793, \9286 );
and \U$6391 ( \15504 , RIdec9e60_761, \9288 );
and \U$6392 ( \15505 , RIdec7160_729, \9290 );
and \U$6393 ( \15506 , RIdeb3660_505, \9292 );
and \U$6394 ( \15507 , RIde94508_313, \9294 );
and \U$6395 ( \15508 , RIe16d268_2619, \9296 );
and \U$6396 ( \15509 , RIe159060_2390, \9298 );
and \U$6397 ( \15510 , RIe142860_2134, \9300 );
and \U$6398 ( \15511 , RIdf37258_2004, \9302 );
and \U$6399 ( \15512 , RIdf2b8b8_1872, \9304 );
and \U$6400 ( \15513 , RIdf1c138_1696, \9306 );
and \U$6401 ( \15514 , RIdeff830_1371, \9308 );
and \U$6402 ( \15515 , RIdee6330_1083, \9310 );
and \U$6403 ( \15516 , RIdedb098_956, \9312 );
and \U$6404 ( \15517 , RIde7a450_186, \9314 );
or \U$6405 ( \15518 , \15454 , \15455 , \15456 , \15457 , \15458 , \15459 , \15460 , \15461 , \15462 , \15463 , \15464 , \15465 , \15466 , \15467 , \15468 , \15469 , \15470 , \15471 , \15472 , \15473 , \15474 , \15475 , \15476 , \15477 , \15478 , \15479 , \15480 , \15481 , \15482 , \15483 , \15484 , \15485 , \15486 , \15487 , \15488 , \15489 , \15490 , \15491 , \15492 , \15493 , \15494 , \15495 , \15496 , \15497 , \15498 , \15499 , \15500 , \15501 , \15502 , \15503 , \15504 , \15505 , \15506 , \15507 , \15508 , \15509 , \15510 , \15511 , \15512 , \15513 , \15514 , \15515 , \15516 , \15517 );
or \U$6406 ( \15519 , \15453 , \15518 );
_DC g2c99 ( \15520_nG2c99 , \15519 , \9323 );
buf \U$6407 ( \15521 , \15520_nG2c99 );
and \U$6408 ( \15522 , RIe19c6f8_3157, \9333 );
and \U$6409 ( \15523 , RIe1999f8_3125, \9335 );
and \U$6410 ( \15524 , RIf1450b8_5245, \9337 );
and \U$6411 ( \15525 , RIe196cf8_3093, \9339 );
and \U$6412 ( \15526 , RIf143fd8_5233, \9341 );
and \U$6413 ( \15527 , RIe193ff8_3061, \9343 );
and \U$6414 ( \15528 , RIe1912f8_3029, \9345 );
and \U$6415 ( \15529 , RIe18e5f8_2997, \9347 );
and \U$6416 ( \15530 , RIe188bf8_2933, \9349 );
and \U$6417 ( \15531 , RIe185ef8_2901, \9351 );
and \U$6418 ( \15532 , RIfe973f8_8065, \9353 );
and \U$6419 ( \15533 , RIe1831f8_2869, \9355 );
and \U$6420 ( \15534 , RIf142958_5217, \9357 );
and \U$6421 ( \15535 , RIe1804f8_2837, \9359 );
and \U$6422 ( \15536 , RIe17d7f8_2805, \9361 );
and \U$6423 ( \15537 , RIe17aaf8_2773, \9363 );
and \U$6424 ( \15538 , RIf141b48_5207, \9365 );
and \U$6425 ( \15539 , RIfc542f0_5980, \9367 );
and \U$6426 ( \15540 , RIfc800a8_6479, \9369 );
and \U$6427 ( \15541 , RIe175260_2710, \9371 );
and \U$6428 ( \15542 , RIfca0bc8_6851, \9373 );
and \U$6429 ( \15543 , RIfc48680_5846, \9375 );
and \U$6430 ( \15544 , RIee3dea0_5163, \9377 );
and \U$6431 ( \15545 , RIfcc6878_7281, \9379 );
and \U$6432 ( \15546 , RIee3ba10_5137, \9381 );
and \U$6433 ( \15547 , RIee3a930_5125, \9383 );
and \U$6434 ( \15548 , RIfe97290_8064, \9385 );
and \U$6435 ( \15549 , RIe172b00_2682, \9387 );
and \U$6436 ( \15550 , RIf16f958_5729, \9389 );
and \U$6437 ( \15551 , RIf16ee18_5721, \9391 );
and \U$6438 ( \15552 , RIf16da68_5707, \9393 );
and \U$6439 ( \15553 , RIf16d360_5702, \9395 );
and \U$6440 ( \15554 , RIfe96e58_8061, \9397 );
and \U$6441 ( \15555 , RIe222a50_4684, \9399 );
and \U$6442 ( \15556 , RIfe96cf0_8060, \9401 );
and \U$6443 ( \15557 , RIe21fd50_4652, \9403 );
and \U$6444 ( \15558 , RIf16a660_5670, \9405 );
and \U$6445 ( \15559 , RIe21d050_4620, \9407 );
and \U$6446 ( \15560 , RIe217650_4556, \9409 );
and \U$6447 ( \15561 , RIe214950_4524, \9411 );
and \U$6448 ( \15562 , RIf169f58_5665, \9413 );
and \U$6449 ( \15563 , RIe211c50_4492, \9415 );
and \U$6450 ( \15564 , RIf168770_5648, \9417 );
and \U$6451 ( \15565 , RIe20ef50_4460, \9419 );
and \U$6452 ( \15566 , RIf1677f8_5637, \9421 );
and \U$6453 ( \15567 , RIe20c250_4428, \9423 );
and \U$6454 ( \15568 , RIe209550_4396, \9425 );
and \U$6455 ( \15569 , RIe206850_4364, \9427 );
and \U$6456 ( \15570 , RIf166880_5626, \9429 );
and \U$6457 ( \15571 , RIf1657a0_5614, \9431 );
and \U$6458 ( \15572 , RIe201dc8_4311, \9433 );
and \U$6459 ( \15573 , RIe2005e0_4294, \9435 );
and \U$6460 ( \15574 , RIfe96b88_8059, \9437 );
and \U$6461 ( \15575 , RIf163b80_5594, \9439 );
and \U$6462 ( \15576 , RIf162c08_5583, \9441 );
and \U$6463 ( \15577 , RIf161420_5566, \9443 );
and \U$6464 ( \15578 , RIf15f530_5544, \9445 );
and \U$6465 ( \15579 , RIf15d7a8_5523, \9447 );
and \U$6466 ( \15580 , RIfe968b8_8057, \9449 );
and \U$6467 ( \15581 , RIfe96a20_8058, \9451 );
and \U$6468 ( \15582 , RIfcb3fc0_7070, \9453 );
and \U$6469 ( \15583 , RIfc7cf70_6444, \9455 );
and \U$6470 ( \15584 , RIfc579c8_6019, \9457 );
and \U$6471 ( \15585 , RIf159590_5476, \9459 );
or \U$6472 ( \15586 , \15522 , \15523 , \15524 , \15525 , \15526 , \15527 , \15528 , \15529 , \15530 , \15531 , \15532 , \15533 , \15534 , \15535 , \15536 , \15537 , \15538 , \15539 , \15540 , \15541 , \15542 , \15543 , \15544 , \15545 , \15546 , \15547 , \15548 , \15549 , \15550 , \15551 , \15552 , \15553 , \15554 , \15555 , \15556 , \15557 , \15558 , \15559 , \15560 , \15561 , \15562 , \15563 , \15564 , \15565 , \15566 , \15567 , \15568 , \15569 , \15570 , \15571 , \15572 , \15573 , \15574 , \15575 , \15576 , \15577 , \15578 , \15579 , \15580 , \15581 , \15582 , \15583 , \15584 , \15585 );
and \U$6473 ( \15587 , RIf1584b0_5464, \9462 );
and \U$6474 ( \15588 , RIf157268_5451, \9464 );
and \U$6475 ( \15589 , RIf1569f8_5445, \9466 );
and \U$6476 ( \15590 , RIfe965e8_8055, \9468 );
and \U$6477 ( \15591 , RIf155d50_5436, \9470 );
and \U$6478 ( \15592 , RIf155210_5428, \9472 );
and \U$6479 ( \15593 , RIf153e60_5414, \9474 );
and \U$6480 ( \15594 , RIfe96750_8056, \9476 );
and \U$6481 ( \15595 , RIf1527e0_5398, \9478 );
and \U$6482 ( \15596 , RIf151430_5384, \9480 );
and \U$6483 ( \15597 , RIfcd2650_7416, \9482 );
and \U$6484 ( \15598 , RIe1f2648_4135, \9484 );
and \U$6485 ( \15599 , RIf14f108_5359, \9486 );
and \U$6486 ( \15600 , RIfc7f298_6469, \9488 );
and \U$6487 ( \15601 , RIf14d4e8_5339, \9490 );
and \U$6488 ( \15602 , RIe1ed350_4076, \9492 );
and \U$6489 ( \15603 , RIe1ea7b8_4045, \9494 );
and \U$6490 ( \15604 , RIe1e7ab8_4013, \9496 );
and \U$6491 ( \15605 , RIe1e4db8_3981, \9498 );
and \U$6492 ( \15606 , RIe1e20b8_3949, \9500 );
and \U$6493 ( \15607 , RIe1df3b8_3917, \9502 );
and \U$6494 ( \15608 , RIe1dc6b8_3885, \9504 );
and \U$6495 ( \15609 , RIe1d99b8_3853, \9506 );
and \U$6496 ( \15610 , RIe1d6cb8_3821, \9508 );
and \U$6497 ( \15611 , RIe1d12b8_3757, \9510 );
and \U$6498 ( \15612 , RIe1ce5b8_3725, \9512 );
and \U$6499 ( \15613 , RIe1cb8b8_3693, \9514 );
and \U$6500 ( \15614 , RIe1c8bb8_3661, \9516 );
and \U$6501 ( \15615 , RIe1c5eb8_3629, \9518 );
and \U$6502 ( \15616 , RIe1c31b8_3597, \9520 );
and \U$6503 ( \15617 , RIe1c04b8_3565, \9522 );
and \U$6504 ( \15618 , RIe1bd7b8_3533, \9524 );
and \U$6505 ( \15619 , RIf14c138_5325, \9526 );
and \U$6506 ( \15620 , RIf14ad88_5311, \9528 );
and \U$6507 ( \15621 , RIe1b8790_3476, \9530 );
and \U$6508 ( \15622 , RIfe96480_8054, \9532 );
and \U$6509 ( \15623 , RIf14a0e0_5302, \9534 );
and \U$6510 ( \15624 , RIf149870_5296, \9536 );
and \U$6511 ( \15625 , RIfe97128_8063, \9538 );
and \U$6512 ( \15626 , RIfe96318_8053, \9540 );
and \U$6513 ( \15627 , RIf148628_5283, \9542 );
and \U$6514 ( \15628 , RIfc58d78_6033, \9544 );
and \U$6515 ( \15629 , RIe1b20e8_3403, \9546 );
and \U$6516 ( \15630 , RIe1b04c8_3383, \9548 );
and \U$6517 ( \15631 , RIf146cd8_5265, \9550 );
and \U$6518 ( \15632 , RIfc591b0_6036, \9552 );
and \U$6519 ( \15633 , RIfe961b0_8052, \9554 );
and \U$6520 ( \15634 , RIfe96fc0_8062, \9556 );
and \U$6521 ( \15635 , RIe1a7af8_3285, \9558 );
and \U$6522 ( \15636 , RIe1a4df8_3253, \9560 );
and \U$6523 ( \15637 , RIe1a20f8_3221, \9562 );
and \U$6524 ( \15638 , RIe19f3f8_3189, \9564 );
and \U$6525 ( \15639 , RIe18b8f8_2965, \9566 );
and \U$6526 ( \15640 , RIe177df8_2741, \9568 );
and \U$6527 ( \15641 , RIe225750_4716, \9570 );
and \U$6528 ( \15642 , RIe21a350_4588, \9572 );
and \U$6529 ( \15643 , RIe203b50_4332, \9574 );
and \U$6530 ( \15644 , RIe1fdbb0_4264, \9576 );
and \U$6531 ( \15645 , RIe1f6f68_4187, \9578 );
and \U$6532 ( \15646 , RIe1efab0_4104, \9580 );
and \U$6533 ( \15647 , RIe1d3fb8_3789, \9582 );
and \U$6534 ( \15648 , RIe1baab8_3501, \9584 );
and \U$6535 ( \15649 , RIe1ad930_3352, \9586 );
and \U$6536 ( \15650 , RIe16ff68_2651, \9588 );
or \U$6537 ( \15651 , \15587 , \15588 , \15589 , \15590 , \15591 , \15592 , \15593 , \15594 , \15595 , \15596 , \15597 , \15598 , \15599 , \15600 , \15601 , \15602 , \15603 , \15604 , \15605 , \15606 , \15607 , \15608 , \15609 , \15610 , \15611 , \15612 , \15613 , \15614 , \15615 , \15616 , \15617 , \15618 , \15619 , \15620 , \15621 , \15622 , \15623 , \15624 , \15625 , \15626 , \15627 , \15628 , \15629 , \15630 , \15631 , \15632 , \15633 , \15634 , \15635 , \15636 , \15637 , \15638 , \15639 , \15640 , \15641 , \15642 , \15643 , \15644 , \15645 , \15646 , \15647 , \15648 , \15649 , \15650 );
or \U$6538 ( \15652 , \15586 , \15651 );
_DC g3dc6 ( \15653_nG3dc6 , \15652 , \9597 );
buf \U$6539 ( \15654 , \15653_nG3dc6 );
xor \U$6540 ( \15655 , \15521 , \15654 );
and \U$6541 ( \15656 , RIdec42f8_696, \9059 );
and \U$6542 ( \15657 , RIdec15f8_664, \9061 );
and \U$6543 ( \15658 , RIfcc6cb0_7284, \9063 );
and \U$6544 ( \15659 , RIdebe8f8_632, \9065 );
and \U$6545 ( \15660 , RIfe93780_8022, \9067 );
and \U$6546 ( \15661 , RIdebbbf8_600, \9069 );
and \U$6547 ( \15662 , RIdeb8ef8_568, \9071 );
and \U$6548 ( \15663 , RIdeb61f8_536, \9073 );
and \U$6549 ( \15664 , RIee1ea00_4807, \9075 );
and \U$6550 ( \15665 , RIdeb07f8_472, \9077 );
and \U$6551 ( \15666 , RIee1e2f8_4802, \9079 );
and \U$6552 ( \15667 , RIdeadaf8_440, \9081 );
and \U$6553 ( \15668 , RIfc5d3c8_6083, \9083 );
and \U$6554 ( \15669 , RIdea7cc0_408, \9085 );
and \U$6555 ( \15670 , RIdea13c0_376, \9087 );
and \U$6556 ( \15671 , RIde9aac0_344, \9089 );
and \U$6557 ( \15672 , RIfc58238_6025, \9091 );
and \U$6558 ( \15673 , RIfcc3b78_7249, \9093 );
and \U$6559 ( \15674 , RIfc7d0d8_6445, \9095 );
and \U$6560 ( \15675 , RIfc59750_6040, \9097 );
and \U$6561 ( \15676 , RIfe93a50_8024, \9099 );
and \U$6562 ( \15677 , RIfe938e8_8023, \9101 );
and \U$6563 ( \15678 , RIde88370_254, \9103 );
and \U$6564 ( \15679 , RIde83e88_233, \9105 );
and \U$6565 ( \15680 , RIfc5f420_6106, \9107 );
and \U$6566 ( \15681 , RIfc976b8_6745, \9109 );
and \U$6567 ( \15682 , RIfc90a70_6668, \9111 );
and \U$6568 ( \15683 , RIfc60500_6118, \9113 );
and \U$6569 ( \15684 , RIee38a40_5103, \9115 );
and \U$6570 ( \15685 , RIe16ab08_2591, \9117 );
and \U$6571 ( \15686 , RIe169488_2575, \9119 );
and \U$6572 ( \15687 , RIe166ff8_2549, \9121 );
and \U$6573 ( \15688 , RIe1642f8_2517, \9123 );
and \U$6574 ( \15689 , RIe1615f8_2485, \9125 );
and \U$6575 ( \15690 , RIee369e8_5080, \9127 );
and \U$6576 ( \15691 , RIe15e8f8_2453, \9129 );
and \U$6577 ( \15692 , RIee35bd8_5070, \9131 );
and \U$6578 ( \15693 , RIe15bbf8_2421, \9133 );
and \U$6579 ( \15694 , RIe1561f8_2357, \9135 );
and \U$6580 ( \15695 , RIe1534f8_2325, \9137 );
and \U$6581 ( \15696 , RIfc3ee28_5741, \9139 );
and \U$6582 ( \15697 , RIe1507f8_2293, \9141 );
and \U$6583 ( \15698 , RIfce6c90_7648, \9143 );
and \U$6584 ( \15699 , RIe14daf8_2261, \9145 );
and \U$6585 ( \15700 , RIfcca7c0_7326, \9147 );
and \U$6586 ( \15701 , RIe14adf8_2229, \9149 );
and \U$6587 ( \15702 , RIe1480f8_2197, \9151 );
and \U$6588 ( \15703 , RIe1453f8_2165, \9153 );
and \U$6589 ( \15704 , RIee33b80_5047, \9155 );
and \U$6590 ( \15705 , RIee32938_5034, \9157 );
and \U$6591 ( \15706 , RIee316f0_5021, \9159 );
and \U$6592 ( \15707 , RIee30bb0_5013, \9161 );
and \U$6593 ( \15708 , RIe1403d0_2108, \9163 );
and \U$6594 ( \15709 , RIfe93618_8021, \9165 );
and \U$6595 ( \15710 , RIdf3bfb0_2059, \9167 );
and \U$6596 ( \15711 , RIfe934b0_8020, \9169 );
and \U$6597 ( \15712 , RIfcd0d00_7398, \9171 );
and \U$6598 ( \15713 , RIee2ecc0_4991, \9173 );
and \U$6599 ( \15714 , RIee2e720_4987, \9175 );
and \U$6600 ( \15715 , RIee2cb00_4967, \9177 );
and \U$6601 ( \15716 , RIfe93bb8_8025, \9179 );
and \U$6602 ( \15717 , RIdf32938_1952, \9181 );
and \U$6603 ( \15718 , RIdf30340_1925, \9183 );
and \U$6604 ( \15719 , RIdf2e450_1903, \9185 );
or \U$6605 ( \15720 , \15656 , \15657 , \15658 , \15659 , \15660 , \15661 , \15662 , \15663 , \15664 , \15665 , \15666 , \15667 , \15668 , \15669 , \15670 , \15671 , \15672 , \15673 , \15674 , \15675 , \15676 , \15677 , \15678 , \15679 , \15680 , \15681 , \15682 , \15683 , \15684 , \15685 , \15686 , \15687 , \15688 , \15689 , \15690 , \15691 , \15692 , \15693 , \15694 , \15695 , \15696 , \15697 , \15698 , \15699 , \15700 , \15701 , \15702 , \15703 , \15704 , \15705 , \15706 , \15707 , \15708 , \15709 , \15710 , \15711 , \15712 , \15713 , \15714 , \15715 , \15716 , \15717 , \15718 , \15719 );
and \U$6606 ( \15721 , RIee2b048_4948, \9188 );
and \U$6607 ( \15722 , RIee29b30_4933, \9190 );
and \U$6608 ( \15723 , RIfc67148_6195, \9192 );
and \U$6609 ( \15724 , RIfc6fb18_6293, \9194 );
and \U$6610 ( \15725 , RIdf29860_1849, \9196 );
and \U$6611 ( \15726 , RIfe931e0_8018, \9198 );
and \U$6612 ( \15727 , RIfe93348_8019, \9200 );
and \U$6613 ( \15728 , RIfe93078_8017, \9202 );
and \U$6614 ( \15729 , RIfc672b0_6196, \9204 );
and \U$6615 ( \15730 , RIfca8788_6939, \9206 );
and \U$6616 ( \15731 , RIdf22510_1767, \9208 );
and \U$6617 ( \15732 , RIfcea7a0_7690, \9210 );
and \U$6618 ( \15733 , RIdf20ff8_1752, \9212 );
and \U$6619 ( \15734 , RIdf1ecd0_1727, \9214 );
and \U$6620 ( \15735 , RIdf1aab8_1680, \9216 );
and \U$6621 ( \15736 , RIfea7c58_8225, \9218 );
and \U$6622 ( \15737 , RIdf15ec8_1626, \9220 );
and \U$6623 ( \15738 , RIdf131c8_1594, \9222 );
and \U$6624 ( \15739 , RIdf104c8_1562, \9224 );
and \U$6625 ( \15740 , RIdf0d7c8_1530, \9226 );
and \U$6626 ( \15741 , RIdf0aac8_1498, \9228 );
and \U$6627 ( \15742 , RIdf07dc8_1466, \9230 );
and \U$6628 ( \15743 , RIdf050c8_1434, \9232 );
and \U$6629 ( \15744 , RIdf023c8_1402, \9234 );
and \U$6630 ( \15745 , RIdefc9c8_1338, \9236 );
and \U$6631 ( \15746 , RIdef9cc8_1306, \9238 );
and \U$6632 ( \15747 , RIdef6fc8_1274, \9240 );
and \U$6633 ( \15748 , RIdef42c8_1242, \9242 );
and \U$6634 ( \15749 , RIdef15c8_1210, \9244 );
and \U$6635 ( \15750 , RIdeee8c8_1178, \9246 );
and \U$6636 ( \15751 , RIdeebbc8_1146, \9248 );
and \U$6637 ( \15752 , RIdee8ec8_1114, \9250 );
and \U$6638 ( \15753 , RIee24f40_4879, \9252 );
and \U$6639 ( \15754 , RIee24130_4869, \9254 );
and \U$6640 ( \15755 , RIee235f0_4861, \9256 );
and \U$6641 ( \15756 , RIee22c18_4854, \9258 );
and \U$6642 ( \15757 , RIfe93d20_8026, \9260 );
and \U$6643 ( \15758 , RIdee1fb0_1035, \9262 );
and \U$6644 ( \15759 , RIdee0228_1014, \9264 );
and \U$6645 ( \15760 , RIdeddc30_987, \9266 );
and \U$6646 ( \15761 , RIfc684f8_6209, \9268 );
and \U$6647 ( \15762 , RIee21ca0_4843, \9270 );
and \U$6648 ( \15763 , RIfc68390_6208, \9272 );
and \U$6649 ( \15764 , RIee20d28_4832, \9274 );
and \U$6650 ( \15765 , RIded8aa0_929, \9276 );
and \U$6651 ( \15766 , RIfe93ff0_8028, \9278 );
and \U$6652 ( \15767 , RIded45b8_880, \9280 );
and \U$6653 ( \15768 , RIfe93e88_8027, \9282 );
and \U$6654 ( \15769 , RIdecf6f8_824, \9284 );
and \U$6655 ( \15770 , RIdecc9f8_792, \9286 );
and \U$6656 ( \15771 , RIdec9cf8_760, \9288 );
and \U$6657 ( \15772 , RIdec6ff8_728, \9290 );
and \U$6658 ( \15773 , RIdeb34f8_504, \9292 );
and \U$6659 ( \15774 , RIde941c0_312, \9294 );
and \U$6660 ( \15775 , RIe16d100_2618, \9296 );
and \U$6661 ( \15776 , RIe158ef8_2389, \9298 );
and \U$6662 ( \15777 , RIe1426f8_2133, \9300 );
and \U$6663 ( \15778 , RIdf370f0_2003, \9302 );
and \U$6664 ( \15779 , RIdf2b750_1871, \9304 );
and \U$6665 ( \15780 , RIdf1bfd0_1695, \9306 );
and \U$6666 ( \15781 , RIdeff6c8_1370, \9308 );
and \U$6667 ( \15782 , RIdee61c8_1082, \9310 );
and \U$6668 ( \15783 , RIdedaf30_955, \9312 );
and \U$6669 ( \15784 , RIde7a108_185, \9314 );
or \U$6670 ( \15785 , \15721 , \15722 , \15723 , \15724 , \15725 , \15726 , \15727 , \15728 , \15729 , \15730 , \15731 , \15732 , \15733 , \15734 , \15735 , \15736 , \15737 , \15738 , \15739 , \15740 , \15741 , \15742 , \15743 , \15744 , \15745 , \15746 , \15747 , \15748 , \15749 , \15750 , \15751 , \15752 , \15753 , \15754 , \15755 , \15756 , \15757 , \15758 , \15759 , \15760 , \15761 , \15762 , \15763 , \15764 , \15765 , \15766 , \15767 , \15768 , \15769 , \15770 , \15771 , \15772 , \15773 , \15774 , \15775 , \15776 , \15777 , \15778 , \15779 , \15780 , \15781 , \15782 , \15783 , \15784 );
or \U$6671 ( \15786 , \15720 , \15785 );
_DC g2d1e ( \15787_nG2d1e , \15786 , \9323 );
buf \U$6672 ( \15788 , \15787_nG2d1e );
and \U$6673 ( \15789 , RIe19c590_3156, \9333 );
and \U$6674 ( \15790 , RIe199890_3124, \9335 );
and \U$6675 ( \15791 , RIf144f50_5244, \9337 );
and \U$6676 ( \15792 , RIe196b90_3092, \9339 );
and \U$6677 ( \15793 , RIfc76058_6365, \9341 );
and \U$6678 ( \15794 , RIe193e90_3060, \9343 );
and \U$6679 ( \15795 , RIe191190_3028, \9345 );
and \U$6680 ( \15796 , RIe18e490_2996, \9347 );
and \U$6681 ( \15797 , RIe188a90_2932, \9349 );
and \U$6682 ( \15798 , RIe185d90_2900, \9351 );
and \U$6683 ( \15799 , RIfccd8f8_7361, \9353 );
and \U$6684 ( \15800 , RIe183090_2868, \9355 );
and \U$6685 ( \15801 , RIfc76e68_6375, \9357 );
and \U$6686 ( \15802 , RIe180390_2836, \9359 );
and \U$6687 ( \15803 , RIe17d690_2804, \9361 );
and \U$6688 ( \15804 , RIe17a990_2772, \9363 );
and \U$6689 ( \15805 , RIf1419e0_5206, \9365 );
and \U$6690 ( \15806 , RIf140630_5192, \9367 );
and \U$6691 ( \15807 , RIe176bb0_2728, \9369 );
and \U$6692 ( \15808 , RIe1750f8_2709, \9371 );
and \U$6693 ( \15809 , RIfcd1840_7406, \9373 );
and \U$6694 ( \15810 , RIfc5f6f0_6108, \9375 );
and \U$6695 ( \15811 , RIee3dd38_5162, \9377 );
and \U$6696 ( \15812 , RIee3cc58_5150, \9379 );
and \U$6697 ( \15813 , RIee3b8a8_5136, \9381 );
and \U$6698 ( \15814 , RIee3a7c8_5124, \9383 );
and \U$6699 ( \15815 , RIee39580_5111, \9385 );
and \U$6700 ( \15816 , RIfea9008_8239, \9387 );
and \U$6701 ( \15817 , RIf16f7f0_5728, \9389 );
and \U$6702 ( \15818 , RIf16ecb0_5720, \9391 );
and \U$6703 ( \15819 , RIf16d900_5706, \9393 );
and \U$6704 ( \15820 , RIfc78ec0_6398, \9395 );
and \U$6705 ( \15821 , RIfcc8060_7298, \9397 );
and \U$6706 ( \15822 , RIe2228e8_4683, \9399 );
and \U$6707 ( \15823 , RIfc5a3f8_6049, \9401 );
and \U$6708 ( \15824 , RIe21fbe8_4651, \9403 );
and \U$6709 ( \15825 , RIfc74000_6342, \9405 );
and \U$6710 ( \15826 , RIe21cee8_4619, \9407 );
and \U$6711 ( \15827 , RIe2174e8_4555, \9409 );
and \U$6712 ( \15828 , RIe2147e8_4523, \9411 );
and \U$6713 ( \15829 , RIfca2c20_6874, \9413 );
and \U$6714 ( \15830 , RIe211ae8_4491, \9415 );
and \U$6715 ( \15831 , RIfca2950_6872, \9417 );
and \U$6716 ( \15832 , RIe20ede8_4459, \9419 );
and \U$6717 ( \15833 , RIfcc24f8_7233, \9421 );
and \U$6718 ( \15834 , RIe20c0e8_4427, \9423 );
and \U$6719 ( \15835 , RIe2093e8_4395, \9425 );
and \U$6720 ( \15836 , RIe2066e8_4363, \9427 );
and \U$6721 ( \15837 , RIfc45110_5808, \9429 );
and \U$6722 ( \15838 , RIfcc6f80_7286, \9431 );
and \U$6723 ( \15839 , RIfe92f10_8016, \9433 );
and \U$6724 ( \15840 , RIfe92970_8012, \9435 );
and \U$6725 ( \15841 , RIf164af8_5605, \9437 );
and \U$6726 ( \15842 , RIf163a18_5593, \9439 );
and \U$6727 ( \15843 , RIf162aa0_5582, \9441 );
and \U$6728 ( \15844 , RIfe92ad8_8013, \9443 );
and \U$6729 ( \15845 , RIf15f3c8_5543, \9445 );
and \U$6730 ( \15846 , RIf15d640_5522, \9447 );
and \U$6731 ( \15847 , RIfe92808_8011, \9449 );
and \U$6732 ( \15848 , RIfe92c40_8014, \9451 );
and \U$6733 ( \15849 , RIfe926a0_8010, \9453 );
and \U$6734 ( \15850 , RIfe92da8_8015, \9455 );
and \U$6735 ( \15851 , RIfe92538_8009, \9457 );
and \U$6736 ( \15852 , RIfcb5a78_7089, \9459 );
or \U$6737 ( \15853 , \15789 , \15790 , \15791 , \15792 , \15793 , \15794 , \15795 , \15796 , \15797 , \15798 , \15799 , \15800 , \15801 , \15802 , \15803 , \15804 , \15805 , \15806 , \15807 , \15808 , \15809 , \15810 , \15811 , \15812 , \15813 , \15814 , \15815 , \15816 , \15817 , \15818 , \15819 , \15820 , \15821 , \15822 , \15823 , \15824 , \15825 , \15826 , \15827 , \15828 , \15829 , \15830 , \15831 , \15832 , \15833 , \15834 , \15835 , \15836 , \15837 , \15838 , \15839 , \15840 , \15841 , \15842 , \15843 , \15844 , \15845 , \15846 , \15847 , \15848 , \15849 , \15850 , \15851 , \15852 );
and \U$6738 ( \15854 , RIf158348_5463, \9462 );
and \U$6739 ( \15855 , RIf157100_5450, \9464 );
and \U$6740 ( \15856 , RIfc53be8_5975, \9466 );
and \U$6741 ( \15857 , RIfec38b8_8345, \9468 );
and \U$6742 ( \15858 , RIfcc5ea0_7274, \9470 );
and \U$6743 ( \15859 , RIf1550a8_5427, \9472 );
and \U$6744 ( \15860 , RIf153cf8_5413, \9474 );
and \U$6745 ( \15861 , RIfec3a20_8346, \9476 );
and \U$6746 ( \15862 , RIf152678_5397, \9478 );
and \U$6747 ( \15863 , RIfec3750_8344, \9480 );
and \U$6748 ( \15864 , RIf14ff18_5369, \9482 );
and \U$6749 ( \15865 , RIfe923d0_8008, \9484 );
and \U$6750 ( \15866 , RIf14efa0_5358, \9486 );
and \U$6751 ( \15867 , RIf14e898_5353, \9488 );
and \U$6752 ( \15868 , RIf14d380_5338, \9490 );
and \U$6753 ( \15869 , RIfe92268_8007, \9492 );
and \U$6754 ( \15870 , RIe1ea650_4044, \9494 );
and \U$6755 ( \15871 , RIe1e7950_4012, \9496 );
and \U$6756 ( \15872 , RIe1e4c50_3980, \9498 );
and \U$6757 ( \15873 , RIe1e1f50_3948, \9500 );
and \U$6758 ( \15874 , RIe1df250_3916, \9502 );
and \U$6759 ( \15875 , RIe1dc550_3884, \9504 );
and \U$6760 ( \15876 , RIe1d9850_3852, \9506 );
and \U$6761 ( \15877 , RIe1d6b50_3820, \9508 );
and \U$6762 ( \15878 , RIe1d1150_3756, \9510 );
and \U$6763 ( \15879 , RIe1ce450_3724, \9512 );
and \U$6764 ( \15880 , RIe1cb750_3692, \9514 );
and \U$6765 ( \15881 , RIe1c8a50_3660, \9516 );
and \U$6766 ( \15882 , RIe1c5d50_3628, \9518 );
and \U$6767 ( \15883 , RIe1c3050_3596, \9520 );
and \U$6768 ( \15884 , RIe1c0350_3564, \9522 );
and \U$6769 ( \15885 , RIe1bd650_3532, \9524 );
and \U$6770 ( \15886 , RIfcda4e0_7506, \9526 );
and \U$6771 ( \15887 , RIfc9d220_6810, \9528 );
and \U$6772 ( \15888 , RIe1b8628_3475, \9530 );
and \U$6773 ( \15889 , RIe1b6738_3453, \9532 );
and \U$6774 ( \15890 , RIfc4f2c8_5923, \9534 );
and \U$6775 ( \15891 , RIfce16c8_7587, \9536 );
and \U$6776 ( \15892 , RIfe91cc8_8003, \9538 );
and \U$6777 ( \15893 , RIfe91e30_8004, \9540 );
and \U$6778 ( \15894 , RIf1484c0_5282, \9542 );
and \U$6779 ( \15895 , RIf147548_5271, \9544 );
and \U$6780 ( \15896 , RIfe91f98_8005, \9546 );
and \U$6781 ( \15897 , RIfe91b60_8002, \9548 );
and \U$6782 ( \15898 , RIf146b70_5264, \9550 );
and \U$6783 ( \15899 , RIfc9f548_6835, \9552 );
and \U$6784 ( \15900 , RIfe92100_8006, \9554 );
and \U$6785 ( \15901 , RIfe919f8_8001, \9556 );
and \U$6786 ( \15902 , RIe1a7990_3284, \9558 );
and \U$6787 ( \15903 , RIe1a4c90_3252, \9560 );
and \U$6788 ( \15904 , RIe1a1f90_3220, \9562 );
and \U$6789 ( \15905 , RIe19f290_3188, \9564 );
and \U$6790 ( \15906 , RIe18b790_2964, \9566 );
and \U$6791 ( \15907 , RIe177c90_2740, \9568 );
and \U$6792 ( \15908 , RIe2255e8_4715, \9570 );
and \U$6793 ( \15909 , RIe21a1e8_4587, \9572 );
and \U$6794 ( \15910 , RIe2039e8_4331, \9574 );
and \U$6795 ( \15911 , RIe1fda48_4263, \9576 );
and \U$6796 ( \15912 , RIe1f6e00_4186, \9578 );
and \U$6797 ( \15913 , RIe1ef948_4103, \9580 );
and \U$6798 ( \15914 , RIe1d3e50_3788, \9582 );
and \U$6799 ( \15915 , RIe1ba950_3500, \9584 );
and \U$6800 ( \15916 , RIe1ad7c8_3351, \9586 );
and \U$6801 ( \15917 , RIe16fe00_2650, \9588 );
or \U$6802 ( \15918 , \15854 , \15855 , \15856 , \15857 , \15858 , \15859 , \15860 , \15861 , \15862 , \15863 , \15864 , \15865 , \15866 , \15867 , \15868 , \15869 , \15870 , \15871 , \15872 , \15873 , \15874 , \15875 , \15876 , \15877 , \15878 , \15879 , \15880 , \15881 , \15882 , \15883 , \15884 , \15885 , \15886 , \15887 , \15888 , \15889 , \15890 , \15891 , \15892 , \15893 , \15894 , \15895 , \15896 , \15897 , \15898 , \15899 , \15900 , \15901 , \15902 , \15903 , \15904 , \15905 , \15906 , \15907 , \15908 , \15909 , \15910 , \15911 , \15912 , \15913 , \15914 , \15915 , \15916 , \15917 );
or \U$6803 ( \15919 , \15853 , \15918 );
_DC g3e4b ( \15920_nG3e4b , \15919 , \9597 );
buf \U$6804 ( \15921 , \15920_nG3e4b );
and \U$6805 ( \15922 , \15788 , \15921 );
and \U$6806 ( \15923 , \14212 , \14345 );
and \U$6807 ( \15924 , \14345 , \14620 );
and \U$6808 ( \15925 , \14212 , \14620 );
or \U$6809 ( \15926 , \15923 , \15924 , \15925 );
and \U$6810 ( \15927 , \15921 , \15926 );
and \U$6811 ( \15928 , \15788 , \15926 );
or \U$6812 ( \15929 , \15922 , \15927 , \15928 );
xor \U$6813 ( \15930 , \15655 , \15929 );
buf g4436 ( \15931_nG4436 , \15930 );
xor \U$6814 ( \15932 , \15788 , \15921 );
xor \U$6815 ( \15933 , \15932 , \15926 );
buf g4439 ( \15934_nG4439 , \15933 );
nand \U$6816 ( \15935 , \15934_nG4439 , \14622_nG443c );
and \U$6817 ( \15936 , \15931_nG4436 , \15935 );
xor \U$6818 ( \15937 , \15934_nG4439 , \14622_nG443c );
not \U$6819 ( \15938 , \15937 );
xor \U$6820 ( \15939 , \15931_nG4436 , \15934_nG4439 );
and \U$6821 ( \15940 , \15938 , \15939 );
and \U$6823 ( \15941 , \15937 , \10694_nG9c0e );
or \U$6824 ( \15942 , 1'b0 , \15941 );
xor \U$6825 ( \15943 , \15936 , \15942 );
xor \U$6826 ( \15944 , \15936 , \15943 );
buf \U$6827 ( \15945 , \15944 );
buf \U$6828 ( \15946 , \15945 );
and \U$6829 ( \15947 , \15388 , \15946 );
and \U$6830 ( \15948 , \15032 , \15048 );
and \U$6831 ( \15949 , \15032 , \15378 );
and \U$6832 ( \15950 , \15048 , \15378 );
or \U$6833 ( \15951 , \15948 , \15949 , \15950 );
buf \U$6834 ( \15952 , \15951 );
and \U$6835 ( \15953 , \15037 , \15039 );
and \U$6836 ( \15954 , \15037 , \15046 );
and \U$6837 ( \15955 , \15039 , \15046 );
or \U$6838 ( \15956 , \15953 , \15954 , \15955 );
buf \U$6839 ( \15957 , \15956 );
and \U$6840 ( \15958 , \14631 , \10995_nG9c0b );
and \U$6841 ( \15959 , \14628 , \11283_nG9c08 );
or \U$6842 ( \15960 , \15958 , \15959 );
xor \U$6843 ( \15961 , \14627 , \15960 );
buf \U$6844 ( \15962 , \15961 );
buf \U$6846 ( \15963 , \15962 );
and \U$6847 ( \15964 , \13370 , \11598_nG9c05 );
and \U$6848 ( \15965 , \13367 , \12470_nG9c02 );
or \U$6849 ( \15966 , \15964 , \15965 );
xor \U$6850 ( \15967 , \13366 , \15966 );
buf \U$6851 ( \15968 , \15967 );
buf \U$6853 ( \15969 , \15968 );
xor \U$6854 ( \15970 , \15963 , \15969 );
buf \U$6855 ( \15971 , \15970 );
and \U$6856 ( \15972 , \15009 , \15015 );
buf \U$6857 ( \15973 , \15972 );
xor \U$6858 ( \15974 , \15971 , \15973 );
and \U$6859 ( \15975 , \12157 , \12801_nG9bff );
and \U$6860 ( \15976 , \12154 , \13705_nG9bfc );
or \U$6861 ( \15977 , \15975 , \15976 );
xor \U$6862 ( \15978 , \12153 , \15977 );
buf \U$6863 ( \15979 , \15978 );
buf \U$6865 ( \15980 , \15979 );
xor \U$6866 ( \15981 , \15974 , \15980 );
buf \U$6867 ( \15982 , \15981 );
xor \U$6868 ( \15983 , \15957 , \15982 );
and \U$6869 ( \15984 , \15017 , \15023 );
and \U$6870 ( \15985 , \15017 , \15030 );
and \U$6871 ( \15986 , \15023 , \15030 );
or \U$6872 ( \15987 , \15984 , \15985 , \15986 );
buf \U$6873 ( \15988 , \15987 );
and \U$6874 ( \15989 , \10421 , \14070_nG9bf9 );
and \U$6875 ( \15990 , \10418 , \14984_nG9bf6 );
or \U$6876 ( \15991 , \15989 , \15990 );
xor \U$6877 ( \15992 , \10417 , \15991 );
buf \U$6878 ( \15993 , \15992 );
buf \U$6880 ( \15994 , \15993 );
xor \U$6881 ( \15995 , \15988 , \15994 );
and \U$6882 ( \15996 , \10707 , \15373_nG9bf3 );
and \U$6883 ( \15997 , \15352 , \15356 );
and \U$6884 ( \15998 , \15356 , \15361 );
and \U$6885 ( \15999 , \15352 , \15361 );
or \U$6886 ( \16000 , \15997 , \15998 , \15999 );
and \U$6887 ( \16001 , \15321 , \10983 );
and \U$6888 ( \16002 , RIdec42f8_696, \9333 );
and \U$6889 ( \16003 , RIdec15f8_664, \9335 );
and \U$6890 ( \16004 , RIfcc6cb0_7284, \9337 );
and \U$6891 ( \16005 , RIdebe8f8_632, \9339 );
and \U$6892 ( \16006 , RIfe93780_8022, \9341 );
and \U$6893 ( \16007 , RIdebbbf8_600, \9343 );
and \U$6894 ( \16008 , RIdeb8ef8_568, \9345 );
and \U$6895 ( \16009 , RIdeb61f8_536, \9347 );
and \U$6896 ( \16010 , RIee1ea00_4807, \9349 );
and \U$6897 ( \16011 , RIdeb07f8_472, \9351 );
and \U$6898 ( \16012 , RIee1e2f8_4802, \9353 );
and \U$6899 ( \16013 , RIdeadaf8_440, \9355 );
and \U$6900 ( \16014 , RIfc5d3c8_6083, \9357 );
and \U$6901 ( \16015 , RIdea7cc0_408, \9359 );
and \U$6902 ( \16016 , RIdea13c0_376, \9361 );
and \U$6903 ( \16017 , RIde9aac0_344, \9363 );
and \U$6904 ( \16018 , RIfc58238_6025, \9365 );
and \U$6905 ( \16019 , RIfcc3b78_7249, \9367 );
and \U$6906 ( \16020 , RIfc7d0d8_6445, \9369 );
and \U$6907 ( \16021 , RIfc59750_6040, \9371 );
and \U$6908 ( \16022 , RIfe93a50_8024, \9373 );
and \U$6909 ( \16023 , RIfe938e8_8023, \9375 );
and \U$6910 ( \16024 , RIde88370_254, \9377 );
and \U$6911 ( \16025 , RIde83e88_233, \9379 );
and \U$6912 ( \16026 , RIfc5f420_6106, \9381 );
and \U$6913 ( \16027 , RIfc976b8_6745, \9383 );
and \U$6914 ( \16028 , RIfc90a70_6668, \9385 );
and \U$6915 ( \16029 , RIfc60500_6118, \9387 );
and \U$6916 ( \16030 , RIee38a40_5103, \9389 );
and \U$6917 ( \16031 , RIe16ab08_2591, \9391 );
and \U$6918 ( \16032 , RIe169488_2575, \9393 );
and \U$6919 ( \16033 , RIe166ff8_2549, \9395 );
and \U$6920 ( \16034 , RIe1642f8_2517, \9397 );
and \U$6921 ( \16035 , RIe1615f8_2485, \9399 );
and \U$6922 ( \16036 , RIee369e8_5080, \9401 );
and \U$6923 ( \16037 , RIe15e8f8_2453, \9403 );
and \U$6924 ( \16038 , RIee35bd8_5070, \9405 );
and \U$6925 ( \16039 , RIe15bbf8_2421, \9407 );
and \U$6926 ( \16040 , RIe1561f8_2357, \9409 );
and \U$6927 ( \16041 , RIe1534f8_2325, \9411 );
and \U$6928 ( \16042 , RIfc3ee28_5741, \9413 );
and \U$6929 ( \16043 , RIe1507f8_2293, \9415 );
and \U$6930 ( \16044 , RIfce6c90_7648, \9417 );
and \U$6931 ( \16045 , RIe14daf8_2261, \9419 );
and \U$6932 ( \16046 , RIfcca7c0_7326, \9421 );
and \U$6933 ( \16047 , RIe14adf8_2229, \9423 );
and \U$6934 ( \16048 , RIe1480f8_2197, \9425 );
and \U$6935 ( \16049 , RIe1453f8_2165, \9427 );
and \U$6936 ( \16050 , RIee33b80_5047, \9429 );
and \U$6937 ( \16051 , RIee32938_5034, \9431 );
and \U$6938 ( \16052 , RIee316f0_5021, \9433 );
and \U$6939 ( \16053 , RIee30bb0_5013, \9435 );
and \U$6940 ( \16054 , RIe1403d0_2108, \9437 );
and \U$6941 ( \16055 , RIfe93618_8021, \9439 );
and \U$6942 ( \16056 , RIdf3bfb0_2059, \9441 );
and \U$6943 ( \16057 , RIfe934b0_8020, \9443 );
and \U$6944 ( \16058 , RIfcd0d00_7398, \9445 );
and \U$6945 ( \16059 , RIee2ecc0_4991, \9447 );
and \U$6946 ( \16060 , RIee2e720_4987, \9449 );
and \U$6947 ( \16061 , RIee2cb00_4967, \9451 );
and \U$6948 ( \16062 , RIfe93bb8_8025, \9453 );
and \U$6949 ( \16063 , RIdf32938_1952, \9455 );
and \U$6950 ( \16064 , RIdf30340_1925, \9457 );
and \U$6951 ( \16065 , RIdf2e450_1903, \9459 );
or \U$6952 ( \16066 , \16002 , \16003 , \16004 , \16005 , \16006 , \16007 , \16008 , \16009 , \16010 , \16011 , \16012 , \16013 , \16014 , \16015 , \16016 , \16017 , \16018 , \16019 , \16020 , \16021 , \16022 , \16023 , \16024 , \16025 , \16026 , \16027 , \16028 , \16029 , \16030 , \16031 , \16032 , \16033 , \16034 , \16035 , \16036 , \16037 , \16038 , \16039 , \16040 , \16041 , \16042 , \16043 , \16044 , \16045 , \16046 , \16047 , \16048 , \16049 , \16050 , \16051 , \16052 , \16053 , \16054 , \16055 , \16056 , \16057 , \16058 , \16059 , \16060 , \16061 , \16062 , \16063 , \16064 , \16065 );
and \U$6953 ( \16067 , RIee2b048_4948, \9462 );
and \U$6954 ( \16068 , RIee29b30_4933, \9464 );
and \U$6955 ( \16069 , RIfc67148_6195, \9466 );
and \U$6956 ( \16070 , RIfc6fb18_6293, \9468 );
and \U$6957 ( \16071 , RIdf29860_1849, \9470 );
and \U$6958 ( \16072 , RIfe931e0_8018, \9472 );
and \U$6959 ( \16073 , RIfe93348_8019, \9474 );
and \U$6960 ( \16074 , RIfe93078_8017, \9476 );
and \U$6961 ( \16075 , RIfc672b0_6196, \9478 );
and \U$6962 ( \16076 , RIfca8788_6939, \9480 );
and \U$6963 ( \16077 , RIdf22510_1767, \9482 );
and \U$6964 ( \16078 , RIfcea7a0_7690, \9484 );
and \U$6965 ( \16079 , RIdf20ff8_1752, \9486 );
and \U$6966 ( \16080 , RIdf1ecd0_1727, \9488 );
and \U$6967 ( \16081 , RIdf1aab8_1680, \9490 );
and \U$6968 ( \16082 , RIfea7c58_8225, \9492 );
and \U$6969 ( \16083 , RIdf15ec8_1626, \9494 );
and \U$6970 ( \16084 , RIdf131c8_1594, \9496 );
and \U$6971 ( \16085 , RIdf104c8_1562, \9498 );
and \U$6972 ( \16086 , RIdf0d7c8_1530, \9500 );
and \U$6973 ( \16087 , RIdf0aac8_1498, \9502 );
and \U$6974 ( \16088 , RIdf07dc8_1466, \9504 );
and \U$6975 ( \16089 , RIdf050c8_1434, \9506 );
and \U$6976 ( \16090 , RIdf023c8_1402, \9508 );
and \U$6977 ( \16091 , RIdefc9c8_1338, \9510 );
and \U$6978 ( \16092 , RIdef9cc8_1306, \9512 );
and \U$6979 ( \16093 , RIdef6fc8_1274, \9514 );
and \U$6980 ( \16094 , RIdef42c8_1242, \9516 );
and \U$6981 ( \16095 , RIdef15c8_1210, \9518 );
and \U$6982 ( \16096 , RIdeee8c8_1178, \9520 );
and \U$6983 ( \16097 , RIdeebbc8_1146, \9522 );
and \U$6984 ( \16098 , RIdee8ec8_1114, \9524 );
and \U$6985 ( \16099 , RIee24f40_4879, \9526 );
and \U$6986 ( \16100 , RIee24130_4869, \9528 );
and \U$6987 ( \16101 , RIee235f0_4861, \9530 );
and \U$6988 ( \16102 , RIee22c18_4854, \9532 );
and \U$6989 ( \16103 , RIfe93d20_8026, \9534 );
and \U$6990 ( \16104 , RIdee1fb0_1035, \9536 );
and \U$6991 ( \16105 , RIdee0228_1014, \9538 );
and \U$6992 ( \16106 , RIdeddc30_987, \9540 );
and \U$6993 ( \16107 , RIfc684f8_6209, \9542 );
and \U$6994 ( \16108 , RIee21ca0_4843, \9544 );
and \U$6995 ( \16109 , RIfc68390_6208, \9546 );
and \U$6996 ( \16110 , RIee20d28_4832, \9548 );
and \U$6997 ( \16111 , RIded8aa0_929, \9550 );
and \U$6998 ( \16112 , RIfe93ff0_8028, \9552 );
and \U$6999 ( \16113 , RIded45b8_880, \9554 );
and \U$7000 ( \16114 , RIfe93e88_8027, \9556 );
and \U$7001 ( \16115 , RIdecf6f8_824, \9558 );
and \U$7002 ( \16116 , RIdecc9f8_792, \9560 );
and \U$7003 ( \16117 , RIdec9cf8_760, \9562 );
and \U$7004 ( \16118 , RIdec6ff8_728, \9564 );
and \U$7005 ( \16119 , RIdeb34f8_504, \9566 );
and \U$7006 ( \16120 , RIde941c0_312, \9568 );
and \U$7007 ( \16121 , RIe16d100_2618, \9570 );
and \U$7008 ( \16122 , RIe158ef8_2389, \9572 );
and \U$7009 ( \16123 , RIe1426f8_2133, \9574 );
and \U$7010 ( \16124 , RIdf370f0_2003, \9576 );
and \U$7011 ( \16125 , RIdf2b750_1871, \9578 );
and \U$7012 ( \16126 , RIdf1bfd0_1695, \9580 );
and \U$7013 ( \16127 , RIdeff6c8_1370, \9582 );
and \U$7014 ( \16128 , RIdee61c8_1082, \9584 );
and \U$7015 ( \16129 , RIdedaf30_955, \9586 );
and \U$7016 ( \16130 , RIde7a108_185, \9588 );
or \U$7017 ( \16131 , \16067 , \16068 , \16069 , \16070 , \16071 , \16072 , \16073 , \16074 , \16075 , \16076 , \16077 , \16078 , \16079 , \16080 , \16081 , \16082 , \16083 , \16084 , \16085 , \16086 , \16087 , \16088 , \16089 , \16090 , \16091 , \16092 , \16093 , \16094 , \16095 , \16096 , \16097 , \16098 , \16099 , \16100 , \16101 , \16102 , \16103 , \16104 , \16105 , \16106 , \16107 , \16108 , \16109 , \16110 , \16111 , \16112 , \16113 , \16114 , \16115 , \16116 , \16117 , \16118 , \16119 , \16120 , \16121 , \16122 , \16123 , \16124 , \16125 , \16126 , \16127 , \16128 , \16129 , \16130 );
or \U$7018 ( \16132 , \16066 , \16131 );
_DC g6595 ( \16133_nG6595 , \16132 , \9597 );
and \U$7019 ( \16134 , RIe19c590_3156, \9059 );
and \U$7020 ( \16135 , RIe199890_3124, \9061 );
and \U$7021 ( \16136 , RIf144f50_5244, \9063 );
and \U$7022 ( \16137 , RIe196b90_3092, \9065 );
and \U$7023 ( \16138 , RIfc76058_6365, \9067 );
and \U$7024 ( \16139 , RIe193e90_3060, \9069 );
and \U$7025 ( \16140 , RIe191190_3028, \9071 );
and \U$7026 ( \16141 , RIe18e490_2996, \9073 );
and \U$7027 ( \16142 , RIe188a90_2932, \9075 );
and \U$7028 ( \16143 , RIe185d90_2900, \9077 );
and \U$7029 ( \16144 , RIfccd8f8_7361, \9079 );
and \U$7030 ( \16145 , RIe183090_2868, \9081 );
and \U$7031 ( \16146 , RIfc76e68_6375, \9083 );
and \U$7032 ( \16147 , RIe180390_2836, \9085 );
and \U$7033 ( \16148 , RIe17d690_2804, \9087 );
and \U$7034 ( \16149 , RIe17a990_2772, \9089 );
and \U$7035 ( \16150 , RIf1419e0_5206, \9091 );
and \U$7036 ( \16151 , RIf140630_5192, \9093 );
and \U$7037 ( \16152 , RIe176bb0_2728, \9095 );
and \U$7038 ( \16153 , RIe1750f8_2709, \9097 );
and \U$7039 ( \16154 , RIfcd1840_7406, \9099 );
and \U$7040 ( \16155 , RIfc5f6f0_6108, \9101 );
and \U$7041 ( \16156 , RIee3dd38_5162, \9103 );
and \U$7042 ( \16157 , RIee3cc58_5150, \9105 );
and \U$7043 ( \16158 , RIee3b8a8_5136, \9107 );
and \U$7044 ( \16159 , RIee3a7c8_5124, \9109 );
and \U$7045 ( \16160 , RIee39580_5111, \9111 );
and \U$7046 ( \16161 , RIfea9008_8239, \9113 );
and \U$7047 ( \16162 , RIf16f7f0_5728, \9115 );
and \U$7048 ( \16163 , RIf16ecb0_5720, \9117 );
and \U$7049 ( \16164 , RIf16d900_5706, \9119 );
and \U$7050 ( \16165 , RIfc78ec0_6398, \9121 );
and \U$7051 ( \16166 , RIfcc8060_7298, \9123 );
and \U$7052 ( \16167 , RIe2228e8_4683, \9125 );
and \U$7053 ( \16168 , RIfc5a3f8_6049, \9127 );
and \U$7054 ( \16169 , RIe21fbe8_4651, \9129 );
and \U$7055 ( \16170 , RIfc74000_6342, \9131 );
and \U$7056 ( \16171 , RIe21cee8_4619, \9133 );
and \U$7057 ( \16172 , RIe2174e8_4555, \9135 );
and \U$7058 ( \16173 , RIe2147e8_4523, \9137 );
and \U$7059 ( \16174 , RIfca2c20_6874, \9139 );
and \U$7060 ( \16175 , RIe211ae8_4491, \9141 );
and \U$7061 ( \16176 , RIfca2950_6872, \9143 );
and \U$7062 ( \16177 , RIe20ede8_4459, \9145 );
and \U$7063 ( \16178 , RIfcc24f8_7233, \9147 );
and \U$7064 ( \16179 , RIe20c0e8_4427, \9149 );
and \U$7065 ( \16180 , RIe2093e8_4395, \9151 );
and \U$7066 ( \16181 , RIe2066e8_4363, \9153 );
and \U$7067 ( \16182 , RIfc45110_5808, \9155 );
and \U$7068 ( \16183 , RIfcc6f80_7286, \9157 );
and \U$7069 ( \16184 , RIfe92f10_8016, \9159 );
and \U$7070 ( \16185 , RIfe92970_8012, \9161 );
and \U$7071 ( \16186 , RIf164af8_5605, \9163 );
and \U$7072 ( \16187 , RIf163a18_5593, \9165 );
and \U$7073 ( \16188 , RIf162aa0_5582, \9167 );
and \U$7074 ( \16189 , RIfe92ad8_8013, \9169 );
and \U$7075 ( \16190 , RIf15f3c8_5543, \9171 );
and \U$7076 ( \16191 , RIf15d640_5522, \9173 );
and \U$7077 ( \16192 , RIfe92808_8011, \9175 );
and \U$7078 ( \16193 , RIfe92c40_8014, \9177 );
and \U$7079 ( \16194 , RIfe926a0_8010, \9179 );
and \U$7080 ( \16195 , RIfe92da8_8015, \9181 );
and \U$7081 ( \16196 , RIfe92538_8009, \9183 );
and \U$7082 ( \16197 , RIfcb5a78_7089, \9185 );
or \U$7083 ( \16198 , \16134 , \16135 , \16136 , \16137 , \16138 , \16139 , \16140 , \16141 , \16142 , \16143 , \16144 , \16145 , \16146 , \16147 , \16148 , \16149 , \16150 , \16151 , \16152 , \16153 , \16154 , \16155 , \16156 , \16157 , \16158 , \16159 , \16160 , \16161 , \16162 , \16163 , \16164 , \16165 , \16166 , \16167 , \16168 , \16169 , \16170 , \16171 , \16172 , \16173 , \16174 , \16175 , \16176 , \16177 , \16178 , \16179 , \16180 , \16181 , \16182 , \16183 , \16184 , \16185 , \16186 , \16187 , \16188 , \16189 , \16190 , \16191 , \16192 , \16193 , \16194 , \16195 , \16196 , \16197 );
and \U$7084 ( \16199 , RIf158348_5463, \9188 );
and \U$7085 ( \16200 , RIf157100_5450, \9190 );
and \U$7086 ( \16201 , RIfc53be8_5975, \9192 );
and \U$7087 ( \16202 , RIfec38b8_8345, \9194 );
and \U$7088 ( \16203 , RIfcc5ea0_7274, \9196 );
and \U$7089 ( \16204 , RIf1550a8_5427, \9198 );
and \U$7090 ( \16205 , RIf153cf8_5413, \9200 );
and \U$7091 ( \16206 , RIfec3a20_8346, \9202 );
and \U$7092 ( \16207 , RIf152678_5397, \9204 );
and \U$7093 ( \16208 , RIfec3750_8344, \9206 );
and \U$7094 ( \16209 , RIf14ff18_5369, \9208 );
and \U$7095 ( \16210 , RIfe923d0_8008, \9210 );
and \U$7096 ( \16211 , RIf14efa0_5358, \9212 );
and \U$7097 ( \16212 , RIf14e898_5353, \9214 );
and \U$7098 ( \16213 , RIf14d380_5338, \9216 );
and \U$7099 ( \16214 , RIfe92268_8007, \9218 );
and \U$7100 ( \16215 , RIe1ea650_4044, \9220 );
and \U$7101 ( \16216 , RIe1e7950_4012, \9222 );
and \U$7102 ( \16217 , RIe1e4c50_3980, \9224 );
and \U$7103 ( \16218 , RIe1e1f50_3948, \9226 );
and \U$7104 ( \16219 , RIe1df250_3916, \9228 );
and \U$7105 ( \16220 , RIe1dc550_3884, \9230 );
and \U$7106 ( \16221 , RIe1d9850_3852, \9232 );
and \U$7107 ( \16222 , RIe1d6b50_3820, \9234 );
and \U$7108 ( \16223 , RIe1d1150_3756, \9236 );
and \U$7109 ( \16224 , RIe1ce450_3724, \9238 );
and \U$7110 ( \16225 , RIe1cb750_3692, \9240 );
and \U$7111 ( \16226 , RIe1c8a50_3660, \9242 );
and \U$7112 ( \16227 , RIe1c5d50_3628, \9244 );
and \U$7113 ( \16228 , RIe1c3050_3596, \9246 );
and \U$7114 ( \16229 , RIe1c0350_3564, \9248 );
and \U$7115 ( \16230 , RIe1bd650_3532, \9250 );
and \U$7116 ( \16231 , RIfcda4e0_7506, \9252 );
and \U$7117 ( \16232 , RIfc9d220_6810, \9254 );
and \U$7118 ( \16233 , RIe1b8628_3475, \9256 );
and \U$7119 ( \16234 , RIe1b6738_3453, \9258 );
and \U$7120 ( \16235 , RIfc4f2c8_5923, \9260 );
and \U$7121 ( \16236 , RIfce16c8_7587, \9262 );
and \U$7122 ( \16237 , RIfe91cc8_8003, \9264 );
and \U$7123 ( \16238 , RIfe91e30_8004, \9266 );
and \U$7124 ( \16239 , RIf1484c0_5282, \9268 );
and \U$7125 ( \16240 , RIf147548_5271, \9270 );
and \U$7126 ( \16241 , RIfe91f98_8005, \9272 );
and \U$7127 ( \16242 , RIfe91b60_8002, \9274 );
and \U$7128 ( \16243 , RIf146b70_5264, \9276 );
and \U$7129 ( \16244 , RIfc9f548_6835, \9278 );
and \U$7130 ( \16245 , RIfe92100_8006, \9280 );
and \U$7131 ( \16246 , RIfe919f8_8001, \9282 );
and \U$7132 ( \16247 , RIe1a7990_3284, \9284 );
and \U$7133 ( \16248 , RIe1a4c90_3252, \9286 );
and \U$7134 ( \16249 , RIe1a1f90_3220, \9288 );
and \U$7135 ( \16250 , RIe19f290_3188, \9290 );
and \U$7136 ( \16251 , RIe18b790_2964, \9292 );
and \U$7137 ( \16252 , RIe177c90_2740, \9294 );
and \U$7138 ( \16253 , RIe2255e8_4715, \9296 );
and \U$7139 ( \16254 , RIe21a1e8_4587, \9298 );
and \U$7140 ( \16255 , RIe2039e8_4331, \9300 );
and \U$7141 ( \16256 , RIe1fda48_4263, \9302 );
and \U$7142 ( \16257 , RIe1f6e00_4186, \9304 );
and \U$7143 ( \16258 , RIe1ef948_4103, \9306 );
and \U$7144 ( \16259 , RIe1d3e50_3788, \9308 );
and \U$7145 ( \16260 , RIe1ba950_3500, \9310 );
and \U$7146 ( \16261 , RIe1ad7c8_3351, \9312 );
and \U$7147 ( \16262 , RIe16fe00_2650, \9314 );
or \U$7148 ( \16263 , \16199 , \16200 , \16201 , \16202 , \16203 , \16204 , \16205 , \16206 , \16207 , \16208 , \16209 , \16210 , \16211 , \16212 , \16213 , \16214 , \16215 , \16216 , \16217 , \16218 , \16219 , \16220 , \16221 , \16222 , \16223 , \16224 , \16225 , \16226 , \16227 , \16228 , \16229 , \16230 , \16231 , \16232 , \16233 , \16234 , \16235 , \16236 , \16237 , \16238 , \16239 , \16240 , \16241 , \16242 , \16243 , \16244 , \16245 , \16246 , \16247 , \16248 , \16249 , \16250 , \16251 , \16252 , \16253 , \16254 , \16255 , \16256 , \16257 , \16258 , \16259 , \16260 , \16261 , \16262 );
or \U$7149 ( \16264 , \16198 , \16263 );
_DC g6596 ( \16265_nG6596 , \16264 , \9323 );
and g6597 ( \16266_nG6597 , \16133_nG6595 , \16265_nG6596 );
buf \U$7150 ( \16267 , \16266_nG6597 );
and \U$7151 ( \16268 , \16267 , \10691 );
nor \U$7152 ( \16269 , \16001 , \16268 );
xnor \U$7153 ( \16270 , \16269 , \10980 );
and \U$7154 ( \16271 , \12769 , \12790 );
and \U$7155 ( \16272 , \13679 , \12461 );
nor \U$7156 ( \16273 , \16271 , \16272 );
xnor \U$7157 ( \16274 , \16273 , \12780 );
xor \U$7158 ( \16275 , \16270 , \16274 );
and \U$7159 ( \16276 , \10988 , \15336 );
and \U$7160 ( \16277 , \11270 , \14963 );
nor \U$7161 ( \16278 , \16276 , \16277 );
xnor \U$7162 ( \16279 , \16278 , \15342 );
xor \U$7163 ( \16280 , \16275 , \16279 );
xor \U$7164 ( \16281 , \16000 , \16280 );
and \U$7165 ( \16282 , \15324 , \15328 );
and \U$7166 ( \16283 , \15328 , \15343 );
and \U$7167 ( \16284 , \15324 , \15343 );
or \U$7168 ( \16285 , \16282 , \16283 , \16284 );
and \U$7169 ( \16286 , \15349 , \15351 );
xor \U$7170 ( \16287 , \16285 , \16286 );
and \U$7171 ( \16288 , \14024 , \11574 );
and \U$7172 ( \16289 , \14950 , \11278 );
nor \U$7173 ( \16290 , \16288 , \16289 );
xnor \U$7174 ( \16291 , \16290 , \11580 );
and \U$7175 ( \16292 , \11586 , \14054 );
and \U$7176 ( \16293 , \12448 , \13692 );
nor \U$7177 ( \16294 , \16292 , \16293 );
xnor \U$7178 ( \16295 , \16294 , \14035 );
xor \U$7179 ( \16296 , \16291 , \16295 );
_DC g4f34 ( \16297_nG4f34 , \16132 , \9597 );
_DC g4fb8 ( \16298_nG4fb8 , \16264 , \9323 );
xor g4fb9 ( \16299_nG4fb9 , \16297_nG4f34 , \16298_nG4fb8 );
buf \U$7180 ( \16300 , \16299_nG4fb9 );
xor \U$7181 ( \16301 , \16300 , \15333 );
and \U$7182 ( \16302 , \10687 , \16301 );
xor \U$7183 ( \16303 , \16296 , \16302 );
xor \U$7184 ( \16304 , \16287 , \16303 );
xor \U$7185 ( \16305 , \16281 , \16304 );
and \U$7186 ( \16306 , \15054 , \15344 );
and \U$7187 ( \16307 , \15344 , \15362 );
and \U$7188 ( \16308 , \15054 , \15362 );
or \U$7189 ( \16309 , \16306 , \16307 , \16308 );
xor \U$7190 ( \16310 , \16305 , \16309 );
and \U$7191 ( \16311 , \15363 , \15367 );
and \U$7192 ( \16312 , \15368 , \15371 );
or \U$7193 ( \16313 , \16311 , \16312 );
xor \U$7194 ( \16314 , \16310 , \16313 );
buf g9bf0 ( \16315_nG9bf0 , \16314 );
and \U$7195 ( \16316 , \10704 , \16315_nG9bf0 );
or \U$7196 ( \16317 , \15996 , \16316 );
xor \U$7197 ( \16318 , \10703 , \16317 );
buf \U$7198 ( \16319 , \16318 );
buf \U$7200 ( \16320 , \16319 );
xor \U$7201 ( \16321 , \15995 , \16320 );
buf \U$7202 ( \16322 , \16321 );
xor \U$7203 ( \16323 , \15983 , \16322 );
buf \U$7204 ( \16324 , \16323 );
xor \U$7205 ( \16325 , \15952 , \16324 );
and \U$7206 ( \16326 , \15006 , \15380 );
and \U$7207 ( \16327 , \15006 , \15386 );
and \U$7208 ( \16328 , \15380 , \15386 );
or \U$7209 ( \16329 , \16326 , \16327 , \16328 );
buf \U$7210 ( \16330 , \16329 );
xor \U$7211 ( \16331 , \16325 , \16330 );
and \U$7212 ( \16332 , \15388 , \16331 );
and \U$7213 ( \16333 , \15946 , \16331 );
or \U$7214 ( \16334 , \15947 , \16332 , \16333 );
and \U$7215 ( \16335 , \15971 , \15973 );
and \U$7216 ( \16336 , \15971 , \15980 );
and \U$7217 ( \16337 , \15973 , \15980 );
or \U$7218 ( \16338 , \16335 , \16336 , \16337 );
buf \U$7219 ( \16339 , \16338 );
and \U$7220 ( \16340 , \10421 , \14984_nG9bf6 );
and \U$7221 ( \16341 , \10418 , \15373_nG9bf3 );
or \U$7222 ( \16342 , \16340 , \16341 );
xor \U$7223 ( \16343 , \10417 , \16342 );
buf \U$7224 ( \16344 , \16343 );
buf \U$7226 ( \16345 , \16344 );
xor \U$7227 ( \16346 , \16339 , \16345 );
and \U$7228 ( \16347 , \10707 , \16315_nG9bf0 );
and \U$7229 ( \16348 , \16285 , \16286 );
and \U$7230 ( \16349 , \16286 , \16303 );
and \U$7231 ( \16350 , \16285 , \16303 );
or \U$7232 ( \16351 , \16348 , \16349 , \16350 );
and \U$7233 ( \16352 , \14950 , \11574 );
and \U$7234 ( \16353 , \15321 , \11278 );
nor \U$7235 ( \16354 , \16352 , \16353 );
xnor \U$7236 ( \16355 , \16354 , \11580 );
not \U$7237 ( \16356 , \16302 );
and \U$7238 ( \16357 , RIdec4460_697, \9333 );
and \U$7239 ( \16358 , RIdec1760_665, \9335 );
and \U$7240 ( \16359 , RIee1fae0_4819, \9337 );
and \U$7241 ( \16360 , RIdebea60_633, \9339 );
and \U$7242 ( \16361 , RIee1f108_4812, \9341 );
and \U$7243 ( \16362 , RIdebbd60_601, \9343 );
and \U$7244 ( \16363 , RIdeb9060_569, \9345 );
and \U$7245 ( \16364 , RIdeb6360_537, \9347 );
and \U$7246 ( \16365 , RIee1eb68_4808, \9349 );
and \U$7247 ( \16366 , RIdeb0960_473, \9351 );
and \U$7248 ( \16367 , RIee1e460_4803, \9353 );
and \U$7249 ( \16368 , RIdeadc60_441, \9355 );
and \U$7250 ( \16369 , RIee1d7b8_4794, \9357 );
and \U$7251 ( \16370 , RIdea8008_409, \9359 );
and \U$7252 ( \16371 , RIdea1708_377, \9361 );
and \U$7253 ( \16372 , RIde9ae08_345, \9363 );
and \U$7254 ( \16373 , RIfe957d8_8045, \9365 );
and \U$7255 ( \16374 , RIfe95508_8043, \9367 );
and \U$7256 ( \16375 , RIfe95670_8044, \9369 );
and \U$7257 ( \16376 , RIee1a7e8_4760, \9371 );
and \U$7258 ( \16377 , RIfe95aa8_8047, \9373 );
and \U$7259 ( \16378 , RIfe95238_8041, \9375 );
and \U$7260 ( \16379 , RIfe95940_8046, \9377 );
and \U$7261 ( \16380 , RIfe953a0_8042, \9379 );
and \U$7262 ( \16381 , RIee1a0e0_4755, \9381 );
and \U$7263 ( \16382 , RIee19ca8_4752, \9383 );
and \U$7264 ( \16383 , RIee19870_4749, \9385 );
and \U$7265 ( \16384 , RIee19438_4746, \9387 );
and \U$7266 ( \16385 , RIee38ba8_5104, \9389 );
and \U$7267 ( \16386 , RIfe95c10_8048, \9391 );
and \U$7268 ( \16387 , RIee384a0_5099, \9393 );
and \U$7269 ( \16388 , RIfea9440_8242, \9395 );
and \U$7270 ( \16389 , RIe164460_2518, \9397 );
and \U$7271 ( \16390 , RIe161760_2486, \9399 );
and \U$7272 ( \16391 , RIfe942c0_8030, \9401 );
and \U$7273 ( \16392 , RIe15ea60_2454, \9403 );
and \U$7274 ( \16393 , RIfe94158_8029, \9405 );
and \U$7275 ( \16394 , RIe15bd60_2422, \9407 );
and \U$7276 ( \16395 , RIe156360_2358, \9409 );
and \U$7277 ( \16396 , RIe153660_2326, \9411 );
and \U$7278 ( \16397 , RIfe94428_8031, \9413 );
and \U$7279 ( \16398 , RIe150960_2294, \9415 );
and \U$7280 ( \16399 , RIfe94590_8032, \9417 );
and \U$7281 ( \16400 , RIe14dc60_2262, \9419 );
and \U$7282 ( \16401 , RIfc5c2e8_6071, \9421 );
and \U$7283 ( \16402 , RIe14af60_2230, \9423 );
and \U$7284 ( \16403 , RIe148260_2198, \9425 );
and \U$7285 ( \16404 , RIe145560_2166, \9427 );
and \U$7286 ( \16405 , RIee33ce8_5048, \9429 );
and \U$7287 ( \16406 , RIee32aa0_5035, \9431 );
and \U$7288 ( \16407 , RIee31858_5022, \9433 );
and \U$7289 ( \16408 , RIfc5d530_6084, \9435 );
and \U$7290 ( \16409 , RIe140538_2109, \9437 );
and \U$7291 ( \16410 , RIdf3e2d8_2084, \9439 );
and \U$7292 ( \16411 , RIdf3c118_2060, \9441 );
and \U$7293 ( \16412 , RIdf39df0_2035, \9443 );
and \U$7294 ( \16413 , RIfcdd780_7542, \9445 );
and \U$7295 ( \16414 , RIee2ee28_4992, \9447 );
and \U$7296 ( \16415 , RIfcc88d0_7304, \9449 );
and \U$7297 ( \16416 , RIee2cc68_4968, \9451 );
and \U$7298 ( \16417 , RIdf34990_1975, \9453 );
and \U$7299 ( \16418 , RIdf32aa0_1953, \9455 );
and \U$7300 ( \16419 , RIdf304a8_1926, \9457 );
and \U$7301 ( \16420 , RIdf2e5b8_1904, \9459 );
or \U$7302 ( \16421 , \16357 , \16358 , \16359 , \16360 , \16361 , \16362 , \16363 , \16364 , \16365 , \16366 , \16367 , \16368 , \16369 , \16370 , \16371 , \16372 , \16373 , \16374 , \16375 , \16376 , \16377 , \16378 , \16379 , \16380 , \16381 , \16382 , \16383 , \16384 , \16385 , \16386 , \16387 , \16388 , \16389 , \16390 , \16391 , \16392 , \16393 , \16394 , \16395 , \16396 , \16397 , \16398 , \16399 , \16400 , \16401 , \16402 , \16403 , \16404 , \16405 , \16406 , \16407 , \16408 , \16409 , \16410 , \16411 , \16412 , \16413 , \16414 , \16415 , \16416 , \16417 , \16418 , \16419 , \16420 );
and \U$7303 ( \16422 , RIee2b1b0_4949, \9462 );
and \U$7304 ( \16423 , RIfe946f8_8033, \9464 );
and \U$7305 ( \16424 , RIfcb2940_7054, \9466 );
and \U$7306 ( \16425 , RIee273d0_4905, \9468 );
and \U$7307 ( \16426 , RIfe949c8_8035, \9470 );
and \U$7308 ( \16427 , RIdf27538_1824, \9472 );
and \U$7309 ( \16428 , RIfe94b30_8036, \9474 );
and \U$7310 ( \16429 , RIfe94860_8034, \9476 );
and \U$7311 ( \16430 , RIee26f98_4902, \9478 );
and \U$7312 ( \16431 , RIee269f8_4898, \9480 );
and \U$7313 ( \16432 , RIee26728_4896, \9482 );
and \U$7314 ( \16433 , RIee26458_4894, \9484 );
and \U$7315 ( \16434 , RIee26188_4892, \9486 );
and \U$7316 ( \16435 , RIfe94c98_8037, \9488 );
and \U$7317 ( \16436 , RIee25d50_4889, \9490 );
and \U$7318 ( \16437 , RIfea9170_8240, \9492 );
and \U$7319 ( \16438 , RIdf16030_1627, \9494 );
and \U$7320 ( \16439 , RIdf13330_1595, \9496 );
and \U$7321 ( \16440 , RIdf10630_1563, \9498 );
and \U$7322 ( \16441 , RIdf0d930_1531, \9500 );
and \U$7323 ( \16442 , RIdf0ac30_1499, \9502 );
and \U$7324 ( \16443 , RIdf07f30_1467, \9504 );
and \U$7325 ( \16444 , RIdf05230_1435, \9506 );
and \U$7326 ( \16445 , RIdf02530_1403, \9508 );
and \U$7327 ( \16446 , RIdefcb30_1339, \9510 );
and \U$7328 ( \16447 , RIdef9e30_1307, \9512 );
and \U$7329 ( \16448 , RIdef7130_1275, \9514 );
and \U$7330 ( \16449 , RIdef4430_1243, \9516 );
and \U$7331 ( \16450 , RIdef1730_1211, \9518 );
and \U$7332 ( \16451 , RIdeeea30_1179, \9520 );
and \U$7333 ( \16452 , RIdeebd30_1147, \9522 );
and \U$7334 ( \16453 , RIdee9030_1115, \9524 );
and \U$7335 ( \16454 , RIee250a8_4880, \9526 );
and \U$7336 ( \16455 , RIee24298_4870, \9528 );
and \U$7337 ( \16456 , RIee23758_4862, \9530 );
and \U$7338 ( \16457 , RIee22d80_4855, \9532 );
and \U$7339 ( \16458 , RIfe950d0_8040, \9534 );
and \U$7340 ( \16459 , RIfe94f68_8039, \9536 );
and \U$7341 ( \16460 , RIfe94e00_8038, \9538 );
and \U$7342 ( \16461 , RIdeddd98_988, \9540 );
and \U$7343 ( \16462 , RIee22ab0_4853, \9542 );
and \U$7344 ( \16463 , RIee21e08_4844, \9544 );
and \U$7345 ( \16464 , RIfca46d8_6893, \9546 );
and \U$7346 ( \16465 , RIfc5dad0_6088, \9548 );
and \U$7347 ( \16466 , RIfeaa250_8252, \9550 );
and \U$7348 ( \16467 , RIfe96048_8051, \9552 );
and \U$7349 ( \16468 , RIfe95d78_8049, \9554 );
and \U$7350 ( \16469 , RIfe95ee0_8050, \9556 );
and \U$7351 ( \16470 , RIdecf860_825, \9558 );
and \U$7352 ( \16471 , RIdeccb60_793, \9560 );
and \U$7353 ( \16472 , RIdec9e60_761, \9562 );
and \U$7354 ( \16473 , RIdec7160_729, \9564 );
and \U$7355 ( \16474 , RIdeb3660_505, \9566 );
and \U$7356 ( \16475 , RIde94508_313, \9568 );
and \U$7357 ( \16476 , RIe16d268_2619, \9570 );
and \U$7358 ( \16477 , RIe159060_2390, \9572 );
and \U$7359 ( \16478 , RIe142860_2134, \9574 );
and \U$7360 ( \16479 , RIdf37258_2004, \9576 );
and \U$7361 ( \16480 , RIdf2b8b8_1872, \9578 );
and \U$7362 ( \16481 , RIdf1c138_1696, \9580 );
and \U$7363 ( \16482 , RIdeff830_1371, \9582 );
and \U$7364 ( \16483 , RIdee6330_1083, \9584 );
and \U$7365 ( \16484 , RIdedb098_956, \9586 );
and \U$7366 ( \16485 , RIde7a450_186, \9588 );
or \U$7367 ( \16486 , \16422 , \16423 , \16424 , \16425 , \16426 , \16427 , \16428 , \16429 , \16430 , \16431 , \16432 , \16433 , \16434 , \16435 , \16436 , \16437 , \16438 , \16439 , \16440 , \16441 , \16442 , \16443 , \16444 , \16445 , \16446 , \16447 , \16448 , \16449 , \16450 , \16451 , \16452 , \16453 , \16454 , \16455 , \16456 , \16457 , \16458 , \16459 , \16460 , \16461 , \16462 , \16463 , \16464 , \16465 , \16466 , \16467 , \16468 , \16469 , \16470 , \16471 , \16472 , \16473 , \16474 , \16475 , \16476 , \16477 , \16478 , \16479 , \16480 , \16481 , \16482 , \16483 , \16484 , \16485 );
or \U$7368 ( \16487 , \16421 , \16486 );
_DC g503d ( \16488_nG503d , \16487 , \9597 );
and \U$7369 ( \16489 , RIe19c6f8_3157, \9059 );
and \U$7370 ( \16490 , RIe1999f8_3125, \9061 );
and \U$7371 ( \16491 , RIf1450b8_5245, \9063 );
and \U$7372 ( \16492 , RIe196cf8_3093, \9065 );
and \U$7373 ( \16493 , RIf143fd8_5233, \9067 );
and \U$7374 ( \16494 , RIe193ff8_3061, \9069 );
and \U$7375 ( \16495 , RIe1912f8_3029, \9071 );
and \U$7376 ( \16496 , RIe18e5f8_2997, \9073 );
and \U$7377 ( \16497 , RIe188bf8_2933, \9075 );
and \U$7378 ( \16498 , RIe185ef8_2901, \9077 );
and \U$7379 ( \16499 , RIfe973f8_8065, \9079 );
and \U$7380 ( \16500 , RIe1831f8_2869, \9081 );
and \U$7381 ( \16501 , RIf142958_5217, \9083 );
and \U$7382 ( \16502 , RIe1804f8_2837, \9085 );
and \U$7383 ( \16503 , RIe17d7f8_2805, \9087 );
and \U$7384 ( \16504 , RIe17aaf8_2773, \9089 );
and \U$7385 ( \16505 , RIf141b48_5207, \9091 );
and \U$7386 ( \16506 , RIfc542f0_5980, \9093 );
and \U$7387 ( \16507 , RIfc800a8_6479, \9095 );
and \U$7388 ( \16508 , RIe175260_2710, \9097 );
and \U$7389 ( \16509 , RIfca0bc8_6851, \9099 );
and \U$7390 ( \16510 , RIfc48680_5846, \9101 );
and \U$7391 ( \16511 , RIee3dea0_5163, \9103 );
and \U$7392 ( \16512 , RIfcc6878_7281, \9105 );
and \U$7393 ( \16513 , RIee3ba10_5137, \9107 );
and \U$7394 ( \16514 , RIee3a930_5125, \9109 );
and \U$7395 ( \16515 , RIfe97290_8064, \9111 );
and \U$7396 ( \16516 , RIe172b00_2682, \9113 );
and \U$7397 ( \16517 , RIf16f958_5729, \9115 );
and \U$7398 ( \16518 , RIf16ee18_5721, \9117 );
and \U$7399 ( \16519 , RIf16da68_5707, \9119 );
and \U$7400 ( \16520 , RIf16d360_5702, \9121 );
and \U$7401 ( \16521 , RIfe96e58_8061, \9123 );
and \U$7402 ( \16522 , RIe222a50_4684, \9125 );
and \U$7403 ( \16523 , RIfe96cf0_8060, \9127 );
and \U$7404 ( \16524 , RIe21fd50_4652, \9129 );
and \U$7405 ( \16525 , RIf16a660_5670, \9131 );
and \U$7406 ( \16526 , RIe21d050_4620, \9133 );
and \U$7407 ( \16527 , RIe217650_4556, \9135 );
and \U$7408 ( \16528 , RIe214950_4524, \9137 );
and \U$7409 ( \16529 , RIf169f58_5665, \9139 );
and \U$7410 ( \16530 , RIe211c50_4492, \9141 );
and \U$7411 ( \16531 , RIf168770_5648, \9143 );
and \U$7412 ( \16532 , RIe20ef50_4460, \9145 );
and \U$7413 ( \16533 , RIf1677f8_5637, \9147 );
and \U$7414 ( \16534 , RIe20c250_4428, \9149 );
and \U$7415 ( \16535 , RIe209550_4396, \9151 );
and \U$7416 ( \16536 , RIe206850_4364, \9153 );
and \U$7417 ( \16537 , RIf166880_5626, \9155 );
and \U$7418 ( \16538 , RIf1657a0_5614, \9157 );
and \U$7419 ( \16539 , RIe201dc8_4311, \9159 );
and \U$7420 ( \16540 , RIe2005e0_4294, \9161 );
and \U$7421 ( \16541 , RIfe96b88_8059, \9163 );
and \U$7422 ( \16542 , RIf163b80_5594, \9165 );
and \U$7423 ( \16543 , RIf162c08_5583, \9167 );
and \U$7424 ( \16544 , RIf161420_5566, \9169 );
and \U$7425 ( \16545 , RIf15f530_5544, \9171 );
and \U$7426 ( \16546 , RIf15d7a8_5523, \9173 );
and \U$7427 ( \16547 , RIfe968b8_8057, \9175 );
and \U$7428 ( \16548 , RIfe96a20_8058, \9177 );
and \U$7429 ( \16549 , RIfcb3fc0_7070, \9179 );
and \U$7430 ( \16550 , RIfc7cf70_6444, \9181 );
and \U$7431 ( \16551 , RIfc579c8_6019, \9183 );
and \U$7432 ( \16552 , RIf159590_5476, \9185 );
or \U$7433 ( \16553 , \16489 , \16490 , \16491 , \16492 , \16493 , \16494 , \16495 , \16496 , \16497 , \16498 , \16499 , \16500 , \16501 , \16502 , \16503 , \16504 , \16505 , \16506 , \16507 , \16508 , \16509 , \16510 , \16511 , \16512 , \16513 , \16514 , \16515 , \16516 , \16517 , \16518 , \16519 , \16520 , \16521 , \16522 , \16523 , \16524 , \16525 , \16526 , \16527 , \16528 , \16529 , \16530 , \16531 , \16532 , \16533 , \16534 , \16535 , \16536 , \16537 , \16538 , \16539 , \16540 , \16541 , \16542 , \16543 , \16544 , \16545 , \16546 , \16547 , \16548 , \16549 , \16550 , \16551 , \16552 );
and \U$7434 ( \16554 , RIf1584b0_5464, \9188 );
and \U$7435 ( \16555 , RIf157268_5451, \9190 );
and \U$7436 ( \16556 , RIf1569f8_5445, \9192 );
and \U$7437 ( \16557 , RIfe965e8_8055, \9194 );
and \U$7438 ( \16558 , RIf155d50_5436, \9196 );
and \U$7439 ( \16559 , RIf155210_5428, \9198 );
and \U$7440 ( \16560 , RIf153e60_5414, \9200 );
and \U$7441 ( \16561 , RIfe96750_8056, \9202 );
and \U$7442 ( \16562 , RIf1527e0_5398, \9204 );
and \U$7443 ( \16563 , RIf151430_5384, \9206 );
and \U$7444 ( \16564 , RIfcd2650_7416, \9208 );
and \U$7445 ( \16565 , RIe1f2648_4135, \9210 );
and \U$7446 ( \16566 , RIf14f108_5359, \9212 );
and \U$7447 ( \16567 , RIfc7f298_6469, \9214 );
and \U$7448 ( \16568 , RIf14d4e8_5339, \9216 );
and \U$7449 ( \16569 , RIe1ed350_4076, \9218 );
and \U$7450 ( \16570 , RIe1ea7b8_4045, \9220 );
and \U$7451 ( \16571 , RIe1e7ab8_4013, \9222 );
and \U$7452 ( \16572 , RIe1e4db8_3981, \9224 );
and \U$7453 ( \16573 , RIe1e20b8_3949, \9226 );
and \U$7454 ( \16574 , RIe1df3b8_3917, \9228 );
and \U$7455 ( \16575 , RIe1dc6b8_3885, \9230 );
and \U$7456 ( \16576 , RIe1d99b8_3853, \9232 );
and \U$7457 ( \16577 , RIe1d6cb8_3821, \9234 );
and \U$7458 ( \16578 , RIe1d12b8_3757, \9236 );
and \U$7459 ( \16579 , RIe1ce5b8_3725, \9238 );
and \U$7460 ( \16580 , RIe1cb8b8_3693, \9240 );
and \U$7461 ( \16581 , RIe1c8bb8_3661, \9242 );
and \U$7462 ( \16582 , RIe1c5eb8_3629, \9244 );
and \U$7463 ( \16583 , RIe1c31b8_3597, \9246 );
and \U$7464 ( \16584 , RIe1c04b8_3565, \9248 );
and \U$7465 ( \16585 , RIe1bd7b8_3533, \9250 );
and \U$7466 ( \16586 , RIf14c138_5325, \9252 );
and \U$7467 ( \16587 , RIf14ad88_5311, \9254 );
and \U$7468 ( \16588 , RIe1b8790_3476, \9256 );
and \U$7469 ( \16589 , RIfe96480_8054, \9258 );
and \U$7470 ( \16590 , RIf14a0e0_5302, \9260 );
and \U$7471 ( \16591 , RIf149870_5296, \9262 );
and \U$7472 ( \16592 , RIfe97128_8063, \9264 );
and \U$7473 ( \16593 , RIfe96318_8053, \9266 );
and \U$7474 ( \16594 , RIf148628_5283, \9268 );
and \U$7475 ( \16595 , RIfc58d78_6033, \9270 );
and \U$7476 ( \16596 , RIe1b20e8_3403, \9272 );
and \U$7477 ( \16597 , RIe1b04c8_3383, \9274 );
and \U$7478 ( \16598 , RIf146cd8_5265, \9276 );
and \U$7479 ( \16599 , RIfc591b0_6036, \9278 );
and \U$7480 ( \16600 , RIfe961b0_8052, \9280 );
and \U$7481 ( \16601 , RIfe96fc0_8062, \9282 );
and \U$7482 ( \16602 , RIe1a7af8_3285, \9284 );
and \U$7483 ( \16603 , RIe1a4df8_3253, \9286 );
and \U$7484 ( \16604 , RIe1a20f8_3221, \9288 );
and \U$7485 ( \16605 , RIe19f3f8_3189, \9290 );
and \U$7486 ( \16606 , RIe18b8f8_2965, \9292 );
and \U$7487 ( \16607 , RIe177df8_2741, \9294 );
and \U$7488 ( \16608 , RIe225750_4716, \9296 );
and \U$7489 ( \16609 , RIe21a350_4588, \9298 );
and \U$7490 ( \16610 , RIe203b50_4332, \9300 );
and \U$7491 ( \16611 , RIe1fdbb0_4264, \9302 );
and \U$7492 ( \16612 , RIe1f6f68_4187, \9304 );
and \U$7493 ( \16613 , RIe1efab0_4104, \9306 );
and \U$7494 ( \16614 , RIe1d3fb8_3789, \9308 );
and \U$7495 ( \16615 , RIe1baab8_3501, \9310 );
and \U$7496 ( \16616 , RIe1ad930_3352, \9312 );
and \U$7497 ( \16617 , RIe16ff68_2651, \9314 );
or \U$7498 ( \16618 , \16554 , \16555 , \16556 , \16557 , \16558 , \16559 , \16560 , \16561 , \16562 , \16563 , \16564 , \16565 , \16566 , \16567 , \16568 , \16569 , \16570 , \16571 , \16572 , \16573 , \16574 , \16575 , \16576 , \16577 , \16578 , \16579 , \16580 , \16581 , \16582 , \16583 , \16584 , \16585 , \16586 , \16587 , \16588 , \16589 , \16590 , \16591 , \16592 , \16593 , \16594 , \16595 , \16596 , \16597 , \16598 , \16599 , \16600 , \16601 , \16602 , \16603 , \16604 , \16605 , \16606 , \16607 , \16608 , \16609 , \16610 , \16611 , \16612 , \16613 , \16614 , \16615 , \16616 , \16617 );
or \U$7499 ( \16619 , \16553 , \16618 );
_DC g50c1 ( \16620_nG50c1 , \16619 , \9323 );
xor g50c2 ( \16621_nG50c2 , \16488_nG503d , \16620_nG50c1 );
buf \U$7500 ( \16622 , \16621_nG50c2 );
and \U$7501 ( \16623 , \16300 , \15333 );
not \U$7502 ( \16624 , \16623 );
and \U$7503 ( \16625 , \16622 , \16624 );
and \U$7504 ( \16626 , \16356 , \16625 );
xor \U$7505 ( \16627 , \16355 , \16626 );
and \U$7506 ( \16628 , \13679 , \12790 );
and \U$7507 ( \16629 , \14024 , \12461 );
nor \U$7508 ( \16630 , \16628 , \16629 );
xnor \U$7509 ( \16631 , \16630 , \12780 );
xor \U$7510 ( \16632 , \16627 , \16631 );
xor \U$7511 ( \16633 , \16622 , \16300 );
not \U$7512 ( \16634 , \16301 );
and \U$7513 ( \16635 , \16633 , \16634 );
and \U$7514 ( \16636 , \10687 , \16635 );
and \U$7515 ( \16637 , \10988 , \16301 );
nor \U$7516 ( \16638 , \16636 , \16637 );
xnor \U$7517 ( \16639 , \16638 , \16625 );
xor \U$7518 ( \16640 , \16632 , \16639 );
xor \U$7519 ( \16641 , \16351 , \16640 );
and \U$7520 ( \16642 , \16291 , \16295 );
and \U$7521 ( \16643 , \16295 , \16302 );
and \U$7522 ( \16644 , \16291 , \16302 );
or \U$7523 ( \16645 , \16642 , \16643 , \16644 );
and \U$7524 ( \16646 , \16270 , \16274 );
and \U$7525 ( \16647 , \16274 , \16279 );
and \U$7526 ( \16648 , \16270 , \16279 );
or \U$7527 ( \16649 , \16646 , \16647 , \16648 );
xor \U$7528 ( \16650 , \16645 , \16649 );
and \U$7529 ( \16651 , \16267 , \10983 );
_DC g6598 ( \16652_nG6598 , \16487 , \9597 );
_DC g6599 ( \16653_nG6599 , \16619 , \9323 );
and g659a ( \16654_nG659a , \16652_nG6598 , \16653_nG6599 );
buf \U$7530 ( \16655 , \16654_nG659a );
and \U$7531 ( \16656 , \16655 , \10691 );
nor \U$7532 ( \16657 , \16651 , \16656 );
xnor \U$7533 ( \16658 , \16657 , \10980 );
and \U$7534 ( \16659 , \12448 , \14054 );
and \U$7535 ( \16660 , \12769 , \13692 );
nor \U$7536 ( \16661 , \16659 , \16660 );
xnor \U$7537 ( \16662 , \16661 , \14035 );
xor \U$7538 ( \16663 , \16658 , \16662 );
and \U$7539 ( \16664 , \11270 , \15336 );
and \U$7540 ( \16665 , \11586 , \14963 );
nor \U$7541 ( \16666 , \16664 , \16665 );
xnor \U$7542 ( \16667 , \16666 , \15342 );
xor \U$7543 ( \16668 , \16663 , \16667 );
xor \U$7544 ( \16669 , \16650 , \16668 );
xor \U$7545 ( \16670 , \16641 , \16669 );
and \U$7546 ( \16671 , \16000 , \16280 );
and \U$7547 ( \16672 , \16280 , \16304 );
and \U$7548 ( \16673 , \16000 , \16304 );
or \U$7549 ( \16674 , \16671 , \16672 , \16673 );
xor \U$7550 ( \16675 , \16670 , \16674 );
and \U$7551 ( \16676 , \16305 , \16309 );
and \U$7552 ( \16677 , \16310 , \16313 );
or \U$7553 ( \16678 , \16676 , \16677 );
xor \U$7554 ( \16679 , \16675 , \16678 );
buf g9bed ( \16680_nG9bed , \16679 );
and \U$7555 ( \16681 , \10704 , \16680_nG9bed );
or \U$7556 ( \16682 , \16347 , \16681 );
xor \U$7557 ( \16683 , \10703 , \16682 );
buf \U$7558 ( \16684 , \16683 );
buf \U$7560 ( \16685 , \16684 );
xor \U$7561 ( \16686 , \16346 , \16685 );
buf \U$7562 ( \16687 , \16686 );
and \U$7563 ( \16688 , \15988 , \15994 );
and \U$7564 ( \16689 , \15988 , \16320 );
and \U$7565 ( \16690 , \15994 , \16320 );
or \U$7566 ( \16691 , \16688 , \16689 , \16690 );
buf \U$7567 ( \16692 , \16691 );
xor \U$7568 ( \16693 , \16687 , \16692 );
and \U$7569 ( \16694 , \15936 , \15943 );
buf \U$7570 ( \16695 , \16694 );
buf \U$7572 ( \16696 , \16695 );
and \U$7573 ( \16697 , \14631 , \11283_nG9c08 );
and \U$7574 ( \16698 , \14628 , \11598_nG9c05 );
or \U$7575 ( \16699 , \16697 , \16698 );
xor \U$7576 ( \16700 , \14627 , \16699 );
buf \U$7577 ( \16701 , \16700 );
buf \U$7579 ( \16702 , \16701 );
xor \U$7580 ( \16703 , \16696 , \16702 );
buf \U$7581 ( \16704 , \16703 );
and \U$7582 ( \16705 , \15940 , \10694_nG9c0e );
and \U$7583 ( \16706 , \15937 , \10995_nG9c0b );
or \U$7584 ( \16707 , \16705 , \16706 );
xor \U$7585 ( \16708 , \15936 , \16707 );
buf \U$7586 ( \16709 , \16708 );
buf \U$7588 ( \16710 , \16709 );
xor \U$7589 ( \16711 , \16704 , \16710 );
and \U$7590 ( \16712 , \13370 , \12470_nG9c02 );
and \U$7591 ( \16713 , \13367 , \12801_nG9bff );
or \U$7592 ( \16714 , \16712 , \16713 );
xor \U$7593 ( \16715 , \13366 , \16714 );
buf \U$7594 ( \16716 , \16715 );
buf \U$7596 ( \16717 , \16716 );
xor \U$7597 ( \16718 , \16711 , \16717 );
buf \U$7598 ( \16719 , \16718 );
and \U$7599 ( \16720 , \15963 , \15969 );
buf \U$7600 ( \16721 , \16720 );
xor \U$7601 ( \16722 , \16719 , \16721 );
and \U$7602 ( \16723 , \12157 , \13705_nG9bfc );
and \U$7603 ( \16724 , \12154 , \14070_nG9bf9 );
or \U$7604 ( \16725 , \16723 , \16724 );
xor \U$7605 ( \16726 , \12153 , \16725 );
buf \U$7606 ( \16727 , \16726 );
buf \U$7608 ( \16728 , \16727 );
xor \U$7609 ( \16729 , \16722 , \16728 );
buf \U$7610 ( \16730 , \16729 );
xor \U$7611 ( \16731 , \16693 , \16730 );
buf \U$7612 ( \16732 , \16731 );
and \U$7613 ( \16733 , \15957 , \15982 );
and \U$7614 ( \16734 , \15957 , \16322 );
and \U$7615 ( \16735 , \15982 , \16322 );
or \U$7616 ( \16736 , \16733 , \16734 , \16735 );
buf \U$7617 ( \16737 , \16736 );
xor \U$7618 ( \16738 , \16732 , \16737 );
and \U$7619 ( \16739 , \15952 , \16324 );
and \U$7620 ( \16740 , \15952 , \16330 );
and \U$7621 ( \16741 , \16324 , \16330 );
or \U$7622 ( \16742 , \16739 , \16740 , \16741 );
buf \U$7623 ( \16743 , \16742 );
xor \U$7624 ( \16744 , \16738 , \16743 );
and \U$7625 ( \16745 , \16334 , \16744 );
and \U$7626 ( \16746 , RIdec4730_699, \9059 );
and \U$7627 ( \16747 , RIdec1a30_667, \9061 );
and \U$7628 ( \16748 , RIfce3f90_7616, \9063 );
and \U$7629 ( \16749 , RIdebed30_635, \9065 );
and \U$7630 ( \16750 , RIfcc3308_7243, \9067 );
and \U$7631 ( \16751 , RIdebc030_603, \9069 );
and \U$7632 ( \16752 , RIdeb9330_571, \9071 );
and \U$7633 ( \16753 , RIdeb6630_539, \9073 );
and \U$7634 ( \16754 , RIfc8c588_6619, \9075 );
and \U$7635 ( \16755 , RIdeb0c30_475, \9077 );
and \U$7636 ( \16756 , RIfc5a998_6053, \9079 );
and \U$7637 ( \16757 , RIdeadf30_443, \9081 );
and \U$7638 ( \16758 , RIfc99b48_6771, \9083 );
and \U$7639 ( \16759 , RIdea8698_411, \9085 );
and \U$7640 ( \16760 , RIdea1d98_379, \9087 );
and \U$7641 ( \16761 , RIde9b498_347, \9089 );
and \U$7642 ( \16762 , RIfc78bf0_6396, \9091 );
and \U$7643 ( \16763 , RIfcbc558_7165, \9093 );
and \U$7644 ( \16764 , RIfca12d0_6856, \9095 );
and \U$7645 ( \16765 , RIfca3fd0_6888, \9097 );
and \U$7646 ( \16766 , RIfec2670_8332, \9099 );
and \U$7647 ( \16767 , RIfec2508_8331, \9101 );
and \U$7648 ( \16768 , RIde88a00_256, \9103 );
and \U$7649 ( \16769 , RIde84518_235, \9105 );
and \U$7650 ( \16770 , RIfcc35d8_7245, \9107 );
and \U$7651 ( \16771 , RIfcb57a8_7087, \9109 );
and \U$7652 ( \16772 , RIfc5a290_6048, \9111 );
and \U$7653 ( \16773 , RIfca3058_6877, \9113 );
and \U$7654 ( \16774 , RIee38e78_5106, \9115 );
and \U$7655 ( \16775 , RIfec27d8_8333, \9117 );
and \U$7656 ( \16776 , RIfca3328_6879, \9119 );
and \U$7657 ( \16777 , RIe1672c8_2551, \9121 );
and \U$7658 ( \16778 , RIe164730_2520, \9123 );
and \U$7659 ( \16779 , RIe161a30_2488, \9125 );
and \U$7660 ( \16780 , RIee36cb8_5082, \9127 );
and \U$7661 ( \16781 , RIe15ed30_2456, \9129 );
and \U$7662 ( \16782 , RIfcc7250_7288, \9131 );
and \U$7663 ( \16783 , RIe15c030_2424, \9133 );
and \U$7664 ( \16784 , RIe156630_2360, \9135 );
and \U$7665 ( \16785 , RIe153930_2328, \9137 );
and \U$7666 ( \16786 , RIfcc7688_7291, \9139 );
and \U$7667 ( \16787 , RIe150c30_2296, \9141 );
and \U$7668 ( \16788 , RIfc8af08_6603, \9143 );
and \U$7669 ( \16789 , RIe14df30_2264, \9145 );
and \U$7670 ( \16790 , RIfc9a250_6776, \9147 );
and \U$7671 ( \16791 , RIe14b230_2232, \9149 );
and \U$7672 ( \16792 , RIe148530_2200, \9151 );
and \U$7673 ( \16793 , RIe145830_2168, \9153 );
and \U$7674 ( \16794 , RIfc9aac0_6782, \9155 );
and \U$7675 ( \16795 , RIfc56bb8_6009, \9157 );
and \U$7676 ( \16796 , RIfca1ca8_6863, \9159 );
and \U$7677 ( \16797 , RIfcec960_7714, \9161 );
and \U$7678 ( \16798 , RIe1406a0_2110, \9163 );
and \U$7679 ( \16799 , RIdf3e440_2085, \9165 );
and \U$7680 ( \16800 , RIdf3c280_2061, \9167 );
and \U$7681 ( \16801 , RIdf39f58_2036, \9169 );
and \U$7682 ( \16802 , RIfc9a958_6781, \9171 );
and \U$7683 ( \16803 , RIee2f0f8_4994, \9173 );
and \U$7684 ( \16804 , RIfcdb458_7517, \9175 );
and \U$7685 ( \16805 , RIee2cf38_4970, \9177 );
and \U$7686 ( \16806 , RIdf34c60_1977, \9179 );
and \U$7687 ( \16807 , RIfec2940_8334, \9181 );
and \U$7688 ( \16808 , RIdf30778_1928, \9183 );
and \U$7689 ( \16809 , RIdf2e888_1906, \9185 );
or \U$7690 ( \16810 , \16746 , \16747 , \16748 , \16749 , \16750 , \16751 , \16752 , \16753 , \16754 , \16755 , \16756 , \16757 , \16758 , \16759 , \16760 , \16761 , \16762 , \16763 , \16764 , \16765 , \16766 , \16767 , \16768 , \16769 , \16770 , \16771 , \16772 , \16773 , \16774 , \16775 , \16776 , \16777 , \16778 , \16779 , \16780 , \16781 , \16782 , \16783 , \16784 , \16785 , \16786 , \16787 , \16788 , \16789 , \16790 , \16791 , \16792 , \16793 , \16794 , \16795 , \16796 , \16797 , \16798 , \16799 , \16800 , \16801 , \16802 , \16803 , \16804 , \16805 , \16806 , \16807 , \16808 , \16809 );
and \U$7691 ( \16811 , RIee2b480_4951, \9188 );
and \U$7692 ( \16812 , RIfec23a0_8330, \9190 );
and \U$7693 ( \16813 , RIee288e8_4920, \9192 );
and \U$7694 ( \16814 , RIfec2238_8329, \9194 );
and \U$7695 ( \16815 , RIdf29b30_1851, \9196 );
and \U$7696 ( \16816 , RIdf27808_1826, \9198 );
and \U$7697 ( \16817 , RIdf25a80_1805, \9200 );
and \U$7698 ( \16818 , RIdf23e60_1785, \9202 );
and \U$7699 ( \16819 , RIfc55100_5990, \9204 );
and \U$7700 ( \16820 , RIfcd9f40_7502, \9206 );
and \U$7701 ( \16821 , RIfc54f98_5989, \9208 );
and \U$7702 ( \16822 , RIfc54cc8_5987, \9210 );
and \U$7703 ( \16823 , RIfc4b218_5877, \9212 );
and \U$7704 ( \16824 , RIdf1efa0_1729, \9214 );
and \U$7705 ( \16825 , RIfcc69e0_7282, \9216 );
and \U$7706 ( \16826 , RIdf18bc8_1658, \9218 );
and \U$7707 ( \16827 , RIdf16300_1629, \9220 );
and \U$7708 ( \16828 , RIdf13600_1597, \9222 );
and \U$7709 ( \16829 , RIdf10900_1565, \9224 );
and \U$7710 ( \16830 , RIdf0dc00_1533, \9226 );
and \U$7711 ( \16831 , RIdf0af00_1501, \9228 );
and \U$7712 ( \16832 , RIdf08200_1469, \9230 );
and \U$7713 ( \16833 , RIdf05500_1437, \9232 );
and \U$7714 ( \16834 , RIdf02800_1405, \9234 );
and \U$7715 ( \16835 , RIdefce00_1341, \9236 );
and \U$7716 ( \16836 , RIdefa100_1309, \9238 );
and \U$7717 ( \16837 , RIdef7400_1277, \9240 );
and \U$7718 ( \16838 , RIdef4700_1245, \9242 );
and \U$7719 ( \16839 , RIdef1a00_1213, \9244 );
and \U$7720 ( \16840 , RIdeeed00_1181, \9246 );
and \U$7721 ( \16841 , RIdeec000_1149, \9248 );
and \U$7722 ( \16842 , RIdee9300_1117, \9250 );
and \U$7723 ( \16843 , RIfce4ad0_7624, \9252 );
and \U$7724 ( \16844 , RIfc9e8a0_6826, \9254 );
and \U$7725 ( \16845 , RIfcc46b8_7257, \9256 );
and \U$7726 ( \16846 , RIfcd4108_7435, \9258 );
and \U$7727 ( \16847 , RIdee4440_1061, \9260 );
and \U$7728 ( \16848 , RIdee2280_1037, \9262 );
and \U$7729 ( \16849 , RIdee0390_1015, \9264 );
and \U$7730 ( \16850 , RIdede068_990, \9266 );
and \U$7731 ( \16851 , RIfcda0a8_7503, \9268 );
and \U$7732 ( \16852 , RIfce54a8_7631, \9270 );
and \U$7733 ( \16853 , RIfca0790_6848, \9272 );
and \U$7734 ( \16854 , RIfc50ee8_5943, \9274 );
and \U$7735 ( \16855 , RIded8d70_931, \9276 );
and \U$7736 ( \16856 , RIded68e0_905, \9278 );
and \U$7737 ( \16857 , RIded4888_882, \9280 );
and \U$7738 ( \16858 , RIded2560_857, \9282 );
and \U$7739 ( \16859 , RIdecfb30_827, \9284 );
and \U$7740 ( \16860 , RIdecce30_795, \9286 );
and \U$7741 ( \16861 , RIdeca130_763, \9288 );
and \U$7742 ( \16862 , RIdec7430_731, \9290 );
and \U$7743 ( \16863 , RIdeb3930_507, \9292 );
and \U$7744 ( \16864 , RIde94b98_315, \9294 );
and \U$7745 ( \16865 , RIe16d538_2621, \9296 );
and \U$7746 ( \16866 , RIe159330_2392, \9298 );
and \U$7747 ( \16867 , RIe142b30_2136, \9300 );
and \U$7748 ( \16868 , RIdf37528_2006, \9302 );
and \U$7749 ( \16869 , RIdf2bb88_1874, \9304 );
and \U$7750 ( \16870 , RIdf1c408_1698, \9306 );
and \U$7751 ( \16871 , RIdeffb00_1373, \9308 );
and \U$7752 ( \16872 , RIdee6600_1085, \9310 );
and \U$7753 ( \16873 , RIdedb368_958, \9312 );
and \U$7754 ( \16874 , RIde7aae0_188, \9314 );
or \U$7755 ( \16875 , \16811 , \16812 , \16813 , \16814 , \16815 , \16816 , \16817 , \16818 , \16819 , \16820 , \16821 , \16822 , \16823 , \16824 , \16825 , \16826 , \16827 , \16828 , \16829 , \16830 , \16831 , \16832 , \16833 , \16834 , \16835 , \16836 , \16837 , \16838 , \16839 , \16840 , \16841 , \16842 , \16843 , \16844 , \16845 , \16846 , \16847 , \16848 , \16849 , \16850 , \16851 , \16852 , \16853 , \16854 , \16855 , \16856 , \16857 , \16858 , \16859 , \16860 , \16861 , \16862 , \16863 , \16864 , \16865 , \16866 , \16867 , \16868 , \16869 , \16870 , \16871 , \16872 , \16873 , \16874 );
or \U$7756 ( \16876 , \16810 , \16875 );
_DC g2b8f ( \16877_nG2b8f , \16876 , \9323 );
buf \U$7757 ( \16878 , \16877_nG2b8f );
and \U$7758 ( \16879 , RIe19c9c8_3159, \9333 );
and \U$7759 ( \16880 , RIe199cc8_3127, \9335 );
and \U$7760 ( \16881 , RIfe8ea28_7967, \9337 );
and \U$7761 ( \16882 , RIe196fc8_3095, \9339 );
and \U$7762 ( \16883 , RIfec20d0_8328, \9341 );
and \U$7763 ( \16884 , RIe1942c8_3063, \9343 );
and \U$7764 ( \16885 , RIe1915c8_3031, \9345 );
and \U$7765 ( \16886 , RIe18e8c8_2999, \9347 );
and \U$7766 ( \16887 , RIe188ec8_2935, \9349 );
and \U$7767 ( \16888 , RIe1861c8_2903, \9351 );
and \U$7768 ( \16889 , RIfc68228_6207, \9353 );
and \U$7769 ( \16890 , RIe1834c8_2871, \9355 );
and \U$7770 ( \16891 , RIfccb5d0_7336, \9357 );
and \U$7771 ( \16892 , RIe1807c8_2839, \9359 );
and \U$7772 ( \16893 , RIe17dac8_2807, \9361 );
and \U$7773 ( \16894 , RIe17adc8_2775, \9363 );
and \U$7774 ( \16895 , RIf141e18_5209, \9365 );
and \U$7775 ( \16896 , RIf140900_5194, \9367 );
and \U$7776 ( \16897 , RIf140090_5188, \9369 );
and \U$7777 ( \16898 , RIe1753c8_2711, \9371 );
and \U$7778 ( \16899 , RIf13f988_5183, \9373 );
and \U$7779 ( \16900 , RIf13ece0_5174, \9375 );
and \U$7780 ( \16901 , RIee3e170_5165, \9377 );
and \U$7781 ( \16902 , RIee3cf28_5152, \9379 );
and \U$7782 ( \16903 , RIee3bce0_5139, \9381 );
and \U$7783 ( \16904 , RIee3ac00_5127, \9383 );
and \U$7784 ( \16905 , RIee39850_5113, \9385 );
and \U$7785 ( \16906 , RIe172dd0_2684, \9387 );
and \U$7786 ( \16907 , RIf16fc28_5731, \9389 );
and \U$7787 ( \16908 , RIf16f0e8_5723, \9391 );
and \U$7788 ( \16909 , RIf16dd38_5709, \9393 );
and \U$7789 ( \16910 , RIfce9120_7674, \9395 );
and \U$7790 ( \16911 , RIfc404a8_5757, \9397 );
and \U$7791 ( \16912 , RIe222d20_4686, \9399 );
and \U$7792 ( \16913 , RIf16b8a8_5683, \9401 );
and \U$7793 ( \16914 , RIe220020_4654, \9403 );
and \U$7794 ( \16915 , RIf16a930_5672, \9405 );
and \U$7795 ( \16916 , RIe21d320_4622, \9407 );
and \U$7796 ( \16917 , RIe217920_4558, \9409 );
and \U$7797 ( \16918 , RIe214c20_4526, \9411 );
and \U$7798 ( \16919 , RIfc5b910_6064, \9413 );
and \U$7799 ( \16920 , RIe211f20_4494, \9415 );
and \U$7800 ( \16921 , RIfe8e8c0_7966, \9417 );
and \U$7801 ( \16922 , RIe20f220_4462, \9419 );
and \U$7802 ( \16923 , RIfe8e758_7965, \9421 );
and \U$7803 ( \16924 , RIe20c520_4430, \9423 );
and \U$7804 ( \16925 , RIe209820_4398, \9425 );
and \U$7805 ( \16926 , RIe206b20_4366, \9427 );
and \U$7806 ( \16927 , RIf166b50_5628, \9429 );
and \U$7807 ( \16928 , RIf165a70_5616, \9431 );
and \U$7808 ( \16929 , RIfe8dd80_7958, \9433 );
and \U$7809 ( \16930 , RIfe8dab0_7956, \9435 );
and \U$7810 ( \16931 , RIf164c60_5606, \9437 );
and \U$7811 ( \16932 , RIf163e50_5596, \9439 );
and \U$7812 ( \16933 , RIf162ed8_5585, \9441 );
and \U$7813 ( \16934 , RIf1616f0_5568, \9443 );
and \U$7814 ( \16935 , RIf15f800_5546, \9445 );
and \U$7815 ( \16936 , RIf15da78_5525, \9447 );
and \U$7816 ( \16937 , RIfe8d948_7955, \9449 );
and \U$7817 ( \16938 , RIfe8dc18_7957, \9451 );
and \U$7818 ( \16939 , RIf15c560_5510, \9453 );
and \U$7819 ( \16940 , RIf15b048_5495, \9455 );
and \U$7820 ( \16941 , RIfc62828_6143, \9457 );
and \U$7821 ( \16942 , RIf159860_5478, \9459 );
or \U$7822 ( \16943 , \16879 , \16880 , \16881 , \16882 , \16883 , \16884 , \16885 , \16886 , \16887 , \16888 , \16889 , \16890 , \16891 , \16892 , \16893 , \16894 , \16895 , \16896 , \16897 , \16898 , \16899 , \16900 , \16901 , \16902 , \16903 , \16904 , \16905 , \16906 , \16907 , \16908 , \16909 , \16910 , \16911 , \16912 , \16913 , \16914 , \16915 , \16916 , \16917 , \16918 , \16919 , \16920 , \16921 , \16922 , \16923 , \16924 , \16925 , \16926 , \16927 , \16928 , \16929 , \16930 , \16931 , \16932 , \16933 , \16934 , \16935 , \16936 , \16937 , \16938 , \16939 , \16940 , \16941 , \16942 );
and \U$7823 ( \16944 , RIf158780_5466, \9462 );
and \U$7824 ( \16945 , RIf157538_5453, \9464 );
and \U$7825 ( \16946 , RIfca6e38_6921, \9466 );
and \U$7826 ( \16947 , RIe1f9b00_4218, \9468 );
and \U$7827 ( \16948 , RIfc61e50_6136, \9470 );
and \U$7828 ( \16949 , RIfc61748_6131, \9472 );
and \U$7829 ( \16950 , RIf154130_5416, \9474 );
and \U$7830 ( \16951 , RIe1f4ad8_4161, \9476 );
and \U$7831 ( \16952 , RIf152ab0_5400, \9478 );
and \U$7832 ( \16953 , RIf151700_5386, \9480 );
and \U$7833 ( \16954 , RIf1501e8_5371, \9482 );
and \U$7834 ( \16955 , RIe1f27b0_4136, \9484 );
and \U$7835 ( \16956 , RIfc60ed8_6125, \9486 );
and \U$7836 ( \16957 , RIfc7b620_6426, \9488 );
and \U$7837 ( \16958 , RIf14d7b8_5341, \9490 );
and \U$7838 ( \16959 , RIe1ed4b8_4077, \9492 );
and \U$7839 ( \16960 , RIe1eaa88_4047, \9494 );
and \U$7840 ( \16961 , RIe1e7d88_4015, \9496 );
and \U$7841 ( \16962 , RIe1e5088_3983, \9498 );
and \U$7842 ( \16963 , RIe1e2388_3951, \9500 );
and \U$7843 ( \16964 , RIe1df688_3919, \9502 );
and \U$7844 ( \16965 , RIe1dc988_3887, \9504 );
and \U$7845 ( \16966 , RIe1d9c88_3855, \9506 );
and \U$7846 ( \16967 , RIe1d6f88_3823, \9508 );
and \U$7847 ( \16968 , RIe1d1588_3759, \9510 );
and \U$7848 ( \16969 , RIe1ce888_3727, \9512 );
and \U$7849 ( \16970 , RIe1cbb88_3695, \9514 );
and \U$7850 ( \16971 , RIe1c8e88_3663, \9516 );
and \U$7851 ( \16972 , RIe1c6188_3631, \9518 );
and \U$7852 ( \16973 , RIe1c3488_3599, \9520 );
and \U$7853 ( \16974 , RIe1c0788_3567, \9522 );
and \U$7854 ( \16975 , RIe1bda88_3535, \9524 );
and \U$7855 ( \16976 , RIfca4de0_6898, \9526 );
and \U$7856 ( \16977 , RIfc5ea48_6099, \9528 );
and \U$7857 ( \16978 , RIe1b8a60_3478, \9530 );
and \U$7858 ( \16979 , RIe1b6a08_3455, \9532 );
and \U$7859 ( \16980 , RIfcbd638_7177, \9534 );
and \U$7860 ( \16981 , RIfc44fa8_5807, \9536 );
and \U$7861 ( \16982 , RIfe8e5f0_7964, \9538 );
and \U$7862 ( \16983 , RIfe8e1b8_7961, \9540 );
and \U$7863 ( \16984 , RIf1488f8_5285, \9542 );
and \U$7864 ( \16985 , RIf147818_5273, \9544 );
and \U$7865 ( \16986 , RIfe8e050_7960, \9546 );
and \U$7866 ( \16987 , RIfe8e488_7963, \9548 );
and \U$7867 ( \16988 , RIf146e40_5266, \9550 );
and \U$7868 ( \16989 , RIf146030_5256, \9552 );
and \U$7869 ( \16990 , RIfe8dee8_7959, \9554 );
and \U$7870 ( \16991 , RIfe8e320_7962, \9556 );
and \U$7871 ( \16992 , RIe1a7dc8_3287, \9558 );
and \U$7872 ( \16993 , RIe1a50c8_3255, \9560 );
and \U$7873 ( \16994 , RIe1a23c8_3223, \9562 );
and \U$7874 ( \16995 , RIe19f6c8_3191, \9564 );
and \U$7875 ( \16996 , RIe18bbc8_2967, \9566 );
and \U$7876 ( \16997 , RIe1780c8_2743, \9568 );
and \U$7877 ( \16998 , RIe225a20_4718, \9570 );
and \U$7878 ( \16999 , RIe21a620_4590, \9572 );
and \U$7879 ( \17000 , RIe203e20_4334, \9574 );
and \U$7880 ( \17001 , RIe1fde80_4266, \9576 );
and \U$7881 ( \17002 , RIe1f7238_4189, \9578 );
and \U$7882 ( \17003 , RIe1efd80_4106, \9580 );
and \U$7883 ( \17004 , RIe1d4288_3791, \9582 );
and \U$7884 ( \17005 , RIe1bad88_3503, \9584 );
and \U$7885 ( \17006 , RIe1adc00_3354, \9586 );
and \U$7886 ( \17007 , RIe170238_2653, \9588 );
or \U$7887 ( \17008 , \16944 , \16945 , \16946 , \16947 , \16948 , \16949 , \16950 , \16951 , \16952 , \16953 , \16954 , \16955 , \16956 , \16957 , \16958 , \16959 , \16960 , \16961 , \16962 , \16963 , \16964 , \16965 , \16966 , \16967 , \16968 , \16969 , \16970 , \16971 , \16972 , \16973 , \16974 , \16975 , \16976 , \16977 , \16978 , \16979 , \16980 , \16981 , \16982 , \16983 , \16984 , \16985 , \16986 , \16987 , \16988 , \16989 , \16990 , \16991 , \16992 , \16993 , \16994 , \16995 , \16996 , \16997 , \16998 , \16999 , \17000 , \17001 , \17002 , \17003 , \17004 , \17005 , \17006 , \17007 );
or \U$7888 ( \17009 , \16943 , \17008 );
_DC g3cbc ( \17010_nG3cbc , \17009 , \9597 );
buf \U$7889 ( \17011 , \17010_nG3cbc );
xor \U$7890 ( \17012 , \16878 , \17011 );
and \U$7891 ( \17013 , RIdec45c8_698, \9059 );
and \U$7892 ( \17014 , RIdec18c8_666, \9061 );
and \U$7893 ( \17015 , RIfce85e0_7666, \9063 );
and \U$7894 ( \17016 , RIdebebc8_634, \9065 );
and \U$7895 ( \17017 , RIfcb8bb0_7124, \9067 );
and \U$7896 ( \17018 , RIdebbec8_602, \9069 );
and \U$7897 ( \17019 , RIdeb91c8_570, \9071 );
and \U$7898 ( \17020 , RIdeb64c8_538, \9073 );
and \U$7899 ( \17021 , RIfc85d78_6545, \9075 );
and \U$7900 ( \17022 , RIdeb0ac8_474, \9077 );
and \U$7901 ( \17023 , RIfc85aa8_6543, \9079 );
and \U$7902 ( \17024 , RIdeaddc8_442, \9081 );
and \U$7903 ( \17025 , RIfc4d3d8_5901, \9083 );
and \U$7904 ( \17026 , RIdea8350_410, \9085 );
and \U$7905 ( \17027 , RIdea1a50_378, \9087 );
and \U$7906 ( \17028 , RIde9b150_346, \9089 );
and \U$7907 ( \17029 , RIfc85ee0_6546, \9091 );
and \U$7908 ( \17030 , RIfc9c9b0_6804, \9093 );
and \U$7909 ( \17031 , RIfce13f8_7585, \9095 );
and \U$7910 ( \17032 , RIfcb8778_7121, \9097 );
and \U$7911 ( \17033 , RIfe8d510_7952, \9099 );
and \U$7912 ( \17034 , RIfe8d3a8_7951, \9101 );
and \U$7913 ( \17035 , RIde886b8_255, \9103 );
and \U$7914 ( \17036 , RIde841d0_234, \9105 );
and \U$7915 ( \17037 , RIde806c0_216, \9107 );
and \U$7916 ( \17038 , RIfcb8070_7116, \9109 );
and \U$7917 ( \17039 , RIfce1128_7583, \9111 );
and \U$7918 ( \17040 , RIfc9c140_6798, \9113 );
and \U$7919 ( \17041 , RIee38d10_5105, \9115 );
and \U$7920 ( \17042 , RIe16ac70_2592, \9117 );
and \U$7921 ( \17043 , RIfc850d0_6536, \9119 );
and \U$7922 ( \17044 , RIe167160_2550, \9121 );
and \U$7923 ( \17045 , RIe1645c8_2519, \9123 );
and \U$7924 ( \17046 , RIe1618c8_2487, \9125 );
and \U$7925 ( \17047 , RIee36b50_5081, \9127 );
and \U$7926 ( \17048 , RIe15ebc8_2455, \9129 );
and \U$7927 ( \17049 , RIee35d40_5071, \9131 );
and \U$7928 ( \17050 , RIe15bec8_2423, \9133 );
and \U$7929 ( \17051 , RIe1564c8_2359, \9135 );
and \U$7930 ( \17052 , RIe1537c8_2327, \9137 );
and \U$7931 ( \17053 , RIfc3ef90_5742, \9139 );
and \U$7932 ( \17054 , RIe150ac8_2295, \9141 );
and \U$7933 ( \17055 , RIfe8d7e0_7954, \9143 );
and \U$7934 ( \17056 , RIe14ddc8_2263, \9145 );
and \U$7935 ( \17057 , RIfce0fc0_7582, \9147 );
and \U$7936 ( \17058 , RIe14b0c8_2231, \9149 );
and \U$7937 ( \17059 , RIe1483c8_2199, \9151 );
and \U$7938 ( \17060 , RIe1456c8_2167, \9153 );
and \U$7939 ( \17061 , RIee33e50_5049, \9155 );
and \U$7940 ( \17062 , RIee32c08_5036, \9157 );
and \U$7941 ( \17063 , RIee319c0_5023, \9159 );
and \U$7942 ( \17064 , RIee30d18_5014, \9161 );
and \U$7943 ( \17065 , RIfe8cf70_7948, \9163 );
and \U$7944 ( \17066 , RIfe8ce08_7947, \9165 );
and \U$7945 ( \17067 , RIfe8d240_7950, \9167 );
and \U$7946 ( \17068 , RIfe8d0d8_7949, \9169 );
and \U$7947 ( \17069 , RIfce9dc8_7683, \9171 );
and \U$7948 ( \17070 , RIee2ef90_4993, \9173 );
and \U$7949 ( \17071 , RIfce51d8_7629, \9175 );
and \U$7950 ( \17072 , RIee2cdd0_4969, \9177 );
and \U$7951 ( \17073 , RIdf34af8_1976, \9179 );
and \U$7952 ( \17074 , RIfe8d678_7953, \9181 );
and \U$7953 ( \17075 , RIdf30610_1927, \9183 );
and \U$7954 ( \17076 , RIdf2e720_1905, \9185 );
or \U$7955 ( \17077 , \17013 , \17014 , \17015 , \17016 , \17017 , \17018 , \17019 , \17020 , \17021 , \17022 , \17023 , \17024 , \17025 , \17026 , \17027 , \17028 , \17029 , \17030 , \17031 , \17032 , \17033 , \17034 , \17035 , \17036 , \17037 , \17038 , \17039 , \17040 , \17041 , \17042 , \17043 , \17044 , \17045 , \17046 , \17047 , \17048 , \17049 , \17050 , \17051 , \17052 , \17053 , \17054 , \17055 , \17056 , \17057 , \17058 , \17059 , \17060 , \17061 , \17062 , \17063 , \17064 , \17065 , \17066 , \17067 , \17068 , \17069 , \17070 , \17071 , \17072 , \17073 , \17074 , \17075 , \17076 );
and \U$7956 ( \17078 , RIee2b318_4950, \9188 );
and \U$7957 ( \17079 , RIee29c98_4934, \9190 );
and \U$7958 ( \17080 , RIee28780_4919, \9192 );
and \U$7959 ( \17081 , RIee27538_4906, \9194 );
and \U$7960 ( \17082 , RIdf299c8_1850, \9196 );
and \U$7961 ( \17083 , RIdf276a0_1825, \9198 );
and \U$7962 ( \17084 , RIdf25918_1804, \9200 );
and \U$7963 ( \17085 , RIdf23cf8_1784, \9202 );
and \U$7964 ( \17086 , RIfc83ff0_6524, \9204 );
and \U$7965 ( \17087 , RIfcb73c8_7107, \9206 );
and \U$7966 ( \17088 , RIfc51320_5946, \9208 );
and \U$7967 ( \17089 , RIfcdaa80_7510, \9210 );
and \U$7968 ( \17090 , RIfc83d20_6522, \9212 );
and \U$7969 ( \17091 , RIdf1ee38_1728, \9214 );
and \U$7970 ( \17092 , RIfc51b90_5952, \9216 );
and \U$7971 ( \17093 , RIdf18a60_1657, \9218 );
and \U$7972 ( \17094 , RIdf16198_1628, \9220 );
and \U$7973 ( \17095 , RIdf13498_1596, \9222 );
and \U$7974 ( \17096 , RIdf10798_1564, \9224 );
and \U$7975 ( \17097 , RIdf0da98_1532, \9226 );
and \U$7976 ( \17098 , RIdf0ad98_1500, \9228 );
and \U$7977 ( \17099 , RIdf08098_1468, \9230 );
and \U$7978 ( \17100 , RIdf05398_1436, \9232 );
and \U$7979 ( \17101 , RIdf02698_1404, \9234 );
and \U$7980 ( \17102 , RIdefcc98_1340, \9236 );
and \U$7981 ( \17103 , RIdef9f98_1308, \9238 );
and \U$7982 ( \17104 , RIdef7298_1276, \9240 );
and \U$7983 ( \17105 , RIdef4598_1244, \9242 );
and \U$7984 ( \17106 , RIdef1898_1212, \9244 );
and \U$7985 ( \17107 , RIdeeeb98_1180, \9246 );
and \U$7986 ( \17108 , RIdeebe98_1148, \9248 );
and \U$7987 ( \17109 , RIdee9198_1116, \9250 );
and \U$7988 ( \17110 , RIee25210_4881, \9252 );
and \U$7989 ( \17111 , RIee24400_4871, \9254 );
and \U$7990 ( \17112 , RIee238c0_4863, \9256 );
and \U$7991 ( \17113 , RIee22ee8_4856, \9258 );
and \U$7992 ( \17114 , RIfe8cca0_7946, \9260 );
and \U$7993 ( \17115 , RIdee2118_1036, \9262 );
and \U$7994 ( \17116 , RIfe8cb38_7945, \9264 );
and \U$7995 ( \17117 , RIdeddf00_989, \9266 );
and \U$7996 ( \17118 , RIfcc5a68_7271, \9268 );
and \U$7997 ( \17119 , RIee21f70_4845, \9270 );
and \U$7998 ( \17120 , RIfcb6cc0_7102, \9272 );
and \U$7999 ( \17121 , RIee20e90_4833, \9274 );
and \U$8000 ( \17122 , RIded8c08_930, \9276 );
and \U$8001 ( \17123 , RIded6778_904, \9278 );
and \U$8002 ( \17124 , RIded4720_881, \9280 );
and \U$8003 ( \17125 , RIded23f8_856, \9282 );
and \U$8004 ( \17126 , RIdecf9c8_826, \9284 );
and \U$8005 ( \17127 , RIdecccc8_794, \9286 );
and \U$8006 ( \17128 , RIdec9fc8_762, \9288 );
and \U$8007 ( \17129 , RIdec72c8_730, \9290 );
and \U$8008 ( \17130 , RIdeb37c8_506, \9292 );
and \U$8009 ( \17131 , RIde94850_314, \9294 );
and \U$8010 ( \17132 , RIe16d3d0_2620, \9296 );
and \U$8011 ( \17133 , RIe1591c8_2391, \9298 );
and \U$8012 ( \17134 , RIe1429c8_2135, \9300 );
and \U$8013 ( \17135 , RIdf373c0_2005, \9302 );
and \U$8014 ( \17136 , RIdf2ba20_1873, \9304 );
and \U$8015 ( \17137 , RIdf1c2a0_1697, \9306 );
and \U$8016 ( \17138 , RIdeff998_1372, \9308 );
and \U$8017 ( \17139 , RIdee6498_1084, \9310 );
and \U$8018 ( \17140 , RIdedb200_957, \9312 );
and \U$8019 ( \17141 , RIde7a798_187, \9314 );
or \U$8020 ( \17142 , \17078 , \17079 , \17080 , \17081 , \17082 , \17083 , \17084 , \17085 , \17086 , \17087 , \17088 , \17089 , \17090 , \17091 , \17092 , \17093 , \17094 , \17095 , \17096 , \17097 , \17098 , \17099 , \17100 , \17101 , \17102 , \17103 , \17104 , \17105 , \17106 , \17107 , \17108 , \17109 , \17110 , \17111 , \17112 , \17113 , \17114 , \17115 , \17116 , \17117 , \17118 , \17119 , \17120 , \17121 , \17122 , \17123 , \17124 , \17125 , \17126 , \17127 , \17128 , \17129 , \17130 , \17131 , \17132 , \17133 , \17134 , \17135 , \17136 , \17137 , \17138 , \17139 , \17140 , \17141 );
or \U$8021 ( \17143 , \17077 , \17142 );
_DC g2c14 ( \17144_nG2c14 , \17143 , \9323 );
buf \U$8022 ( \17145 , \17144_nG2c14 );
and \U$8023 ( \17146 , RIe19c860_3158, \9333 );
and \U$8024 ( \17147 , RIe199b60_3126, \9335 );
and \U$8025 ( \17148 , RIf145220_5246, \9337 );
and \U$8026 ( \17149 , RIe196e60_3094, \9339 );
and \U$8027 ( \17150 , RIf144140_5234, \9341 );
and \U$8028 ( \17151 , RIe194160_3062, \9343 );
and \U$8029 ( \17152 , RIe191460_3030, \9345 );
and \U$8030 ( \17153 , RIe18e760_2998, \9347 );
and \U$8031 ( \17154 , RIe188d60_2934, \9349 );
and \U$8032 ( \17155 , RIe186060_2902, \9351 );
and \U$8033 ( \17156 , RIf1431c8_5223, \9353 );
and \U$8034 ( \17157 , RIe183360_2870, \9355 );
and \U$8035 ( \17158 , RIf142ac0_5218, \9357 );
and \U$8036 ( \17159 , RIe180660_2838, \9359 );
and \U$8037 ( \17160 , RIe17d960_2806, \9361 );
and \U$8038 ( \17161 , RIe17ac60_2774, \9363 );
and \U$8039 ( \17162 , RIf141cb0_5208, \9365 );
and \U$8040 ( \17163 , RIf140798_5193, \9367 );
and \U$8041 ( \17164 , RIf13ff28_5187, \9369 );
and \U$8042 ( \17165 , RIfe8be90_7936, \9371 );
and \U$8043 ( \17166 , RIfceb880_7702, \9373 );
and \U$8044 ( \17167 , RIf13eb78_5173, \9375 );
and \U$8045 ( \17168 , RIee3e008_5164, \9377 );
and \U$8046 ( \17169 , RIee3cdc0_5151, \9379 );
and \U$8047 ( \17170 , RIee3bb78_5138, \9381 );
and \U$8048 ( \17171 , RIee3aa98_5126, \9383 );
and \U$8049 ( \17172 , RIee396e8_5112, \9385 );
and \U$8050 ( \17173 , RIe172c68_2683, \9387 );
and \U$8051 ( \17174 , RIf16fac0_5730, \9389 );
and \U$8052 ( \17175 , RIf16ef80_5722, \9391 );
and \U$8053 ( \17176 , RIf16dbd0_5708, \9393 );
and \U$8054 ( \17177 , RIfcc4af0_7260, \9395 );
and \U$8055 ( \17178 , RIf16c820_5694, \9397 );
and \U$8056 ( \17179 , RIe222bb8_4685, \9399 );
and \U$8057 ( \17180 , RIf16b740_5682, \9401 );
and \U$8058 ( \17181 , RIe21feb8_4653, \9403 );
and \U$8059 ( \17182 , RIf16a7c8_5671, \9405 );
and \U$8060 ( \17183 , RIe21d1b8_4621, \9407 );
and \U$8061 ( \17184 , RIe2177b8_4557, \9409 );
and \U$8062 ( \17185 , RIe214ab8_4525, \9411 );
and \U$8063 ( \17186 , RIfe8c430_7940, \9413 );
and \U$8064 ( \17187 , RIe211db8_4493, \9415 );
and \U$8065 ( \17188 , RIf1688d8_5649, \9417 );
and \U$8066 ( \17189 , RIe20f0b8_4461, \9419 );
and \U$8067 ( \17190 , RIf167960_5638, \9421 );
and \U$8068 ( \17191 , RIe20c3b8_4429, \9423 );
and \U$8069 ( \17192 , RIe2096b8_4397, \9425 );
and \U$8070 ( \17193 , RIe2069b8_4365, \9427 );
and \U$8071 ( \17194 , RIf1669e8_5627, \9429 );
and \U$8072 ( \17195 , RIf165908_5615, \9431 );
and \U$8073 ( \17196 , RIfe8c9d0_7944, \9433 );
and \U$8074 ( \17197 , RIfe8c700_7942, \9435 );
and \U$8075 ( \17198 , RIfc9c578_6801, \9437 );
and \U$8076 ( \17199 , RIf163ce8_5595, \9439 );
and \U$8077 ( \17200 , RIf162d70_5584, \9441 );
and \U$8078 ( \17201 , RIf161588_5567, \9443 );
and \U$8079 ( \17202 , RIf15f698_5545, \9445 );
and \U$8080 ( \17203 , RIf15d910_5524, \9447 );
and \U$8081 ( \17204 , RIfe8c598_7941, \9449 );
and \U$8082 ( \17205 , RIfe8c868_7943, \9451 );
and \U$8083 ( \17206 , RIf15c3f8_5509, \9453 );
and \U$8084 ( \17207 , RIf15aee0_5494, \9455 );
and \U$8085 ( \17208 , RIf15a0d0_5484, \9457 );
and \U$8086 ( \17209 , RIf1596f8_5477, \9459 );
or \U$8087 ( \17210 , \17146 , \17147 , \17148 , \17149 , \17150 , \17151 , \17152 , \17153 , \17154 , \17155 , \17156 , \17157 , \17158 , \17159 , \17160 , \17161 , \17162 , \17163 , \17164 , \17165 , \17166 , \17167 , \17168 , \17169 , \17170 , \17171 , \17172 , \17173 , \17174 , \17175 , \17176 , \17177 , \17178 , \17179 , \17180 , \17181 , \17182 , \17183 , \17184 , \17185 , \17186 , \17187 , \17188 , \17189 , \17190 , \17191 , \17192 , \17193 , \17194 , \17195 , \17196 , \17197 , \17198 , \17199 , \17200 , \17201 , \17202 , \17203 , \17204 , \17205 , \17206 , \17207 , \17208 , \17209 );
and \U$8088 ( \17211 , RIf158618_5465, \9462 );
and \U$8089 ( \17212 , RIf1573d0_5452, \9464 );
and \U$8090 ( \17213 , RIf156b60_5446, \9466 );
and \U$8091 ( \17214 , RIfec1f68_8327, \9468 );
and \U$8092 ( \17215 , RIf155eb8_5437, \9470 );
and \U$8093 ( \17216 , RIf155378_5429, \9472 );
and \U$8094 ( \17217 , RIf153fc8_5415, \9474 );
and \U$8095 ( \17218 , RIfe8bff8_7937, \9476 );
and \U$8096 ( \17219 , RIf152948_5399, \9478 );
and \U$8097 ( \17220 , RIf151598_5385, \9480 );
and \U$8098 ( \17221 , RIf150080_5370, \9482 );
and \U$8099 ( \17222 , RIfe8c2c8_7939, \9484 );
and \U$8100 ( \17223 , RIf14f270_5360, \9486 );
and \U$8101 ( \17224 , RIfc503a8_5935, \9488 );
and \U$8102 ( \17225 , RIf14d650_5340, \9490 );
and \U$8103 ( \17226 , RIfe8c160_7938, \9492 );
and \U$8104 ( \17227 , RIe1ea920_4046, \9494 );
and \U$8105 ( \17228 , RIe1e7c20_4014, \9496 );
and \U$8106 ( \17229 , RIe1e4f20_3982, \9498 );
and \U$8107 ( \17230 , RIe1e2220_3950, \9500 );
and \U$8108 ( \17231 , RIe1df520_3918, \9502 );
and \U$8109 ( \17232 , RIe1dc820_3886, \9504 );
and \U$8110 ( \17233 , RIe1d9b20_3854, \9506 );
and \U$8111 ( \17234 , RIe1d6e20_3822, \9508 );
and \U$8112 ( \17235 , RIe1d1420_3758, \9510 );
and \U$8113 ( \17236 , RIe1ce720_3726, \9512 );
and \U$8114 ( \17237 , RIe1cba20_3694, \9514 );
and \U$8115 ( \17238 , RIe1c8d20_3662, \9516 );
and \U$8116 ( \17239 , RIe1c6020_3630, \9518 );
and \U$8117 ( \17240 , RIe1c3320_3598, \9520 );
and \U$8118 ( \17241 , RIe1c0620_3566, \9522 );
and \U$8119 ( \17242 , RIe1bd920_3534, \9524 );
and \U$8120 ( \17243 , RIf14c2a0_5326, \9526 );
and \U$8121 ( \17244 , RIf14aef0_5312, \9528 );
and \U$8122 ( \17245 , RIe1b88f8_3477, \9530 );
and \U$8123 ( \17246 , RIe1b68a0_3454, \9532 );
and \U$8124 ( \17247 , RIfcd4db0_7444, \9534 );
and \U$8125 ( \17248 , RIfc4ebc0_5918, \9536 );
and \U$8126 ( \17249 , RIfec1e00_8326, \9538 );
and \U$8127 ( \17250 , RIfe8bd28_7935, \9540 );
and \U$8128 ( \17251 , RIf148790_5284, \9542 );
and \U$8129 ( \17252 , RIf1476b0_5272, \9544 );
and \U$8130 ( \17253 , RIfe8ba58_7933, \9546 );
and \U$8131 ( \17254 , RIfec1b30_8324, \9548 );
and \U$8132 ( \17255 , RIfc4e788_5915, \9550 );
and \U$8133 ( \17256 , RIfcb8e80_7126, \9552 );
and \U$8134 ( \17257 , RIfe8bbc0_7934, \9554 );
and \U$8135 ( \17258 , RIfec1c98_8325, \9556 );
and \U$8136 ( \17259 , RIe1a7c60_3286, \9558 );
and \U$8137 ( \17260 , RIe1a4f60_3254, \9560 );
and \U$8138 ( \17261 , RIe1a2260_3222, \9562 );
and \U$8139 ( \17262 , RIe19f560_3190, \9564 );
and \U$8140 ( \17263 , RIe18ba60_2966, \9566 );
and \U$8141 ( \17264 , RIe177f60_2742, \9568 );
and \U$8142 ( \17265 , RIe2258b8_4717, \9570 );
and \U$8143 ( \17266 , RIe21a4b8_4589, \9572 );
and \U$8144 ( \17267 , RIe203cb8_4333, \9574 );
and \U$8145 ( \17268 , RIe1fdd18_4265, \9576 );
and \U$8146 ( \17269 , RIe1f70d0_4188, \9578 );
and \U$8147 ( \17270 , RIe1efc18_4105, \9580 );
and \U$8148 ( \17271 , RIe1d4120_3790, \9582 );
and \U$8149 ( \17272 , RIe1bac20_3502, \9584 );
and \U$8150 ( \17273 , RIe1ada98_3353, \9586 );
and \U$8151 ( \17274 , RIe1700d0_2652, \9588 );
or \U$8152 ( \17275 , \17211 , \17212 , \17213 , \17214 , \17215 , \17216 , \17217 , \17218 , \17219 , \17220 , \17221 , \17222 , \17223 , \17224 , \17225 , \17226 , \17227 , \17228 , \17229 , \17230 , \17231 , \17232 , \17233 , \17234 , \17235 , \17236 , \17237 , \17238 , \17239 , \17240 , \17241 , \17242 , \17243 , \17244 , \17245 , \17246 , \17247 , \17248 , \17249 , \17250 , \17251 , \17252 , \17253 , \17254 , \17255 , \17256 , \17257 , \17258 , \17259 , \17260 , \17261 , \17262 , \17263 , \17264 , \17265 , \17266 , \17267 , \17268 , \17269 , \17270 , \17271 , \17272 , \17273 , \17274 );
or \U$8153 ( \17276 , \17210 , \17275 );
_DC g3d41 ( \17277_nG3d41 , \17276 , \9597 );
buf \U$8154 ( \17278 , \17277_nG3d41 );
and \U$8155 ( \17279 , \17145 , \17278 );
and \U$8156 ( \17280 , \15521 , \15654 );
and \U$8157 ( \17281 , \15654 , \15929 );
and \U$8158 ( \17282 , \15521 , \15929 );
or \U$8159 ( \17283 , \17280 , \17281 , \17282 );
and \U$8160 ( \17284 , \17278 , \17283 );
and \U$8161 ( \17285 , \17145 , \17283 );
or \U$8162 ( \17286 , \17279 , \17284 , \17285 );
xor \U$8163 ( \17287 , \17012 , \17286 );
buf g4430 ( \17288_nG4430 , \17287 );
xor \U$8164 ( \17289 , \17145 , \17278 );
xor \U$8165 ( \17290 , \17289 , \17283 );
buf g4433 ( \17291_nG4433 , \17290 );
nand \U$8166 ( \17292 , \17291_nG4433 , \15931_nG4436 );
and \U$8167 ( \17293 , \17288_nG4430 , \17292 );
xor \U$8168 ( \17294 , \17291_nG4433 , \15931_nG4436 );
not \U$8169 ( \17295 , \17294 );
xor \U$8170 ( \17296 , \17288_nG4430 , \17291_nG4433 );
and \U$8171 ( \17297 , \17295 , \17296 );
and \U$8173 ( \17298 , \17294 , \10694_nG9c0e );
or \U$8174 ( \17299 , 1'b0 , \17298 );
xor \U$8175 ( \17300 , \17293 , \17299 );
xor \U$8176 ( \17301 , \17293 , \17300 );
buf \U$8177 ( \17302 , \17301 );
buf \U$8178 ( \17303 , \17302 );
and \U$8179 ( \17304 , \16745 , \17303 );
and \U$8180 ( \17305 , \16719 , \16721 );
and \U$8181 ( \17306 , \16719 , \16728 );
and \U$8182 ( \17307 , \16721 , \16728 );
or \U$8183 ( \17308 , \17305 , \17306 , \17307 );
buf \U$8184 ( \17309 , \17308 );
and \U$8185 ( \17310 , \15940 , \10995_nG9c0b );
and \U$8186 ( \17311 , \15937 , \11283_nG9c08 );
or \U$8187 ( \17312 , \17310 , \17311 );
xor \U$8188 ( \17313 , \15936 , \17312 );
buf \U$8189 ( \17314 , \17313 );
buf \U$8191 ( \17315 , \17314 );
and \U$8192 ( \17316 , \14631 , \11598_nG9c05 );
and \U$8193 ( \17317 , \14628 , \12470_nG9c02 );
or \U$8194 ( \17318 , \17316 , \17317 );
xor \U$8195 ( \17319 , \14627 , \17318 );
buf \U$8196 ( \17320 , \17319 );
buf \U$8198 ( \17321 , \17320 );
xor \U$8199 ( \17322 , \17315 , \17321 );
buf \U$8200 ( \17323 , \17322 );
and \U$8201 ( \17324 , \16696 , \16702 );
buf \U$8202 ( \17325 , \17324 );
xor \U$8203 ( \17326 , \17323 , \17325 );
and \U$8204 ( \17327 , \13370 , \12801_nG9bff );
and \U$8205 ( \17328 , \13367 , \13705_nG9bfc );
or \U$8206 ( \17329 , \17327 , \17328 );
xor \U$8207 ( \17330 , \13366 , \17329 );
buf \U$8208 ( \17331 , \17330 );
buf \U$8210 ( \17332 , \17331 );
xor \U$8211 ( \17333 , \17326 , \17332 );
buf \U$8212 ( \17334 , \17333 );
xor \U$8213 ( \17335 , \17309 , \17334 );
and \U$8214 ( \17336 , \10707 , \16680_nG9bed );
and \U$8215 ( \17337 , \16351 , \16640 );
and \U$8216 ( \17338 , \16640 , \16669 );
and \U$8217 ( \17339 , \16351 , \16669 );
or \U$8218 ( \17340 , \17337 , \17338 , \17339 );
and \U$8219 ( \17341 , \16645 , \16649 );
and \U$8220 ( \17342 , \16649 , \16668 );
and \U$8221 ( \17343 , \16645 , \16668 );
or \U$8222 ( \17344 , \17341 , \17342 , \17343 );
and \U$8223 ( \17345 , \16658 , \16662 );
and \U$8224 ( \17346 , \16662 , \16667 );
and \U$8225 ( \17347 , \16658 , \16667 );
or \U$8226 ( \17348 , \17345 , \17346 , \17347 );
and \U$8227 ( \17349 , \16355 , \16626 );
xor \U$8228 ( \17350 , \17348 , \17349 );
and \U$8229 ( \17351 , \14024 , \12790 );
and \U$8230 ( \17352 , \14950 , \12461 );
nor \U$8231 ( \17353 , \17351 , \17352 );
xnor \U$8232 ( \17354 , \17353 , \12780 );
xor \U$8233 ( \17355 , \17350 , \17354 );
xor \U$8234 ( \17356 , \17344 , \17355 );
and \U$8235 ( \17357 , \16627 , \16631 );
and \U$8236 ( \17358 , \16631 , \16639 );
and \U$8237 ( \17359 , \16627 , \16639 );
or \U$8238 ( \17360 , \17357 , \17358 , \17359 );
and \U$8239 ( \17361 , \16655 , \10983 );
and \U$8240 ( \17362 , RIdec45c8_698, \9333 );
and \U$8241 ( \17363 , RIdec18c8_666, \9335 );
and \U$8242 ( \17364 , RIfce85e0_7666, \9337 );
and \U$8243 ( \17365 , RIdebebc8_634, \9339 );
and \U$8244 ( \17366 , RIfcb8bb0_7124, \9341 );
and \U$8245 ( \17367 , RIdebbec8_602, \9343 );
and \U$8246 ( \17368 , RIdeb91c8_570, \9345 );
and \U$8247 ( \17369 , RIdeb64c8_538, \9347 );
and \U$8248 ( \17370 , RIfc85d78_6545, \9349 );
and \U$8249 ( \17371 , RIdeb0ac8_474, \9351 );
and \U$8250 ( \17372 , RIfc85aa8_6543, \9353 );
and \U$8251 ( \17373 , RIdeaddc8_442, \9355 );
and \U$8252 ( \17374 , RIfc4d3d8_5901, \9357 );
and \U$8253 ( \17375 , RIdea8350_410, \9359 );
and \U$8254 ( \17376 , RIdea1a50_378, \9361 );
and \U$8255 ( \17377 , RIde9b150_346, \9363 );
and \U$8256 ( \17378 , RIfc85ee0_6546, \9365 );
and \U$8257 ( \17379 , RIfc9c9b0_6804, \9367 );
and \U$8258 ( \17380 , RIfce13f8_7585, \9369 );
and \U$8259 ( \17381 , RIfcb8778_7121, \9371 );
and \U$8260 ( \17382 , RIfe8d510_7952, \9373 );
and \U$8261 ( \17383 , RIfe8d3a8_7951, \9375 );
and \U$8262 ( \17384 , RIde886b8_255, \9377 );
and \U$8263 ( \17385 , RIde841d0_234, \9379 );
and \U$8264 ( \17386 , RIde806c0_216, \9381 );
and \U$8265 ( \17387 , RIfcb8070_7116, \9383 );
and \U$8266 ( \17388 , RIfce1128_7583, \9385 );
and \U$8267 ( \17389 , RIfc9c140_6798, \9387 );
and \U$8268 ( \17390 , RIee38d10_5105, \9389 );
and \U$8269 ( \17391 , RIe16ac70_2592, \9391 );
and \U$8270 ( \17392 , RIfc850d0_6536, \9393 );
and \U$8271 ( \17393 , RIe167160_2550, \9395 );
and \U$8272 ( \17394 , RIe1645c8_2519, \9397 );
and \U$8273 ( \17395 , RIe1618c8_2487, \9399 );
and \U$8274 ( \17396 , RIee36b50_5081, \9401 );
and \U$8275 ( \17397 , RIe15ebc8_2455, \9403 );
and \U$8276 ( \17398 , RIee35d40_5071, \9405 );
and \U$8277 ( \17399 , RIe15bec8_2423, \9407 );
and \U$8278 ( \17400 , RIe1564c8_2359, \9409 );
and \U$8279 ( \17401 , RIe1537c8_2327, \9411 );
and \U$8280 ( \17402 , RIfc3ef90_5742, \9413 );
and \U$8281 ( \17403 , RIe150ac8_2295, \9415 );
and \U$8282 ( \17404 , RIfe8d7e0_7954, \9417 );
and \U$8283 ( \17405 , RIe14ddc8_2263, \9419 );
and \U$8284 ( \17406 , RIfce0fc0_7582, \9421 );
and \U$8285 ( \17407 , RIe14b0c8_2231, \9423 );
and \U$8286 ( \17408 , RIe1483c8_2199, \9425 );
and \U$8287 ( \17409 , RIe1456c8_2167, \9427 );
and \U$8288 ( \17410 , RIee33e50_5049, \9429 );
and \U$8289 ( \17411 , RIee32c08_5036, \9431 );
and \U$8290 ( \17412 , RIee319c0_5023, \9433 );
and \U$8291 ( \17413 , RIee30d18_5014, \9435 );
and \U$8292 ( \17414 , RIfe8cf70_7948, \9437 );
and \U$8293 ( \17415 , RIfe8ce08_7947, \9439 );
and \U$8294 ( \17416 , RIfe8d240_7950, \9441 );
and \U$8295 ( \17417 , RIfe8d0d8_7949, \9443 );
and \U$8296 ( \17418 , RIfce9dc8_7683, \9445 );
and \U$8297 ( \17419 , RIee2ef90_4993, \9447 );
and \U$8298 ( \17420 , RIfce51d8_7629, \9449 );
and \U$8299 ( \17421 , RIee2cdd0_4969, \9451 );
and \U$8300 ( \17422 , RIdf34af8_1976, \9453 );
and \U$8301 ( \17423 , RIfe8d678_7953, \9455 );
and \U$8302 ( \17424 , RIdf30610_1927, \9457 );
and \U$8303 ( \17425 , RIdf2e720_1905, \9459 );
or \U$8304 ( \17426 , \17362 , \17363 , \17364 , \17365 , \17366 , \17367 , \17368 , \17369 , \17370 , \17371 , \17372 , \17373 , \17374 , \17375 , \17376 , \17377 , \17378 , \17379 , \17380 , \17381 , \17382 , \17383 , \17384 , \17385 , \17386 , \17387 , \17388 , \17389 , \17390 , \17391 , \17392 , \17393 , \17394 , \17395 , \17396 , \17397 , \17398 , \17399 , \17400 , \17401 , \17402 , \17403 , \17404 , \17405 , \17406 , \17407 , \17408 , \17409 , \17410 , \17411 , \17412 , \17413 , \17414 , \17415 , \17416 , \17417 , \17418 , \17419 , \17420 , \17421 , \17422 , \17423 , \17424 , \17425 );
and \U$8305 ( \17427 , RIee2b318_4950, \9462 );
and \U$8306 ( \17428 , RIee29c98_4934, \9464 );
and \U$8307 ( \17429 , RIee28780_4919, \9466 );
and \U$8308 ( \17430 , RIee27538_4906, \9468 );
and \U$8309 ( \17431 , RIdf299c8_1850, \9470 );
and \U$8310 ( \17432 , RIdf276a0_1825, \9472 );
and \U$8311 ( \17433 , RIdf25918_1804, \9474 );
and \U$8312 ( \17434 , RIdf23cf8_1784, \9476 );
and \U$8313 ( \17435 , RIfc83ff0_6524, \9478 );
and \U$8314 ( \17436 , RIfcb73c8_7107, \9480 );
and \U$8315 ( \17437 , RIfc51320_5946, \9482 );
and \U$8316 ( \17438 , RIfcdaa80_7510, \9484 );
and \U$8317 ( \17439 , RIfc83d20_6522, \9486 );
and \U$8318 ( \17440 , RIdf1ee38_1728, \9488 );
and \U$8319 ( \17441 , RIfc51b90_5952, \9490 );
and \U$8320 ( \17442 , RIdf18a60_1657, \9492 );
and \U$8321 ( \17443 , RIdf16198_1628, \9494 );
and \U$8322 ( \17444 , RIdf13498_1596, \9496 );
and \U$8323 ( \17445 , RIdf10798_1564, \9498 );
and \U$8324 ( \17446 , RIdf0da98_1532, \9500 );
and \U$8325 ( \17447 , RIdf0ad98_1500, \9502 );
and \U$8326 ( \17448 , RIdf08098_1468, \9504 );
and \U$8327 ( \17449 , RIdf05398_1436, \9506 );
and \U$8328 ( \17450 , RIdf02698_1404, \9508 );
and \U$8329 ( \17451 , RIdefcc98_1340, \9510 );
and \U$8330 ( \17452 , RIdef9f98_1308, \9512 );
and \U$8331 ( \17453 , RIdef7298_1276, \9514 );
and \U$8332 ( \17454 , RIdef4598_1244, \9516 );
and \U$8333 ( \17455 , RIdef1898_1212, \9518 );
and \U$8334 ( \17456 , RIdeeeb98_1180, \9520 );
and \U$8335 ( \17457 , RIdeebe98_1148, \9522 );
and \U$8336 ( \17458 , RIdee9198_1116, \9524 );
and \U$8337 ( \17459 , RIee25210_4881, \9526 );
and \U$8338 ( \17460 , RIee24400_4871, \9528 );
and \U$8339 ( \17461 , RIee238c0_4863, \9530 );
and \U$8340 ( \17462 , RIee22ee8_4856, \9532 );
and \U$8341 ( \17463 , RIfe8cca0_7946, \9534 );
and \U$8342 ( \17464 , RIdee2118_1036, \9536 );
and \U$8343 ( \17465 , RIfe8cb38_7945, \9538 );
and \U$8344 ( \17466 , RIdeddf00_989, \9540 );
and \U$8345 ( \17467 , RIfcc5a68_7271, \9542 );
and \U$8346 ( \17468 , RIee21f70_4845, \9544 );
and \U$8347 ( \17469 , RIfcb6cc0_7102, \9546 );
and \U$8348 ( \17470 , RIee20e90_4833, \9548 );
and \U$8349 ( \17471 , RIded8c08_930, \9550 );
and \U$8350 ( \17472 , RIded6778_904, \9552 );
and \U$8351 ( \17473 , RIded4720_881, \9554 );
and \U$8352 ( \17474 , RIded23f8_856, \9556 );
and \U$8353 ( \17475 , RIdecf9c8_826, \9558 );
and \U$8354 ( \17476 , RIdecccc8_794, \9560 );
and \U$8355 ( \17477 , RIdec9fc8_762, \9562 );
and \U$8356 ( \17478 , RIdec72c8_730, \9564 );
and \U$8357 ( \17479 , RIdeb37c8_506, \9566 );
and \U$8358 ( \17480 , RIde94850_314, \9568 );
and \U$8359 ( \17481 , RIe16d3d0_2620, \9570 );
and \U$8360 ( \17482 , RIe1591c8_2391, \9572 );
and \U$8361 ( \17483 , RIe1429c8_2135, \9574 );
and \U$8362 ( \17484 , RIdf373c0_2005, \9576 );
and \U$8363 ( \17485 , RIdf2ba20_1873, \9578 );
and \U$8364 ( \17486 , RIdf1c2a0_1697, \9580 );
and \U$8365 ( \17487 , RIdeff998_1372, \9582 );
and \U$8366 ( \17488 , RIdee6498_1084, \9584 );
and \U$8367 ( \17489 , RIdedb200_957, \9586 );
and \U$8368 ( \17490 , RIde7a798_187, \9588 );
or \U$8369 ( \17491 , \17427 , \17428 , \17429 , \17430 , \17431 , \17432 , \17433 , \17434 , \17435 , \17436 , \17437 , \17438 , \17439 , \17440 , \17441 , \17442 , \17443 , \17444 , \17445 , \17446 , \17447 , \17448 , \17449 , \17450 , \17451 , \17452 , \17453 , \17454 , \17455 , \17456 , \17457 , \17458 , \17459 , \17460 , \17461 , \17462 , \17463 , \17464 , \17465 , \17466 , \17467 , \17468 , \17469 , \17470 , \17471 , \17472 , \17473 , \17474 , \17475 , \17476 , \17477 , \17478 , \17479 , \17480 , \17481 , \17482 , \17483 , \17484 , \17485 , \17486 , \17487 , \17488 , \17489 , \17490 );
or \U$8370 ( \17492 , \17426 , \17491 );
_DC g659b ( \17493_nG659b , \17492 , \9597 );
and \U$8371 ( \17494 , RIe19c860_3158, \9059 );
and \U$8372 ( \17495 , RIe199b60_3126, \9061 );
and \U$8373 ( \17496 , RIf145220_5246, \9063 );
and \U$8374 ( \17497 , RIe196e60_3094, \9065 );
and \U$8375 ( \17498 , RIf144140_5234, \9067 );
and \U$8376 ( \17499 , RIe194160_3062, \9069 );
and \U$8377 ( \17500 , RIe191460_3030, \9071 );
and \U$8378 ( \17501 , RIe18e760_2998, \9073 );
and \U$8379 ( \17502 , RIe188d60_2934, \9075 );
and \U$8380 ( \17503 , RIe186060_2902, \9077 );
and \U$8381 ( \17504 , RIf1431c8_5223, \9079 );
and \U$8382 ( \17505 , RIe183360_2870, \9081 );
and \U$8383 ( \17506 , RIf142ac0_5218, \9083 );
and \U$8384 ( \17507 , RIe180660_2838, \9085 );
and \U$8385 ( \17508 , RIe17d960_2806, \9087 );
and \U$8386 ( \17509 , RIe17ac60_2774, \9089 );
and \U$8387 ( \17510 , RIf141cb0_5208, \9091 );
and \U$8388 ( \17511 , RIf140798_5193, \9093 );
and \U$8389 ( \17512 , RIf13ff28_5187, \9095 );
and \U$8390 ( \17513 , RIfe8be90_7936, \9097 );
and \U$8391 ( \17514 , RIfceb880_7702, \9099 );
and \U$8392 ( \17515 , RIf13eb78_5173, \9101 );
and \U$8393 ( \17516 , RIee3e008_5164, \9103 );
and \U$8394 ( \17517 , RIee3cdc0_5151, \9105 );
and \U$8395 ( \17518 , RIee3bb78_5138, \9107 );
and \U$8396 ( \17519 , RIee3aa98_5126, \9109 );
and \U$8397 ( \17520 , RIee396e8_5112, \9111 );
and \U$8398 ( \17521 , RIe172c68_2683, \9113 );
and \U$8399 ( \17522 , RIf16fac0_5730, \9115 );
and \U$8400 ( \17523 , RIf16ef80_5722, \9117 );
and \U$8401 ( \17524 , RIf16dbd0_5708, \9119 );
and \U$8402 ( \17525 , RIfcc4af0_7260, \9121 );
and \U$8403 ( \17526 , RIf16c820_5694, \9123 );
and \U$8404 ( \17527 , RIe222bb8_4685, \9125 );
and \U$8405 ( \17528 , RIf16b740_5682, \9127 );
and \U$8406 ( \17529 , RIe21feb8_4653, \9129 );
and \U$8407 ( \17530 , RIf16a7c8_5671, \9131 );
and \U$8408 ( \17531 , RIe21d1b8_4621, \9133 );
and \U$8409 ( \17532 , RIe2177b8_4557, \9135 );
and \U$8410 ( \17533 , RIe214ab8_4525, \9137 );
and \U$8411 ( \17534 , RIfe8c430_7940, \9139 );
and \U$8412 ( \17535 , RIe211db8_4493, \9141 );
and \U$8413 ( \17536 , RIf1688d8_5649, \9143 );
and \U$8414 ( \17537 , RIe20f0b8_4461, \9145 );
and \U$8415 ( \17538 , RIf167960_5638, \9147 );
and \U$8416 ( \17539 , RIe20c3b8_4429, \9149 );
and \U$8417 ( \17540 , RIe2096b8_4397, \9151 );
and \U$8418 ( \17541 , RIe2069b8_4365, \9153 );
and \U$8419 ( \17542 , RIf1669e8_5627, \9155 );
and \U$8420 ( \17543 , RIf165908_5615, \9157 );
and \U$8421 ( \17544 , RIfe8c9d0_7944, \9159 );
and \U$8422 ( \17545 , RIfe8c700_7942, \9161 );
and \U$8423 ( \17546 , RIfc9c578_6801, \9163 );
and \U$8424 ( \17547 , RIf163ce8_5595, \9165 );
and \U$8425 ( \17548 , RIf162d70_5584, \9167 );
and \U$8426 ( \17549 , RIf161588_5567, \9169 );
and \U$8427 ( \17550 , RIf15f698_5545, \9171 );
and \U$8428 ( \17551 , RIf15d910_5524, \9173 );
and \U$8429 ( \17552 , RIfe8c598_7941, \9175 );
and \U$8430 ( \17553 , RIfe8c868_7943, \9177 );
and \U$8431 ( \17554 , RIf15c3f8_5509, \9179 );
and \U$8432 ( \17555 , RIf15aee0_5494, \9181 );
and \U$8433 ( \17556 , RIf15a0d0_5484, \9183 );
and \U$8434 ( \17557 , RIf1596f8_5477, \9185 );
or \U$8435 ( \17558 , \17494 , \17495 , \17496 , \17497 , \17498 , \17499 , \17500 , \17501 , \17502 , \17503 , \17504 , \17505 , \17506 , \17507 , \17508 , \17509 , \17510 , \17511 , \17512 , \17513 , \17514 , \17515 , \17516 , \17517 , \17518 , \17519 , \17520 , \17521 , \17522 , \17523 , \17524 , \17525 , \17526 , \17527 , \17528 , \17529 , \17530 , \17531 , \17532 , \17533 , \17534 , \17535 , \17536 , \17537 , \17538 , \17539 , \17540 , \17541 , \17542 , \17543 , \17544 , \17545 , \17546 , \17547 , \17548 , \17549 , \17550 , \17551 , \17552 , \17553 , \17554 , \17555 , \17556 , \17557 );
and \U$8436 ( \17559 , RIf158618_5465, \9188 );
and \U$8437 ( \17560 , RIf1573d0_5452, \9190 );
and \U$8438 ( \17561 , RIf156b60_5446, \9192 );
and \U$8439 ( \17562 , RIfec1f68_8327, \9194 );
and \U$8440 ( \17563 , RIf155eb8_5437, \9196 );
and \U$8441 ( \17564 , RIf155378_5429, \9198 );
and \U$8442 ( \17565 , RIf153fc8_5415, \9200 );
and \U$8443 ( \17566 , RIfe8bff8_7937, \9202 );
and \U$8444 ( \17567 , RIf152948_5399, \9204 );
and \U$8445 ( \17568 , RIf151598_5385, \9206 );
and \U$8446 ( \17569 , RIf150080_5370, \9208 );
and \U$8447 ( \17570 , RIfe8c2c8_7939, \9210 );
and \U$8448 ( \17571 , RIf14f270_5360, \9212 );
and \U$8449 ( \17572 , RIfc503a8_5935, \9214 );
and \U$8450 ( \17573 , RIf14d650_5340, \9216 );
and \U$8451 ( \17574 , RIfe8c160_7938, \9218 );
and \U$8452 ( \17575 , RIe1ea920_4046, \9220 );
and \U$8453 ( \17576 , RIe1e7c20_4014, \9222 );
and \U$8454 ( \17577 , RIe1e4f20_3982, \9224 );
and \U$8455 ( \17578 , RIe1e2220_3950, \9226 );
and \U$8456 ( \17579 , RIe1df520_3918, \9228 );
and \U$8457 ( \17580 , RIe1dc820_3886, \9230 );
and \U$8458 ( \17581 , RIe1d9b20_3854, \9232 );
and \U$8459 ( \17582 , RIe1d6e20_3822, \9234 );
and \U$8460 ( \17583 , RIe1d1420_3758, \9236 );
and \U$8461 ( \17584 , RIe1ce720_3726, \9238 );
and \U$8462 ( \17585 , RIe1cba20_3694, \9240 );
and \U$8463 ( \17586 , RIe1c8d20_3662, \9242 );
and \U$8464 ( \17587 , RIe1c6020_3630, \9244 );
and \U$8465 ( \17588 , RIe1c3320_3598, \9246 );
and \U$8466 ( \17589 , RIe1c0620_3566, \9248 );
and \U$8467 ( \17590 , RIe1bd920_3534, \9250 );
and \U$8468 ( \17591 , RIf14c2a0_5326, \9252 );
and \U$8469 ( \17592 , RIf14aef0_5312, \9254 );
and \U$8470 ( \17593 , RIe1b88f8_3477, \9256 );
and \U$8471 ( \17594 , RIe1b68a0_3454, \9258 );
and \U$8472 ( \17595 , RIfcd4db0_7444, \9260 );
and \U$8473 ( \17596 , RIfc4ebc0_5918, \9262 );
and \U$8474 ( \17597 , RIfec1e00_8326, \9264 );
and \U$8475 ( \17598 , RIfe8bd28_7935, \9266 );
and \U$8476 ( \17599 , RIf148790_5284, \9268 );
and \U$8477 ( \17600 , RIf1476b0_5272, \9270 );
and \U$8478 ( \17601 , RIfe8ba58_7933, \9272 );
and \U$8479 ( \17602 , RIfec1b30_8324, \9274 );
and \U$8480 ( \17603 , RIfc4e788_5915, \9276 );
and \U$8481 ( \17604 , RIfcb8e80_7126, \9278 );
and \U$8482 ( \17605 , RIfe8bbc0_7934, \9280 );
and \U$8483 ( \17606 , RIfec1c98_8325, \9282 );
and \U$8484 ( \17607 , RIe1a7c60_3286, \9284 );
and \U$8485 ( \17608 , RIe1a4f60_3254, \9286 );
and \U$8486 ( \17609 , RIe1a2260_3222, \9288 );
and \U$8487 ( \17610 , RIe19f560_3190, \9290 );
and \U$8488 ( \17611 , RIe18ba60_2966, \9292 );
and \U$8489 ( \17612 , RIe177f60_2742, \9294 );
and \U$8490 ( \17613 , RIe2258b8_4717, \9296 );
and \U$8491 ( \17614 , RIe21a4b8_4589, \9298 );
and \U$8492 ( \17615 , RIe203cb8_4333, \9300 );
and \U$8493 ( \17616 , RIe1fdd18_4265, \9302 );
and \U$8494 ( \17617 , RIe1f70d0_4188, \9304 );
and \U$8495 ( \17618 , RIe1efc18_4105, \9306 );
and \U$8496 ( \17619 , RIe1d4120_3790, \9308 );
and \U$8497 ( \17620 , RIe1bac20_3502, \9310 );
and \U$8498 ( \17621 , RIe1ada98_3353, \9312 );
and \U$8499 ( \17622 , RIe1700d0_2652, \9314 );
or \U$8500 ( \17623 , \17559 , \17560 , \17561 , \17562 , \17563 , \17564 , \17565 , \17566 , \17567 , \17568 , \17569 , \17570 , \17571 , \17572 , \17573 , \17574 , \17575 , \17576 , \17577 , \17578 , \17579 , \17580 , \17581 , \17582 , \17583 , \17584 , \17585 , \17586 , \17587 , \17588 , \17589 , \17590 , \17591 , \17592 , \17593 , \17594 , \17595 , \17596 , \17597 , \17598 , \17599 , \17600 , \17601 , \17602 , \17603 , \17604 , \17605 , \17606 , \17607 , \17608 , \17609 , \17610 , \17611 , \17612 , \17613 , \17614 , \17615 , \17616 , \17617 , \17618 , \17619 , \17620 , \17621 , \17622 );
or \U$8501 ( \17624 , \17558 , \17623 );
_DC g659c ( \17625_nG659c , \17624 , \9323 );
and g659d ( \17626_nG659d , \17493_nG659b , \17625_nG659c );
buf \U$8502 ( \17627 , \17626_nG659d );
and \U$8503 ( \17628 , \17627 , \10691 );
nor \U$8504 ( \17629 , \17361 , \17628 );
xnor \U$8505 ( \17630 , \17629 , \10980 );
and \U$8506 ( \17631 , \11586 , \15336 );
and \U$8507 ( \17632 , \12448 , \14963 );
nor \U$8508 ( \17633 , \17631 , \17632 );
xnor \U$8509 ( \17634 , \17633 , \15342 );
xor \U$8510 ( \17635 , \17630 , \17634 );
and \U$8511 ( \17636 , \10988 , \16635 );
and \U$8512 ( \17637 , \11270 , \16301 );
nor \U$8513 ( \17638 , \17636 , \17637 );
xnor \U$8514 ( \17639 , \17638 , \16625 );
xor \U$8515 ( \17640 , \17635 , \17639 );
xor \U$8516 ( \17641 , \17360 , \17640 );
and \U$8517 ( \17642 , \15321 , \11574 );
and \U$8518 ( \17643 , \16267 , \11278 );
nor \U$8519 ( \17644 , \17642 , \17643 );
xnor \U$8520 ( \17645 , \17644 , \11580 );
and \U$8521 ( \17646 , \12769 , \14054 );
and \U$8522 ( \17647 , \13679 , \13692 );
nor \U$8523 ( \17648 , \17646 , \17647 );
xnor \U$8524 ( \17649 , \17648 , \14035 );
xor \U$8525 ( \17650 , \17645 , \17649 );
_DC g5146 ( \17651_nG5146 , \17492 , \9597 );
_DC g51ca ( \17652_nG51ca , \17624 , \9323 );
xor g51cb ( \17653_nG51cb , \17651_nG5146 , \17652_nG51ca );
buf \U$8526 ( \17654 , \17653_nG51cb );
xor \U$8527 ( \17655 , \17654 , \16622 );
and \U$8528 ( \17656 , \10687 , \17655 );
xor \U$8529 ( \17657 , \17650 , \17656 );
xor \U$8530 ( \17658 , \17641 , \17657 );
xor \U$8531 ( \17659 , \17356 , \17658 );
xor \U$8532 ( \17660 , \17340 , \17659 );
and \U$8533 ( \17661 , \16670 , \16674 );
and \U$8534 ( \17662 , \16675 , \16678 );
or \U$8535 ( \17663 , \17661 , \17662 );
xor \U$8536 ( \17664 , \17660 , \17663 );
buf g9bea ( \17665_nG9bea , \17664 );
and \U$8537 ( \17666 , \10704 , \17665_nG9bea );
or \U$8538 ( \17667 , \17336 , \17666 );
xor \U$8539 ( \17668 , \10703 , \17667 );
buf \U$8540 ( \17669 , \17668 );
buf \U$8542 ( \17670 , \17669 );
xor \U$8543 ( \17671 , \17335 , \17670 );
buf \U$8544 ( \17672 , \17671 );
and \U$8545 ( \17673 , \16339 , \16345 );
and \U$8546 ( \17674 , \16339 , \16685 );
and \U$8547 ( \17675 , \16345 , \16685 );
or \U$8548 ( \17676 , \17673 , \17674 , \17675 );
buf \U$8549 ( \17677 , \17676 );
xor \U$8550 ( \17678 , \17672 , \17677 );
and \U$8551 ( \17679 , \16704 , \16710 );
and \U$8552 ( \17680 , \16704 , \16717 );
and \U$8553 ( \17681 , \16710 , \16717 );
or \U$8554 ( \17682 , \17679 , \17680 , \17681 );
buf \U$8555 ( \17683 , \17682 );
and \U$8556 ( \17684 , \12157 , \14070_nG9bf9 );
and \U$8557 ( \17685 , \12154 , \14984_nG9bf6 );
or \U$8558 ( \17686 , \17684 , \17685 );
xor \U$8559 ( \17687 , \12153 , \17686 );
buf \U$8560 ( \17688 , \17687 );
buf \U$8562 ( \17689 , \17688 );
xor \U$8563 ( \17690 , \17683 , \17689 );
and \U$8564 ( \17691 , \10421 , \15373_nG9bf3 );
and \U$8565 ( \17692 , \10418 , \16315_nG9bf0 );
or \U$8566 ( \17693 , \17691 , \17692 );
xor \U$8567 ( \17694 , \10417 , \17693 );
buf \U$8568 ( \17695 , \17694 );
buf \U$8570 ( \17696 , \17695 );
xor \U$8571 ( \17697 , \17690 , \17696 );
buf \U$8572 ( \17698 , \17697 );
xor \U$8573 ( \17699 , \17678 , \17698 );
buf \U$8574 ( \17700 , \17699 );
and \U$8575 ( \17701 , \16687 , \16692 );
and \U$8576 ( \17702 , \16687 , \16730 );
and \U$8577 ( \17703 , \16692 , \16730 );
or \U$8578 ( \17704 , \17701 , \17702 , \17703 );
buf \U$8579 ( \17705 , \17704 );
xor \U$8580 ( \17706 , \17700 , \17705 );
and \U$8581 ( \17707 , \16732 , \16737 );
and \U$8582 ( \17708 , \16732 , \16743 );
and \U$8583 ( \17709 , \16737 , \16743 );
or \U$8584 ( \17710 , \17707 , \17708 , \17709 );
buf \U$8585 ( \17711 , \17710 );
xor \U$8586 ( \17712 , \17706 , \17711 );
and \U$8587 ( \17713 , \16745 , \17712 );
and \U$8588 ( \17714 , \17303 , \17712 );
or \U$8589 ( \17715 , \17304 , \17713 , \17714 );
and \U$8590 ( \17716 , \17309 , \17334 );
and \U$8591 ( \17717 , \17309 , \17670 );
and \U$8592 ( \17718 , \17334 , \17670 );
or \U$8593 ( \17719 , \17716 , \17717 , \17718 );
buf \U$8594 ( \17720 , \17719 );
and \U$8595 ( \17721 , \17683 , \17689 );
and \U$8596 ( \17722 , \17683 , \17696 );
and \U$8597 ( \17723 , \17689 , \17696 );
or \U$8598 ( \17724 , \17721 , \17722 , \17723 );
buf \U$8599 ( \17725 , \17724 );
and \U$8600 ( \17726 , \17293 , \17300 );
buf \U$8601 ( \17727 , \17726 );
buf \U$8603 ( \17728 , \17727 );
and \U$8604 ( \17729 , \15940 , \11283_nG9c08 );
and \U$8605 ( \17730 , \15937 , \11598_nG9c05 );
or \U$8606 ( \17731 , \17729 , \17730 );
xor \U$8607 ( \17732 , \15936 , \17731 );
buf \U$8608 ( \17733 , \17732 );
buf \U$8610 ( \17734 , \17733 );
xor \U$8611 ( \17735 , \17728 , \17734 );
buf \U$8612 ( \17736 , \17735 );
and \U$8613 ( \17737 , \17297 , \10694_nG9c0e );
and \U$8614 ( \17738 , \17294 , \10995_nG9c0b );
or \U$8615 ( \17739 , \17737 , \17738 );
xor \U$8616 ( \17740 , \17293 , \17739 );
buf \U$8617 ( \17741 , \17740 );
buf \U$8619 ( \17742 , \17741 );
xor \U$8620 ( \17743 , \17736 , \17742 );
and \U$8621 ( \17744 , \14631 , \12470_nG9c02 );
and \U$8622 ( \17745 , \14628 , \12801_nG9bff );
or \U$8623 ( \17746 , \17744 , \17745 );
xor \U$8624 ( \17747 , \14627 , \17746 );
buf \U$8625 ( \17748 , \17747 );
buf \U$8627 ( \17749 , \17748 );
xor \U$8628 ( \17750 , \17743 , \17749 );
buf \U$8629 ( \17751 , \17750 );
and \U$8630 ( \17752 , \17315 , \17321 );
buf \U$8631 ( \17753 , \17752 );
xor \U$8632 ( \17754 , \17751 , \17753 );
and \U$8633 ( \17755 , \13370 , \13705_nG9bfc );
and \U$8634 ( \17756 , \13367 , \14070_nG9bf9 );
or \U$8635 ( \17757 , \17755 , \17756 );
xor \U$8636 ( \17758 , \13366 , \17757 );
buf \U$8637 ( \17759 , \17758 );
buf \U$8639 ( \17760 , \17759 );
xor \U$8640 ( \17761 , \17754 , \17760 );
buf \U$8641 ( \17762 , \17761 );
xor \U$8642 ( \17763 , \17725 , \17762 );
and \U$8643 ( \17764 , \10707 , \17665_nG9bea );
and \U$8644 ( \17765 , \17360 , \17640 );
and \U$8645 ( \17766 , \17640 , \17657 );
and \U$8646 ( \17767 , \17360 , \17657 );
or \U$8647 ( \17768 , \17765 , \17766 , \17767 );
and \U$8648 ( \17769 , \17627 , \10983 );
and \U$8649 ( \17770 , RIdec4730_699, \9333 );
and \U$8650 ( \17771 , RIdec1a30_667, \9335 );
and \U$8651 ( \17772 , RIfce3f90_7616, \9337 );
and \U$8652 ( \17773 , RIdebed30_635, \9339 );
and \U$8653 ( \17774 , RIfcc3308_7243, \9341 );
and \U$8654 ( \17775 , RIdebc030_603, \9343 );
and \U$8655 ( \17776 , RIdeb9330_571, \9345 );
and \U$8656 ( \17777 , RIdeb6630_539, \9347 );
and \U$8657 ( \17778 , RIfc8c588_6619, \9349 );
and \U$8658 ( \17779 , RIdeb0c30_475, \9351 );
and \U$8659 ( \17780 , RIfc5a998_6053, \9353 );
and \U$8660 ( \17781 , RIdeadf30_443, \9355 );
and \U$8661 ( \17782 , RIfc99b48_6771, \9357 );
and \U$8662 ( \17783 , RIdea8698_411, \9359 );
and \U$8663 ( \17784 , RIdea1d98_379, \9361 );
and \U$8664 ( \17785 , RIde9b498_347, \9363 );
and \U$8665 ( \17786 , RIfc78bf0_6396, \9365 );
and \U$8666 ( \17787 , RIfcbc558_7165, \9367 );
and \U$8667 ( \17788 , RIfca12d0_6856, \9369 );
and \U$8668 ( \17789 , RIfca3fd0_6888, \9371 );
and \U$8669 ( \17790 , RIfec2670_8332, \9373 );
and \U$8670 ( \17791 , RIfec2508_8331, \9375 );
and \U$8671 ( \17792 , RIde88a00_256, \9377 );
and \U$8672 ( \17793 , RIde84518_235, \9379 );
and \U$8673 ( \17794 , RIfcc35d8_7245, \9381 );
and \U$8674 ( \17795 , RIfcb57a8_7087, \9383 );
and \U$8675 ( \17796 , RIfc5a290_6048, \9385 );
and \U$8676 ( \17797 , RIfca3058_6877, \9387 );
and \U$8677 ( \17798 , RIee38e78_5106, \9389 );
and \U$8678 ( \17799 , RIfec27d8_8333, \9391 );
and \U$8679 ( \17800 , RIfca3328_6879, \9393 );
and \U$8680 ( \17801 , RIe1672c8_2551, \9395 );
and \U$8681 ( \17802 , RIe164730_2520, \9397 );
and \U$8682 ( \17803 , RIe161a30_2488, \9399 );
and \U$8683 ( \17804 , RIee36cb8_5082, \9401 );
and \U$8684 ( \17805 , RIe15ed30_2456, \9403 );
and \U$8685 ( \17806 , RIfcc7250_7288, \9405 );
and \U$8686 ( \17807 , RIe15c030_2424, \9407 );
and \U$8687 ( \17808 , RIe156630_2360, \9409 );
and \U$8688 ( \17809 , RIe153930_2328, \9411 );
and \U$8689 ( \17810 , RIfcc7688_7291, \9413 );
and \U$8690 ( \17811 , RIe150c30_2296, \9415 );
and \U$8691 ( \17812 , RIfc8af08_6603, \9417 );
and \U$8692 ( \17813 , RIe14df30_2264, \9419 );
and \U$8693 ( \17814 , RIfc9a250_6776, \9421 );
and \U$8694 ( \17815 , RIe14b230_2232, \9423 );
and \U$8695 ( \17816 , RIe148530_2200, \9425 );
and \U$8696 ( \17817 , RIe145830_2168, \9427 );
and \U$8697 ( \17818 , RIfc9aac0_6782, \9429 );
and \U$8698 ( \17819 , RIfc56bb8_6009, \9431 );
and \U$8699 ( \17820 , RIfca1ca8_6863, \9433 );
and \U$8700 ( \17821 , RIfcec960_7714, \9435 );
and \U$8701 ( \17822 , RIe1406a0_2110, \9437 );
and \U$8702 ( \17823 , RIdf3e440_2085, \9439 );
and \U$8703 ( \17824 , RIdf3c280_2061, \9441 );
and \U$8704 ( \17825 , RIdf39f58_2036, \9443 );
and \U$8705 ( \17826 , RIfc9a958_6781, \9445 );
and \U$8706 ( \17827 , RIee2f0f8_4994, \9447 );
and \U$8707 ( \17828 , RIfcdb458_7517, \9449 );
and \U$8708 ( \17829 , RIee2cf38_4970, \9451 );
and \U$8709 ( \17830 , RIdf34c60_1977, \9453 );
and \U$8710 ( \17831 , RIfec2940_8334, \9455 );
and \U$8711 ( \17832 , RIdf30778_1928, \9457 );
and \U$8712 ( \17833 , RIdf2e888_1906, \9459 );
or \U$8713 ( \17834 , \17770 , \17771 , \17772 , \17773 , \17774 , \17775 , \17776 , \17777 , \17778 , \17779 , \17780 , \17781 , \17782 , \17783 , \17784 , \17785 , \17786 , \17787 , \17788 , \17789 , \17790 , \17791 , \17792 , \17793 , \17794 , \17795 , \17796 , \17797 , \17798 , \17799 , \17800 , \17801 , \17802 , \17803 , \17804 , \17805 , \17806 , \17807 , \17808 , \17809 , \17810 , \17811 , \17812 , \17813 , \17814 , \17815 , \17816 , \17817 , \17818 , \17819 , \17820 , \17821 , \17822 , \17823 , \17824 , \17825 , \17826 , \17827 , \17828 , \17829 , \17830 , \17831 , \17832 , \17833 );
and \U$8714 ( \17835 , RIee2b480_4951, \9462 );
and \U$8715 ( \17836 , RIfec23a0_8330, \9464 );
and \U$8716 ( \17837 , RIee288e8_4920, \9466 );
and \U$8717 ( \17838 , RIfec2238_8329, \9468 );
and \U$8718 ( \17839 , RIdf29b30_1851, \9470 );
and \U$8719 ( \17840 , RIdf27808_1826, \9472 );
and \U$8720 ( \17841 , RIdf25a80_1805, \9474 );
and \U$8721 ( \17842 , RIdf23e60_1785, \9476 );
and \U$8722 ( \17843 , RIfc55100_5990, \9478 );
and \U$8723 ( \17844 , RIfcd9f40_7502, \9480 );
and \U$8724 ( \17845 , RIfc54f98_5989, \9482 );
and \U$8725 ( \17846 , RIfc54cc8_5987, \9484 );
and \U$8726 ( \17847 , RIfc4b218_5877, \9486 );
and \U$8727 ( \17848 , RIdf1efa0_1729, \9488 );
and \U$8728 ( \17849 , RIfcc69e0_7282, \9490 );
and \U$8729 ( \17850 , RIdf18bc8_1658, \9492 );
and \U$8730 ( \17851 , RIdf16300_1629, \9494 );
and \U$8731 ( \17852 , RIdf13600_1597, \9496 );
and \U$8732 ( \17853 , RIdf10900_1565, \9498 );
and \U$8733 ( \17854 , RIdf0dc00_1533, \9500 );
and \U$8734 ( \17855 , RIdf0af00_1501, \9502 );
and \U$8735 ( \17856 , RIdf08200_1469, \9504 );
and \U$8736 ( \17857 , RIdf05500_1437, \9506 );
and \U$8737 ( \17858 , RIdf02800_1405, \9508 );
and \U$8738 ( \17859 , RIdefce00_1341, \9510 );
and \U$8739 ( \17860 , RIdefa100_1309, \9512 );
and \U$8740 ( \17861 , RIdef7400_1277, \9514 );
and \U$8741 ( \17862 , RIdef4700_1245, \9516 );
and \U$8742 ( \17863 , RIdef1a00_1213, \9518 );
and \U$8743 ( \17864 , RIdeeed00_1181, \9520 );
and \U$8744 ( \17865 , RIdeec000_1149, \9522 );
and \U$8745 ( \17866 , RIdee9300_1117, \9524 );
and \U$8746 ( \17867 , RIfce4ad0_7624, \9526 );
and \U$8747 ( \17868 , RIfc9e8a0_6826, \9528 );
and \U$8748 ( \17869 , RIfcc46b8_7257, \9530 );
and \U$8749 ( \17870 , RIfcd4108_7435, \9532 );
and \U$8750 ( \17871 , RIdee4440_1061, \9534 );
and \U$8751 ( \17872 , RIdee2280_1037, \9536 );
and \U$8752 ( \17873 , RIdee0390_1015, \9538 );
and \U$8753 ( \17874 , RIdede068_990, \9540 );
and \U$8754 ( \17875 , RIfcda0a8_7503, \9542 );
and \U$8755 ( \17876 , RIfce54a8_7631, \9544 );
and \U$8756 ( \17877 , RIfca0790_6848, \9546 );
and \U$8757 ( \17878 , RIfc50ee8_5943, \9548 );
and \U$8758 ( \17879 , RIded8d70_931, \9550 );
and \U$8759 ( \17880 , RIded68e0_905, \9552 );
and \U$8760 ( \17881 , RIded4888_882, \9554 );
and \U$8761 ( \17882 , RIded2560_857, \9556 );
and \U$8762 ( \17883 , RIdecfb30_827, \9558 );
and \U$8763 ( \17884 , RIdecce30_795, \9560 );
and \U$8764 ( \17885 , RIdeca130_763, \9562 );
and \U$8765 ( \17886 , RIdec7430_731, \9564 );
and \U$8766 ( \17887 , RIdeb3930_507, \9566 );
and \U$8767 ( \17888 , RIde94b98_315, \9568 );
and \U$8768 ( \17889 , RIe16d538_2621, \9570 );
and \U$8769 ( \17890 , RIe159330_2392, \9572 );
and \U$8770 ( \17891 , RIe142b30_2136, \9574 );
and \U$8771 ( \17892 , RIdf37528_2006, \9576 );
and \U$8772 ( \17893 , RIdf2bb88_1874, \9578 );
and \U$8773 ( \17894 , RIdf1c408_1698, \9580 );
and \U$8774 ( \17895 , RIdeffb00_1373, \9582 );
and \U$8775 ( \17896 , RIdee6600_1085, \9584 );
and \U$8776 ( \17897 , RIdedb368_958, \9586 );
and \U$8777 ( \17898 , RIde7aae0_188, \9588 );
or \U$8778 ( \17899 , \17835 , \17836 , \17837 , \17838 , \17839 , \17840 , \17841 , \17842 , \17843 , \17844 , \17845 , \17846 , \17847 , \17848 , \17849 , \17850 , \17851 , \17852 , \17853 , \17854 , \17855 , \17856 , \17857 , \17858 , \17859 , \17860 , \17861 , \17862 , \17863 , \17864 , \17865 , \17866 , \17867 , \17868 , \17869 , \17870 , \17871 , \17872 , \17873 , \17874 , \17875 , \17876 , \17877 , \17878 , \17879 , \17880 , \17881 , \17882 , \17883 , \17884 , \17885 , \17886 , \17887 , \17888 , \17889 , \17890 , \17891 , \17892 , \17893 , \17894 , \17895 , \17896 , \17897 , \17898 );
or \U$8779 ( \17900 , \17834 , \17899 );
_DC g659e ( \17901_nG659e , \17900 , \9597 );
and \U$8780 ( \17902 , RIe19c9c8_3159, \9059 );
and \U$8781 ( \17903 , RIe199cc8_3127, \9061 );
and \U$8782 ( \17904 , RIfe8ea28_7967, \9063 );
and \U$8783 ( \17905 , RIe196fc8_3095, \9065 );
and \U$8784 ( \17906 , RIfec20d0_8328, \9067 );
and \U$8785 ( \17907 , RIe1942c8_3063, \9069 );
and \U$8786 ( \17908 , RIe1915c8_3031, \9071 );
and \U$8787 ( \17909 , RIe18e8c8_2999, \9073 );
and \U$8788 ( \17910 , RIe188ec8_2935, \9075 );
and \U$8789 ( \17911 , RIe1861c8_2903, \9077 );
and \U$8790 ( \17912 , RIfc68228_6207, \9079 );
and \U$8791 ( \17913 , RIe1834c8_2871, \9081 );
and \U$8792 ( \17914 , RIfccb5d0_7336, \9083 );
and \U$8793 ( \17915 , RIe1807c8_2839, \9085 );
and \U$8794 ( \17916 , RIe17dac8_2807, \9087 );
and \U$8795 ( \17917 , RIe17adc8_2775, \9089 );
and \U$8796 ( \17918 , RIf141e18_5209, \9091 );
and \U$8797 ( \17919 , RIf140900_5194, \9093 );
and \U$8798 ( \17920 , RIf140090_5188, \9095 );
and \U$8799 ( \17921 , RIe1753c8_2711, \9097 );
and \U$8800 ( \17922 , RIf13f988_5183, \9099 );
and \U$8801 ( \17923 , RIf13ece0_5174, \9101 );
and \U$8802 ( \17924 , RIee3e170_5165, \9103 );
and \U$8803 ( \17925 , RIee3cf28_5152, \9105 );
and \U$8804 ( \17926 , RIee3bce0_5139, \9107 );
and \U$8805 ( \17927 , RIee3ac00_5127, \9109 );
and \U$8806 ( \17928 , RIee39850_5113, \9111 );
and \U$8807 ( \17929 , RIe172dd0_2684, \9113 );
and \U$8808 ( \17930 , RIf16fc28_5731, \9115 );
and \U$8809 ( \17931 , RIf16f0e8_5723, \9117 );
and \U$8810 ( \17932 , RIf16dd38_5709, \9119 );
and \U$8811 ( \17933 , RIfce9120_7674, \9121 );
and \U$8812 ( \17934 , RIfc404a8_5757, \9123 );
and \U$8813 ( \17935 , RIe222d20_4686, \9125 );
and \U$8814 ( \17936 , RIf16b8a8_5683, \9127 );
and \U$8815 ( \17937 , RIe220020_4654, \9129 );
and \U$8816 ( \17938 , RIf16a930_5672, \9131 );
and \U$8817 ( \17939 , RIe21d320_4622, \9133 );
and \U$8818 ( \17940 , RIe217920_4558, \9135 );
and \U$8819 ( \17941 , RIe214c20_4526, \9137 );
and \U$8820 ( \17942 , RIfc5b910_6064, \9139 );
and \U$8821 ( \17943 , RIe211f20_4494, \9141 );
and \U$8822 ( \17944 , RIfe8e8c0_7966, \9143 );
and \U$8823 ( \17945 , RIe20f220_4462, \9145 );
and \U$8824 ( \17946 , RIfe8e758_7965, \9147 );
and \U$8825 ( \17947 , RIe20c520_4430, \9149 );
and \U$8826 ( \17948 , RIe209820_4398, \9151 );
and \U$8827 ( \17949 , RIe206b20_4366, \9153 );
and \U$8828 ( \17950 , RIf166b50_5628, \9155 );
and \U$8829 ( \17951 , RIf165a70_5616, \9157 );
and \U$8830 ( \17952 , RIfe8dd80_7958, \9159 );
and \U$8831 ( \17953 , RIfe8dab0_7956, \9161 );
and \U$8832 ( \17954 , RIf164c60_5606, \9163 );
and \U$8833 ( \17955 , RIf163e50_5596, \9165 );
and \U$8834 ( \17956 , RIf162ed8_5585, \9167 );
and \U$8835 ( \17957 , RIf1616f0_5568, \9169 );
and \U$8836 ( \17958 , RIf15f800_5546, \9171 );
and \U$8837 ( \17959 , RIf15da78_5525, \9173 );
and \U$8838 ( \17960 , RIfe8d948_7955, \9175 );
and \U$8839 ( \17961 , RIfe8dc18_7957, \9177 );
and \U$8840 ( \17962 , RIf15c560_5510, \9179 );
and \U$8841 ( \17963 , RIf15b048_5495, \9181 );
and \U$8842 ( \17964 , RIfc62828_6143, \9183 );
and \U$8843 ( \17965 , RIf159860_5478, \9185 );
or \U$8844 ( \17966 , \17902 , \17903 , \17904 , \17905 , \17906 , \17907 , \17908 , \17909 , \17910 , \17911 , \17912 , \17913 , \17914 , \17915 , \17916 , \17917 , \17918 , \17919 , \17920 , \17921 , \17922 , \17923 , \17924 , \17925 , \17926 , \17927 , \17928 , \17929 , \17930 , \17931 , \17932 , \17933 , \17934 , \17935 , \17936 , \17937 , \17938 , \17939 , \17940 , \17941 , \17942 , \17943 , \17944 , \17945 , \17946 , \17947 , \17948 , \17949 , \17950 , \17951 , \17952 , \17953 , \17954 , \17955 , \17956 , \17957 , \17958 , \17959 , \17960 , \17961 , \17962 , \17963 , \17964 , \17965 );
and \U$8845 ( \17967 , RIf158780_5466, \9188 );
and \U$8846 ( \17968 , RIf157538_5453, \9190 );
and \U$8847 ( \17969 , RIfca6e38_6921, \9192 );
and \U$8848 ( \17970 , RIe1f9b00_4218, \9194 );
and \U$8849 ( \17971 , RIfc61e50_6136, \9196 );
and \U$8850 ( \17972 , RIfc61748_6131, \9198 );
and \U$8851 ( \17973 , RIf154130_5416, \9200 );
and \U$8852 ( \17974 , RIe1f4ad8_4161, \9202 );
and \U$8853 ( \17975 , RIf152ab0_5400, \9204 );
and \U$8854 ( \17976 , RIf151700_5386, \9206 );
and \U$8855 ( \17977 , RIf1501e8_5371, \9208 );
and \U$8856 ( \17978 , RIe1f27b0_4136, \9210 );
and \U$8857 ( \17979 , RIfc60ed8_6125, \9212 );
and \U$8858 ( \17980 , RIfc7b620_6426, \9214 );
and \U$8859 ( \17981 , RIf14d7b8_5341, \9216 );
and \U$8860 ( \17982 , RIe1ed4b8_4077, \9218 );
and \U$8861 ( \17983 , RIe1eaa88_4047, \9220 );
and \U$8862 ( \17984 , RIe1e7d88_4015, \9222 );
and \U$8863 ( \17985 , RIe1e5088_3983, \9224 );
and \U$8864 ( \17986 , RIe1e2388_3951, \9226 );
and \U$8865 ( \17987 , RIe1df688_3919, \9228 );
and \U$8866 ( \17988 , RIe1dc988_3887, \9230 );
and \U$8867 ( \17989 , RIe1d9c88_3855, \9232 );
and \U$8868 ( \17990 , RIe1d6f88_3823, \9234 );
and \U$8869 ( \17991 , RIe1d1588_3759, \9236 );
and \U$8870 ( \17992 , RIe1ce888_3727, \9238 );
and \U$8871 ( \17993 , RIe1cbb88_3695, \9240 );
and \U$8872 ( \17994 , RIe1c8e88_3663, \9242 );
and \U$8873 ( \17995 , RIe1c6188_3631, \9244 );
and \U$8874 ( \17996 , RIe1c3488_3599, \9246 );
and \U$8875 ( \17997 , RIe1c0788_3567, \9248 );
and \U$8876 ( \17998 , RIe1bda88_3535, \9250 );
and \U$8877 ( \17999 , RIfca4de0_6898, \9252 );
and \U$8878 ( \18000 , RIfc5ea48_6099, \9254 );
and \U$8879 ( \18001 , RIe1b8a60_3478, \9256 );
and \U$8880 ( \18002 , RIe1b6a08_3455, \9258 );
and \U$8881 ( \18003 , RIfcbd638_7177, \9260 );
and \U$8882 ( \18004 , RIfc44fa8_5807, \9262 );
and \U$8883 ( \18005 , RIfe8e5f0_7964, \9264 );
and \U$8884 ( \18006 , RIfe8e1b8_7961, \9266 );
and \U$8885 ( \18007 , RIf1488f8_5285, \9268 );
and \U$8886 ( \18008 , RIf147818_5273, \9270 );
and \U$8887 ( \18009 , RIfe8e050_7960, \9272 );
and \U$8888 ( \18010 , RIfe8e488_7963, \9274 );
and \U$8889 ( \18011 , RIf146e40_5266, \9276 );
and \U$8890 ( \18012 , RIf146030_5256, \9278 );
and \U$8891 ( \18013 , RIfe8dee8_7959, \9280 );
and \U$8892 ( \18014 , RIfe8e320_7962, \9282 );
and \U$8893 ( \18015 , RIe1a7dc8_3287, \9284 );
and \U$8894 ( \18016 , RIe1a50c8_3255, \9286 );
and \U$8895 ( \18017 , RIe1a23c8_3223, \9288 );
and \U$8896 ( \18018 , RIe19f6c8_3191, \9290 );
and \U$8897 ( \18019 , RIe18bbc8_2967, \9292 );
and \U$8898 ( \18020 , RIe1780c8_2743, \9294 );
and \U$8899 ( \18021 , RIe225a20_4718, \9296 );
and \U$8900 ( \18022 , RIe21a620_4590, \9298 );
and \U$8901 ( \18023 , RIe203e20_4334, \9300 );
and \U$8902 ( \18024 , RIe1fde80_4266, \9302 );
and \U$8903 ( \18025 , RIe1f7238_4189, \9304 );
and \U$8904 ( \18026 , RIe1efd80_4106, \9306 );
and \U$8905 ( \18027 , RIe1d4288_3791, \9308 );
and \U$8906 ( \18028 , RIe1bad88_3503, \9310 );
and \U$8907 ( \18029 , RIe1adc00_3354, \9312 );
and \U$8908 ( \18030 , RIe170238_2653, \9314 );
or \U$8909 ( \18031 , \17967 , \17968 , \17969 , \17970 , \17971 , \17972 , \17973 , \17974 , \17975 , \17976 , \17977 , \17978 , \17979 , \17980 , \17981 , \17982 , \17983 , \17984 , \17985 , \17986 , \17987 , \17988 , \17989 , \17990 , \17991 , \17992 , \17993 , \17994 , \17995 , \17996 , \17997 , \17998 , \17999 , \18000 , \18001 , \18002 , \18003 , \18004 , \18005 , \18006 , \18007 , \18008 , \18009 , \18010 , \18011 , \18012 , \18013 , \18014 , \18015 , \18016 , \18017 , \18018 , \18019 , \18020 , \18021 , \18022 , \18023 , \18024 , \18025 , \18026 , \18027 , \18028 , \18029 , \18030 );
or \U$8910 ( \18032 , \17966 , \18031 );
_DC g659f ( \18033_nG659f , \18032 , \9323 );
and g65a0 ( \18034_nG65a0 , \17901_nG659e , \18033_nG659f );
buf \U$8911 ( \18035 , \18034_nG65a0 );
and \U$8912 ( \18036 , \18035 , \10691 );
nor \U$8913 ( \18037 , \17769 , \18036 );
xnor \U$8914 ( \18038 , \18037 , \10980 );
not \U$8915 ( \18039 , \17656 );
_DC g524f ( \18040_nG524f , \17900 , \9597 );
_DC g52d3 ( \18041_nG52d3 , \18032 , \9323 );
xor g52d4 ( \18042_nG52d4 , \18040_nG524f , \18041_nG52d3 );
buf \U$8916 ( \18043 , \18042_nG52d4 );
and \U$8917 ( \18044 , \17654 , \16622 );
not \U$8918 ( \18045 , \18044 );
and \U$8919 ( \18046 , \18043 , \18045 );
and \U$8920 ( \18047 , \18039 , \18046 );
xor \U$8921 ( \18048 , \18038 , \18047 );
and \U$8922 ( \18049 , \17630 , \17634 );
and \U$8923 ( \18050 , \17634 , \17639 );
and \U$8924 ( \18051 , \17630 , \17639 );
or \U$8925 ( \18052 , \18049 , \18050 , \18051 );
xor \U$8926 ( \18053 , \18048 , \18052 );
and \U$8927 ( \18054 , \17645 , \17649 );
and \U$8928 ( \18055 , \17649 , \17656 );
and \U$8929 ( \18056 , \17645 , \17656 );
or \U$8930 ( \18057 , \18054 , \18055 , \18056 );
xor \U$8931 ( \18058 , \18053 , \18057 );
xor \U$8932 ( \18059 , \17768 , \18058 );
and \U$8933 ( \18060 , \17348 , \17349 );
and \U$8934 ( \18061 , \17349 , \17354 );
and \U$8935 ( \18062 , \17348 , \17354 );
or \U$8936 ( \18063 , \18060 , \18061 , \18062 );
and \U$8937 ( \18064 , \16267 , \11574 );
and \U$8938 ( \18065 , \16655 , \11278 );
nor \U$8939 ( \18066 , \18064 , \18065 );
xnor \U$8940 ( \18067 , \18066 , \11580 );
and \U$8941 ( \18068 , \13679 , \14054 );
and \U$8942 ( \18069 , \14024 , \13692 );
nor \U$8943 ( \18070 , \18068 , \18069 );
xnor \U$8944 ( \18071 , \18070 , \14035 );
xor \U$8945 ( \18072 , \18067 , \18071 );
and \U$8946 ( \18073 , \12448 , \15336 );
and \U$8947 ( \18074 , \12769 , \14963 );
nor \U$8948 ( \18075 , \18073 , \18074 );
xnor \U$8949 ( \18076 , \18075 , \15342 );
xor \U$8950 ( \18077 , \18072 , \18076 );
xor \U$8951 ( \18078 , \18063 , \18077 );
and \U$8952 ( \18079 , \14950 , \12790 );
and \U$8953 ( \18080 , \15321 , \12461 );
nor \U$8954 ( \18081 , \18079 , \18080 );
xnor \U$8955 ( \18082 , \18081 , \12780 );
and \U$8956 ( \18083 , \11270 , \16635 );
and \U$8957 ( \18084 , \11586 , \16301 );
nor \U$8958 ( \18085 , \18083 , \18084 );
xnor \U$8959 ( \18086 , \18085 , \16625 );
xor \U$8960 ( \18087 , \18082 , \18086 );
xor \U$8961 ( \18088 , \18043 , \17654 );
not \U$8962 ( \18089 , \17655 );
and \U$8963 ( \18090 , \18088 , \18089 );
and \U$8964 ( \18091 , \10687 , \18090 );
and \U$8965 ( \18092 , \10988 , \17655 );
nor \U$8966 ( \18093 , \18091 , \18092 );
xnor \U$8967 ( \18094 , \18093 , \18046 );
xor \U$8968 ( \18095 , \18087 , \18094 );
xor \U$8969 ( \18096 , \18078 , \18095 );
xor \U$8970 ( \18097 , \18059 , \18096 );
and \U$8971 ( \18098 , \17344 , \17355 );
and \U$8972 ( \18099 , \17355 , \17658 );
and \U$8973 ( \18100 , \17344 , \17658 );
or \U$8974 ( \18101 , \18098 , \18099 , \18100 );
xor \U$8975 ( \18102 , \18097 , \18101 );
and \U$8976 ( \18103 , \17340 , \17659 );
and \U$8977 ( \18104 , \17660 , \17663 );
or \U$8978 ( \18105 , \18103 , \18104 );
xor \U$8979 ( \18106 , \18102 , \18105 );
buf g9be7 ( \18107_nG9be7 , \18106 );
and \U$8980 ( \18108 , \10704 , \18107_nG9be7 );
or \U$8981 ( \18109 , \17764 , \18108 );
xor \U$8982 ( \18110 , \10703 , \18109 );
buf \U$8983 ( \18111 , \18110 );
buf \U$8985 ( \18112 , \18111 );
xor \U$8986 ( \18113 , \17763 , \18112 );
buf \U$8987 ( \18114 , \18113 );
xor \U$8988 ( \18115 , \17720 , \18114 );
and \U$8989 ( \18116 , \17323 , \17325 );
and \U$8990 ( \18117 , \17323 , \17332 );
and \U$8991 ( \18118 , \17325 , \17332 );
or \U$8992 ( \18119 , \18116 , \18117 , \18118 );
buf \U$8993 ( \18120 , \18119 );
and \U$8994 ( \18121 , \12157 , \14984_nG9bf6 );
and \U$8995 ( \18122 , \12154 , \15373_nG9bf3 );
or \U$8996 ( \18123 , \18121 , \18122 );
xor \U$8997 ( \18124 , \12153 , \18123 );
buf \U$8998 ( \18125 , \18124 );
buf \U$9000 ( \18126 , \18125 );
xor \U$9001 ( \18127 , \18120 , \18126 );
and \U$9002 ( \18128 , \10421 , \16315_nG9bf0 );
and \U$9003 ( \18129 , \10418 , \16680_nG9bed );
or \U$9004 ( \18130 , \18128 , \18129 );
xor \U$9005 ( \18131 , \10417 , \18130 );
buf \U$9006 ( \18132 , \18131 );
buf \U$9008 ( \18133 , \18132 );
xor \U$9009 ( \18134 , \18127 , \18133 );
buf \U$9010 ( \18135 , \18134 );
xor \U$9011 ( \18136 , \18115 , \18135 );
buf \U$9012 ( \18137 , \18136 );
and \U$9013 ( \18138 , \17672 , \17677 );
and \U$9014 ( \18139 , \17672 , \17698 );
and \U$9015 ( \18140 , \17677 , \17698 );
or \U$9016 ( \18141 , \18138 , \18139 , \18140 );
buf \U$9017 ( \18142 , \18141 );
xor \U$9018 ( \18143 , \18137 , \18142 );
and \U$9019 ( \18144 , \17700 , \17705 );
and \U$9020 ( \18145 , \17700 , \17711 );
and \U$9021 ( \18146 , \17705 , \17711 );
or \U$9022 ( \18147 , \18144 , \18145 , \18146 );
buf \U$9023 ( \18148 , \18147 );
xor \U$9024 ( \18149 , \18143 , \18148 );
and \U$9025 ( \18150 , \17715 , \18149 );
and \U$9026 ( \18151 , RIdec4a00_701, \9059 );
and \U$9027 ( \18152 , RIdec1d00_669, \9061 );
and \U$9028 ( \18153 , RIfcad7b0_6996, \9063 );
and \U$9029 ( \18154 , RIdebf000_637, \9065 );
and \U$9030 ( \18155 , RIfc64cb8_6169, \9067 );
and \U$9031 ( \18156 , RIdebc300_605, \9069 );
and \U$9032 ( \18157 , RIdeb9600_573, \9071 );
and \U$9033 ( \18158 , RIdeb6900_541, \9073 );
and \U$9034 ( \18159 , RIfc6f9b0_6292, \9075 );
and \U$9035 ( \18160 , RIdeb0f00_477, \9077 );
and \U$9036 ( \18161 , RIfc657f8_6177, \9079 );
and \U$9037 ( \18162 , RIdeae200_445, \9081 );
and \U$9038 ( \18163 , RIfce69c0_7646, \9083 );
and \U$9039 ( \18164 , RIdea8d28_413, \9085 );
and \U$9040 ( \18165 , RIdea2428_381, \9087 );
and \U$9041 ( \18166 , RIde9bb28_349, \9089 );
and \U$9042 ( \18167 , RIfc6fc80_6294, \9091 );
and \U$9043 ( \18168 , RIee1b760_4771, \9093 );
and \U$9044 ( \18169 , RIfca8080_6934, \9095 );
and \U$9045 ( \18170 , RIfe8b8f0_7932, \9097 );
and \U$9046 ( \18171 , RIde90020_292, \9099 );
and \U$9047 ( \18172 , RIde8c510_274, \9101 );
and \U$9048 ( \18173 , RIde89090_258, \9103 );
and \U$9049 ( \18174 , RIde84ba8_237, \9105 );
and \U$9050 ( \18175 , RIfc65ac8_6179, \9107 );
and \U$9051 ( \18176 , RIfcad210_6992, \9109 );
and \U$9052 ( \18177 , RIfcce168_7367, \9111 );
and \U$9053 ( \18178 , RIfcce2d0_7368, \9113 );
and \U$9054 ( \18179 , RIfc51488_5947, \9115 );
and \U$9055 ( \18180 , RIe16af40_2594, \9117 );
and \U$9056 ( \18181 , RIfc65c30_6180, \9119 );
and \U$9057 ( \18182 , RIe167598_2553, \9121 );
and \U$9058 ( \18183 , RIe164a00_2522, \9123 );
and \U$9059 ( \18184 , RIe161d00_2490, \9125 );
and \U$9060 ( \18185 , RIfc66e78_6193, \9127 );
and \U$9061 ( \18186 , RIe15f000_2458, \9129 );
and \U$9062 ( \18187 , RIfc6e498_6277, \9131 );
and \U$9063 ( \18188 , RIe15c300_2426, \9133 );
and \U$9064 ( \18189 , RIe156900_2362, \9135 );
and \U$9065 ( \18190 , RIe153c00_2330, \9137 );
and \U$9066 ( \18191 , RIfc6e330_6276, \9139 );
and \U$9067 ( \18192 , RIe150f00_2298, \9141 );
and \U$9068 ( \18193 , RIfccda60_7362, \9143 );
and \U$9069 ( \18194 , RIe14e200_2266, \9145 );
and \U$9070 ( \18195 , RIfc6e1c8_6275, \9147 );
and \U$9071 ( \18196 , RIe14b500_2234, \9149 );
and \U$9072 ( \18197 , RIe148800_2202, \9151 );
and \U$9073 ( \18198 , RIe145b00_2170, \9153 );
and \U$9074 ( \18199 , RIee33fb8_5050, \9155 );
and \U$9075 ( \18200 , RIee32d70_5037, \9157 );
and \U$9076 ( \18201 , RIee31c90_5025, \9159 );
and \U$9077 ( \18202 , RIee30fe8_5016, \9161 );
and \U$9078 ( \18203 , RIfea8630_8232, \9163 );
and \U$9079 ( \18204 , RIdf3e5a8_2086, \9165 );
and \U$9080 ( \18205 , RIdf3c550_2063, \9167 );
and \U$9081 ( \18206 , RIfea8798_8233, \9169 );
and \U$9082 ( \18207 , RIfc6e060_6274, \9171 );
and \U$9083 ( \18208 , RIfcac6d0_6984, \9173 );
and \U$9084 ( \18209 , RIfc56078_6001, \9175 );
and \U$9085 ( \18210 , RIfc6e600_6278, \9177 );
and \U$9086 ( \18211 , RIdf34dc8_1978, \9179 );
and \U$9087 ( \18212 , RIdf32d70_1955, \9181 );
and \U$9088 ( \18213 , RIfea84c8_8231, \9183 );
and \U$9089 ( \18214 , RIdf2eb58_1908, \9185 );
or \U$9090 ( \18215 , \18151 , \18152 , \18153 , \18154 , \18155 , \18156 , \18157 , \18158 , \18159 , \18160 , \18161 , \18162 , \18163 , \18164 , \18165 , \18166 , \18167 , \18168 , \18169 , \18170 , \18171 , \18172 , \18173 , \18174 , \18175 , \18176 , \18177 , \18178 , \18179 , \18180 , \18181 , \18182 , \18183 , \18184 , \18185 , \18186 , \18187 , \18188 , \18189 , \18190 , \18191 , \18192 , \18193 , \18194 , \18195 , \18196 , \18197 , \18198 , \18199 , \18200 , \18201 , \18202 , \18203 , \18204 , \18205 , \18206 , \18207 , \18208 , \18209 , \18210 , \18211 , \18212 , \18213 , \18214 );
and \U$9091 ( \18216 , RIee2b750_4953, \9188 );
and \U$9092 ( \18217 , RIfc6ee70_6284, \9190 );
and \U$9093 ( \18218 , RIfc6efd8_6285, \9192 );
and \U$9094 ( \18219 , RIee27808_4908, \9194 );
and \U$9095 ( \18220 , RIfe8b788_7931, \9196 );
and \U$9096 ( \18221 , RIdf27ad8_1828, \9198 );
and \U$9097 ( \18222 , RIdf25d50_1807, \9200 );
and \U$9098 ( \18223 , RIdf24130_1787, \9202 );
and \U$9099 ( \18224 , RIfc66608_6187, \9204 );
and \U$9100 ( \18225 , RIfccde98_7365, \9206 );
and \U$9101 ( \18226 , RIfc66a40_6190, \9208 );
and \U$9102 ( \18227 , RIfc668d8_6189, \9210 );
and \U$9103 ( \18228 , RIfcacf40_6990, \9212 );
and \U$9104 ( \18229 , RIfeaaef8_8261, \9214 );
and \U$9105 ( \18230 , RIfc6e8d0_6280, \9216 );
and \U$9106 ( \18231 , RIdf18d30_1659, \9218 );
and \U$9107 ( \18232 , RIdf165d0_1631, \9220 );
and \U$9108 ( \18233 , RIdf138d0_1599, \9222 );
and \U$9109 ( \18234 , RIdf10bd0_1567, \9224 );
and \U$9110 ( \18235 , RIdf0ded0_1535, \9226 );
and \U$9111 ( \18236 , RIdf0b1d0_1503, \9228 );
and \U$9112 ( \18237 , RIdf084d0_1471, \9230 );
and \U$9113 ( \18238 , RIdf057d0_1439, \9232 );
and \U$9114 ( \18239 , RIdf02ad0_1407, \9234 );
and \U$9115 ( \18240 , RIdefd0d0_1343, \9236 );
and \U$9116 ( \18241 , RIdefa3d0_1311, \9238 );
and \U$9117 ( \18242 , RIdef76d0_1279, \9240 );
and \U$9118 ( \18243 , RIdef49d0_1247, \9242 );
and \U$9119 ( \18244 , RIdef1cd0_1215, \9244 );
and \U$9120 ( \18245 , RIdeeefd0_1183, \9246 );
and \U$9121 ( \18246 , RIdeec2d0_1151, \9248 );
and \U$9122 ( \18247 , RIdee95d0_1119, \9250 );
and \U$9123 ( \18248 , RIfc6dc28_6271, \9252 );
and \U$9124 ( \18249 , RIfc67c88_6203, \9254 );
and \U$9125 ( \18250 , RIfccb300_7334, \9256 );
and \U$9126 ( \18251 , RIfccd4c0_7358, \9258 );
and \U$9127 ( \18252 , RIfea81f8_8229, \9260 );
and \U$9128 ( \18253 , RIfea8360_8230, \9262 );
and \U$9129 ( \18254 , RIdee04f8_1016, \9264 );
and \U$9130 ( \18255 , RIdede338_992, \9266 );
and \U$9131 ( \18256 , RIfc6def8_6273, \9268 );
and \U$9132 ( \18257 , RIfcac130_6980, \9270 );
and \U$9133 ( \18258 , RIfc67b20_6202, \9272 );
and \U$9134 ( \18259 , RIfc67df0_6204, \9274 );
and \U$9135 ( \18260 , RIded9040_933, \9276 );
and \U$9136 ( \18261 , RIded6a48_906, \9278 );
and \U$9137 ( \18262 , RIded4b58_884, \9280 );
and \U$9138 ( \18263 , RIded26c8_858, \9282 );
and \U$9139 ( \18264 , RIdecfe00_829, \9284 );
and \U$9140 ( \18265 , RIdecd100_797, \9286 );
and \U$9141 ( \18266 , RIdeca400_765, \9288 );
and \U$9142 ( \18267 , RIdec7700_733, \9290 );
and \U$9143 ( \18268 , RIdeb3c00_509, \9292 );
and \U$9144 ( \18269 , RIde95228_317, \9294 );
and \U$9145 ( \18270 , RIe16d808_2623, \9296 );
and \U$9146 ( \18271 , RIe159600_2394, \9298 );
and \U$9147 ( \18272 , RIe142e00_2138, \9300 );
and \U$9148 ( \18273 , RIdf377f8_2008, \9302 );
and \U$9149 ( \18274 , RIdf2be58_1876, \9304 );
and \U$9150 ( \18275 , RIdf1c6d8_1700, \9306 );
and \U$9151 ( \18276 , RIdeffdd0_1375, \9308 );
and \U$9152 ( \18277 , RIdee68d0_1087, \9310 );
and \U$9153 ( \18278 , RIdedb638_960, \9312 );
and \U$9154 ( \18279 , RIde7b170_190, \9314 );
or \U$9155 ( \18280 , \18216 , \18217 , \18218 , \18219 , \18220 , \18221 , \18222 , \18223 , \18224 , \18225 , \18226 , \18227 , \18228 , \18229 , \18230 , \18231 , \18232 , \18233 , \18234 , \18235 , \18236 , \18237 , \18238 , \18239 , \18240 , \18241 , \18242 , \18243 , \18244 , \18245 , \18246 , \18247 , \18248 , \18249 , \18250 , \18251 , \18252 , \18253 , \18254 , \18255 , \18256 , \18257 , \18258 , \18259 , \18260 , \18261 , \18262 , \18263 , \18264 , \18265 , \18266 , \18267 , \18268 , \18269 , \18270 , \18271 , \18272 , \18273 , \18274 , \18275 , \18276 , \18277 , \18278 , \18279 );
or \U$9156 ( \18281 , \18215 , \18280 );
_DC g2a85 ( \18282_nG2a85 , \18281 , \9323 );
buf \U$9157 ( \18283 , \18282_nG2a85 );
and \U$9158 ( \18284 , RIe19cc98_3161, \9333 );
and \U$9159 ( \18285 , RIe199f98_3129, \9335 );
and \U$9160 ( \18286 , RIfc73088_6331, \9337 );
and \U$9161 ( \18287 , RIe197298_3097, \9339 );
and \U$9162 ( \18288 , RIf1442a8_5235, \9341 );
and \U$9163 ( \18289 , RIe194598_3065, \9343 );
and \U$9164 ( \18290 , RIe191898_3033, \9345 );
and \U$9165 ( \18291 , RIe18eb98_3001, \9347 );
and \U$9166 ( \18292 , RIe189198_2937, \9349 );
and \U$9167 ( \18293 , RIe186498_2905, \9351 );
and \U$9168 ( \18294 , RIfc72278_6321, \9353 );
and \U$9169 ( \18295 , RIe183798_2873, \9355 );
and \U$9170 ( \18296 , RIfc61ce8_6135, \9357 );
and \U$9171 ( \18297 , RIe180a98_2841, \9359 );
and \U$9172 ( \18298 , RIe17dd98_2809, \9361 );
and \U$9173 ( \18299 , RIe17b098_2777, \9363 );
and \U$9174 ( \18300 , RIfcaf268_7015, \9365 );
and \U$9175 ( \18301 , RIfca6a00_6918, \9367 );
and \U$9176 ( \18302 , RIfcc9b18_7317, \9369 );
and \U$9177 ( \18303 , RIe175530_2712, \9371 );
and \U$9178 ( \18304 , RIfc72818_6325, \9373 );
and \U$9179 ( \18305 , RIfc726b0_6324, \9375 );
and \U$9180 ( \18306 , RIfccf7e8_7383, \9377 );
and \U$9181 ( \18307 , RIfc72548_6323, \9379 );
and \U$9182 ( \18308 , RIee3be48_5140, \9381 );
and \U$9183 ( \18309 , RIee3ad68_5128, \9383 );
and \U$9184 ( \18310 , RIfc71fa8_6319, \9385 );
and \U$9185 ( \18311 , RIe1730a0_2686, \9387 );
and \U$9186 ( \18312 , RIfcaef98_7013, \9389 );
and \U$9187 ( \18313 , RIfccf518_7381, \9391 );
and \U$9188 ( \18314 , RIfc71e40_6318, \9393 );
and \U$9189 ( \18315 , RIfc62120_6138, \9395 );
and \U$9190 ( \18316 , RIfe8b350_7928, \9397 );
and \U$9191 ( \18317 , RIe222ff0_4688, \9399 );
and \U$9192 ( \18318 , RIfcc9f50_7320, \9401 );
and \U$9193 ( \18319 , RIe2202f0_4656, \9403 );
and \U$9194 ( \18320 , RIfc4a570_5868, \9405 );
and \U$9195 ( \18321 , RIe21d5f0_4624, \9407 );
and \U$9196 ( \18322 , RIe217bf0_4560, \9409 );
and \U$9197 ( \18323 , RIe214ef0_4528, \9411 );
and \U$9198 ( \18324 , RIfccf3b0_7380, \9413 );
and \U$9199 ( \18325 , RIe2121f0_4496, \9415 );
and \U$9200 ( \18326 , RIf168ba8_5651, \9417 );
and \U$9201 ( \18327 , RIe20f4f0_4464, \9419 );
and \U$9202 ( \18328 , RIfc71300_6310, \9421 );
and \U$9203 ( \18329 , RIe20c7f0_4432, \9423 );
and \U$9204 ( \18330 , RIe209af0_4400, \9425 );
and \U$9205 ( \18331 , RIe206df0_4368, \9427 );
and \U$9206 ( \18332 , RIfc718a0_6314, \9429 );
and \U$9207 ( \18333 , RIfc71a08_6315, \9431 );
and \U$9208 ( \18334 , RIe202098_4313, \9433 );
and \U$9209 ( \18335 , RIfe8b1e8_7927, \9435 );
and \U$9210 ( \18336 , RIfc715d0_6312, \9437 );
and \U$9211 ( \18337 , RIfce6588_7643, \9439 );
and \U$9212 ( \18338 , RIfc62c60_6146, \9441 );
and \U$9213 ( \18339 , RIf161858_5569, \9443 );
and \U$9214 ( \18340 , RIf15fad0_5548, \9445 );
and \U$9215 ( \18341 , RIf15dbe0_5526, \9447 );
and \U$9216 ( \18342 , RIe1fc698_4249, \9449 );
and \U$9217 ( \18343 , RIfe8b4b8_7929, \9451 );
and \U$9218 ( \18344 , RIfcae5c0_7006, \9453 );
and \U$9219 ( \18345 , RIfc63098_6149, \9455 );
and \U$9220 ( \18346 , RIfc63200_6150, \9457 );
and \U$9221 ( \18347 , RIfc71198_6309, \9459 );
or \U$9222 ( \18348 , \18284 , \18285 , \18286 , \18287 , \18288 , \18289 , \18290 , \18291 , \18292 , \18293 , \18294 , \18295 , \18296 , \18297 , \18298 , \18299 , \18300 , \18301 , \18302 , \18303 , \18304 , \18305 , \18306 , \18307 , \18308 , \18309 , \18310 , \18311 , \18312 , \18313 , \18314 , \18315 , \18316 , \18317 , \18318 , \18319 , \18320 , \18321 , \18322 , \18323 , \18324 , \18325 , \18326 , \18327 , \18328 , \18329 , \18330 , \18331 , \18332 , \18333 , \18334 , \18335 , \18336 , \18337 , \18338 , \18339 , \18340 , \18341 , \18342 , \18343 , \18344 , \18345 , \18346 , \18347 );
and \U$9223 ( \18349 , RIf158a50_5468, \9462 );
and \U$9224 ( \18350 , RIf1576a0_5454, \9464 );
and \U$9225 ( \18351 , RIfcdc808_7531, \9466 );
and \U$9226 ( \18352 , RIfe8b620_7930, \9468 );
and \U$9227 ( \18353 , RIfc634d0_6152, \9470 );
and \U$9228 ( \18354 , RIfcceb40_7374, \9472 );
and \U$9229 ( \18355 , RIf154400_5418, \9474 );
and \U$9230 ( \18356 , RIe1f4da8_4163, \9476 );
and \U$9231 ( \18357 , RIf152c18_5401, \9478 );
and \U$9232 ( \18358 , RIf151868_5387, \9480 );
and \U$9233 ( \18359 , RIfc4d108_5899, \9482 );
and \U$9234 ( \18360 , RIe1f2a80_4138, \9484 );
and \U$9235 ( \18361 , RIfc70a90_6304, \9486 );
and \U$9236 ( \18362 , RIfc63bd8_6157, \9488 );
and \U$9237 ( \18363 , RIfca7810_6928, \9490 );
and \U$9238 ( \18364 , RIe1ed788_4079, \9492 );
and \U$9239 ( \18365 , RIe1ead58_4049, \9494 );
and \U$9240 ( \18366 , RIe1e8058_4017, \9496 );
and \U$9241 ( \18367 , RIe1e5358_3985, \9498 );
and \U$9242 ( \18368 , RIe1e2658_3953, \9500 );
and \U$9243 ( \18369 , RIe1df958_3921, \9502 );
and \U$9244 ( \18370 , RIe1dcc58_3889, \9504 );
and \U$9245 ( \18371 , RIe1d9f58_3857, \9506 );
and \U$9246 ( \18372 , RIe1d7258_3825, \9508 );
and \U$9247 ( \18373 , RIe1d1858_3761, \9510 );
and \U$9248 ( \18374 , RIe1ceb58_3729, \9512 );
and \U$9249 ( \18375 , RIe1cbe58_3697, \9514 );
and \U$9250 ( \18376 , RIe1c9158_3665, \9516 );
and \U$9251 ( \18377 , RIe1c6458_3633, \9518 );
and \U$9252 ( \18378 , RIe1c3758_3601, \9520 );
and \U$9253 ( \18379 , RIe1c0a58_3569, \9522 );
and \U$9254 ( \18380 , RIe1bdd58_3537, \9524 );
and \U$9255 ( \18381 , RIf14c408_5327, \9526 );
and \U$9256 ( \18382 , RIf14b1c0_5314, \9528 );
and \U$9257 ( \18383 , RIe1b8d30_3480, \9530 );
and \U$9258 ( \18384 , RIe1b6cd8_3457, \9532 );
and \U$9259 ( \18385 , RIfc707c0_6302, \9534 );
and \U$9260 ( \18386 , RIfca7c48_6931, \9536 );
and \U$9261 ( \18387 , RIe1b4de8_3435, \9538 );
and \U$9262 ( \18388 , RIe1b3a38_3421, \9540 );
and \U$9263 ( \18389 , RIfc70220_6298, \9542 );
and \U$9264 ( \18390 , RIfcce870_7372, \9544 );
and \U$9265 ( \18391 , RIe1b23b8_3405, \9546 );
and \U$9266 ( \18392 , RIe1b0630_3384, \9548 );
and \U$9267 ( \18393 , RIfc645b0_6164, \9550 );
and \U$9268 ( \18394 , RIfc700b8_6297, \9552 );
and \U$9269 ( \18395 , RIfeaac28_8259, \9554 );
and \U$9270 ( \18396 , RIe1aa690_3316, \9556 );
and \U$9271 ( \18397 , RIe1a8098_3289, \9558 );
and \U$9272 ( \18398 , RIe1a5398_3257, \9560 );
and \U$9273 ( \18399 , RIe1a2698_3225, \9562 );
and \U$9274 ( \18400 , RIe19f998_3193, \9564 );
and \U$9275 ( \18401 , RIe18be98_2969, \9566 );
and \U$9276 ( \18402 , RIe178398_2745, \9568 );
and \U$9277 ( \18403 , RIe225cf0_4720, \9570 );
and \U$9278 ( \18404 , RIe21a8f0_4592, \9572 );
and \U$9279 ( \18405 , RIe2040f0_4336, \9574 );
and \U$9280 ( \18406 , RIe1fe150_4268, \9576 );
and \U$9281 ( \18407 , RIe1f7508_4191, \9578 );
and \U$9282 ( \18408 , RIe1f0050_4108, \9580 );
and \U$9283 ( \18409 , RIe1d4558_3793, \9582 );
and \U$9284 ( \18410 , RIe1bb058_3505, \9584 );
and \U$9285 ( \18411 , RIe1aded0_3356, \9586 );
and \U$9286 ( \18412 , RIe170508_2655, \9588 );
or \U$9287 ( \18413 , \18349 , \18350 , \18351 , \18352 , \18353 , \18354 , \18355 , \18356 , \18357 , \18358 , \18359 , \18360 , \18361 , \18362 , \18363 , \18364 , \18365 , \18366 , \18367 , \18368 , \18369 , \18370 , \18371 , \18372 , \18373 , \18374 , \18375 , \18376 , \18377 , \18378 , \18379 , \18380 , \18381 , \18382 , \18383 , \18384 , \18385 , \18386 , \18387 , \18388 , \18389 , \18390 , \18391 , \18392 , \18393 , \18394 , \18395 , \18396 , \18397 , \18398 , \18399 , \18400 , \18401 , \18402 , \18403 , \18404 , \18405 , \18406 , \18407 , \18408 , \18409 , \18410 , \18411 , \18412 );
or \U$9288 ( \18414 , \18348 , \18413 );
_DC g3bb2 ( \18415_nG3bb2 , \18414 , \9597 );
buf \U$9289 ( \18416 , \18415_nG3bb2 );
xor \U$9290 ( \18417 , \18283 , \18416 );
and \U$9291 ( \18418 , RIdec4898_700, \9059 );
and \U$9292 ( \18419 , RIdec1b98_668, \9061 );
and \U$9293 ( \18420 , RIfc661d0_6184, \9063 );
and \U$9294 ( \18421 , RIdebee98_636, \9065 );
and \U$9295 ( \18422 , RIfce6b28_7647, \9067 );
and \U$9296 ( \18423 , RIdebc198_604, \9069 );
and \U$9297 ( \18424 , RIdeb9498_572, \9071 );
and \U$9298 ( \18425 , RIdeb6798_540, \9073 );
and \U$9299 ( \18426 , RIfc40d18_5763, \9075 );
and \U$9300 ( \18427 , RIdeb0d98_476, \9077 );
and \U$9301 ( \18428 , RIfcad648_6995, \9079 );
and \U$9302 ( \18429 , RIdeae098_444, \9081 );
and \U$9303 ( \18430 , RIfcaa510_6960, \9083 );
and \U$9304 ( \18431 , RIdea89e0_412, \9085 );
and \U$9305 ( \18432 , RIdea20e0_380, \9087 );
and \U$9306 ( \18433 , RIde9b7e0_348, \9089 );
and \U$9307 ( \18434 , RIfcab320_6970, \9091 );
and \U$9308 ( \18435 , RIfca8350_6936, \9093 );
and \U$9309 ( \18436 , RIfc6f6e0_6290, \9095 );
and \U$9310 ( \18437 , RIfcaa240_6958, \9097 );
and \U$9311 ( \18438 , RIde8fcd8_291, \9099 );
and \U$9312 ( \18439 , RIfe8aae0_7922, \9101 );
and \U$9313 ( \18440 , RIde88d48_257, \9103 );
and \U$9314 ( \18441 , RIde84860_236, \9105 );
and \U$9315 ( \18442 , RIde80a08_217, \9107 );
and \U$9316 ( \18443 , RIfc64718_6165, \9109 );
and \U$9317 ( \18444 , RIfcae020_7002, \9111 );
and \U$9318 ( \18445 , RIfcadeb8_7001, \9113 );
and \U$9319 ( \18446 , RIee38fe0_5107, \9115 );
and \U$9320 ( \18447 , RIe16add8_2593, \9117 );
and \U$9321 ( \18448 , RIe1695f0_2576, \9119 );
and \U$9322 ( \18449 , RIe167430_2552, \9121 );
and \U$9323 ( \18450 , RIe164898_2521, \9123 );
and \U$9324 ( \18451 , RIe161b98_2489, \9125 );
and \U$9325 ( \18452 , RIfe8a3d8_7917, \9127 );
and \U$9326 ( \18453 , RIe15ee98_2457, \9129 );
and \U$9327 ( \18454 , RIfe8a270_7916, \9131 );
and \U$9328 ( \18455 , RIe15c198_2425, \9133 );
and \U$9329 ( \18456 , RIe156798_2361, \9135 );
and \U$9330 ( \18457 , RIe153a98_2329, \9137 );
and \U$9331 ( \18458 , RIfc3f0f8_5743, \9139 );
and \U$9332 ( \18459 , RIe150d98_2297, \9141 );
and \U$9333 ( \18460 , RIfcab050_6968, \9143 );
and \U$9334 ( \18461 , RIe14e098_2265, \9145 );
and \U$9335 ( \18462 , RIfcca658_7325, \9147 );
and \U$9336 ( \18463 , RIe14b398_2233, \9149 );
and \U$9337 ( \18464 , RIe148698_2201, \9151 );
and \U$9338 ( \18465 , RIe145998_2169, \9153 );
and \U$9339 ( \18466 , RIfe8a810_7920, \9155 );
and \U$9340 ( \18467 , RIfe8a6a8_7919, \9157 );
and \U$9341 ( \18468 , RIee31b28_5024, \9159 );
and \U$9342 ( \18469 , RIee30e80_5015, \9161 );
and \U$9343 ( \18470 , RIe140808_2111, \9163 );
and \U$9344 ( \18471 , RIfe8a540_7918, \9165 );
and \U$9345 ( \18472 , RIdf3c3e8_2062, \9167 );
and \U$9346 ( \18473 , RIdf3a0c0_2037, \9169 );
and \U$9347 ( \18474 , RIfc6b1f8_6241, \9171 );
and \U$9348 ( \18475 , RIee2f260_4995, \9173 );
and \U$9349 ( \18476 , RIfc70d60_6306, \9175 );
and \U$9350 ( \18477 , RIee2d0a0_4971, \9177 );
and \U$9351 ( \18478 , RIfe8a978_7921, \9179 );
and \U$9352 ( \18479 , RIdf32c08_1954, \9181 );
and \U$9353 ( \18480 , RIdf308e0_1929, \9183 );
and \U$9354 ( \18481 , RIdf2e9f0_1907, \9185 );
or \U$9355 ( \18482 , \18418 , \18419 , \18420 , \18421 , \18422 , \18423 , \18424 , \18425 , \18426 , \18427 , \18428 , \18429 , \18430 , \18431 , \18432 , \18433 , \18434 , \18435 , \18436 , \18437 , \18438 , \18439 , \18440 , \18441 , \18442 , \18443 , \18444 , \18445 , \18446 , \18447 , \18448 , \18449 , \18450 , \18451 , \18452 , \18453 , \18454 , \18455 , \18456 , \18457 , \18458 , \18459 , \18460 , \18461 , \18462 , \18463 , \18464 , \18465 , \18466 , \18467 , \18468 , \18469 , \18470 , \18471 , \18472 , \18473 , \18474 , \18475 , \18476 , \18477 , \18478 , \18479 , \18480 , \18481 );
and \U$9356 ( \18483 , RIee2b5e8_4952, \9188 );
and \U$9357 ( \18484 , RIee29e00_4935, \9190 );
and \U$9358 ( \18485 , RIee28a50_4921, \9192 );
and \U$9359 ( \18486 , RIee276a0_4907, \9194 );
and \U$9360 ( \18487 , RIdf29c98_1852, \9196 );
and \U$9361 ( \18488 , RIdf27970_1827, \9198 );
and \U$9362 ( \18489 , RIdf25be8_1806, \9200 );
and \U$9363 ( \18490 , RIdf23fc8_1786, \9202 );
and \U$9364 ( \18491 , RIfc6aaf0_6236, \9204 );
and \U$9365 ( \18492 , RIfc6ac58_6237, \9206 );
and \U$9366 ( \18493 , RIdf22678_1768, \9208 );
and \U$9367 ( \18494 , RIfcdd4b0_7540, \9210 );
and \U$9368 ( \18495 , RIdf21160_1753, \9212 );
and \U$9369 ( \18496 , RIdf1f108_1730, \9214 );
and \U$9370 ( \18497 , RIdf1ac20_1681, \9216 );
and \U$9371 ( \18498 , RIfeaa7f0_8256, \9218 );
and \U$9372 ( \18499 , RIdf16468_1630, \9220 );
and \U$9373 ( \18500 , RIdf13768_1598, \9222 );
and \U$9374 ( \18501 , RIdf10a68_1566, \9224 );
and \U$9375 ( \18502 , RIdf0dd68_1534, \9226 );
and \U$9376 ( \18503 , RIdf0b068_1502, \9228 );
and \U$9377 ( \18504 , RIdf08368_1470, \9230 );
and \U$9378 ( \18505 , RIdf05668_1438, \9232 );
and \U$9379 ( \18506 , RIdf02968_1406, \9234 );
and \U$9380 ( \18507 , RIdefcf68_1342, \9236 );
and \U$9381 ( \18508 , RIdefa268_1310, \9238 );
and \U$9382 ( \18509 , RIdef7568_1278, \9240 );
and \U$9383 ( \18510 , RIdef4868_1246, \9242 );
and \U$9384 ( \18511 , RIdef1b68_1214, \9244 );
and \U$9385 ( \18512 , RIdeeee68_1182, \9246 );
and \U$9386 ( \18513 , RIdeec168_1150, \9248 );
and \U$9387 ( \18514 , RIdee9468_1118, \9250 );
and \U$9388 ( \18515 , RIee25378_4882, \9252 );
and \U$9389 ( \18516 , RIee24568_4872, \9254 );
and \U$9390 ( \18517 , RIee23a28_4864, \9256 );
and \U$9391 ( \18518 , RIee23050_4857, \9258 );
and \U$9392 ( \18519 , RIfe8adb0_7924, \9260 );
and \U$9393 ( \18520 , RIdee23e8_1038, \9262 );
and \U$9394 ( \18521 , RIfe8ac48_7923, \9264 );
and \U$9395 ( \18522 , RIdede1d0_991, \9266 );
and \U$9396 ( \18523 , RIfca5650_6904, \9268 );
and \U$9397 ( \18524 , RIee220d8_4846, \9270 );
and \U$9398 ( \18525 , RIfceeb20_7738, \9272 );
and \U$9399 ( \18526 , RIee20ff8_4834, \9274 );
and \U$9400 ( \18527 , RIded8ed8_932, \9276 );
and \U$9401 ( \18528 , RIfe8af18_7925, \9278 );
and \U$9402 ( \18529 , RIded49f0_883, \9280 );
and \U$9403 ( \18530 , RIfe8b080_7926, \9282 );
and \U$9404 ( \18531 , RIdecfc98_828, \9284 );
and \U$9405 ( \18532 , RIdeccf98_796, \9286 );
and \U$9406 ( \18533 , RIdeca298_764, \9288 );
and \U$9407 ( \18534 , RIdec7598_732, \9290 );
and \U$9408 ( \18535 , RIdeb3a98_508, \9292 );
and \U$9409 ( \18536 , RIde94ee0_316, \9294 );
and \U$9410 ( \18537 , RIe16d6a0_2622, \9296 );
and \U$9411 ( \18538 , RIe159498_2393, \9298 );
and \U$9412 ( \18539 , RIe142c98_2137, \9300 );
and \U$9413 ( \18540 , RIdf37690_2007, \9302 );
and \U$9414 ( \18541 , RIdf2bcf0_1875, \9304 );
and \U$9415 ( \18542 , RIdf1c570_1699, \9306 );
and \U$9416 ( \18543 , RIdeffc68_1374, \9308 );
and \U$9417 ( \18544 , RIdee6768_1086, \9310 );
and \U$9418 ( \18545 , RIdedb4d0_959, \9312 );
and \U$9419 ( \18546 , RIde7ae28_189, \9314 );
or \U$9420 ( \18547 , \18483 , \18484 , \18485 , \18486 , \18487 , \18488 , \18489 , \18490 , \18491 , \18492 , \18493 , \18494 , \18495 , \18496 , \18497 , \18498 , \18499 , \18500 , \18501 , \18502 , \18503 , \18504 , \18505 , \18506 , \18507 , \18508 , \18509 , \18510 , \18511 , \18512 , \18513 , \18514 , \18515 , \18516 , \18517 , \18518 , \18519 , \18520 , \18521 , \18522 , \18523 , \18524 , \18525 , \18526 , \18527 , \18528 , \18529 , \18530 , \18531 , \18532 , \18533 , \18534 , \18535 , \18536 , \18537 , \18538 , \18539 , \18540 , \18541 , \18542 , \18543 , \18544 , \18545 , \18546 );
or \U$9421 ( \18548 , \18482 , \18547 );
_DC g2b0a ( \18549_nG2b0a , \18548 , \9323 );
buf \U$9422 ( \18550 , \18549_nG2b0a );
and \U$9423 ( \18551 , RIe19cb30_3160, \9333 );
and \U$9424 ( \18552 , RIe199e30_3128, \9335 );
and \U$9425 ( \18553 , RIf145388_5247, \9337 );
and \U$9426 ( \18554 , RIe197130_3096, \9339 );
and \U$9427 ( \18555 , RIfe8a108_7915, \9341 );
and \U$9428 ( \18556 , RIe194430_3064, \9343 );
and \U$9429 ( \18557 , RIe191730_3032, \9345 );
and \U$9430 ( \18558 , RIe18ea30_3000, \9347 );
and \U$9431 ( \18559 , RIe189030_2936, \9349 );
and \U$9432 ( \18560 , RIe186330_2904, \9351 );
and \U$9433 ( \18561 , RIfc6c878_6257, \9353 );
and \U$9434 ( \18562 , RIe183630_2872, \9355 );
and \U$9435 ( \18563 , RIfcabcf8_6977, \9357 );
and \U$9436 ( \18564 , RIe180930_2840, \9359 );
and \U$9437 ( \18565 , RIe17dc30_2808, \9361 );
and \U$9438 ( \18566 , RIe17af30_2776, \9363 );
and \U$9439 ( \18567 , RIfcccc50_7352, \9365 );
and \U$9440 ( \18568 , RIfcccdb8_7353, \9367 );
and \U$9441 ( \18569 , RIe176d18_2729, \9369 );
and \U$9442 ( \18570 , RIfea7af0_8224, \9371 );
and \U$9443 ( \18571 , RIfe89fa0_7914, \9373 );
and \U$9444 ( \18572 , RIfe89e38_7913, \9375 );
and \U$9445 ( \18573 , RIfcdd078_7537, \9377 );
and \U$9446 ( \18574 , RIfccb738_7337, \9379 );
and \U$9447 ( \18575 , RIfca9868_6951, \9381 );
and \U$9448 ( \18576 , RIfcabb90_6976, \9383 );
and \U$9449 ( \18577 , RIfca99d0_6952, \9385 );
and \U$9450 ( \18578 , RIe172f38_2685, \9387 );
and \U$9451 ( \18579 , RIf16fd90_5732, \9389 );
and \U$9452 ( \18580 , RIf16f250_5724, \9391 );
and \U$9453 ( \18581 , RIfc6c440_6254, \9393 );
and \U$9454 ( \18582 , RIfcaba28_6975, \9395 );
and \U$9455 ( \18583 , RIfc40610_5758, \9397 );
and \U$9456 ( \18584 , RIe222e88_4687, \9399 );
and \U$9457 ( \18585 , RIfc5d260_6082, \9401 );
and \U$9458 ( \18586 , RIe220188_4655, \9403 );
and \U$9459 ( \18587 , RIfcab758_6973, \9405 );
and \U$9460 ( \18588 , RIe21d488_4623, \9407 );
and \U$9461 ( \18589 , RIe217a88_4559, \9409 );
and \U$9462 ( \18590 , RIe214d88_4527, \9411 );
and \U$9463 ( \18591 , RIfe892f8_7905, \9413 );
and \U$9464 ( \18592 , RIe212088_4495, \9415 );
and \U$9465 ( \18593 , RIf168a40_5650, \9417 );
and \U$9466 ( \18594 , RIe20f388_4463, \9419 );
and \U$9467 ( \18595 , RIf167ac8_5639, \9421 );
and \U$9468 ( \18596 , RIe20c688_4431, \9423 );
and \U$9469 ( \18597 , RIe209988_4399, \9425 );
and \U$9470 ( \18598 , RIe206c88_4367, \9427 );
and \U$9471 ( \18599 , RIfc6c2d8_6253, \9429 );
and \U$9472 ( \18600 , RIfceec88_7739, \9431 );
and \U$9473 ( \18601 , RIe201f30_4312, \9433 );
and \U$9474 ( \18602 , RIe200748_4295, \9435 );
and \U$9475 ( \18603 , RIf164dc8_5607, \9437 );
and \U$9476 ( \18604 , RIf163fb8_5597, \9439 );
and \U$9477 ( \18605 , RIf163040_5586, \9441 );
and \U$9478 ( \18606 , RIfe895c8_7907, \9443 );
and \U$9479 ( \18607 , RIf15f968_5547, \9445 );
and \U$9480 ( \18608 , RIfe89898_7909, \9447 );
and \U$9481 ( \18609 , RIfe89460_7906, \9449 );
and \U$9482 ( \18610 , RIe1fb5b8_4237, \9451 );
and \U$9483 ( \18611 , RIf15c6c8_5511, \9453 );
and \U$9484 ( \18612 , RIfe89730_7908, \9455 );
and \U$9485 ( \18613 , RIf15a238_5485, \9457 );
and \U$9486 ( \18614 , RIf1599c8_5479, \9459 );
or \U$9487 ( \18615 , \18551 , \18552 , \18553 , \18554 , \18555 , \18556 , \18557 , \18558 , \18559 , \18560 , \18561 , \18562 , \18563 , \18564 , \18565 , \18566 , \18567 , \18568 , \18569 , \18570 , \18571 , \18572 , \18573 , \18574 , \18575 , \18576 , \18577 , \18578 , \18579 , \18580 , \18581 , \18582 , \18583 , \18584 , \18585 , \18586 , \18587 , \18588 , \18589 , \18590 , \18591 , \18592 , \18593 , \18594 , \18595 , \18596 , \18597 , \18598 , \18599 , \18600 , \18601 , \18602 , \18603 , \18604 , \18605 , \18606 , \18607 , \18608 , \18609 , \18610 , \18611 , \18612 , \18613 , \18614 );
and \U$9488 ( \18616 , RIf1588e8_5467, \9462 );
and \U$9489 ( \18617 , RIfe89cd0_7912, \9464 );
and \U$9490 ( \18618 , RIfc5ba78_6065, \9466 );
and \U$9491 ( \18619 , RIe1f9c68_4219, \9468 );
and \U$9492 ( \18620 , RIfc5bd48_6067, \9470 );
and \U$9493 ( \18621 , RIf1554e0_5430, \9472 );
and \U$9494 ( \18622 , RIf154298_5417, \9474 );
and \U$9495 ( \18623 , RIe1f4c40_4162, \9476 );
and \U$9496 ( \18624 , RIfe89b68_7911, \9478 );
and \U$9497 ( \18625 , RIfe89a00_7910, \9480 );
and \U$9498 ( \18626 , RIf150350_5372, \9482 );
and \U$9499 ( \18627 , RIe1f2918_4137, \9484 );
and \U$9500 ( \18628 , RIf14f3d8_5361, \9486 );
and \U$9501 ( \18629 , RIfccc818_7349, \9488 );
and \U$9502 ( \18630 , RIf14d920_5342, \9490 );
and \U$9503 ( \18631 , RIe1ed620_4078, \9492 );
and \U$9504 ( \18632 , RIe1eabf0_4048, \9494 );
and \U$9505 ( \18633 , RIe1e7ef0_4016, \9496 );
and \U$9506 ( \18634 , RIe1e51f0_3984, \9498 );
and \U$9507 ( \18635 , RIe1e24f0_3952, \9500 );
and \U$9508 ( \18636 , RIe1df7f0_3920, \9502 );
and \U$9509 ( \18637 , RIe1dcaf0_3888, \9504 );
and \U$9510 ( \18638 , RIe1d9df0_3856, \9506 );
and \U$9511 ( \18639 , RIe1d70f0_3824, \9508 );
and \U$9512 ( \18640 , RIe1d16f0_3760, \9510 );
and \U$9513 ( \18641 , RIe1ce9f0_3728, \9512 );
and \U$9514 ( \18642 , RIe1cbcf0_3696, \9514 );
and \U$9515 ( \18643 , RIe1c8ff0_3664, \9516 );
and \U$9516 ( \18644 , RIe1c62f0_3632, \9518 );
and \U$9517 ( \18645 , RIe1c35f0_3600, \9520 );
and \U$9518 ( \18646 , RIe1c08f0_3568, \9522 );
and \U$9519 ( \18647 , RIe1bdbf0_3536, \9524 );
and \U$9520 ( \18648 , RIfc680c0_6206, \9526 );
and \U$9521 ( \18649 , RIf14b058_5313, \9528 );
and \U$9522 ( \18650 , RIe1b8bc8_3479, \9530 );
and \U$9523 ( \18651 , RIe1b6b70_3456, \9532 );
and \U$9524 ( \18652 , RIfcac298_6981, \9534 );
and \U$9525 ( \18653 , RIf1499d8_5297, \9536 );
and \U$9526 ( \18654 , RIfe89190_7904, \9538 );
and \U$9527 ( \18655 , RIfec19c8_8323, \9540 );
and \U$9528 ( \18656 , RIf148a60_5286, \9542 );
and \U$9529 ( \18657 , RIfccdd30_7364, \9544 );
and \U$9530 ( \18658 , RIe1b2250_3404, \9546 );
and \U$9531 ( \18659 , RIfec1860_8322, \9548 );
and \U$9532 ( \18660 , RIfc6e768_6279, \9550 );
and \U$9533 ( \18661 , RIfc54728_5983, \9552 );
and \U$9534 ( \18662 , RIe1abfe0_3334, \9554 );
and \U$9535 ( \18663 , RIe1aa528_3315, \9556 );
and \U$9536 ( \18664 , RIe1a7f30_3288, \9558 );
and \U$9537 ( \18665 , RIe1a5230_3256, \9560 );
and \U$9538 ( \18666 , RIe1a2530_3224, \9562 );
and \U$9539 ( \18667 , RIe19f830_3192, \9564 );
and \U$9540 ( \18668 , RIe18bd30_2968, \9566 );
and \U$9541 ( \18669 , RIe178230_2744, \9568 );
and \U$9542 ( \18670 , RIe225b88_4719, \9570 );
and \U$9543 ( \18671 , RIe21a788_4591, \9572 );
and \U$9544 ( \18672 , RIe203f88_4335, \9574 );
and \U$9545 ( \18673 , RIe1fdfe8_4267, \9576 );
and \U$9546 ( \18674 , RIe1f73a0_4190, \9578 );
and \U$9547 ( \18675 , RIe1efee8_4107, \9580 );
and \U$9548 ( \18676 , RIe1d43f0_3792, \9582 );
and \U$9549 ( \18677 , RIe1baef0_3504, \9584 );
and \U$9550 ( \18678 , RIe1add68_3355, \9586 );
and \U$9551 ( \18679 , RIe1703a0_2654, \9588 );
or \U$9552 ( \18680 , \18616 , \18617 , \18618 , \18619 , \18620 , \18621 , \18622 , \18623 , \18624 , \18625 , \18626 , \18627 , \18628 , \18629 , \18630 , \18631 , \18632 , \18633 , \18634 , \18635 , \18636 , \18637 , \18638 , \18639 , \18640 , \18641 , \18642 , \18643 , \18644 , \18645 , \18646 , \18647 , \18648 , \18649 , \18650 , \18651 , \18652 , \18653 , \18654 , \18655 , \18656 , \18657 , \18658 , \18659 , \18660 , \18661 , \18662 , \18663 , \18664 , \18665 , \18666 , \18667 , \18668 , \18669 , \18670 , \18671 , \18672 , \18673 , \18674 , \18675 , \18676 , \18677 , \18678 , \18679 );
or \U$9553 ( \18681 , \18615 , \18680 );
_DC g3c37 ( \18682_nG3c37 , \18681 , \9597 );
buf \U$9554 ( \18683 , \18682_nG3c37 );
and \U$9555 ( \18684 , \18550 , \18683 );
and \U$9556 ( \18685 , \16878 , \17011 );
and \U$9557 ( \18686 , \17011 , \17286 );
and \U$9558 ( \18687 , \16878 , \17286 );
or \U$9559 ( \18688 , \18685 , \18686 , \18687 );
and \U$9560 ( \18689 , \18683 , \18688 );
and \U$9561 ( \18690 , \18550 , \18688 );
or \U$9562 ( \18691 , \18684 , \18689 , \18690 );
xor \U$9563 ( \18692 , \18417 , \18691 );
buf g442a ( \18693_nG442a , \18692 );
xor \U$9564 ( \18694 , \18550 , \18683 );
xor \U$9565 ( \18695 , \18694 , \18688 );
buf g442d ( \18696_nG442d , \18695 );
nand \U$9566 ( \18697 , \18696_nG442d , \17288_nG4430 );
and \U$9567 ( \18698 , \18693_nG442a , \18697 );
xor \U$9568 ( \18699 , \18696_nG442d , \17288_nG4430 );
not \U$9569 ( \18700 , \18699 );
xor \U$9570 ( \18701 , \18693_nG442a , \18696_nG442d );
and \U$9571 ( \18702 , \18700 , \18701 );
and \U$9573 ( \18703 , \18699 , \10694_nG9c0e );
or \U$9574 ( \18704 , 1'b0 , \18703 );
xor \U$9575 ( \18705 , \18698 , \18704 );
xor \U$9576 ( \18706 , \18698 , \18705 );
buf \U$9577 ( \18707 , \18706 );
buf \U$9578 ( \18708 , \18707 );
and \U$9579 ( \18709 , \18150 , \18708 );
and \U$9580 ( \18710 , \18137 , \18142 );
and \U$9581 ( \18711 , \18137 , \18148 );
and \U$9582 ( \18712 , \18142 , \18148 );
or \U$9583 ( \18713 , \18710 , \18711 , \18712 );
buf \U$9584 ( \18714 , \18713 );
and \U$9585 ( \18715 , \17725 , \17762 );
and \U$9586 ( \18716 , \17725 , \18112 );
and \U$9587 ( \18717 , \17762 , \18112 );
or \U$9588 ( \18718 , \18715 , \18716 , \18717 );
buf \U$9589 ( \18719 , \18718 );
and \U$9590 ( \18720 , \17297 , \10995_nG9c0b );
and \U$9591 ( \18721 , \17294 , \11283_nG9c08 );
or \U$9592 ( \18722 , \18720 , \18721 );
xor \U$9593 ( \18723 , \17293 , \18722 );
buf \U$9594 ( \18724 , \18723 );
buf \U$9596 ( \18725 , \18724 );
and \U$9597 ( \18726 , \15940 , \11598_nG9c05 );
and \U$9598 ( \18727 , \15937 , \12470_nG9c02 );
or \U$9599 ( \18728 , \18726 , \18727 );
xor \U$9600 ( \18729 , \15936 , \18728 );
buf \U$9601 ( \18730 , \18729 );
buf \U$9603 ( \18731 , \18730 );
xor \U$9604 ( \18732 , \18725 , \18731 );
buf \U$9605 ( \18733 , \18732 );
and \U$9606 ( \18734 , \17728 , \17734 );
buf \U$9607 ( \18735 , \18734 );
xor \U$9608 ( \18736 , \18733 , \18735 );
and \U$9609 ( \18737 , \14631 , \12801_nG9bff );
and \U$9610 ( \18738 , \14628 , \13705_nG9bfc );
or \U$9611 ( \18739 , \18737 , \18738 );
xor \U$9612 ( \18740 , \14627 , \18739 );
buf \U$9613 ( \18741 , \18740 );
buf \U$9615 ( \18742 , \18741 );
xor \U$9616 ( \18743 , \18736 , \18742 );
buf \U$9617 ( \18744 , \18743 );
and \U$9618 ( \18745 , \10421 , \16680_nG9bed );
and \U$9619 ( \18746 , \10418 , \17665_nG9bea );
or \U$9620 ( \18747 , \18745 , \18746 );
xor \U$9621 ( \18748 , \10417 , \18747 );
buf \U$9622 ( \18749 , \18748 );
buf \U$9624 ( \18750 , \18749 );
xor \U$9625 ( \18751 , \18744 , \18750 );
and \U$9626 ( \18752 , \10707 , \18107_nG9be7 );
and \U$9627 ( \18753 , \18063 , \18077 );
and \U$9628 ( \18754 , \18077 , \18095 );
and \U$9629 ( \18755 , \18063 , \18095 );
or \U$9630 ( \18756 , \18753 , \18754 , \18755 );
and \U$9631 ( \18757 , \18067 , \18071 );
and \U$9632 ( \18758 , \18071 , \18076 );
and \U$9633 ( \18759 , \18067 , \18076 );
or \U$9634 ( \18760 , \18757 , \18758 , \18759 );
and \U$9635 ( \18761 , \18082 , \18086 );
and \U$9636 ( \18762 , \18086 , \18094 );
and \U$9637 ( \18763 , \18082 , \18094 );
or \U$9638 ( \18764 , \18761 , \18762 , \18763 );
xor \U$9639 ( \18765 , \18760 , \18764 );
and \U$9640 ( \18766 , \18035 , \10983 );
and \U$9641 ( \18767 , RIdec4898_700, \9333 );
and \U$9642 ( \18768 , RIdec1b98_668, \9335 );
and \U$9643 ( \18769 , RIfc661d0_6184, \9337 );
and \U$9644 ( \18770 , RIdebee98_636, \9339 );
and \U$9645 ( \18771 , RIfce6b28_7647, \9341 );
and \U$9646 ( \18772 , RIdebc198_604, \9343 );
and \U$9647 ( \18773 , RIdeb9498_572, \9345 );
and \U$9648 ( \18774 , RIdeb6798_540, \9347 );
and \U$9649 ( \18775 , RIfc40d18_5763, \9349 );
and \U$9650 ( \18776 , RIdeb0d98_476, \9351 );
and \U$9651 ( \18777 , RIfcad648_6995, \9353 );
and \U$9652 ( \18778 , RIdeae098_444, \9355 );
and \U$9653 ( \18779 , RIfcaa510_6960, \9357 );
and \U$9654 ( \18780 , RIdea89e0_412, \9359 );
and \U$9655 ( \18781 , RIdea20e0_380, \9361 );
and \U$9656 ( \18782 , RIde9b7e0_348, \9363 );
and \U$9657 ( \18783 , RIfcab320_6970, \9365 );
and \U$9658 ( \18784 , RIfca8350_6936, \9367 );
and \U$9659 ( \18785 , RIfc6f6e0_6290, \9369 );
and \U$9660 ( \18786 , RIfcaa240_6958, \9371 );
and \U$9661 ( \18787 , RIde8fcd8_291, \9373 );
and \U$9662 ( \18788 , RIfe8aae0_7922, \9375 );
and \U$9663 ( \18789 , RIde88d48_257, \9377 );
and \U$9664 ( \18790 , RIde84860_236, \9379 );
and \U$9665 ( \18791 , RIde80a08_217, \9381 );
and \U$9666 ( \18792 , RIfc64718_6165, \9383 );
and \U$9667 ( \18793 , RIfcae020_7002, \9385 );
and \U$9668 ( \18794 , RIfcadeb8_7001, \9387 );
and \U$9669 ( \18795 , RIee38fe0_5107, \9389 );
and \U$9670 ( \18796 , RIe16add8_2593, \9391 );
and \U$9671 ( \18797 , RIe1695f0_2576, \9393 );
and \U$9672 ( \18798 , RIe167430_2552, \9395 );
and \U$9673 ( \18799 , RIe164898_2521, \9397 );
and \U$9674 ( \18800 , RIe161b98_2489, \9399 );
and \U$9675 ( \18801 , RIfe8a3d8_7917, \9401 );
and \U$9676 ( \18802 , RIe15ee98_2457, \9403 );
and \U$9677 ( \18803 , RIfe8a270_7916, \9405 );
and \U$9678 ( \18804 , RIe15c198_2425, \9407 );
and \U$9679 ( \18805 , RIe156798_2361, \9409 );
and \U$9680 ( \18806 , RIe153a98_2329, \9411 );
and \U$9681 ( \18807 , RIfc3f0f8_5743, \9413 );
and \U$9682 ( \18808 , RIe150d98_2297, \9415 );
and \U$9683 ( \18809 , RIfcab050_6968, \9417 );
and \U$9684 ( \18810 , RIe14e098_2265, \9419 );
and \U$9685 ( \18811 , RIfcca658_7325, \9421 );
and \U$9686 ( \18812 , RIe14b398_2233, \9423 );
and \U$9687 ( \18813 , RIe148698_2201, \9425 );
and \U$9688 ( \18814 , RIe145998_2169, \9427 );
and \U$9689 ( \18815 , RIfe8a810_7920, \9429 );
and \U$9690 ( \18816 , RIfe8a6a8_7919, \9431 );
and \U$9691 ( \18817 , RIee31b28_5024, \9433 );
and \U$9692 ( \18818 , RIee30e80_5015, \9435 );
and \U$9693 ( \18819 , RIe140808_2111, \9437 );
and \U$9694 ( \18820 , RIfe8a540_7918, \9439 );
and \U$9695 ( \18821 , RIdf3c3e8_2062, \9441 );
and \U$9696 ( \18822 , RIdf3a0c0_2037, \9443 );
and \U$9697 ( \18823 , RIfc6b1f8_6241, \9445 );
and \U$9698 ( \18824 , RIee2f260_4995, \9447 );
and \U$9699 ( \18825 , RIfc70d60_6306, \9449 );
and \U$9700 ( \18826 , RIee2d0a0_4971, \9451 );
and \U$9701 ( \18827 , RIfe8a978_7921, \9453 );
and \U$9702 ( \18828 , RIdf32c08_1954, \9455 );
and \U$9703 ( \18829 , RIdf308e0_1929, \9457 );
and \U$9704 ( \18830 , RIdf2e9f0_1907, \9459 );
or \U$9705 ( \18831 , \18767 , \18768 , \18769 , \18770 , \18771 , \18772 , \18773 , \18774 , \18775 , \18776 , \18777 , \18778 , \18779 , \18780 , \18781 , \18782 , \18783 , \18784 , \18785 , \18786 , \18787 , \18788 , \18789 , \18790 , \18791 , \18792 , \18793 , \18794 , \18795 , \18796 , \18797 , \18798 , \18799 , \18800 , \18801 , \18802 , \18803 , \18804 , \18805 , \18806 , \18807 , \18808 , \18809 , \18810 , \18811 , \18812 , \18813 , \18814 , \18815 , \18816 , \18817 , \18818 , \18819 , \18820 , \18821 , \18822 , \18823 , \18824 , \18825 , \18826 , \18827 , \18828 , \18829 , \18830 );
and \U$9706 ( \18832 , RIee2b5e8_4952, \9462 );
and \U$9707 ( \18833 , RIee29e00_4935, \9464 );
and \U$9708 ( \18834 , RIee28a50_4921, \9466 );
and \U$9709 ( \18835 , RIee276a0_4907, \9468 );
and \U$9710 ( \18836 , RIdf29c98_1852, \9470 );
and \U$9711 ( \18837 , RIdf27970_1827, \9472 );
and \U$9712 ( \18838 , RIdf25be8_1806, \9474 );
and \U$9713 ( \18839 , RIdf23fc8_1786, \9476 );
and \U$9714 ( \18840 , RIfc6aaf0_6236, \9478 );
and \U$9715 ( \18841 , RIfc6ac58_6237, \9480 );
and \U$9716 ( \18842 , RIdf22678_1768, \9482 );
and \U$9717 ( \18843 , RIfcdd4b0_7540, \9484 );
and \U$9718 ( \18844 , RIdf21160_1753, \9486 );
and \U$9719 ( \18845 , RIdf1f108_1730, \9488 );
and \U$9720 ( \18846 , RIdf1ac20_1681, \9490 );
and \U$9721 ( \18847 , RIfeaa7f0_8256, \9492 );
and \U$9722 ( \18848 , RIdf16468_1630, \9494 );
and \U$9723 ( \18849 , RIdf13768_1598, \9496 );
and \U$9724 ( \18850 , RIdf10a68_1566, \9498 );
and \U$9725 ( \18851 , RIdf0dd68_1534, \9500 );
and \U$9726 ( \18852 , RIdf0b068_1502, \9502 );
and \U$9727 ( \18853 , RIdf08368_1470, \9504 );
and \U$9728 ( \18854 , RIdf05668_1438, \9506 );
and \U$9729 ( \18855 , RIdf02968_1406, \9508 );
and \U$9730 ( \18856 , RIdefcf68_1342, \9510 );
and \U$9731 ( \18857 , RIdefa268_1310, \9512 );
and \U$9732 ( \18858 , RIdef7568_1278, \9514 );
and \U$9733 ( \18859 , RIdef4868_1246, \9516 );
and \U$9734 ( \18860 , RIdef1b68_1214, \9518 );
and \U$9735 ( \18861 , RIdeeee68_1182, \9520 );
and \U$9736 ( \18862 , RIdeec168_1150, \9522 );
and \U$9737 ( \18863 , RIdee9468_1118, \9524 );
and \U$9738 ( \18864 , RIee25378_4882, \9526 );
and \U$9739 ( \18865 , RIee24568_4872, \9528 );
and \U$9740 ( \18866 , RIee23a28_4864, \9530 );
and \U$9741 ( \18867 , RIee23050_4857, \9532 );
and \U$9742 ( \18868 , RIfe8adb0_7924, \9534 );
and \U$9743 ( \18869 , RIdee23e8_1038, \9536 );
and \U$9744 ( \18870 , RIfe8ac48_7923, \9538 );
and \U$9745 ( \18871 , RIdede1d0_991, \9540 );
and \U$9746 ( \18872 , RIfca5650_6904, \9542 );
and \U$9747 ( \18873 , RIee220d8_4846, \9544 );
and \U$9748 ( \18874 , RIfceeb20_7738, \9546 );
and \U$9749 ( \18875 , RIee20ff8_4834, \9548 );
and \U$9750 ( \18876 , RIded8ed8_932, \9550 );
and \U$9751 ( \18877 , RIfe8af18_7925, \9552 );
and \U$9752 ( \18878 , RIded49f0_883, \9554 );
and \U$9753 ( \18879 , RIfe8b080_7926, \9556 );
and \U$9754 ( \18880 , RIdecfc98_828, \9558 );
and \U$9755 ( \18881 , RIdeccf98_796, \9560 );
and \U$9756 ( \18882 , RIdeca298_764, \9562 );
and \U$9757 ( \18883 , RIdec7598_732, \9564 );
and \U$9758 ( \18884 , RIdeb3a98_508, \9566 );
and \U$9759 ( \18885 , RIde94ee0_316, \9568 );
and \U$9760 ( \18886 , RIe16d6a0_2622, \9570 );
and \U$9761 ( \18887 , RIe159498_2393, \9572 );
and \U$9762 ( \18888 , RIe142c98_2137, \9574 );
and \U$9763 ( \18889 , RIdf37690_2007, \9576 );
and \U$9764 ( \18890 , RIdf2bcf0_1875, \9578 );
and \U$9765 ( \18891 , RIdf1c570_1699, \9580 );
and \U$9766 ( \18892 , RIdeffc68_1374, \9582 );
and \U$9767 ( \18893 , RIdee6768_1086, \9584 );
and \U$9768 ( \18894 , RIdedb4d0_959, \9586 );
and \U$9769 ( \18895 , RIde7ae28_189, \9588 );
or \U$9770 ( \18896 , \18832 , \18833 , \18834 , \18835 , \18836 , \18837 , \18838 , \18839 , \18840 , \18841 , \18842 , \18843 , \18844 , \18845 , \18846 , \18847 , \18848 , \18849 , \18850 , \18851 , \18852 , \18853 , \18854 , \18855 , \18856 , \18857 , \18858 , \18859 , \18860 , \18861 , \18862 , \18863 , \18864 , \18865 , \18866 , \18867 , \18868 , \18869 , \18870 , \18871 , \18872 , \18873 , \18874 , \18875 , \18876 , \18877 , \18878 , \18879 , \18880 , \18881 , \18882 , \18883 , \18884 , \18885 , \18886 , \18887 , \18888 , \18889 , \18890 , \18891 , \18892 , \18893 , \18894 , \18895 );
or \U$9771 ( \18897 , \18831 , \18896 );
_DC g65a1 ( \18898_nG65a1 , \18897 , \9597 );
and \U$9772 ( \18899 , RIe19cb30_3160, \9059 );
and \U$9773 ( \18900 , RIe199e30_3128, \9061 );
and \U$9774 ( \18901 , RIf145388_5247, \9063 );
and \U$9775 ( \18902 , RIe197130_3096, \9065 );
and \U$9776 ( \18903 , RIfe8a108_7915, \9067 );
and \U$9777 ( \18904 , RIe194430_3064, \9069 );
and \U$9778 ( \18905 , RIe191730_3032, \9071 );
and \U$9779 ( \18906 , RIe18ea30_3000, \9073 );
and \U$9780 ( \18907 , RIe189030_2936, \9075 );
and \U$9781 ( \18908 , RIe186330_2904, \9077 );
and \U$9782 ( \18909 , RIfc6c878_6257, \9079 );
and \U$9783 ( \18910 , RIe183630_2872, \9081 );
and \U$9784 ( \18911 , RIfcabcf8_6977, \9083 );
and \U$9785 ( \18912 , RIe180930_2840, \9085 );
and \U$9786 ( \18913 , RIe17dc30_2808, \9087 );
and \U$9787 ( \18914 , RIe17af30_2776, \9089 );
and \U$9788 ( \18915 , RIfcccc50_7352, \9091 );
and \U$9789 ( \18916 , RIfcccdb8_7353, \9093 );
and \U$9790 ( \18917 , RIe176d18_2729, \9095 );
and \U$9791 ( \18918 , RIfea7af0_8224, \9097 );
and \U$9792 ( \18919 , RIfe89fa0_7914, \9099 );
and \U$9793 ( \18920 , RIfe89e38_7913, \9101 );
and \U$9794 ( \18921 , RIfcdd078_7537, \9103 );
and \U$9795 ( \18922 , RIfccb738_7337, \9105 );
and \U$9796 ( \18923 , RIfca9868_6951, \9107 );
and \U$9797 ( \18924 , RIfcabb90_6976, \9109 );
and \U$9798 ( \18925 , RIfca99d0_6952, \9111 );
and \U$9799 ( \18926 , RIe172f38_2685, \9113 );
and \U$9800 ( \18927 , RIf16fd90_5732, \9115 );
and \U$9801 ( \18928 , RIf16f250_5724, \9117 );
and \U$9802 ( \18929 , RIfc6c440_6254, \9119 );
and \U$9803 ( \18930 , RIfcaba28_6975, \9121 );
and \U$9804 ( \18931 , RIfc40610_5758, \9123 );
and \U$9805 ( \18932 , RIe222e88_4687, \9125 );
and \U$9806 ( \18933 , RIfc5d260_6082, \9127 );
and \U$9807 ( \18934 , RIe220188_4655, \9129 );
and \U$9808 ( \18935 , RIfcab758_6973, \9131 );
and \U$9809 ( \18936 , RIe21d488_4623, \9133 );
and \U$9810 ( \18937 , RIe217a88_4559, \9135 );
and \U$9811 ( \18938 , RIe214d88_4527, \9137 );
and \U$9812 ( \18939 , RIfe892f8_7905, \9139 );
and \U$9813 ( \18940 , RIe212088_4495, \9141 );
and \U$9814 ( \18941 , RIf168a40_5650, \9143 );
and \U$9815 ( \18942 , RIe20f388_4463, \9145 );
and \U$9816 ( \18943 , RIf167ac8_5639, \9147 );
and \U$9817 ( \18944 , RIe20c688_4431, \9149 );
and \U$9818 ( \18945 , RIe209988_4399, \9151 );
and \U$9819 ( \18946 , RIe206c88_4367, \9153 );
and \U$9820 ( \18947 , RIfc6c2d8_6253, \9155 );
and \U$9821 ( \18948 , RIfceec88_7739, \9157 );
and \U$9822 ( \18949 , RIe201f30_4312, \9159 );
and \U$9823 ( \18950 , RIe200748_4295, \9161 );
and \U$9824 ( \18951 , RIf164dc8_5607, \9163 );
and \U$9825 ( \18952 , RIf163fb8_5597, \9165 );
and \U$9826 ( \18953 , RIf163040_5586, \9167 );
and \U$9827 ( \18954 , RIfe895c8_7907, \9169 );
and \U$9828 ( \18955 , RIf15f968_5547, \9171 );
and \U$9829 ( \18956 , RIfe89898_7909, \9173 );
and \U$9830 ( \18957 , RIfe89460_7906, \9175 );
and \U$9831 ( \18958 , RIe1fb5b8_4237, \9177 );
and \U$9832 ( \18959 , RIf15c6c8_5511, \9179 );
and \U$9833 ( \18960 , RIfe89730_7908, \9181 );
and \U$9834 ( \18961 , RIf15a238_5485, \9183 );
and \U$9835 ( \18962 , RIf1599c8_5479, \9185 );
or \U$9836 ( \18963 , \18899 , \18900 , \18901 , \18902 , \18903 , \18904 , \18905 , \18906 , \18907 , \18908 , \18909 , \18910 , \18911 , \18912 , \18913 , \18914 , \18915 , \18916 , \18917 , \18918 , \18919 , \18920 , \18921 , \18922 , \18923 , \18924 , \18925 , \18926 , \18927 , \18928 , \18929 , \18930 , \18931 , \18932 , \18933 , \18934 , \18935 , \18936 , \18937 , \18938 , \18939 , \18940 , \18941 , \18942 , \18943 , \18944 , \18945 , \18946 , \18947 , \18948 , \18949 , \18950 , \18951 , \18952 , \18953 , \18954 , \18955 , \18956 , \18957 , \18958 , \18959 , \18960 , \18961 , \18962 );
and \U$9837 ( \18964 , RIf1588e8_5467, \9188 );
and \U$9838 ( \18965 , RIfe89cd0_7912, \9190 );
and \U$9839 ( \18966 , RIfc5ba78_6065, \9192 );
and \U$9840 ( \18967 , RIe1f9c68_4219, \9194 );
and \U$9841 ( \18968 , RIfc5bd48_6067, \9196 );
and \U$9842 ( \18969 , RIf1554e0_5430, \9198 );
and \U$9843 ( \18970 , RIf154298_5417, \9200 );
and \U$9844 ( \18971 , RIe1f4c40_4162, \9202 );
and \U$9845 ( \18972 , RIfe89b68_7911, \9204 );
and \U$9846 ( \18973 , RIfe89a00_7910, \9206 );
and \U$9847 ( \18974 , RIf150350_5372, \9208 );
and \U$9848 ( \18975 , RIe1f2918_4137, \9210 );
and \U$9849 ( \18976 , RIf14f3d8_5361, \9212 );
and \U$9850 ( \18977 , RIfccc818_7349, \9214 );
and \U$9851 ( \18978 , RIf14d920_5342, \9216 );
and \U$9852 ( \18979 , RIe1ed620_4078, \9218 );
and \U$9853 ( \18980 , RIe1eabf0_4048, \9220 );
and \U$9854 ( \18981 , RIe1e7ef0_4016, \9222 );
and \U$9855 ( \18982 , RIe1e51f0_3984, \9224 );
and \U$9856 ( \18983 , RIe1e24f0_3952, \9226 );
and \U$9857 ( \18984 , RIe1df7f0_3920, \9228 );
and \U$9858 ( \18985 , RIe1dcaf0_3888, \9230 );
and \U$9859 ( \18986 , RIe1d9df0_3856, \9232 );
and \U$9860 ( \18987 , RIe1d70f0_3824, \9234 );
and \U$9861 ( \18988 , RIe1d16f0_3760, \9236 );
and \U$9862 ( \18989 , RIe1ce9f0_3728, \9238 );
and \U$9863 ( \18990 , RIe1cbcf0_3696, \9240 );
and \U$9864 ( \18991 , RIe1c8ff0_3664, \9242 );
and \U$9865 ( \18992 , RIe1c62f0_3632, \9244 );
and \U$9866 ( \18993 , RIe1c35f0_3600, \9246 );
and \U$9867 ( \18994 , RIe1c08f0_3568, \9248 );
and \U$9868 ( \18995 , RIe1bdbf0_3536, \9250 );
and \U$9869 ( \18996 , RIfc680c0_6206, \9252 );
and \U$9870 ( \18997 , RIf14b058_5313, \9254 );
and \U$9871 ( \18998 , RIe1b8bc8_3479, \9256 );
and \U$9872 ( \18999 , RIe1b6b70_3456, \9258 );
and \U$9873 ( \19000 , RIfcac298_6981, \9260 );
and \U$9874 ( \19001 , RIf1499d8_5297, \9262 );
and \U$9875 ( \19002 , RIfe89190_7904, \9264 );
and \U$9876 ( \19003 , RIfec19c8_8323, \9266 );
and \U$9877 ( \19004 , RIf148a60_5286, \9268 );
and \U$9878 ( \19005 , RIfccdd30_7364, \9270 );
and \U$9879 ( \19006 , RIe1b2250_3404, \9272 );
and \U$9880 ( \19007 , RIfec1860_8322, \9274 );
and \U$9881 ( \19008 , RIfc6e768_6279, \9276 );
and \U$9882 ( \19009 , RIfc54728_5983, \9278 );
and \U$9883 ( \19010 , RIe1abfe0_3334, \9280 );
and \U$9884 ( \19011 , RIe1aa528_3315, \9282 );
and \U$9885 ( \19012 , RIe1a7f30_3288, \9284 );
and \U$9886 ( \19013 , RIe1a5230_3256, \9286 );
and \U$9887 ( \19014 , RIe1a2530_3224, \9288 );
and \U$9888 ( \19015 , RIe19f830_3192, \9290 );
and \U$9889 ( \19016 , RIe18bd30_2968, \9292 );
and \U$9890 ( \19017 , RIe178230_2744, \9294 );
and \U$9891 ( \19018 , RIe225b88_4719, \9296 );
and \U$9892 ( \19019 , RIe21a788_4591, \9298 );
and \U$9893 ( \19020 , RIe203f88_4335, \9300 );
and \U$9894 ( \19021 , RIe1fdfe8_4267, \9302 );
and \U$9895 ( \19022 , RIe1f73a0_4190, \9304 );
and \U$9896 ( \19023 , RIe1efee8_4107, \9306 );
and \U$9897 ( \19024 , RIe1d43f0_3792, \9308 );
and \U$9898 ( \19025 , RIe1baef0_3504, \9310 );
and \U$9899 ( \19026 , RIe1add68_3355, \9312 );
and \U$9900 ( \19027 , RIe1703a0_2654, \9314 );
or \U$9901 ( \19028 , \18964 , \18965 , \18966 , \18967 , \18968 , \18969 , \18970 , \18971 , \18972 , \18973 , \18974 , \18975 , \18976 , \18977 , \18978 , \18979 , \18980 , \18981 , \18982 , \18983 , \18984 , \18985 , \18986 , \18987 , \18988 , \18989 , \18990 , \18991 , \18992 , \18993 , \18994 , \18995 , \18996 , \18997 , \18998 , \18999 , \19000 , \19001 , \19002 , \19003 , \19004 , \19005 , \19006 , \19007 , \19008 , \19009 , \19010 , \19011 , \19012 , \19013 , \19014 , \19015 , \19016 , \19017 , \19018 , \19019 , \19020 , \19021 , \19022 , \19023 , \19024 , \19025 , \19026 , \19027 );
or \U$9902 ( \19029 , \18963 , \19028 );
_DC g65a2 ( \19030_nG65a2 , \19029 , \9323 );
and g65a3 ( \19031_nG65a3 , \18898_nG65a1 , \19030_nG65a2 );
buf \U$9903 ( \19032 , \19031_nG65a3 );
and \U$9904 ( \19033 , \19032 , \10691 );
nor \U$9905 ( \19034 , \18766 , \19033 );
xnor \U$9906 ( \19035 , \19034 , \10980 );
and \U$9907 ( \19036 , \16655 , \11574 );
and \U$9908 ( \19037 , \17627 , \11278 );
nor \U$9909 ( \19038 , \19036 , \19037 );
xnor \U$9910 ( \19039 , \19038 , \11580 );
xor \U$9911 ( \19040 , \19035 , \19039 );
_DC g5358 ( \19041_nG5358 , \18897 , \9597 );
_DC g53dc ( \19042_nG53dc , \19029 , \9323 );
xor g53dd ( \19043_nG53dd , \19041_nG5358 , \19042_nG53dc );
buf \U$9912 ( \19044 , \19043_nG53dd );
xor \U$9913 ( \19045 , \19044 , \18043 );
and \U$9914 ( \19046 , \10687 , \19045 );
xor \U$9915 ( \19047 , \19040 , \19046 );
xor \U$9916 ( \19048 , \18765 , \19047 );
xor \U$9917 ( \19049 , \18756 , \19048 );
and \U$9918 ( \19050 , \18048 , \18052 );
and \U$9919 ( \19051 , \18052 , \18057 );
and \U$9920 ( \19052 , \18048 , \18057 );
or \U$9921 ( \19053 , \19050 , \19051 , \19052 );
and \U$9922 ( \19054 , \15321 , \12790 );
and \U$9923 ( \19055 , \16267 , \12461 );
nor \U$9924 ( \19056 , \19054 , \19055 );
xnor \U$9925 ( \19057 , \19056 , \12780 );
and \U$9926 ( \19058 , \14024 , \14054 );
and \U$9927 ( \19059 , \14950 , \13692 );
nor \U$9928 ( \19060 , \19058 , \19059 );
xnor \U$9929 ( \19061 , \19060 , \14035 );
xor \U$9930 ( \19062 , \19057 , \19061 );
and \U$9931 ( \19063 , \12769 , \15336 );
and \U$9932 ( \19064 , \13679 , \14963 );
nor \U$9933 ( \19065 , \19063 , \19064 );
xnor \U$9934 ( \19066 , \19065 , \15342 );
xor \U$9935 ( \19067 , \19062 , \19066 );
xor \U$9936 ( \19068 , \19053 , \19067 );
and \U$9937 ( \19069 , \18038 , \18047 );
and \U$9938 ( \19070 , \11586 , \16635 );
and \U$9939 ( \19071 , \12448 , \16301 );
nor \U$9940 ( \19072 , \19070 , \19071 );
xnor \U$9941 ( \19073 , \19072 , \16625 );
xor \U$9942 ( \19074 , \19069 , \19073 );
and \U$9943 ( \19075 , \10988 , \18090 );
and \U$9944 ( \19076 , \11270 , \17655 );
nor \U$9945 ( \19077 , \19075 , \19076 );
xnor \U$9946 ( \19078 , \19077 , \18046 );
xor \U$9947 ( \19079 , \19074 , \19078 );
xor \U$9948 ( \19080 , \19068 , \19079 );
xor \U$9949 ( \19081 , \19049 , \19080 );
and \U$9950 ( \19082 , \17768 , \18058 );
and \U$9951 ( \19083 , \18058 , \18096 );
and \U$9952 ( \19084 , \17768 , \18096 );
or \U$9953 ( \19085 , \19082 , \19083 , \19084 );
xor \U$9954 ( \19086 , \19081 , \19085 );
and \U$9955 ( \19087 , \18097 , \18101 );
and \U$9956 ( \19088 , \18102 , \18105 );
or \U$9957 ( \19089 , \19087 , \19088 );
xor \U$9958 ( \19090 , \19086 , \19089 );
buf g9be4 ( \19091_nG9be4 , \19090 );
and \U$9959 ( \19092 , \10704 , \19091_nG9be4 );
or \U$9960 ( \19093 , \18752 , \19092 );
xor \U$9961 ( \19094 , \10703 , \19093 );
buf \U$9962 ( \19095 , \19094 );
buf \U$9964 ( \19096 , \19095 );
xor \U$9965 ( \19097 , \18751 , \19096 );
buf \U$9966 ( \19098 , \19097 );
xor \U$9967 ( \19099 , \18719 , \19098 );
and \U$9968 ( \19100 , \18120 , \18126 );
and \U$9969 ( \19101 , \18120 , \18133 );
and \U$9970 ( \19102 , \18126 , \18133 );
or \U$9971 ( \19103 , \19100 , \19101 , \19102 );
buf \U$9972 ( \19104 , \19103 );
and \U$9973 ( \19105 , \17736 , \17742 );
and \U$9974 ( \19106 , \17736 , \17749 );
and \U$9975 ( \19107 , \17742 , \17749 );
or \U$9976 ( \19108 , \19105 , \19106 , \19107 );
buf \U$9977 ( \19109 , \19108 );
and \U$9978 ( \19110 , \13370 , \14070_nG9bf9 );
and \U$9979 ( \19111 , \13367 , \14984_nG9bf6 );
or \U$9980 ( \19112 , \19110 , \19111 );
xor \U$9981 ( \19113 , \13366 , \19112 );
buf \U$9982 ( \19114 , \19113 );
buf \U$9984 ( \19115 , \19114 );
xor \U$9985 ( \19116 , \19109 , \19115 );
and \U$9986 ( \19117 , \12157 , \15373_nG9bf3 );
and \U$9987 ( \19118 , \12154 , \16315_nG9bf0 );
or \U$9988 ( \19119 , \19117 , \19118 );
xor \U$9989 ( \19120 , \12153 , \19119 );
buf \U$9990 ( \19121 , \19120 );
buf \U$9992 ( \19122 , \19121 );
xor \U$9993 ( \19123 , \19116 , \19122 );
buf \U$9994 ( \19124 , \19123 );
xor \U$9995 ( \19125 , \19104 , \19124 );
and \U$9996 ( \19126 , \17751 , \17753 );
and \U$9997 ( \19127 , \17751 , \17760 );
and \U$9998 ( \19128 , \17753 , \17760 );
or \U$9999 ( \19129 , \19126 , \19127 , \19128 );
buf \U$10000 ( \19130 , \19129 );
xor \U$10001 ( \19131 , \19125 , \19130 );
buf \U$10002 ( \19132 , \19131 );
xor \U$10003 ( \19133 , \19099 , \19132 );
buf \U$10004 ( \19134 , \19133 );
xor \U$10005 ( \19135 , \18714 , \19134 );
and \U$10006 ( \19136 , \17720 , \18114 );
and \U$10007 ( \19137 , \17720 , \18135 );
and \U$10008 ( \19138 , \18114 , \18135 );
or \U$10009 ( \19139 , \19136 , \19137 , \19138 );
buf \U$10010 ( \19140 , \19139 );
xor \U$10011 ( \19141 , \19135 , \19140 );
and \U$10012 ( \19142 , \18150 , \19141 );
and \U$10013 ( \19143 , \18708 , \19141 );
or \U$10014 ( \19144 , \18709 , \19142 , \19143 );
and \U$10015 ( \19145 , \18714 , \19134 );
and \U$10016 ( \19146 , \18714 , \19140 );
and \U$10017 ( \19147 , \19134 , \19140 );
or \U$10018 ( \19148 , \19145 , \19146 , \19147 );
buf \U$10019 ( \19149 , \19148 );
and \U$10020 ( \19150 , \19104 , \19124 );
and \U$10021 ( \19151 , \19104 , \19130 );
and \U$10022 ( \19152 , \19124 , \19130 );
or \U$10023 ( \19153 , \19150 , \19151 , \19152 );
buf \U$10024 ( \19154 , \19153 );
and \U$10025 ( \19155 , \19109 , \19115 );
and \U$10026 ( \19156 , \19109 , \19122 );
and \U$10027 ( \19157 , \19115 , \19122 );
or \U$10028 ( \19158 , \19155 , \19156 , \19157 );
buf \U$10029 ( \19159 , \19158 );
and \U$10030 ( \19160 , \18725 , \18731 );
buf \U$10031 ( \19161 , \19160 );
and \U$10032 ( \19162 , \14631 , \13705_nG9bfc );
and \U$10033 ( \19163 , \14628 , \14070_nG9bf9 );
or \U$10034 ( \19164 , \19162 , \19163 );
xor \U$10035 ( \19165 , \14627 , \19164 );
buf \U$10036 ( \19166 , \19165 );
buf \U$10038 ( \19167 , \19166 );
xor \U$10039 ( \19168 , \19161 , \19167 );
and \U$10040 ( \19169 , \13370 , \14984_nG9bf6 );
and \U$10041 ( \19170 , \13367 , \15373_nG9bf3 );
or \U$10042 ( \19171 , \19169 , \19170 );
xor \U$10043 ( \19172 , \13366 , \19171 );
buf \U$10044 ( \19173 , \19172 );
buf \U$10046 ( \19174 , \19173 );
xor \U$10047 ( \19175 , \19168 , \19174 );
buf \U$10048 ( \19176 , \19175 );
xor \U$10049 ( \19177 , \19159 , \19176 );
and \U$10050 ( \19178 , \10421 , \17665_nG9bea );
and \U$10051 ( \19179 , \10418 , \18107_nG9be7 );
or \U$10052 ( \19180 , \19178 , \19179 );
xor \U$10053 ( \19181 , \10417 , \19180 );
buf \U$10054 ( \19182 , \19181 );
buf \U$10056 ( \19183 , \19182 );
xor \U$10057 ( \19184 , \19177 , \19183 );
buf \U$10058 ( \19185 , \19184 );
xor \U$10059 ( \19186 , \19154 , \19185 );
and \U$10060 ( \19187 , \18744 , \18750 );
and \U$10061 ( \19188 , \18744 , \19096 );
and \U$10062 ( \19189 , \18750 , \19096 );
or \U$10063 ( \19190 , \19187 , \19188 , \19189 );
buf \U$10064 ( \19191 , \19190 );
and \U$10065 ( \19192 , \18733 , \18735 );
and \U$10066 ( \19193 , \18733 , \18742 );
and \U$10067 ( \19194 , \18735 , \18742 );
or \U$10068 ( \19195 , \19192 , \19193 , \19194 );
buf \U$10069 ( \19196 , \19195 );
and \U$10070 ( \19197 , \18698 , \18705 );
buf \U$10071 ( \19198 , \19197 );
buf \U$10073 ( \19199 , \19198 );
and \U$10074 ( \19200 , \17297 , \11283_nG9c08 );
and \U$10075 ( \19201 , \17294 , \11598_nG9c05 );
or \U$10076 ( \19202 , \19200 , \19201 );
xor \U$10077 ( \19203 , \17293 , \19202 );
buf \U$10078 ( \19204 , \19203 );
buf \U$10080 ( \19205 , \19204 );
xor \U$10081 ( \19206 , \19199 , \19205 );
buf \U$10082 ( \19207 , \19206 );
and \U$10083 ( \19208 , \18702 , \10694_nG9c0e );
and \U$10084 ( \19209 , \18699 , \10995_nG9c0b );
or \U$10085 ( \19210 , \19208 , \19209 );
xor \U$10086 ( \19211 , \18698 , \19210 );
buf \U$10087 ( \19212 , \19211 );
buf \U$10089 ( \19213 , \19212 );
xor \U$10090 ( \19214 , \19207 , \19213 );
and \U$10091 ( \19215 , \15940 , \12470_nG9c02 );
and \U$10092 ( \19216 , \15937 , \12801_nG9bff );
or \U$10093 ( \19217 , \19215 , \19216 );
xor \U$10094 ( \19218 , \15936 , \19217 );
buf \U$10095 ( \19219 , \19218 );
buf \U$10097 ( \19220 , \19219 );
xor \U$10098 ( \19221 , \19214 , \19220 );
buf \U$10099 ( \19222 , \19221 );
xor \U$10100 ( \19223 , \19196 , \19222 );
and \U$10101 ( \19224 , \12157 , \16315_nG9bf0 );
and \U$10102 ( \19225 , \12154 , \16680_nG9bed );
or \U$10103 ( \19226 , \19224 , \19225 );
xor \U$10104 ( \19227 , \12153 , \19226 );
buf \U$10105 ( \19228 , \19227 );
buf \U$10107 ( \19229 , \19228 );
xor \U$10108 ( \19230 , \19223 , \19229 );
buf \U$10109 ( \19231 , \19230 );
xor \U$10110 ( \19232 , \19191 , \19231 );
and \U$10111 ( \19233 , \10707 , \19091_nG9be4 );
and \U$10112 ( \19234 , \19053 , \19067 );
and \U$10113 ( \19235 , \19067 , \19079 );
and \U$10114 ( \19236 , \19053 , \19079 );
or \U$10115 ( \19237 , \19234 , \19235 , \19236 );
and \U$10116 ( \19238 , \19057 , \19061 );
and \U$10117 ( \19239 , \19061 , \19066 );
and \U$10118 ( \19240 , \19057 , \19066 );
or \U$10119 ( \19241 , \19238 , \19239 , \19240 );
and \U$10120 ( \19242 , \16267 , \12790 );
and \U$10121 ( \19243 , \16655 , \12461 );
nor \U$10122 ( \19244 , \19242 , \19243 );
xnor \U$10123 ( \19245 , \19244 , \12780 );
and \U$10124 ( \19246 , \13679 , \15336 );
and \U$10125 ( \19247 , \14024 , \14963 );
nor \U$10126 ( \19248 , \19246 , \19247 );
xnor \U$10127 ( \19249 , \19248 , \15342 );
xor \U$10128 ( \19250 , \19245 , \19249 );
and \U$10129 ( \19251 , \12448 , \16635 );
and \U$10130 ( \19252 , \12769 , \16301 );
nor \U$10131 ( \19253 , \19251 , \19252 );
xnor \U$10132 ( \19254 , \19253 , \16625 );
xor \U$10133 ( \19255 , \19250 , \19254 );
xor \U$10134 ( \19256 , \19241 , \19255 );
and \U$10135 ( \19257 , \17627 , \11574 );
and \U$10136 ( \19258 , \18035 , \11278 );
nor \U$10137 ( \19259 , \19257 , \19258 );
xnor \U$10138 ( \19260 , \19259 , \11580 );
and \U$10139 ( \19261 , \14950 , \14054 );
and \U$10140 ( \19262 , \15321 , \13692 );
nor \U$10141 ( \19263 , \19261 , \19262 );
xnor \U$10142 ( \19264 , \19263 , \14035 );
xor \U$10143 ( \19265 , \19260 , \19264 );
and \U$10144 ( \19266 , RIdec4a00_701, \9333 );
and \U$10145 ( \19267 , RIdec1d00_669, \9335 );
and \U$10146 ( \19268 , RIfcad7b0_6996, \9337 );
and \U$10147 ( \19269 , RIdebf000_637, \9339 );
and \U$10148 ( \19270 , RIfc64cb8_6169, \9341 );
and \U$10149 ( \19271 , RIdebc300_605, \9343 );
and \U$10150 ( \19272 , RIdeb9600_573, \9345 );
and \U$10151 ( \19273 , RIdeb6900_541, \9347 );
and \U$10152 ( \19274 , RIfc6f9b0_6292, \9349 );
and \U$10153 ( \19275 , RIdeb0f00_477, \9351 );
and \U$10154 ( \19276 , RIfc657f8_6177, \9353 );
and \U$10155 ( \19277 , RIdeae200_445, \9355 );
and \U$10156 ( \19278 , RIfce69c0_7646, \9357 );
and \U$10157 ( \19279 , RIdea8d28_413, \9359 );
and \U$10158 ( \19280 , RIdea2428_381, \9361 );
and \U$10159 ( \19281 , RIde9bb28_349, \9363 );
and \U$10160 ( \19282 , RIfc6fc80_6294, \9365 );
and \U$10161 ( \19283 , RIee1b760_4771, \9367 );
and \U$10162 ( \19284 , RIfca8080_6934, \9369 );
and \U$10163 ( \19285 , RIfe8b8f0_7932, \9371 );
and \U$10164 ( \19286 , RIde90020_292, \9373 );
and \U$10165 ( \19287 , RIde8c510_274, \9375 );
and \U$10166 ( \19288 , RIde89090_258, \9377 );
and \U$10167 ( \19289 , RIde84ba8_237, \9379 );
and \U$10168 ( \19290 , RIfc65ac8_6179, \9381 );
and \U$10169 ( \19291 , RIfcad210_6992, \9383 );
and \U$10170 ( \19292 , RIfcce168_7367, \9385 );
and \U$10171 ( \19293 , RIfcce2d0_7368, \9387 );
and \U$10172 ( \19294 , RIfc51488_5947, \9389 );
and \U$10173 ( \19295 , RIe16af40_2594, \9391 );
and \U$10174 ( \19296 , RIfc65c30_6180, \9393 );
and \U$10175 ( \19297 , RIe167598_2553, \9395 );
and \U$10176 ( \19298 , RIe164a00_2522, \9397 );
and \U$10177 ( \19299 , RIe161d00_2490, \9399 );
and \U$10178 ( \19300 , RIfc66e78_6193, \9401 );
and \U$10179 ( \19301 , RIe15f000_2458, \9403 );
and \U$10180 ( \19302 , RIfc6e498_6277, \9405 );
and \U$10181 ( \19303 , RIe15c300_2426, \9407 );
and \U$10182 ( \19304 , RIe156900_2362, \9409 );
and \U$10183 ( \19305 , RIe153c00_2330, \9411 );
and \U$10184 ( \19306 , RIfc6e330_6276, \9413 );
and \U$10185 ( \19307 , RIe150f00_2298, \9415 );
and \U$10186 ( \19308 , RIfccda60_7362, \9417 );
and \U$10187 ( \19309 , RIe14e200_2266, \9419 );
and \U$10188 ( \19310 , RIfc6e1c8_6275, \9421 );
and \U$10189 ( \19311 , RIe14b500_2234, \9423 );
and \U$10190 ( \19312 , RIe148800_2202, \9425 );
and \U$10191 ( \19313 , RIe145b00_2170, \9427 );
and \U$10192 ( \19314 , RIee33fb8_5050, \9429 );
and \U$10193 ( \19315 , RIee32d70_5037, \9431 );
and \U$10194 ( \19316 , RIee31c90_5025, \9433 );
and \U$10195 ( \19317 , RIee30fe8_5016, \9435 );
and \U$10196 ( \19318 , RIfea8630_8232, \9437 );
and \U$10197 ( \19319 , RIdf3e5a8_2086, \9439 );
and \U$10198 ( \19320 , RIdf3c550_2063, \9441 );
and \U$10199 ( \19321 , RIfea8798_8233, \9443 );
and \U$10200 ( \19322 , RIfc6e060_6274, \9445 );
and \U$10201 ( \19323 , RIfcac6d0_6984, \9447 );
and \U$10202 ( \19324 , RIfc56078_6001, \9449 );
and \U$10203 ( \19325 , RIfc6e600_6278, \9451 );
and \U$10204 ( \19326 , RIdf34dc8_1978, \9453 );
and \U$10205 ( \19327 , RIdf32d70_1955, \9455 );
and \U$10206 ( \19328 , RIfea84c8_8231, \9457 );
and \U$10207 ( \19329 , RIdf2eb58_1908, \9459 );
or \U$10208 ( \19330 , \19266 , \19267 , \19268 , \19269 , \19270 , \19271 , \19272 , \19273 , \19274 , \19275 , \19276 , \19277 , \19278 , \19279 , \19280 , \19281 , \19282 , \19283 , \19284 , \19285 , \19286 , \19287 , \19288 , \19289 , \19290 , \19291 , \19292 , \19293 , \19294 , \19295 , \19296 , \19297 , \19298 , \19299 , \19300 , \19301 , \19302 , \19303 , \19304 , \19305 , \19306 , \19307 , \19308 , \19309 , \19310 , \19311 , \19312 , \19313 , \19314 , \19315 , \19316 , \19317 , \19318 , \19319 , \19320 , \19321 , \19322 , \19323 , \19324 , \19325 , \19326 , \19327 , \19328 , \19329 );
and \U$10209 ( \19331 , RIee2b750_4953, \9462 );
and \U$10210 ( \19332 , RIfc6ee70_6284, \9464 );
and \U$10211 ( \19333 , RIfc6efd8_6285, \9466 );
and \U$10212 ( \19334 , RIee27808_4908, \9468 );
and \U$10213 ( \19335 , RIfe8b788_7931, \9470 );
and \U$10214 ( \19336 , RIdf27ad8_1828, \9472 );
and \U$10215 ( \19337 , RIdf25d50_1807, \9474 );
and \U$10216 ( \19338 , RIdf24130_1787, \9476 );
and \U$10217 ( \19339 , RIfc66608_6187, \9478 );
and \U$10218 ( \19340 , RIfccde98_7365, \9480 );
and \U$10219 ( \19341 , RIfc66a40_6190, \9482 );
and \U$10220 ( \19342 , RIfc668d8_6189, \9484 );
and \U$10221 ( \19343 , RIfcacf40_6990, \9486 );
and \U$10222 ( \19344 , RIfeaaef8_8261, \9488 );
and \U$10223 ( \19345 , RIfc6e8d0_6280, \9490 );
and \U$10224 ( \19346 , RIdf18d30_1659, \9492 );
and \U$10225 ( \19347 , RIdf165d0_1631, \9494 );
and \U$10226 ( \19348 , RIdf138d0_1599, \9496 );
and \U$10227 ( \19349 , RIdf10bd0_1567, \9498 );
and \U$10228 ( \19350 , RIdf0ded0_1535, \9500 );
and \U$10229 ( \19351 , RIdf0b1d0_1503, \9502 );
and \U$10230 ( \19352 , RIdf084d0_1471, \9504 );
and \U$10231 ( \19353 , RIdf057d0_1439, \9506 );
and \U$10232 ( \19354 , RIdf02ad0_1407, \9508 );
and \U$10233 ( \19355 , RIdefd0d0_1343, \9510 );
and \U$10234 ( \19356 , RIdefa3d0_1311, \9512 );
and \U$10235 ( \19357 , RIdef76d0_1279, \9514 );
and \U$10236 ( \19358 , RIdef49d0_1247, \9516 );
and \U$10237 ( \19359 , RIdef1cd0_1215, \9518 );
and \U$10238 ( \19360 , RIdeeefd0_1183, \9520 );
and \U$10239 ( \19361 , RIdeec2d0_1151, \9522 );
and \U$10240 ( \19362 , RIdee95d0_1119, \9524 );
and \U$10241 ( \19363 , RIfc6dc28_6271, \9526 );
and \U$10242 ( \19364 , RIfc67c88_6203, \9528 );
and \U$10243 ( \19365 , RIfccb300_7334, \9530 );
and \U$10244 ( \19366 , RIfccd4c0_7358, \9532 );
and \U$10245 ( \19367 , RIfea81f8_8229, \9534 );
and \U$10246 ( \19368 , RIfea8360_8230, \9536 );
and \U$10247 ( \19369 , RIdee04f8_1016, \9538 );
and \U$10248 ( \19370 , RIdede338_992, \9540 );
and \U$10249 ( \19371 , RIfc6def8_6273, \9542 );
and \U$10250 ( \19372 , RIfcac130_6980, \9544 );
and \U$10251 ( \19373 , RIfc67b20_6202, \9546 );
and \U$10252 ( \19374 , RIfc67df0_6204, \9548 );
and \U$10253 ( \19375 , RIded9040_933, \9550 );
and \U$10254 ( \19376 , RIded6a48_906, \9552 );
and \U$10255 ( \19377 , RIded4b58_884, \9554 );
and \U$10256 ( \19378 , RIded26c8_858, \9556 );
and \U$10257 ( \19379 , RIdecfe00_829, \9558 );
and \U$10258 ( \19380 , RIdecd100_797, \9560 );
and \U$10259 ( \19381 , RIdeca400_765, \9562 );
and \U$10260 ( \19382 , RIdec7700_733, \9564 );
and \U$10261 ( \19383 , RIdeb3c00_509, \9566 );
and \U$10262 ( \19384 , RIde95228_317, \9568 );
and \U$10263 ( \19385 , RIe16d808_2623, \9570 );
and \U$10264 ( \19386 , RIe159600_2394, \9572 );
and \U$10265 ( \19387 , RIe142e00_2138, \9574 );
and \U$10266 ( \19388 , RIdf377f8_2008, \9576 );
and \U$10267 ( \19389 , RIdf2be58_1876, \9578 );
and \U$10268 ( \19390 , RIdf1c6d8_1700, \9580 );
and \U$10269 ( \19391 , RIdeffdd0_1375, \9582 );
and \U$10270 ( \19392 , RIdee68d0_1087, \9584 );
and \U$10271 ( \19393 , RIdedb638_960, \9586 );
and \U$10272 ( \19394 , RIde7b170_190, \9588 );
or \U$10273 ( \19395 , \19331 , \19332 , \19333 , \19334 , \19335 , \19336 , \19337 , \19338 , \19339 , \19340 , \19341 , \19342 , \19343 , \19344 , \19345 , \19346 , \19347 , \19348 , \19349 , \19350 , \19351 , \19352 , \19353 , \19354 , \19355 , \19356 , \19357 , \19358 , \19359 , \19360 , \19361 , \19362 , \19363 , \19364 , \19365 , \19366 , \19367 , \19368 , \19369 , \19370 , \19371 , \19372 , \19373 , \19374 , \19375 , \19376 , \19377 , \19378 , \19379 , \19380 , \19381 , \19382 , \19383 , \19384 , \19385 , \19386 , \19387 , \19388 , \19389 , \19390 , \19391 , \19392 , \19393 , \19394 );
or \U$10274 ( \19396 , \19330 , \19395 );
_DC g5461 ( \19397_nG5461 , \19396 , \9597 );
and \U$10275 ( \19398 , RIe19cc98_3161, \9059 );
and \U$10276 ( \19399 , RIe199f98_3129, \9061 );
and \U$10277 ( \19400 , RIfc73088_6331, \9063 );
and \U$10278 ( \19401 , RIe197298_3097, \9065 );
and \U$10279 ( \19402 , RIf1442a8_5235, \9067 );
and \U$10280 ( \19403 , RIe194598_3065, \9069 );
and \U$10281 ( \19404 , RIe191898_3033, \9071 );
and \U$10282 ( \19405 , RIe18eb98_3001, \9073 );
and \U$10283 ( \19406 , RIe189198_2937, \9075 );
and \U$10284 ( \19407 , RIe186498_2905, \9077 );
and \U$10285 ( \19408 , RIfc72278_6321, \9079 );
and \U$10286 ( \19409 , RIe183798_2873, \9081 );
and \U$10287 ( \19410 , RIfc61ce8_6135, \9083 );
and \U$10288 ( \19411 , RIe180a98_2841, \9085 );
and \U$10289 ( \19412 , RIe17dd98_2809, \9087 );
and \U$10290 ( \19413 , RIe17b098_2777, \9089 );
and \U$10291 ( \19414 , RIfcaf268_7015, \9091 );
and \U$10292 ( \19415 , RIfca6a00_6918, \9093 );
and \U$10293 ( \19416 , RIfcc9b18_7317, \9095 );
and \U$10294 ( \19417 , RIe175530_2712, \9097 );
and \U$10295 ( \19418 , RIfc72818_6325, \9099 );
and \U$10296 ( \19419 , RIfc726b0_6324, \9101 );
and \U$10297 ( \19420 , RIfccf7e8_7383, \9103 );
and \U$10298 ( \19421 , RIfc72548_6323, \9105 );
and \U$10299 ( \19422 , RIee3be48_5140, \9107 );
and \U$10300 ( \19423 , RIee3ad68_5128, \9109 );
and \U$10301 ( \19424 , RIfc71fa8_6319, \9111 );
and \U$10302 ( \19425 , RIe1730a0_2686, \9113 );
and \U$10303 ( \19426 , RIfcaef98_7013, \9115 );
and \U$10304 ( \19427 , RIfccf518_7381, \9117 );
and \U$10305 ( \19428 , RIfc71e40_6318, \9119 );
and \U$10306 ( \19429 , RIfc62120_6138, \9121 );
and \U$10307 ( \19430 , RIfe8b350_7928, \9123 );
and \U$10308 ( \19431 , RIe222ff0_4688, \9125 );
and \U$10309 ( \19432 , RIfcc9f50_7320, \9127 );
and \U$10310 ( \19433 , RIe2202f0_4656, \9129 );
and \U$10311 ( \19434 , RIfc4a570_5868, \9131 );
and \U$10312 ( \19435 , RIe21d5f0_4624, \9133 );
and \U$10313 ( \19436 , RIe217bf0_4560, \9135 );
and \U$10314 ( \19437 , RIe214ef0_4528, \9137 );
and \U$10315 ( \19438 , RIfccf3b0_7380, \9139 );
and \U$10316 ( \19439 , RIe2121f0_4496, \9141 );
and \U$10317 ( \19440 , RIf168ba8_5651, \9143 );
and \U$10318 ( \19441 , RIe20f4f0_4464, \9145 );
and \U$10319 ( \19442 , RIfc71300_6310, \9147 );
and \U$10320 ( \19443 , RIe20c7f0_4432, \9149 );
and \U$10321 ( \19444 , RIe209af0_4400, \9151 );
and \U$10322 ( \19445 , RIe206df0_4368, \9153 );
and \U$10323 ( \19446 , RIfc718a0_6314, \9155 );
and \U$10324 ( \19447 , RIfc71a08_6315, \9157 );
and \U$10325 ( \19448 , RIe202098_4313, \9159 );
and \U$10326 ( \19449 , RIfe8b1e8_7927, \9161 );
and \U$10327 ( \19450 , RIfc715d0_6312, \9163 );
and \U$10328 ( \19451 , RIfce6588_7643, \9165 );
and \U$10329 ( \19452 , RIfc62c60_6146, \9167 );
and \U$10330 ( \19453 , RIf161858_5569, \9169 );
and \U$10331 ( \19454 , RIf15fad0_5548, \9171 );
and \U$10332 ( \19455 , RIf15dbe0_5526, \9173 );
and \U$10333 ( \19456 , RIe1fc698_4249, \9175 );
and \U$10334 ( \19457 , RIfe8b4b8_7929, \9177 );
and \U$10335 ( \19458 , RIfcae5c0_7006, \9179 );
and \U$10336 ( \19459 , RIfc63098_6149, \9181 );
and \U$10337 ( \19460 , RIfc63200_6150, \9183 );
and \U$10338 ( \19461 , RIfc71198_6309, \9185 );
or \U$10339 ( \19462 , \19398 , \19399 , \19400 , \19401 , \19402 , \19403 , \19404 , \19405 , \19406 , \19407 , \19408 , \19409 , \19410 , \19411 , \19412 , \19413 , \19414 , \19415 , \19416 , \19417 , \19418 , \19419 , \19420 , \19421 , \19422 , \19423 , \19424 , \19425 , \19426 , \19427 , \19428 , \19429 , \19430 , \19431 , \19432 , \19433 , \19434 , \19435 , \19436 , \19437 , \19438 , \19439 , \19440 , \19441 , \19442 , \19443 , \19444 , \19445 , \19446 , \19447 , \19448 , \19449 , \19450 , \19451 , \19452 , \19453 , \19454 , \19455 , \19456 , \19457 , \19458 , \19459 , \19460 , \19461 );
and \U$10340 ( \19463 , RIf158a50_5468, \9188 );
and \U$10341 ( \19464 , RIf1576a0_5454, \9190 );
and \U$10342 ( \19465 , RIfcdc808_7531, \9192 );
and \U$10343 ( \19466 , RIfe8b620_7930, \9194 );
and \U$10344 ( \19467 , RIfc634d0_6152, \9196 );
and \U$10345 ( \19468 , RIfcceb40_7374, \9198 );
and \U$10346 ( \19469 , RIf154400_5418, \9200 );
and \U$10347 ( \19470 , RIe1f4da8_4163, \9202 );
and \U$10348 ( \19471 , RIf152c18_5401, \9204 );
and \U$10349 ( \19472 , RIf151868_5387, \9206 );
and \U$10350 ( \19473 , RIfc4d108_5899, \9208 );
and \U$10351 ( \19474 , RIe1f2a80_4138, \9210 );
and \U$10352 ( \19475 , RIfc70a90_6304, \9212 );
and \U$10353 ( \19476 , RIfc63bd8_6157, \9214 );
and \U$10354 ( \19477 , RIfca7810_6928, \9216 );
and \U$10355 ( \19478 , RIe1ed788_4079, \9218 );
and \U$10356 ( \19479 , RIe1ead58_4049, \9220 );
and \U$10357 ( \19480 , RIe1e8058_4017, \9222 );
and \U$10358 ( \19481 , RIe1e5358_3985, \9224 );
and \U$10359 ( \19482 , RIe1e2658_3953, \9226 );
and \U$10360 ( \19483 , RIe1df958_3921, \9228 );
and \U$10361 ( \19484 , RIe1dcc58_3889, \9230 );
and \U$10362 ( \19485 , RIe1d9f58_3857, \9232 );
and \U$10363 ( \19486 , RIe1d7258_3825, \9234 );
and \U$10364 ( \19487 , RIe1d1858_3761, \9236 );
and \U$10365 ( \19488 , RIe1ceb58_3729, \9238 );
and \U$10366 ( \19489 , RIe1cbe58_3697, \9240 );
and \U$10367 ( \19490 , RIe1c9158_3665, \9242 );
and \U$10368 ( \19491 , RIe1c6458_3633, \9244 );
and \U$10369 ( \19492 , RIe1c3758_3601, \9246 );
and \U$10370 ( \19493 , RIe1c0a58_3569, \9248 );
and \U$10371 ( \19494 , RIe1bdd58_3537, \9250 );
and \U$10372 ( \19495 , RIf14c408_5327, \9252 );
and \U$10373 ( \19496 , RIf14b1c0_5314, \9254 );
and \U$10374 ( \19497 , RIe1b8d30_3480, \9256 );
and \U$10375 ( \19498 , RIe1b6cd8_3457, \9258 );
and \U$10376 ( \19499 , RIfc707c0_6302, \9260 );
and \U$10377 ( \19500 , RIfca7c48_6931, \9262 );
and \U$10378 ( \19501 , RIe1b4de8_3435, \9264 );
and \U$10379 ( \19502 , RIe1b3a38_3421, \9266 );
and \U$10380 ( \19503 , RIfc70220_6298, \9268 );
and \U$10381 ( \19504 , RIfcce870_7372, \9270 );
and \U$10382 ( \19505 , RIe1b23b8_3405, \9272 );
and \U$10383 ( \19506 , RIe1b0630_3384, \9274 );
and \U$10384 ( \19507 , RIfc645b0_6164, \9276 );
and \U$10385 ( \19508 , RIfc700b8_6297, \9278 );
and \U$10386 ( \19509 , RIfeaac28_8259, \9280 );
and \U$10387 ( \19510 , RIe1aa690_3316, \9282 );
and \U$10388 ( \19511 , RIe1a8098_3289, \9284 );
and \U$10389 ( \19512 , RIe1a5398_3257, \9286 );
and \U$10390 ( \19513 , RIe1a2698_3225, \9288 );
and \U$10391 ( \19514 , RIe19f998_3193, \9290 );
and \U$10392 ( \19515 , RIe18be98_2969, \9292 );
and \U$10393 ( \19516 , RIe178398_2745, \9294 );
and \U$10394 ( \19517 , RIe225cf0_4720, \9296 );
and \U$10395 ( \19518 , RIe21a8f0_4592, \9298 );
and \U$10396 ( \19519 , RIe2040f0_4336, \9300 );
and \U$10397 ( \19520 , RIe1fe150_4268, \9302 );
and \U$10398 ( \19521 , RIe1f7508_4191, \9304 );
and \U$10399 ( \19522 , RIe1f0050_4108, \9306 );
and \U$10400 ( \19523 , RIe1d4558_3793, \9308 );
and \U$10401 ( \19524 , RIe1bb058_3505, \9310 );
and \U$10402 ( \19525 , RIe1aded0_3356, \9312 );
and \U$10403 ( \19526 , RIe170508_2655, \9314 );
or \U$10404 ( \19527 , \19463 , \19464 , \19465 , \19466 , \19467 , \19468 , \19469 , \19470 , \19471 , \19472 , \19473 , \19474 , \19475 , \19476 , \19477 , \19478 , \19479 , \19480 , \19481 , \19482 , \19483 , \19484 , \19485 , \19486 , \19487 , \19488 , \19489 , \19490 , \19491 , \19492 , \19493 , \19494 , \19495 , \19496 , \19497 , \19498 , \19499 , \19500 , \19501 , \19502 , \19503 , \19504 , \19505 , \19506 , \19507 , \19508 , \19509 , \19510 , \19511 , \19512 , \19513 , \19514 , \19515 , \19516 , \19517 , \19518 , \19519 , \19520 , \19521 , \19522 , \19523 , \19524 , \19525 , \19526 );
or \U$10405 ( \19528 , \19462 , \19527 );
_DC g54e5 ( \19529_nG54e5 , \19528 , \9323 );
xor g54e6 ( \19530_nG54e6 , \19397_nG5461 , \19529_nG54e5 );
buf \U$10406 ( \19531 , \19530_nG54e6 );
xor \U$10407 ( \19532 , \19531 , \19044 );
not \U$10408 ( \19533 , \19045 );
and \U$10409 ( \19534 , \19532 , \19533 );
and \U$10410 ( \19535 , \10687 , \19534 );
and \U$10411 ( \19536 , \10988 , \19045 );
nor \U$10412 ( \19537 , \19535 , \19536 );
and \U$10413 ( \19538 , \19044 , \18043 );
not \U$10414 ( \19539 , \19538 );
and \U$10415 ( \19540 , \19531 , \19539 );
xnor \U$10416 ( \19541 , \19537 , \19540 );
xor \U$10417 ( \19542 , \19265 , \19541 );
xor \U$10418 ( \19543 , \19256 , \19542 );
xor \U$10419 ( \19544 , \19237 , \19543 );
and \U$10420 ( \19545 , \19069 , \19073 );
and \U$10421 ( \19546 , \19073 , \19078 );
and \U$10422 ( \19547 , \19069 , \19078 );
or \U$10423 ( \19548 , \19545 , \19546 , \19547 );
and \U$10424 ( \19549 , \18760 , \18764 );
and \U$10425 ( \19550 , \18764 , \19047 );
and \U$10426 ( \19551 , \18760 , \19047 );
or \U$10427 ( \19552 , \19549 , \19550 , \19551 );
xor \U$10428 ( \19553 , \19548 , \19552 );
and \U$10429 ( \19554 , \19032 , \10983 );
_DC g65a4 ( \19555_nG65a4 , \19396 , \9597 );
_DC g65a5 ( \19556_nG65a5 , \19528 , \9323 );
and g65a6 ( \19557_nG65a6 , \19555_nG65a4 , \19556_nG65a5 );
buf \U$10430 ( \19558 , \19557_nG65a6 );
and \U$10431 ( \19559 , \19558 , \10691 );
nor \U$10432 ( \19560 , \19554 , \19559 );
xnor \U$10433 ( \19561 , \19560 , \10980 );
not \U$10434 ( \19562 , \19046 );
and \U$10435 ( \19563 , \19562 , \19540 );
xor \U$10436 ( \19564 , \19561 , \19563 );
and \U$10437 ( \19565 , \19035 , \19039 );
and \U$10438 ( \19566 , \19039 , \19046 );
and \U$10439 ( \19567 , \19035 , \19046 );
or \U$10440 ( \19568 , \19565 , \19566 , \19567 );
xor \U$10441 ( \19569 , \19564 , \19568 );
and \U$10442 ( \19570 , \11270 , \18090 );
and \U$10443 ( \19571 , \11586 , \17655 );
nor \U$10444 ( \19572 , \19570 , \19571 );
xnor \U$10445 ( \19573 , \19572 , \18046 );
xor \U$10446 ( \19574 , \19569 , \19573 );
xor \U$10447 ( \19575 , \19553 , \19574 );
xor \U$10448 ( \19576 , \19544 , \19575 );
and \U$10449 ( \19577 , \18756 , \19048 );
and \U$10450 ( \19578 , \19048 , \19080 );
and \U$10451 ( \19579 , \18756 , \19080 );
or \U$10452 ( \19580 , \19577 , \19578 , \19579 );
xor \U$10453 ( \19581 , \19576 , \19580 );
and \U$10454 ( \19582 , \19081 , \19085 );
and \U$10455 ( \19583 , \19086 , \19089 );
or \U$10456 ( \19584 , \19582 , \19583 );
xor \U$10457 ( \19585 , \19581 , \19584 );
buf g9be1 ( \19586_nG9be1 , \19585 );
and \U$10458 ( \19587 , \10704 , \19586_nG9be1 );
or \U$10459 ( \19588 , \19233 , \19587 );
xor \U$10460 ( \19589 , \10703 , \19588 );
buf \U$10461 ( \19590 , \19589 );
buf \U$10463 ( \19591 , \19590 );
xor \U$10464 ( \19592 , \19232 , \19591 );
buf \U$10465 ( \19593 , \19592 );
xor \U$10466 ( \19594 , \19186 , \19593 );
buf \U$10467 ( \19595 , \19594 );
xor \U$10468 ( \19596 , \19149 , \19595 );
and \U$10469 ( \19597 , \18719 , \19098 );
and \U$10470 ( \19598 , \18719 , \19132 );
and \U$10471 ( \19599 , \19098 , \19132 );
or \U$10472 ( \19600 , \19597 , \19598 , \19599 );
buf \U$10473 ( \19601 , \19600 );
xor \U$10474 ( \19602 , \19596 , \19601 );
and \U$10475 ( \19603 , \19144 , \19602 );
and \U$10476 ( \19604 , RIdec4cd0_703, \9059 );
and \U$10477 ( \19605 , RIdec1fd0_671, \9061 );
and \U$10478 ( \19606 , RIfc7b4b8_6425, \9063 );
and \U$10479 ( \19607 , RIdebf2d0_639, \9065 );
and \U$10480 ( \19608 , RIfc7b1e8_6423, \9067 );
and \U$10481 ( \19609 , RIdebc5d0_607, \9069 );
and \U$10482 ( \19610 , RIdeb98d0_575, \9071 );
and \U$10483 ( \19611 , RIdeb6bd0_543, \9073 );
and \U$10484 ( \19612 , RIfe83358_7837, \9075 );
and \U$10485 ( \19613 , RIdeb11d0_479, \9077 );
and \U$10486 ( \19614 , RIee1e5c8_4804, \9079 );
and \U$10487 ( \19615 , RIdeae4d0_447, \9081 );
and \U$10488 ( \19616 , RIfc437c0_5790, \9083 );
and \U$10489 ( \19617 , RIdea93b8_415, \9085 );
and \U$10490 ( \19618 , RIdea2ab8_383, \9087 );
and \U$10491 ( \19619 , RIde9c1b8_351, \9089 );
and \U$10492 ( \19620 , RIfc90ea8_6671, \9091 );
and \U$10493 ( \19621 , RIfc7af18_6421, \9093 );
and \U$10494 ( \19622 , RIfe83088_7835, \9095 );
and \U$10495 ( \19623 , RIee1a950_4761, \9097 );
and \U$10496 ( \19624 , RIde906b0_294, \9099 );
and \U$10497 ( \19625 , RIde8cba0_276, \9101 );
and \U$10498 ( \19626 , RIfe82f20_7834, \9103 );
and \U$10499 ( \19627 , RIfe82db8_7833, \9105 );
and \U$10500 ( \19628 , RIee1a248_4756, \9107 );
and \U$10501 ( \19629 , RIfe831f0_7836, \9109 );
and \U$10502 ( \19630 , RIfcc2390_7232, \9111 );
and \U$10503 ( \19631 , RIee195a0_4747, \9113 );
and \U$10504 ( \19632 , RIfcbe718_7189, \9115 );
and \U$10505 ( \19633 , RIfea9e18_8249, \9117 );
and \U$10506 ( \19634 , RIfc43220_5786, \9119 );
and \U$10507 ( \19635 , RIe167868_2555, \9121 );
and \U$10508 ( \19636 , RIe164cd0_2524, \9123 );
and \U$10509 ( \19637 , RIe161fd0_2492, \9125 );
and \U$10510 ( \19638 , RIee36f88_5084, \9127 );
and \U$10511 ( \19639 , RIe15f2d0_2460, \9129 );
and \U$10512 ( \19640 , RIee35ea8_5072, \9131 );
and \U$10513 ( \19641 , RIe15c5d0_2428, \9133 );
and \U$10514 ( \19642 , RIe156bd0_2364, \9135 );
and \U$10515 ( \19643 , RIe153ed0_2332, \9137 );
and \U$10516 ( \19644 , RIfe83628_7839, \9139 );
and \U$10517 ( \19645 , RIe1511d0_2300, \9141 );
and \U$10518 ( \19646 , RIfebfda8_8303, \9143 );
and \U$10519 ( \19647 , RIe14e4d0_2268, \9145 );
and \U$10520 ( \19648 , RIfebfc40_8302, \9147 );
and \U$10521 ( \19649 , RIe14b7d0_2236, \9149 );
and \U$10522 ( \19650 , RIe148ad0_2204, \9151 );
and \U$10523 ( \19651 , RIe145dd0_2172, \9153 );
and \U$10524 ( \19652 , RIee34120_5051, \9155 );
and \U$10525 ( \19653 , RIee32ed8_5038, \9157 );
and \U$10526 ( \19654 , RIee31df8_5026, \9159 );
and \U$10527 ( \19655 , RIfcc1f58_7229, \9161 );
and \U$10528 ( \19656 , RIe140ad8_2113, \9163 );
and \U$10529 ( \19657 , RIdf3e878_2088, \9165 );
and \U$10530 ( \19658 , RIfe834c0_7838, \9167 );
and \U$10531 ( \19659 , RIdf3a390_2039, \9169 );
and \U$10532 ( \19660 , RIfc5a6c8_6051, \9171 );
and \U$10533 ( \19661 , RIfc91e20_6682, \9173 );
and \U$10534 ( \19662 , RIee2e888_4988, \9175 );
and \U$10535 ( \19663 , RIfc96a10_6736, \9177 );
and \U$10536 ( \19664 , RIdf35098_1980, \9179 );
and \U$10537 ( \19665 , RIfeab600_8266, \9181 );
and \U$10538 ( \19666 , RIdf30bb0_1931, \9183 );
and \U$10539 ( \19667 , RIfeab768_8267, \9185 );
or \U$10540 ( \19668 , \19604 , \19605 , \19606 , \19607 , \19608 , \19609 , \19610 , \19611 , \19612 , \19613 , \19614 , \19615 , \19616 , \19617 , \19618 , \19619 , \19620 , \19621 , \19622 , \19623 , \19624 , \19625 , \19626 , \19627 , \19628 , \19629 , \19630 , \19631 , \19632 , \19633 , \19634 , \19635 , \19636 , \19637 , \19638 , \19639 , \19640 , \19641 , \19642 , \19643 , \19644 , \19645 , \19646 , \19647 , \19648 , \19649 , \19650 , \19651 , \19652 , \19653 , \19654 , \19655 , \19656 , \19657 , \19658 , \19659 , \19660 , \19661 , \19662 , \19663 , \19664 , \19665 , \19666 , \19667 );
and \U$10541 ( \19669 , RIfcbe9e8_7191, \9188 );
and \U$10542 ( \19670 , RIfc79fa0_6410, \9190 );
and \U$10543 ( \19671 , RIfc96740_6734, \9192 );
and \U$10544 ( \19672 , RIfc92258_6685, \9194 );
and \U$10545 ( \19673 , RIfea7118_8217, \9196 );
and \U$10546 ( \19674 , RIfea95a8_8243, \9198 );
and \U$10547 ( \19675 , RIdf26020_1809, \9200 );
and \U$10548 ( \19676 , RIdf24400_1789, \9202 );
and \U$10549 ( \19677 , RIfc79a00_6406, \9204 );
and \U$10550 ( \19678 , RIfc5add0_6056, \9206 );
and \U$10551 ( \19679 , RIfce5d18_7637, \9208 );
and \U$10552 ( \19680 , RIfc92690_6688, \9210 );
and \U$10553 ( \19681 , RIfce3018_7605, \9212 );
and \U$10554 ( \19682 , RIdf1f270_1731, \9214 );
and \U$10555 ( \19683 , RIfc79730_6404, \9216 );
and \U$10556 ( \19684 , RIdf19000_1661, \9218 );
and \U$10557 ( \19685 , RIdf168a0_1633, \9220 );
and \U$10558 ( \19686 , RIdf13ba0_1601, \9222 );
and \U$10559 ( \19687 , RIdf10ea0_1569, \9224 );
and \U$10560 ( \19688 , RIdf0e1a0_1537, \9226 );
and \U$10561 ( \19689 , RIdf0b4a0_1505, \9228 );
and \U$10562 ( \19690 , RIdf087a0_1473, \9230 );
and \U$10563 ( \19691 , RIdf05aa0_1441, \9232 );
and \U$10564 ( \19692 , RIdf02da0_1409, \9234 );
and \U$10565 ( \19693 , RIdefd3a0_1345, \9236 );
and \U$10566 ( \19694 , RIdefa6a0_1313, \9238 );
and \U$10567 ( \19695 , RIdef79a0_1281, \9240 );
and \U$10568 ( \19696 , RIdef4ca0_1249, \9242 );
and \U$10569 ( \19697 , RIdef1fa0_1217, \9244 );
and \U$10570 ( \19698 , RIdeef2a0_1185, \9246 );
and \U$10571 ( \19699 , RIdeec5a0_1153, \9248 );
and \U$10572 ( \19700 , RIdee98a0_1121, \9250 );
and \U$10573 ( \19701 , RIfc5b7a8_6063, \9252 );
and \U$10574 ( \19702 , RIfc5b640_6062, \9254 );
and \U$10575 ( \19703 , RIfc931d0_6696, \9256 );
and \U$10576 ( \19704 , RIfcecac8_7715, \9258 );
and \U$10577 ( \19705 , RIdee4710_1063, \9260 );
and \U$10578 ( \19706 , RIdee26b8_1040, \9262 );
and \U$10579 ( \19707 , RIdee07c8_1018, \9264 );
and \U$10580 ( \19708 , RIdede4a0_993, \9266 );
and \U$10581 ( \19709 , RIfcbf0f0_7196, \9268 );
and \U$10582 ( \19710 , RIfcbf528_7199, \9270 );
and \U$10583 ( \19711 , RIfc792f8_6401, \9272 );
and \U$10584 ( \19712 , RIfc93068_6695, \9274 );
and \U$10585 ( \19713 , RIded91a8_934, \9276 );
and \U$10586 ( \19714 , RIded6d18_908, \9278 );
and \U$10587 ( \19715 , RIded4e28_886, \9280 );
and \U$10588 ( \19716 , RIded2998_860, \9282 );
and \U$10589 ( \19717 , RIded00d0_831, \9284 );
and \U$10590 ( \19718 , RIdecd3d0_799, \9286 );
and \U$10591 ( \19719 , RIdeca6d0_767, \9288 );
and \U$10592 ( \19720 , RIdec79d0_735, \9290 );
and \U$10593 ( \19721 , RIdeb3ed0_511, \9292 );
and \U$10594 ( \19722 , RIde958b8_319, \9294 );
and \U$10595 ( \19723 , RIe16dad8_2625, \9296 );
and \U$10596 ( \19724 , RIe1598d0_2396, \9298 );
and \U$10597 ( \19725 , RIe1430d0_2140, \9300 );
and \U$10598 ( \19726 , RIdf37ac8_2010, \9302 );
and \U$10599 ( \19727 , RIdf2c128_1878, \9304 );
and \U$10600 ( \19728 , RIdf1c9a8_1702, \9306 );
and \U$10601 ( \19729 , RIdf000a0_1377, \9308 );
and \U$10602 ( \19730 , RIdee6ba0_1089, \9310 );
and \U$10603 ( \19731 , RIdedb908_962, \9312 );
and \U$10604 ( \19732 , RIde7b800_192, \9314 );
or \U$10605 ( \19733 , \19669 , \19670 , \19671 , \19672 , \19673 , \19674 , \19675 , \19676 , \19677 , \19678 , \19679 , \19680 , \19681 , \19682 , \19683 , \19684 , \19685 , \19686 , \19687 , \19688 , \19689 , \19690 , \19691 , \19692 , \19693 , \19694 , \19695 , \19696 , \19697 , \19698 , \19699 , \19700 , \19701 , \19702 , \19703 , \19704 , \19705 , \19706 , \19707 , \19708 , \19709 , \19710 , \19711 , \19712 , \19713 , \19714 , \19715 , \19716 , \19717 , \19718 , \19719 , \19720 , \19721 , \19722 , \19723 , \19724 , \19725 , \19726 , \19727 , \19728 , \19729 , \19730 , \19731 , \19732 );
or \U$10606 ( \19734 , \19668 , \19733 );
_DC g297b ( \19735_nG297b , \19734 , \9323 );
buf \U$10607 ( \19736 , \19735_nG297b );
and \U$10608 ( \19737 , RIe19cf68_3163, \9333 );
and \U$10609 ( \19738 , RIe19a268_3131, \9335 );
and \U$10610 ( \19739 , RIfc8d7d0_6632, \9337 );
and \U$10611 ( \19740 , RIe197568_3099, \9339 );
and \U$10612 ( \19741 , RIfc561e0_6002, \9341 );
and \U$10613 ( \19742 , RIe194868_3067, \9343 );
and \U$10614 ( \19743 , RIe191b68_3035, \9345 );
and \U$10615 ( \19744 , RIe18ee68_3003, \9347 );
and \U$10616 ( \19745 , RIe189468_2939, \9349 );
and \U$10617 ( \19746 , RIe186768_2907, \9351 );
and \U$10618 ( \19747 , RIf143330_5224, \9353 );
and \U$10619 ( \19748 , RIe183a68_2875, \9355 );
and \U$10620 ( \19749 , RIfc7d948_6451, \9357 );
and \U$10621 ( \19750 , RIe180d68_2843, \9359 );
and \U$10622 ( \19751 , RIe17e068_2811, \9361 );
and \U$10623 ( \19752 , RIe17b368_2779, \9363 );
and \U$10624 ( \19753 , RIfc564b0_6004, \9365 );
and \U$10625 ( \19754 , RIfcd6700_7462, \9367 );
and \U$10626 ( \19755 , RIfc461f0_5820, \9369 );
and \U$10627 ( \19756 , RIe175698_2713, \9371 );
and \U$10628 ( \19757 , RIfc46088_5819, \9373 );
and \U$10629 ( \19758 , RIfc45f20_5818, \9375 );
and \U$10630 ( \19759 , RIfc7dc18_6453, \9377 );
and \U$10631 ( \19760 , RIfcd69d0_7464, \9379 );
and \U$10632 ( \19761 , RIfc98630_6756, \9381 );
and \U$10633 ( \19762 , RIfcc2a98_7237, \9383 );
and \U$10634 ( \19763 , RIfc7d510_6448, \9385 );
and \U$10635 ( \19764 , RIe173208_2687, \9387 );
and \U$10636 ( \19765 , RIfc8e478_6641, \9389 );
and \U$10637 ( \19766 , RIfc45ae8_5815, \9391 );
and \U$10638 ( \19767 , RIfc8e8b0_6644, \9393 );
and \U$10639 ( \19768 , RIfc45980_5814, \9395 );
and \U$10640 ( \19769 , RIfe82ae8_7831, \9397 );
and \U$10641 ( \19770 , RIe2232c0_4690, \9399 );
and \U$10642 ( \19771 , RIf16ba10_5684, \9401 );
and \U$10643 ( \19772 , RIe2205c0_4658, \9403 );
and \U$10644 ( \19773 , RIfcd24e8_7415, \9405 );
and \U$10645 ( \19774 , RIe21d8c0_4626, \9407 );
and \U$10646 ( \19775 , RIe217ec0_4562, \9409 );
and \U$10647 ( \19776 , RIe2151c0_4530, \9411 );
and \U$10648 ( \19777 , RIfebf268_8295, \9413 );
and \U$10649 ( \19778 , RIe2124c0_4498, \9415 );
and \U$10650 ( \19779 , RIf168d10_5652, \9417 );
and \U$10651 ( \19780 , RIe20f7c0_4466, \9419 );
and \U$10652 ( \19781 , RIfc7d240_6446, \9421 );
and \U$10653 ( \19782 , RIe20cac0_4434, \9423 );
and \U$10654 ( \19783 , RIe209dc0_4402, \9425 );
and \U$10655 ( \19784 , RIe2070c0_4370, \9427 );
and \U$10656 ( \19785 , RIf166e20_5630, \9429 );
and \U$10657 ( \19786 , RIfebf6a0_8298, \9431 );
and \U$10658 ( \19787 , RIfebf808_8299, \9433 );
and \U$10659 ( \19788 , RIfebf538_8297, \9435 );
and \U$10660 ( \19789 , RIfc8eb80_6646, \9437 );
and \U$10661 ( \19790 , RIf164120_5598, \9439 );
and \U$10662 ( \19791 , RIfc453e0_5810, \9441 );
and \U$10663 ( \19792 , RIf161b28_5571, \9443 );
and \U$10664 ( \19793 , RIf15fc38_5549, \9445 );
and \U$10665 ( \19794 , RIf15dd48_5527, \9447 );
and \U$10666 ( \19795 , RIe1fc968_4251, \9449 );
and \U$10667 ( \19796 , RIe1fb888_4239, \9451 );
and \U$10668 ( \19797 , RIfebf3d0_8296, \9453 );
and \U$10669 ( \19798 , RIf15b318_5497, \9455 );
and \U$10670 ( \19799 , RIfca2518_6869, \9457 );
and \U$10671 ( \19800 , RIfc8f120_6650, \9459 );
or \U$10672 ( \19801 , \19737 , \19738 , \19739 , \19740 , \19741 , \19742 , \19743 , \19744 , \19745 , \19746 , \19747 , \19748 , \19749 , \19750 , \19751 , \19752 , \19753 , \19754 , \19755 , \19756 , \19757 , \19758 , \19759 , \19760 , \19761 , \19762 , \19763 , \19764 , \19765 , \19766 , \19767 , \19768 , \19769 , \19770 , \19771 , \19772 , \19773 , \19774 , \19775 , \19776 , \19777 , \19778 , \19779 , \19780 , \19781 , \19782 , \19783 , \19784 , \19785 , \19786 , \19787 , \19788 , \19789 , \19790 , \19791 , \19792 , \19793 , \19794 , \19795 , \19796 , \19797 , \19798 , \19799 , \19800 );
and \U$10673 ( \19802 , RIfebfad8_8301, \9462 );
and \U$10674 ( \19803 , RIfebf970_8300, \9464 );
and \U$10675 ( \19804 , RIfc7cca0_6442, \9466 );
and \U$10676 ( \19805 , RIe1f9dd0_4220, \9468 );
and \U$10677 ( \19806 , RIfe82c50_7832, \9470 );
and \U$10678 ( \19807 , RIf155648_5431, \9472 );
and \U$10679 ( \19808 , RIfc8f288_6651, \9474 );
and \U$10680 ( \19809 , RIe1f4f10_4164, \9476 );
and \U$10681 ( \19810 , RIf152d80_5402, \9478 );
and \U$10682 ( \19811 , RIfc8f828_6655, \9480 );
and \U$10683 ( \19812 , RIfcb3b88_7067, \9482 );
and \U$10684 ( \19813 , RIe1f2d50_4140, \9484 );
and \U$10685 ( \19814 , RIfc445d0_5800, \9486 );
and \U$10686 ( \19815 , RIfc8faf8_6657, \9488 );
and \U$10687 ( \19816 , RIf14da88_5343, \9490 );
and \U$10688 ( \19817 , RIe1eda58_4081, \9492 );
and \U$10689 ( \19818 , RIe1eb028_4051, \9494 );
and \U$10690 ( \19819 , RIe1e8328_4019, \9496 );
and \U$10691 ( \19820 , RIe1e5628_3987, \9498 );
and \U$10692 ( \19821 , RIe1e2928_3955, \9500 );
and \U$10693 ( \19822 , RIe1dfc28_3923, \9502 );
and \U$10694 ( \19823 , RIe1dcf28_3891, \9504 );
and \U$10695 ( \19824 , RIe1da228_3859, \9506 );
and \U$10696 ( \19825 , RIe1d7528_3827, \9508 );
and \U$10697 ( \19826 , RIe1d1b28_3763, \9510 );
and \U$10698 ( \19827 , RIe1cee28_3731, \9512 );
and \U$10699 ( \19828 , RIe1cc128_3699, \9514 );
and \U$10700 ( \19829 , RIe1c9428_3667, \9516 );
and \U$10701 ( \19830 , RIe1c6728_3635, \9518 );
and \U$10702 ( \19831 , RIe1c3a28_3603, \9520 );
and \U$10703 ( \19832 , RIe1c0d28_3571, \9522 );
and \U$10704 ( \19833 , RIe1be028_3539, \9524 );
and \U$10705 ( \19834 , RIfc7bff8_6433, \9526 );
and \U$10706 ( \19835 , RIfc44030_5796, \9528 );
and \U$10707 ( \19836 , RIe1b9000_3482, \9530 );
and \U$10708 ( \19837 , RIe1b6fa8_3459, \9532 );
and \U$10709 ( \19838 , RIfcbdd40_7182, \9534 );
and \U$10710 ( \19839 , RIfc8ff30_6660, \9536 );
and \U$10711 ( \19840 , RIe1b50b8_3437, \9538 );
and \U$10712 ( \19841 , RIe1b3d08_3423, \9540 );
and \U$10713 ( \19842 , RIfcbe178_7185, \9542 );
and \U$10714 ( \19843 , RIfc43d60_5794, \9544 );
and \U$10715 ( \19844 , RIe1b2520_3406, \9546 );
and \U$10716 ( \19845 , RIe1b0798_3385, \9548 );
and \U$10717 ( \19846 , RIfcdb5c0_7518, \9550 );
and \U$10718 ( \19847 , RIfc7ba58_6429, \9552 );
and \U$10719 ( \19848 , RIe1ac148_3335, \9554 );
and \U$10720 ( \19849 , RIe1aa960_3318, \9556 );
and \U$10721 ( \19850 , RIe1a8368_3291, \9558 );
and \U$10722 ( \19851 , RIe1a5668_3259, \9560 );
and \U$10723 ( \19852 , RIe1a2968_3227, \9562 );
and \U$10724 ( \19853 , RIe19fc68_3195, \9564 );
and \U$10725 ( \19854 , RIe18c168_2971, \9566 );
and \U$10726 ( \19855 , RIe178668_2747, \9568 );
and \U$10727 ( \19856 , RIe225fc0_4722, \9570 );
and \U$10728 ( \19857 , RIe21abc0_4594, \9572 );
and \U$10729 ( \19858 , RIe2043c0_4338, \9574 );
and \U$10730 ( \19859 , RIe1fe420_4270, \9576 );
and \U$10731 ( \19860 , RIe1f77d8_4193, \9578 );
and \U$10732 ( \19861 , RIe1f0320_4110, \9580 );
and \U$10733 ( \19862 , RIe1d4828_3795, \9582 );
and \U$10734 ( \19863 , RIe1bb328_3507, \9584 );
and \U$10735 ( \19864 , RIe1ae1a0_3358, \9586 );
and \U$10736 ( \19865 , RIe1707d8_2657, \9588 );
or \U$10737 ( \19866 , \19802 , \19803 , \19804 , \19805 , \19806 , \19807 , \19808 , \19809 , \19810 , \19811 , \19812 , \19813 , \19814 , \19815 , \19816 , \19817 , \19818 , \19819 , \19820 , \19821 , \19822 , \19823 , \19824 , \19825 , \19826 , \19827 , \19828 , \19829 , \19830 , \19831 , \19832 , \19833 , \19834 , \19835 , \19836 , \19837 , \19838 , \19839 , \19840 , \19841 , \19842 , \19843 , \19844 , \19845 , \19846 , \19847 , \19848 , \19849 , \19850 , \19851 , \19852 , \19853 , \19854 , \19855 , \19856 , \19857 , \19858 , \19859 , \19860 , \19861 , \19862 , \19863 , \19864 , \19865 );
or \U$10738 ( \19867 , \19801 , \19866 );
_DC g3aa8 ( \19868_nG3aa8 , \19867 , \9597 );
buf \U$10739 ( \19869 , \19868_nG3aa8 );
xor \U$10740 ( \19870 , \19736 , \19869 );
and \U$10741 ( \19871 , RIdec4b68_702, \9059 );
and \U$10742 ( \19872 , RIdec1e68_670, \9061 );
and \U$10743 ( \19873 , RIfc5df08_6091, \9063 );
and \U$10744 ( \19874 , RIdebf168_638, \9065 );
and \U$10745 ( \19875 , RIfce6df8_7649, \9067 );
and \U$10746 ( \19876 , RIdebc468_606, \9069 );
and \U$10747 ( \19877 , RIdeb9768_574, \9071 );
and \U$10748 ( \19878 , RIdeb6a68_542, \9073 );
and \U$10749 ( \19879 , RIfc75ef0_6364, \9075 );
and \U$10750 ( \19880 , RIdeb1068_478, \9077 );
and \U$10751 ( \19881 , RIfcc12b0_7220, \9079 );
and \U$10752 ( \19882 , RIdeae368_446, \9081 );
and \U$10753 ( \19883 , RIfc5e340_6094, \9083 );
and \U$10754 ( \19884 , RIdea9070_414, \9085 );
and \U$10755 ( \19885 , RIdea2770_382, \9087 );
and \U$10756 ( \19886 , RIde9be70_350, \9089 );
and \U$10757 ( \19887 , RIfced4a0_7722, \9091 );
and \U$10758 ( \19888 , RIfcc1418_7221, \9093 );
and \U$10759 ( \19889 , RIfc95930_6724, \9095 );
and \U$10760 ( \19890 , RIfcec0f0_7708, \9097 );
and \U$10761 ( \19891 , RIde90368_293, \9099 );
and \U$10762 ( \19892 , RIde8c858_275, \9101 );
and \U$10763 ( \19893 , RIde893d8_259, \9103 );
and \U$10764 ( \19894 , RIde84ef0_238, \9105 );
and \U$10765 ( \19895 , RIde80d50_218, \9107 );
and \U$10766 ( \19896 , RIfc95a98_6725, \9109 );
and \U$10767 ( \19897 , RIfced068_7719, \9111 );
and \U$10768 ( \19898 , RIfced1d0_7720, \9113 );
and \U$10769 ( \19899 , RIfcedfe0_7730, \9115 );
and \U$10770 ( \19900 , RIe16b0a8_2595, \9117 );
and \U$10771 ( \19901 , RIe169758_2577, \9119 );
and \U$10772 ( \19902 , RIe167700_2554, \9121 );
and \U$10773 ( \19903 , RIe164b68_2523, \9123 );
and \U$10774 ( \19904 , RIe161e68_2491, \9125 );
and \U$10775 ( \19905 , RIee36e20_5083, \9127 );
and \U$10776 ( \19906 , RIe15f168_2459, \9129 );
and \U$10777 ( \19907 , RIfc426e0_5778, \9131 );
and \U$10778 ( \19908 , RIe15c468_2427, \9133 );
and \U$10779 ( \19909 , RIe156a68_2363, \9135 );
and \U$10780 ( \19910 , RIe153d68_2331, \9137 );
and \U$10781 ( \19911 , RIfe82818_7829, \9139 );
and \U$10782 ( \19912 , RIe151068_2299, \9141 );
and \U$10783 ( \19913 , RIee34c60_5059, \9143 );
and \U$10784 ( \19914 , RIe14e368_2267, \9145 );
and \U$10785 ( \19915 , RIfc5f9c0_6110, \9147 );
and \U$10786 ( \19916 , RIe14b668_2235, \9149 );
and \U$10787 ( \19917 , RIe148968_2203, \9151 );
and \U$10788 ( \19918 , RIe145c68_2171, \9153 );
and \U$10789 ( \19919 , RIfccfef0_7388, \9155 );
and \U$10790 ( \19920 , RIfca57b8_6905, \9157 );
and \U$10791 ( \19921 , RIfc600c8_6115, \9159 );
and \U$10792 ( \19922 , RIfcafda8_7023, \9161 );
and \U$10793 ( \19923 , RIe140970_2112, \9163 );
and \U$10794 ( \19924 , RIdf3e710_2087, \9165 );
and \U$10795 ( \19925 , RIdf3c6b8_2064, \9167 );
and \U$10796 ( \19926 , RIdf3a228_2038, \9169 );
and \U$10797 ( \19927 , RIfc5fc90_6112, \9171 );
and \U$10798 ( \19928 , RIee2f3c8_4996, \9173 );
and \U$10799 ( \19929 , RIfc742d0_6344, \9175 );
and \U$10800 ( \19930 , RIee2d208_4972, \9177 );
and \U$10801 ( \19931 , RIdf34f30_1979, \9179 );
and \U$10802 ( \19932 , RIfebf100_8294, \9181 );
and \U$10803 ( \19933 , RIdf30a48_1930, \9183 );
and \U$10804 ( \19934 , RIdf2ecc0_1909, \9185 );
or \U$10805 ( \19935 , \19871 , \19872 , \19873 , \19874 , \19875 , \19876 , \19877 , \19878 , \19879 , \19880 , \19881 , \19882 , \19883 , \19884 , \19885 , \19886 , \19887 , \19888 , \19889 , \19890 , \19891 , \19892 , \19893 , \19894 , \19895 , \19896 , \19897 , \19898 , \19899 , \19900 , \19901 , \19902 , \19903 , \19904 , \19905 , \19906 , \19907 , \19908 , \19909 , \19910 , \19911 , \19912 , \19913 , \19914 , \19915 , \19916 , \19917 , \19918 , \19919 , \19920 , \19921 , \19922 , \19923 , \19924 , \19925 , \19926 , \19927 , \19928 , \19929 , \19930 , \19931 , \19932 , \19933 , \19934 );
and \U$10806 ( \19936 , RIfcb08e8_7031, \9188 );
and \U$10807 ( \19937 , RIfcee418_7733, \9190 );
and \U$10808 ( \19938 , RIfc95ed0_6728, \9192 );
and \U$10809 ( \19939 , RIfcdef68_7559, \9194 );
and \U$10810 ( \19940 , RIdf29e00_1853, \9196 );
and \U$10811 ( \19941 , RIdf27c40_1829, \9198 );
and \U$10812 ( \19942 , RIdf25eb8_1808, \9200 );
and \U$10813 ( \19943 , RIdf24298_1788, \9202 );
and \U$10814 ( \19944 , RIfc5ed18_6101, \9204 );
and \U$10815 ( \19945 , RIfcee850_7736, \9206 );
and \U$10816 ( \19946 , RIdf227e0_1769, \9208 );
and \U$10817 ( \19947 , RIfc5efe8_6103, \9210 );
and \U$10818 ( \19948 , RIdf212c8_1754, \9212 );
and \U$10819 ( \19949 , RIfeaa520_8254, \9214 );
and \U$10820 ( \19950 , RIdf1ad88_1682, \9216 );
and \U$10821 ( \19951 , RIdf18e98_1660, \9218 );
and \U$10822 ( \19952 , RIdf16738_1632, \9220 );
and \U$10823 ( \19953 , RIdf13a38_1600, \9222 );
and \U$10824 ( \19954 , RIdf10d38_1568, \9224 );
and \U$10825 ( \19955 , RIdf0e038_1536, \9226 );
and \U$10826 ( \19956 , RIdf0b338_1504, \9228 );
and \U$10827 ( \19957 , RIdf08638_1472, \9230 );
and \U$10828 ( \19958 , RIdf05938_1440, \9232 );
and \U$10829 ( \19959 , RIdf02c38_1408, \9234 );
and \U$10830 ( \19960 , RIdefd238_1344, \9236 );
and \U$10831 ( \19961 , RIdefa538_1312, \9238 );
and \U$10832 ( \19962 , RIdef7838_1280, \9240 );
and \U$10833 ( \19963 , RIdef4b38_1248, \9242 );
and \U$10834 ( \19964 , RIdef1e38_1216, \9244 );
and \U$10835 ( \19965 , RIdeef138_1184, \9246 );
and \U$10836 ( \19966 , RIdeec438_1152, \9248 );
and \U$10837 ( \19967 , RIdee9738_1120, \9250 );
and \U$10838 ( \19968 , RIfcc96e0_7314, \9252 );
and \U$10839 ( \19969 , RIfccfd88_7387, \9254 );
and \U$10840 ( \19970 , RIfc60aa0_6122, \9256 );
and \U$10841 ( \19971 , RIfca5ec0_6910, \9258 );
and \U$10842 ( \19972 , RIdee45a8_1062, \9260 );
and \U$10843 ( \19973 , RIdee2550_1039, \9262 );
and \U$10844 ( \19974 , RIdee0660_1017, \9264 );
and \U$10845 ( \19975 , RIfe826b0_7828, \9266 );
and \U$10846 ( \19976 , RIfcdeb30_7556, \9268 );
and \U$10847 ( \19977 , RIfc73bc8_6339, \9270 );
and \U$10848 ( \19978 , RIfca5bf0_6908, \9272 );
and \U$10849 ( \19979 , RIfc73a60_6338, \9274 );
and \U$10850 ( \19980 , RIfe82980_7830, \9276 );
and \U$10851 ( \19981 , RIded6bb0_907, \9278 );
and \U$10852 ( \19982 , RIded4cc0_885, \9280 );
and \U$10853 ( \19983 , RIded2830_859, \9282 );
and \U$10854 ( \19984 , RIdecff68_830, \9284 );
and \U$10855 ( \19985 , RIdecd268_798, \9286 );
and \U$10856 ( \19986 , RIdeca568_766, \9288 );
and \U$10857 ( \19987 , RIdec7868_734, \9290 );
and \U$10858 ( \19988 , RIdeb3d68_510, \9292 );
and \U$10859 ( \19989 , RIde95570_318, \9294 );
and \U$10860 ( \19990 , RIe16d970_2624, \9296 );
and \U$10861 ( \19991 , RIe159768_2395, \9298 );
and \U$10862 ( \19992 , RIe142f68_2139, \9300 );
and \U$10863 ( \19993 , RIdf37960_2009, \9302 );
and \U$10864 ( \19994 , RIdf2bfc0_1877, \9304 );
and \U$10865 ( \19995 , RIdf1c840_1701, \9306 );
and \U$10866 ( \19996 , RIdefff38_1376, \9308 );
and \U$10867 ( \19997 , RIdee6a38_1088, \9310 );
and \U$10868 ( \19998 , RIdedb7a0_961, \9312 );
and \U$10869 ( \19999 , RIde7b4b8_191, \9314 );
or \U$10870 ( \20000 , \19936 , \19937 , \19938 , \19939 , \19940 , \19941 , \19942 , \19943 , \19944 , \19945 , \19946 , \19947 , \19948 , \19949 , \19950 , \19951 , \19952 , \19953 , \19954 , \19955 , \19956 , \19957 , \19958 , \19959 , \19960 , \19961 , \19962 , \19963 , \19964 , \19965 , \19966 , \19967 , \19968 , \19969 , \19970 , \19971 , \19972 , \19973 , \19974 , \19975 , \19976 , \19977 , \19978 , \19979 , \19980 , \19981 , \19982 , \19983 , \19984 , \19985 , \19986 , \19987 , \19988 , \19989 , \19990 , \19991 , \19992 , \19993 , \19994 , \19995 , \19996 , \19997 , \19998 , \19999 );
or \U$10871 ( \20001 , \19935 , \20000 );
_DC g2a00 ( \20002_nG2a00 , \20001 , \9323 );
buf \U$10872 ( \20003 , \20002_nG2a00 );
and \U$10873 ( \20004 , RIe19ce00_3162, \9333 );
and \U$10874 ( \20005 , RIe19a100_3130, \9335 );
and \U$10875 ( \20006 , RIfce96c0_7678, \9337 );
and \U$10876 ( \20007 , RIe197400_3098, \9339 );
and \U$10877 ( \20008 , RIf144410_5236, \9341 );
and \U$10878 ( \20009 , RIe194700_3066, \9343 );
and \U$10879 ( \20010 , RIe191a00_3034, \9345 );
and \U$10880 ( \20011 , RIe18ed00_3002, \9347 );
and \U$10881 ( \20012 , RIe189300_2938, \9349 );
and \U$10882 ( \20013 , RIe186600_2906, \9351 );
and \U$10883 ( \20014 , RIfebee30_8292, \9353 );
and \U$10884 ( \20015 , RIe183900_2874, \9355 );
and \U$10885 ( \20016 , RIfcdbcc8_7523, \9357 );
and \U$10886 ( \20017 , RIe180c00_2842, \9359 );
and \U$10887 ( \20018 , RIe17df00_2810, \9361 );
and \U$10888 ( \20019 , RIe17b200_2778, \9363 );
and \U$10889 ( \20020 , RIf141f80_5210, \9365 );
and \U$10890 ( \20021 , RIfce7398_7653, \9367 );
and \U$10891 ( \20022 , RIfcb1e00_7046, \9369 );
and \U$10892 ( \20023 , RIfe82548_7827, \9371 );
and \U$10893 ( \20024 , RIfca42a0_6890, \9373 );
and \U$10894 ( \20025 , RIfcbff00_7206, \9375 );
and \U$10895 ( \20026 , RIfcaaee8_6967, \9377 );
and \U$10896 ( \20027 , RIee3d090_5153, \9379 );
and \U$10897 ( \20028 , RIfc5c180_6070, \9381 );
and \U$10898 ( \20029 , RIfce35b8_7609, \9383 );
and \U$10899 ( \20030 , RIee399b8_5114, \9385 );
and \U$10900 ( \20031 , RIfea8a68_8235, \9387 );
and \U$10901 ( \20032 , RIf16fef8_5733, \9389 );
and \U$10902 ( \20033 , RIfebecc8_8291, \9391 );
and \U$10903 ( \20034 , RIfc5c450_6072, \9393 );
and \U$10904 ( \20035 , RIfce9288_7675, \9395 );
and \U$10905 ( \20036 , RIfc40778_5759, \9397 );
and \U$10906 ( \20037 , RIe223158_4689, \9399 );
and \U$10907 ( \20038 , RIfce77d0_7656, \9401 );
and \U$10908 ( \20039 , RIe220458_4657, \9403 );
and \U$10909 ( \20040 , RIfce24d8_7597, \9405 );
and \U$10910 ( \20041 , RIe21d758_4625, \9407 );
and \U$10911 ( \20042 , RIe217d58_4561, \9409 );
and \U$10912 ( \20043 , RIe215058_4529, \9411 );
and \U$10913 ( \20044 , RIfce8a18_7669, \9413 );
and \U$10914 ( \20045 , RIe212358_4497, \9415 );
and \U$10915 ( \20046 , RIfce1998_7589, \9417 );
and \U$10916 ( \20047 , RIe20f658_4465, \9419 );
and \U$10917 ( \20048 , RIfc77840_6382, \9421 );
and \U$10918 ( \20049 , RIe20c958_4433, \9423 );
and \U$10919 ( \20050 , RIe209c58_4401, \9425 );
and \U$10920 ( \20051 , RIe206f58_4369, \9427 );
and \U$10921 ( \20052 , RIf166cb8_5629, \9429 );
and \U$10922 ( \20053 , RIf165bd8_5617, \9431 );
and \U$10923 ( \20054 , RIfe81fa8_7823, \9433 );
and \U$10924 ( \20055 , RIfe81e40_7822, \9435 );
and \U$10925 ( \20056 , RIfc5c888_6075, \9437 );
and \U$10926 ( \20057 , RIfceb178_7697, \9439 );
and \U$10927 ( \20058 , RIf1631a8_5587, \9441 );
and \U$10928 ( \20059 , RIf1619c0_5570, \9443 );
and \U$10929 ( \20060 , RIfccf248_7379, \9445 );
and \U$10930 ( \20061 , RIfc77570_6380, \9447 );
and \U$10931 ( \20062 , RIe1fc800_4250, \9449 );
and \U$10932 ( \20063 , RIe1fb720_4238, \9451 );
and \U$10933 ( \20064 , RIf15c830_5512, \9453 );
and \U$10934 ( \20065 , RIf15b1b0_5496, \9455 );
and \U$10935 ( \20066 , RIfcd0fd0_7400, \9457 );
and \U$10936 ( \20067 , RIfccc6b0_7348, \9459 );
or \U$10937 ( \20068 , \20004 , \20005 , \20006 , \20007 , \20008 , \20009 , \20010 , \20011 , \20012 , \20013 , \20014 , \20015 , \20016 , \20017 , \20018 , \20019 , \20020 , \20021 , \20022 , \20023 , \20024 , \20025 , \20026 , \20027 , \20028 , \20029 , \20030 , \20031 , \20032 , \20033 , \20034 , \20035 , \20036 , \20037 , \20038 , \20039 , \20040 , \20041 , \20042 , \20043 , \20044 , \20045 , \20046 , \20047 , \20048 , \20049 , \20050 , \20051 , \20052 , \20053 , \20054 , \20055 , \20056 , \20057 , \20058 , \20059 , \20060 , \20061 , \20062 , \20063 , \20064 , \20065 , \20066 , \20067 );
and \U$10938 ( \20069 , RIf158bb8_5469, \9462 );
and \U$10939 ( \20070 , RIf157808_5455, \9464 );
and \U$10940 ( \20071 , RIfc5d0f8_6081, \9466 );
and \U$10941 ( \20072 , RIfebef98_8293, \9468 );
and \U$10942 ( \20073 , RIfcc8a38_7305, \9470 );
and \U$10943 ( \20074 , RIfcd7ab0_7476, \9472 );
and \U$10944 ( \20075 , RIfcb1428_7039, \9474 );
and \U$10945 ( \20076 , RIfeaa0e8_8251, \9476 );
and \U$10946 ( \20077 , RIfccc548_7347, \9478 );
and \U$10947 ( \20078 , RIfce3450_7608, \9480 );
and \U$10948 ( \20079 , RIf1504b8_5373, \9482 );
and \U$10949 ( \20080 , RIe1f2be8_4139, \9484 );
and \U$10950 ( \20081 , RIf14f540_5362, \9486 );
and \U$10951 ( \20082 , RIfc772a0_6378, \9488 );
and \U$10952 ( \20083 , RIfcec258_7709, \9490 );
and \U$10953 ( \20084 , RIe1ed8f0_4080, \9492 );
and \U$10954 ( \20085 , RIe1eaec0_4050, \9494 );
and \U$10955 ( \20086 , RIe1e81c0_4018, \9496 );
and \U$10956 ( \20087 , RIe1e54c0_3986, \9498 );
and \U$10957 ( \20088 , RIe1e27c0_3954, \9500 );
and \U$10958 ( \20089 , RIe1dfac0_3922, \9502 );
and \U$10959 ( \20090 , RIe1dcdc0_3890, \9504 );
and \U$10960 ( \20091 , RIe1da0c0_3858, \9506 );
and \U$10961 ( \20092 , RIe1d73c0_3826, \9508 );
and \U$10962 ( \20093 , RIe1d19c0_3762, \9510 );
and \U$10963 ( \20094 , RIe1cecc0_3730, \9512 );
and \U$10964 ( \20095 , RIe1cbfc0_3698, \9514 );
and \U$10965 ( \20096 , RIe1c92c0_3666, \9516 );
and \U$10966 ( \20097 , RIe1c65c0_3634, \9518 );
and \U$10967 ( \20098 , RIe1c38c0_3602, \9520 );
and \U$10968 ( \20099 , RIe1c0bc0_3570, \9522 );
and \U$10969 ( \20100 , RIe1bdec0_3538, \9524 );
and \U$10970 ( \20101 , RIf14c570_5328, \9526 );
and \U$10971 ( \20102 , RIf14b328_5315, \9528 );
and \U$10972 ( \20103 , RIe1b8e98_3481, \9530 );
and \U$10973 ( \20104 , RIe1b6e40_3458, \9532 );
and \U$10974 ( \20105 , RIfc76760_6370, \9534 );
and \U$10975 ( \20106 , RIfc94b20_6714, \9536 );
and \U$10976 ( \20107 , RIe1b4f50_3436, \9538 );
and \U$10977 ( \20108 , RIe1b3ba0_3422, \9540 );
and \U$10978 ( \20109 , RIfcec3c0_7710, \9542 );
and \U$10979 ( \20110 , RIfceb010_7696, \9544 );
and \U$10980 ( \20111 , RIfe823e0_7826, \9546 );
and \U$10981 ( \20112 , RIfe82110_7824, \9548 );
and \U$10982 ( \20113 , RIfcdd8e8_7543, \9550 );
and \U$10983 ( \20114 , RIfcc0ba8_7215, \9552 );
and \U$10984 ( \20115 , RIfe82278_7825, \9554 );
and \U$10985 ( \20116 , RIe1aa7f8_3317, \9556 );
and \U$10986 ( \20117 , RIe1a8200_3290, \9558 );
and \U$10987 ( \20118 , RIe1a5500_3258, \9560 );
and \U$10988 ( \20119 , RIe1a2800_3226, \9562 );
and \U$10989 ( \20120 , RIe19fb00_3194, \9564 );
and \U$10990 ( \20121 , RIe18c000_2970, \9566 );
and \U$10991 ( \20122 , RIe178500_2746, \9568 );
and \U$10992 ( \20123 , RIe225e58_4721, \9570 );
and \U$10993 ( \20124 , RIe21aa58_4593, \9572 );
and \U$10994 ( \20125 , RIe204258_4337, \9574 );
and \U$10995 ( \20126 , RIe1fe2b8_4269, \9576 );
and \U$10996 ( \20127 , RIe1f7670_4192, \9578 );
and \U$10997 ( \20128 , RIe1f01b8_4109, \9580 );
and \U$10998 ( \20129 , RIe1d46c0_3794, \9582 );
and \U$10999 ( \20130 , RIe1bb1c0_3506, \9584 );
and \U$11000 ( \20131 , RIe1ae038_3357, \9586 );
and \U$11001 ( \20132 , RIe170670_2656, \9588 );
or \U$11002 ( \20133 , \20069 , \20070 , \20071 , \20072 , \20073 , \20074 , \20075 , \20076 , \20077 , \20078 , \20079 , \20080 , \20081 , \20082 , \20083 , \20084 , \20085 , \20086 , \20087 , \20088 , \20089 , \20090 , \20091 , \20092 , \20093 , \20094 , \20095 , \20096 , \20097 , \20098 , \20099 , \20100 , \20101 , \20102 , \20103 , \20104 , \20105 , \20106 , \20107 , \20108 , \20109 , \20110 , \20111 , \20112 , \20113 , \20114 , \20115 , \20116 , \20117 , \20118 , \20119 , \20120 , \20121 , \20122 , \20123 , \20124 , \20125 , \20126 , \20127 , \20128 , \20129 , \20130 , \20131 , \20132 );
or \U$11003 ( \20134 , \20068 , \20133 );
_DC g3b2d ( \20135_nG3b2d , \20134 , \9597 );
buf \U$11004 ( \20136 , \20135_nG3b2d );
and \U$11005 ( \20137 , \20003 , \20136 );
and \U$11006 ( \20138 , \18283 , \18416 );
and \U$11007 ( \20139 , \18416 , \18691 );
and \U$11008 ( \20140 , \18283 , \18691 );
or \U$11009 ( \20141 , \20138 , \20139 , \20140 );
and \U$11010 ( \20142 , \20136 , \20141 );
and \U$11011 ( \20143 , \20003 , \20141 );
or \U$11012 ( \20144 , \20137 , \20142 , \20143 );
xor \U$11013 ( \20145 , \19870 , \20144 );
buf g4424 ( \20146_nG4424 , \20145 );
xor \U$11014 ( \20147 , \20003 , \20136 );
xor \U$11015 ( \20148 , \20147 , \20141 );
buf g4427 ( \20149_nG4427 , \20148 );
nand \U$11016 ( \20150 , \20149_nG4427 , \18693_nG442a );
and \U$11017 ( \20151 , \20146_nG4424 , \20150 );
xor \U$11018 ( \20152 , \20149_nG4427 , \18693_nG442a );
not \U$11019 ( \20153 , \20152 );
xor \U$11020 ( \20154 , \20146_nG4424 , \20149_nG4427 );
and \U$11021 ( \20155 , \20153 , \20154 );
and \U$11023 ( \20156 , \20152 , \10694_nG9c0e );
or \U$11024 ( \20157 , 1'b0 , \20156 );
xor \U$11025 ( \20158 , \20151 , \20157 );
xor \U$11026 ( \20159 , \20151 , \20158 );
buf \U$11027 ( \20160 , \20159 );
buf \U$11028 ( \20161 , \20160 );
and \U$11029 ( \20162 , \19603 , \20161 );
and \U$11030 ( \20163 , \19149 , \19595 );
and \U$11031 ( \20164 , \19149 , \19601 );
and \U$11032 ( \20165 , \19595 , \19601 );
or \U$11033 ( \20166 , \20163 , \20164 , \20165 );
buf \U$11034 ( \20167 , \20166 );
and \U$11035 ( \20168 , \19154 , \19185 );
and \U$11036 ( \20169 , \19154 , \19593 );
and \U$11037 ( \20170 , \19185 , \19593 );
or \U$11038 ( \20171 , \20168 , \20169 , \20170 );
buf \U$11039 ( \20172 , \20171 );
xor \U$11040 ( \20173 , \20167 , \20172 );
and \U$11041 ( \20174 , \19191 , \19231 );
and \U$11042 ( \20175 , \19191 , \19591 );
and \U$11043 ( \20176 , \19231 , \19591 );
or \U$11044 ( \20177 , \20174 , \20175 , \20176 );
buf \U$11045 ( \20178 , \20177 );
and \U$11046 ( \20179 , \19159 , \19176 );
and \U$11047 ( \20180 , \19159 , \19183 );
and \U$11048 ( \20181 , \19176 , \19183 );
or \U$11049 ( \20182 , \20179 , \20180 , \20181 );
buf \U$11050 ( \20183 , \20182 );
and \U$11051 ( \20184 , \19161 , \19167 );
and \U$11052 ( \20185 , \19161 , \19174 );
and \U$11053 ( \20186 , \19167 , \19174 );
or \U$11054 ( \20187 , \20184 , \20185 , \20186 );
buf \U$11055 ( \20188 , \20187 );
and \U$11056 ( \20189 , \19199 , \19205 );
buf \U$11057 ( \20190 , \20189 );
and \U$11058 ( \20191 , \18702 , \10995_nG9c0b );
and \U$11059 ( \20192 , \18699 , \11283_nG9c08 );
or \U$11060 ( \20193 , \20191 , \20192 );
xor \U$11061 ( \20194 , \18698 , \20193 );
buf \U$11062 ( \20195 , \20194 );
buf \U$11064 ( \20196 , \20195 );
and \U$11065 ( \20197 , \17297 , \11598_nG9c05 );
and \U$11066 ( \20198 , \17294 , \12470_nG9c02 );
or \U$11067 ( \20199 , \20197 , \20198 );
xor \U$11068 ( \20200 , \17293 , \20199 );
buf \U$11069 ( \20201 , \20200 );
buf \U$11071 ( \20202 , \20201 );
xor \U$11072 ( \20203 , \20196 , \20202 );
buf \U$11073 ( \20204 , \20203 );
xor \U$11074 ( \20205 , \20190 , \20204 );
and \U$11075 ( \20206 , \15940 , \12801_nG9bff );
and \U$11076 ( \20207 , \15937 , \13705_nG9bfc );
or \U$11077 ( \20208 , \20206 , \20207 );
xor \U$11078 ( \20209 , \15936 , \20208 );
buf \U$11079 ( \20210 , \20209 );
buf \U$11081 ( \20211 , \20210 );
xor \U$11082 ( \20212 , \20205 , \20211 );
buf \U$11083 ( \20213 , \20212 );
xor \U$11084 ( \20214 , \20188 , \20213 );
and \U$11085 ( \20215 , \12157 , \16680_nG9bed );
and \U$11086 ( \20216 , \12154 , \17665_nG9bea );
or \U$11087 ( \20217 , \20215 , \20216 );
xor \U$11088 ( \20218 , \12153 , \20217 );
buf \U$11089 ( \20219 , \20218 );
buf \U$11091 ( \20220 , \20219 );
xor \U$11092 ( \20221 , \20214 , \20220 );
buf \U$11093 ( \20222 , \20221 );
xor \U$11094 ( \20223 , \20183 , \20222 );
and \U$11095 ( \20224 , \19196 , \19222 );
and \U$11096 ( \20225 , \19196 , \19229 );
and \U$11097 ( \20226 , \19222 , \19229 );
or \U$11098 ( \20227 , \20224 , \20225 , \20226 );
buf \U$11099 ( \20228 , \20227 );
xor \U$11100 ( \20229 , \20223 , \20228 );
buf \U$11101 ( \20230 , \20229 );
xor \U$11102 ( \20231 , \20178 , \20230 );
and \U$11103 ( \20232 , \19207 , \19213 );
and \U$11104 ( \20233 , \19207 , \19220 );
and \U$11105 ( \20234 , \19213 , \19220 );
or \U$11106 ( \20235 , \20232 , \20233 , \20234 );
buf \U$11107 ( \20236 , \20235 );
and \U$11108 ( \20237 , \14631 , \14070_nG9bf9 );
and \U$11109 ( \20238 , \14628 , \14984_nG9bf6 );
or \U$11110 ( \20239 , \20237 , \20238 );
xor \U$11111 ( \20240 , \14627 , \20239 );
buf \U$11112 ( \20241 , \20240 );
buf \U$11114 ( \20242 , \20241 );
xor \U$11115 ( \20243 , \20236 , \20242 );
and \U$11116 ( \20244 , \13370 , \15373_nG9bf3 );
and \U$11117 ( \20245 , \13367 , \16315_nG9bf0 );
or \U$11118 ( \20246 , \20244 , \20245 );
xor \U$11119 ( \20247 , \13366 , \20246 );
buf \U$11120 ( \20248 , \20247 );
buf \U$11122 ( \20249 , \20248 );
xor \U$11123 ( \20250 , \20243 , \20249 );
buf \U$11124 ( \20251 , \20250 );
and \U$11125 ( \20252 , \10421 , \18107_nG9be7 );
and \U$11126 ( \20253 , \10418 , \19091_nG9be4 );
or \U$11127 ( \20254 , \20252 , \20253 );
xor \U$11128 ( \20255 , \10417 , \20254 );
buf \U$11129 ( \20256 , \20255 );
buf \U$11131 ( \20257 , \20256 );
xor \U$11132 ( \20258 , \20251 , \20257 );
and \U$11133 ( \20259 , \10707 , \19586_nG9be1 );
and \U$11134 ( \20260 , \19548 , \19552 );
and \U$11135 ( \20261 , \19552 , \19574 );
and \U$11136 ( \20262 , \19548 , \19574 );
or \U$11137 ( \20263 , \20260 , \20261 , \20262 );
and \U$11138 ( \20264 , \15321 , \14054 );
and \U$11139 ( \20265 , \16267 , \13692 );
nor \U$11140 ( \20266 , \20264 , \20265 );
xnor \U$11141 ( \20267 , \20266 , \14035 );
and \U$11142 ( \20268 , \14024 , \15336 );
and \U$11143 ( \20269 , \14950 , \14963 );
nor \U$11144 ( \20270 , \20268 , \20269 );
xnor \U$11145 ( \20271 , \20270 , \15342 );
xor \U$11146 ( \20272 , \20267 , \20271 );
and \U$11147 ( \20273 , \10988 , \19534 );
and \U$11148 ( \20274 , \11270 , \19045 );
nor \U$11149 ( \20275 , \20273 , \20274 );
xnor \U$11150 ( \20276 , \20275 , \19540 );
xor \U$11151 ( \20277 , \20272 , \20276 );
and \U$11152 ( \20278 , \19558 , \10983 );
and \U$11153 ( \20279 , RIdec4b68_702, \9333 );
and \U$11154 ( \20280 , RIdec1e68_670, \9335 );
and \U$11155 ( \20281 , RIfc5df08_6091, \9337 );
and \U$11156 ( \20282 , RIdebf168_638, \9339 );
and \U$11157 ( \20283 , RIfce6df8_7649, \9341 );
and \U$11158 ( \20284 , RIdebc468_606, \9343 );
and \U$11159 ( \20285 , RIdeb9768_574, \9345 );
and \U$11160 ( \20286 , RIdeb6a68_542, \9347 );
and \U$11161 ( \20287 , RIfc75ef0_6364, \9349 );
and \U$11162 ( \20288 , RIdeb1068_478, \9351 );
and \U$11163 ( \20289 , RIfcc12b0_7220, \9353 );
and \U$11164 ( \20290 , RIdeae368_446, \9355 );
and \U$11165 ( \20291 , RIfc5e340_6094, \9357 );
and \U$11166 ( \20292 , RIdea9070_414, \9359 );
and \U$11167 ( \20293 , RIdea2770_382, \9361 );
and \U$11168 ( \20294 , RIde9be70_350, \9363 );
and \U$11169 ( \20295 , RIfced4a0_7722, \9365 );
and \U$11170 ( \20296 , RIfcc1418_7221, \9367 );
and \U$11171 ( \20297 , RIfc95930_6724, \9369 );
and \U$11172 ( \20298 , RIfcec0f0_7708, \9371 );
and \U$11173 ( \20299 , RIde90368_293, \9373 );
and \U$11174 ( \20300 , RIde8c858_275, \9375 );
and \U$11175 ( \20301 , RIde893d8_259, \9377 );
and \U$11176 ( \20302 , RIde84ef0_238, \9379 );
and \U$11177 ( \20303 , RIde80d50_218, \9381 );
and \U$11178 ( \20304 , RIfc95a98_6725, \9383 );
and \U$11179 ( \20305 , RIfced068_7719, \9385 );
and \U$11180 ( \20306 , RIfced1d0_7720, \9387 );
and \U$11181 ( \20307 , RIfcedfe0_7730, \9389 );
and \U$11182 ( \20308 , RIe16b0a8_2595, \9391 );
and \U$11183 ( \20309 , RIe169758_2577, \9393 );
and \U$11184 ( \20310 , RIe167700_2554, \9395 );
and \U$11185 ( \20311 , RIe164b68_2523, \9397 );
and \U$11186 ( \20312 , RIe161e68_2491, \9399 );
and \U$11187 ( \20313 , RIee36e20_5083, \9401 );
and \U$11188 ( \20314 , RIe15f168_2459, \9403 );
and \U$11189 ( \20315 , RIfc426e0_5778, \9405 );
and \U$11190 ( \20316 , RIe15c468_2427, \9407 );
and \U$11191 ( \20317 , RIe156a68_2363, \9409 );
and \U$11192 ( \20318 , RIe153d68_2331, \9411 );
and \U$11193 ( \20319 , RIfe82818_7829, \9413 );
and \U$11194 ( \20320 , RIe151068_2299, \9415 );
and \U$11195 ( \20321 , RIee34c60_5059, \9417 );
and \U$11196 ( \20322 , RIe14e368_2267, \9419 );
and \U$11197 ( \20323 , RIfc5f9c0_6110, \9421 );
and \U$11198 ( \20324 , RIe14b668_2235, \9423 );
and \U$11199 ( \20325 , RIe148968_2203, \9425 );
and \U$11200 ( \20326 , RIe145c68_2171, \9427 );
and \U$11201 ( \20327 , RIfccfef0_7388, \9429 );
and \U$11202 ( \20328 , RIfca57b8_6905, \9431 );
and \U$11203 ( \20329 , RIfc600c8_6115, \9433 );
and \U$11204 ( \20330 , RIfcafda8_7023, \9435 );
and \U$11205 ( \20331 , RIe140970_2112, \9437 );
and \U$11206 ( \20332 , RIdf3e710_2087, \9439 );
and \U$11207 ( \20333 , RIdf3c6b8_2064, \9441 );
and \U$11208 ( \20334 , RIdf3a228_2038, \9443 );
and \U$11209 ( \20335 , RIfc5fc90_6112, \9445 );
and \U$11210 ( \20336 , RIee2f3c8_4996, \9447 );
and \U$11211 ( \20337 , RIfc742d0_6344, \9449 );
and \U$11212 ( \20338 , RIee2d208_4972, \9451 );
and \U$11213 ( \20339 , RIdf34f30_1979, \9453 );
and \U$11214 ( \20340 , RIfebf100_8294, \9455 );
and \U$11215 ( \20341 , RIdf30a48_1930, \9457 );
and \U$11216 ( \20342 , RIdf2ecc0_1909, \9459 );
or \U$11217 ( \20343 , \20279 , \20280 , \20281 , \20282 , \20283 , \20284 , \20285 , \20286 , \20287 , \20288 , \20289 , \20290 , \20291 , \20292 , \20293 , \20294 , \20295 , \20296 , \20297 , \20298 , \20299 , \20300 , \20301 , \20302 , \20303 , \20304 , \20305 , \20306 , \20307 , \20308 , \20309 , \20310 , \20311 , \20312 , \20313 , \20314 , \20315 , \20316 , \20317 , \20318 , \20319 , \20320 , \20321 , \20322 , \20323 , \20324 , \20325 , \20326 , \20327 , \20328 , \20329 , \20330 , \20331 , \20332 , \20333 , \20334 , \20335 , \20336 , \20337 , \20338 , \20339 , \20340 , \20341 , \20342 );
and \U$11218 ( \20344 , RIfcb08e8_7031, \9462 );
and \U$11219 ( \20345 , RIfcee418_7733, \9464 );
and \U$11220 ( \20346 , RIfc95ed0_6728, \9466 );
and \U$11221 ( \20347 , RIfcdef68_7559, \9468 );
and \U$11222 ( \20348 , RIdf29e00_1853, \9470 );
and \U$11223 ( \20349 , RIdf27c40_1829, \9472 );
and \U$11224 ( \20350 , RIdf25eb8_1808, \9474 );
and \U$11225 ( \20351 , RIdf24298_1788, \9476 );
and \U$11226 ( \20352 , RIfc5ed18_6101, \9478 );
and \U$11227 ( \20353 , RIfcee850_7736, \9480 );
and \U$11228 ( \20354 , RIdf227e0_1769, \9482 );
and \U$11229 ( \20355 , RIfc5efe8_6103, \9484 );
and \U$11230 ( \20356 , RIdf212c8_1754, \9486 );
and \U$11231 ( \20357 , RIfeaa520_8254, \9488 );
and \U$11232 ( \20358 , RIdf1ad88_1682, \9490 );
and \U$11233 ( \20359 , RIdf18e98_1660, \9492 );
and \U$11234 ( \20360 , RIdf16738_1632, \9494 );
and \U$11235 ( \20361 , RIdf13a38_1600, \9496 );
and \U$11236 ( \20362 , RIdf10d38_1568, \9498 );
and \U$11237 ( \20363 , RIdf0e038_1536, \9500 );
and \U$11238 ( \20364 , RIdf0b338_1504, \9502 );
and \U$11239 ( \20365 , RIdf08638_1472, \9504 );
and \U$11240 ( \20366 , RIdf05938_1440, \9506 );
and \U$11241 ( \20367 , RIdf02c38_1408, \9508 );
and \U$11242 ( \20368 , RIdefd238_1344, \9510 );
and \U$11243 ( \20369 , RIdefa538_1312, \9512 );
and \U$11244 ( \20370 , RIdef7838_1280, \9514 );
and \U$11245 ( \20371 , RIdef4b38_1248, \9516 );
and \U$11246 ( \20372 , RIdef1e38_1216, \9518 );
and \U$11247 ( \20373 , RIdeef138_1184, \9520 );
and \U$11248 ( \20374 , RIdeec438_1152, \9522 );
and \U$11249 ( \20375 , RIdee9738_1120, \9524 );
and \U$11250 ( \20376 , RIfcc96e0_7314, \9526 );
and \U$11251 ( \20377 , RIfccfd88_7387, \9528 );
and \U$11252 ( \20378 , RIfc60aa0_6122, \9530 );
and \U$11253 ( \20379 , RIfca5ec0_6910, \9532 );
and \U$11254 ( \20380 , RIdee45a8_1062, \9534 );
and \U$11255 ( \20381 , RIdee2550_1039, \9536 );
and \U$11256 ( \20382 , RIdee0660_1017, \9538 );
and \U$11257 ( \20383 , RIfe826b0_7828, \9540 );
and \U$11258 ( \20384 , RIfcdeb30_7556, \9542 );
and \U$11259 ( \20385 , RIfc73bc8_6339, \9544 );
and \U$11260 ( \20386 , RIfca5bf0_6908, \9546 );
and \U$11261 ( \20387 , RIfc73a60_6338, \9548 );
and \U$11262 ( \20388 , RIfe82980_7830, \9550 );
and \U$11263 ( \20389 , RIded6bb0_907, \9552 );
and \U$11264 ( \20390 , RIded4cc0_885, \9554 );
and \U$11265 ( \20391 , RIded2830_859, \9556 );
and \U$11266 ( \20392 , RIdecff68_830, \9558 );
and \U$11267 ( \20393 , RIdecd268_798, \9560 );
and \U$11268 ( \20394 , RIdeca568_766, \9562 );
and \U$11269 ( \20395 , RIdec7868_734, \9564 );
and \U$11270 ( \20396 , RIdeb3d68_510, \9566 );
and \U$11271 ( \20397 , RIde95570_318, \9568 );
and \U$11272 ( \20398 , RIe16d970_2624, \9570 );
and \U$11273 ( \20399 , RIe159768_2395, \9572 );
and \U$11274 ( \20400 , RIe142f68_2139, \9574 );
and \U$11275 ( \20401 , RIdf37960_2009, \9576 );
and \U$11276 ( \20402 , RIdf2bfc0_1877, \9578 );
and \U$11277 ( \20403 , RIdf1c840_1701, \9580 );
and \U$11278 ( \20404 , RIdefff38_1376, \9582 );
and \U$11279 ( \20405 , RIdee6a38_1088, \9584 );
and \U$11280 ( \20406 , RIdedb7a0_961, \9586 );
and \U$11281 ( \20407 , RIde7b4b8_191, \9588 );
or \U$11282 ( \20408 , \20344 , \20345 , \20346 , \20347 , \20348 , \20349 , \20350 , \20351 , \20352 , \20353 , \20354 , \20355 , \20356 , \20357 , \20358 , \20359 , \20360 , \20361 , \20362 , \20363 , \20364 , \20365 , \20366 , \20367 , \20368 , \20369 , \20370 , \20371 , \20372 , \20373 , \20374 , \20375 , \20376 , \20377 , \20378 , \20379 , \20380 , \20381 , \20382 , \20383 , \20384 , \20385 , \20386 , \20387 , \20388 , \20389 , \20390 , \20391 , \20392 , \20393 , \20394 , \20395 , \20396 , \20397 , \20398 , \20399 , \20400 , \20401 , \20402 , \20403 , \20404 , \20405 , \20406 , \20407 );
or \U$11283 ( \20409 , \20343 , \20408 );
_DC g65a7 ( \20410_nG65a7 , \20409 , \9597 );
and \U$11284 ( \20411 , RIe19ce00_3162, \9059 );
and \U$11285 ( \20412 , RIe19a100_3130, \9061 );
and \U$11286 ( \20413 , RIfce96c0_7678, \9063 );
and \U$11287 ( \20414 , RIe197400_3098, \9065 );
and \U$11288 ( \20415 , RIf144410_5236, \9067 );
and \U$11289 ( \20416 , RIe194700_3066, \9069 );
and \U$11290 ( \20417 , RIe191a00_3034, \9071 );
and \U$11291 ( \20418 , RIe18ed00_3002, \9073 );
and \U$11292 ( \20419 , RIe189300_2938, \9075 );
and \U$11293 ( \20420 , RIe186600_2906, \9077 );
and \U$11294 ( \20421 , RIfebee30_8292, \9079 );
and \U$11295 ( \20422 , RIe183900_2874, \9081 );
and \U$11296 ( \20423 , RIfcdbcc8_7523, \9083 );
and \U$11297 ( \20424 , RIe180c00_2842, \9085 );
and \U$11298 ( \20425 , RIe17df00_2810, \9087 );
and \U$11299 ( \20426 , RIe17b200_2778, \9089 );
and \U$11300 ( \20427 , RIf141f80_5210, \9091 );
and \U$11301 ( \20428 , RIfce7398_7653, \9093 );
and \U$11302 ( \20429 , RIfcb1e00_7046, \9095 );
and \U$11303 ( \20430 , RIfe82548_7827, \9097 );
and \U$11304 ( \20431 , RIfca42a0_6890, \9099 );
and \U$11305 ( \20432 , RIfcbff00_7206, \9101 );
and \U$11306 ( \20433 , RIfcaaee8_6967, \9103 );
and \U$11307 ( \20434 , RIee3d090_5153, \9105 );
and \U$11308 ( \20435 , RIfc5c180_6070, \9107 );
and \U$11309 ( \20436 , RIfce35b8_7609, \9109 );
and \U$11310 ( \20437 , RIee399b8_5114, \9111 );
and \U$11311 ( \20438 , RIfea8a68_8235, \9113 );
and \U$11312 ( \20439 , RIf16fef8_5733, \9115 );
and \U$11313 ( \20440 , RIfebecc8_8291, \9117 );
and \U$11314 ( \20441 , RIfc5c450_6072, \9119 );
and \U$11315 ( \20442 , RIfce9288_7675, \9121 );
and \U$11316 ( \20443 , RIfc40778_5759, \9123 );
and \U$11317 ( \20444 , RIe223158_4689, \9125 );
and \U$11318 ( \20445 , RIfce77d0_7656, \9127 );
and \U$11319 ( \20446 , RIe220458_4657, \9129 );
and \U$11320 ( \20447 , RIfce24d8_7597, \9131 );
and \U$11321 ( \20448 , RIe21d758_4625, \9133 );
and \U$11322 ( \20449 , RIe217d58_4561, \9135 );
and \U$11323 ( \20450 , RIe215058_4529, \9137 );
and \U$11324 ( \20451 , RIfce8a18_7669, \9139 );
and \U$11325 ( \20452 , RIe212358_4497, \9141 );
and \U$11326 ( \20453 , RIfce1998_7589, \9143 );
and \U$11327 ( \20454 , RIe20f658_4465, \9145 );
and \U$11328 ( \20455 , RIfc77840_6382, \9147 );
and \U$11329 ( \20456 , RIe20c958_4433, \9149 );
and \U$11330 ( \20457 , RIe209c58_4401, \9151 );
and \U$11331 ( \20458 , RIe206f58_4369, \9153 );
and \U$11332 ( \20459 , RIf166cb8_5629, \9155 );
and \U$11333 ( \20460 , RIf165bd8_5617, \9157 );
and \U$11334 ( \20461 , RIfe81fa8_7823, \9159 );
and \U$11335 ( \20462 , RIfe81e40_7822, \9161 );
and \U$11336 ( \20463 , RIfc5c888_6075, \9163 );
and \U$11337 ( \20464 , RIfceb178_7697, \9165 );
and \U$11338 ( \20465 , RIf1631a8_5587, \9167 );
and \U$11339 ( \20466 , RIf1619c0_5570, \9169 );
and \U$11340 ( \20467 , RIfccf248_7379, \9171 );
and \U$11341 ( \20468 , RIfc77570_6380, \9173 );
and \U$11342 ( \20469 , RIe1fc800_4250, \9175 );
and \U$11343 ( \20470 , RIe1fb720_4238, \9177 );
and \U$11344 ( \20471 , RIf15c830_5512, \9179 );
and \U$11345 ( \20472 , RIf15b1b0_5496, \9181 );
and \U$11346 ( \20473 , RIfcd0fd0_7400, \9183 );
and \U$11347 ( \20474 , RIfccc6b0_7348, \9185 );
or \U$11348 ( \20475 , \20411 , \20412 , \20413 , \20414 , \20415 , \20416 , \20417 , \20418 , \20419 , \20420 , \20421 , \20422 , \20423 , \20424 , \20425 , \20426 , \20427 , \20428 , \20429 , \20430 , \20431 , \20432 , \20433 , \20434 , \20435 , \20436 , \20437 , \20438 , \20439 , \20440 , \20441 , \20442 , \20443 , \20444 , \20445 , \20446 , \20447 , \20448 , \20449 , \20450 , \20451 , \20452 , \20453 , \20454 , \20455 , \20456 , \20457 , \20458 , \20459 , \20460 , \20461 , \20462 , \20463 , \20464 , \20465 , \20466 , \20467 , \20468 , \20469 , \20470 , \20471 , \20472 , \20473 , \20474 );
and \U$11349 ( \20476 , RIf158bb8_5469, \9188 );
and \U$11350 ( \20477 , RIf157808_5455, \9190 );
and \U$11351 ( \20478 , RIfc5d0f8_6081, \9192 );
and \U$11352 ( \20479 , RIfebef98_8293, \9194 );
and \U$11353 ( \20480 , RIfcc8a38_7305, \9196 );
and \U$11354 ( \20481 , RIfcd7ab0_7476, \9198 );
and \U$11355 ( \20482 , RIfcb1428_7039, \9200 );
and \U$11356 ( \20483 , RIfeaa0e8_8251, \9202 );
and \U$11357 ( \20484 , RIfccc548_7347, \9204 );
and \U$11358 ( \20485 , RIfce3450_7608, \9206 );
and \U$11359 ( \20486 , RIf1504b8_5373, \9208 );
and \U$11360 ( \20487 , RIe1f2be8_4139, \9210 );
and \U$11361 ( \20488 , RIf14f540_5362, \9212 );
and \U$11362 ( \20489 , RIfc772a0_6378, \9214 );
and \U$11363 ( \20490 , RIfcec258_7709, \9216 );
and \U$11364 ( \20491 , RIe1ed8f0_4080, \9218 );
and \U$11365 ( \20492 , RIe1eaec0_4050, \9220 );
and \U$11366 ( \20493 , RIe1e81c0_4018, \9222 );
and \U$11367 ( \20494 , RIe1e54c0_3986, \9224 );
and \U$11368 ( \20495 , RIe1e27c0_3954, \9226 );
and \U$11369 ( \20496 , RIe1dfac0_3922, \9228 );
and \U$11370 ( \20497 , RIe1dcdc0_3890, \9230 );
and \U$11371 ( \20498 , RIe1da0c0_3858, \9232 );
and \U$11372 ( \20499 , RIe1d73c0_3826, \9234 );
and \U$11373 ( \20500 , RIe1d19c0_3762, \9236 );
and \U$11374 ( \20501 , RIe1cecc0_3730, \9238 );
and \U$11375 ( \20502 , RIe1cbfc0_3698, \9240 );
and \U$11376 ( \20503 , RIe1c92c0_3666, \9242 );
and \U$11377 ( \20504 , RIe1c65c0_3634, \9244 );
and \U$11378 ( \20505 , RIe1c38c0_3602, \9246 );
and \U$11379 ( \20506 , RIe1c0bc0_3570, \9248 );
and \U$11380 ( \20507 , RIe1bdec0_3538, \9250 );
and \U$11381 ( \20508 , RIf14c570_5328, \9252 );
and \U$11382 ( \20509 , RIf14b328_5315, \9254 );
and \U$11383 ( \20510 , RIe1b8e98_3481, \9256 );
and \U$11384 ( \20511 , RIe1b6e40_3458, \9258 );
and \U$11385 ( \20512 , RIfc76760_6370, \9260 );
and \U$11386 ( \20513 , RIfc94b20_6714, \9262 );
and \U$11387 ( \20514 , RIe1b4f50_3436, \9264 );
and \U$11388 ( \20515 , RIe1b3ba0_3422, \9266 );
and \U$11389 ( \20516 , RIfcec3c0_7710, \9268 );
and \U$11390 ( \20517 , RIfceb010_7696, \9270 );
and \U$11391 ( \20518 , RIfe823e0_7826, \9272 );
and \U$11392 ( \20519 , RIfe82110_7824, \9274 );
and \U$11393 ( \20520 , RIfcdd8e8_7543, \9276 );
and \U$11394 ( \20521 , RIfcc0ba8_7215, \9278 );
and \U$11395 ( \20522 , RIfe82278_7825, \9280 );
and \U$11396 ( \20523 , RIe1aa7f8_3317, \9282 );
and \U$11397 ( \20524 , RIe1a8200_3290, \9284 );
and \U$11398 ( \20525 , RIe1a5500_3258, \9286 );
and \U$11399 ( \20526 , RIe1a2800_3226, \9288 );
and \U$11400 ( \20527 , RIe19fb00_3194, \9290 );
and \U$11401 ( \20528 , RIe18c000_2970, \9292 );
and \U$11402 ( \20529 , RIe178500_2746, \9294 );
and \U$11403 ( \20530 , RIe225e58_4721, \9296 );
and \U$11404 ( \20531 , RIe21aa58_4593, \9298 );
and \U$11405 ( \20532 , RIe204258_4337, \9300 );
and \U$11406 ( \20533 , RIe1fe2b8_4269, \9302 );
and \U$11407 ( \20534 , RIe1f7670_4192, \9304 );
and \U$11408 ( \20535 , RIe1f01b8_4109, \9306 );
and \U$11409 ( \20536 , RIe1d46c0_3794, \9308 );
and \U$11410 ( \20537 , RIe1bb1c0_3506, \9310 );
and \U$11411 ( \20538 , RIe1ae038_3357, \9312 );
and \U$11412 ( \20539 , RIe170670_2656, \9314 );
or \U$11413 ( \20540 , \20476 , \20477 , \20478 , \20479 , \20480 , \20481 , \20482 , \20483 , \20484 , \20485 , \20486 , \20487 , \20488 , \20489 , \20490 , \20491 , \20492 , \20493 , \20494 , \20495 , \20496 , \20497 , \20498 , \20499 , \20500 , \20501 , \20502 , \20503 , \20504 , \20505 , \20506 , \20507 , \20508 , \20509 , \20510 , \20511 , \20512 , \20513 , \20514 , \20515 , \20516 , \20517 , \20518 , \20519 , \20520 , \20521 , \20522 , \20523 , \20524 , \20525 , \20526 , \20527 , \20528 , \20529 , \20530 , \20531 , \20532 , \20533 , \20534 , \20535 , \20536 , \20537 , \20538 , \20539 );
or \U$11414 ( \20541 , \20475 , \20540 );
_DC g65a8 ( \20542_nG65a8 , \20541 , \9323 );
and g65a9 ( \20543_nG65a9 , \20410_nG65a7 , \20542_nG65a8 );
buf \U$11415 ( \20544 , \20543_nG65a9 );
and \U$11416 ( \20545 , \20544 , \10691 );
nor \U$11417 ( \20546 , \20278 , \20545 );
xnor \U$11418 ( \20547 , \20546 , \10980 );
and \U$11419 ( \20548 , \18035 , \11574 );
and \U$11420 ( \20549 , \19032 , \11278 );
nor \U$11421 ( \20550 , \20548 , \20549 );
xnor \U$11422 ( \20551 , \20550 , \11580 );
xor \U$11423 ( \20552 , \20547 , \20551 );
_DC g556a ( \20553_nG556a , \20409 , \9597 );
_DC g55ee ( \20554_nG55ee , \20541 , \9323 );
xor g55ef ( \20555_nG55ef , \20553_nG556a , \20554_nG55ee );
buf \U$11424 ( \20556 , \20555_nG55ef );
xor \U$11425 ( \20557 , \20556 , \19531 );
and \U$11426 ( \20558 , \10687 , \20557 );
xor \U$11427 ( \20559 , \20552 , \20558 );
xor \U$11428 ( \20560 , \20277 , \20559 );
and \U$11429 ( \20561 , \16655 , \12790 );
and \U$11430 ( \20562 , \17627 , \12461 );
nor \U$11431 ( \20563 , \20561 , \20562 );
xnor \U$11432 ( \20564 , \20563 , \12780 );
and \U$11433 ( \20565 , \12769 , \16635 );
and \U$11434 ( \20566 , \13679 , \16301 );
nor \U$11435 ( \20567 , \20565 , \20566 );
xnor \U$11436 ( \20568 , \20567 , \16625 );
xor \U$11437 ( \20569 , \20564 , \20568 );
and \U$11438 ( \20570 , \11586 , \18090 );
and \U$11439 ( \20571 , \12448 , \17655 );
nor \U$11440 ( \20572 , \20570 , \20571 );
xnor \U$11441 ( \20573 , \20572 , \18046 );
xor \U$11442 ( \20574 , \20569 , \20573 );
xor \U$11443 ( \20575 , \20560 , \20574 );
xor \U$11444 ( \20576 , \20263 , \20575 );
and \U$11445 ( \20577 , \19564 , \19568 );
and \U$11446 ( \20578 , \19568 , \19573 );
and \U$11447 ( \20579 , \19564 , \19573 );
or \U$11448 ( \20580 , \20577 , \20578 , \20579 );
and \U$11449 ( \20581 , \19241 , \19255 );
and \U$11450 ( \20582 , \19255 , \19542 );
and \U$11451 ( \20583 , \19241 , \19542 );
or \U$11452 ( \20584 , \20581 , \20582 , \20583 );
xor \U$11453 ( \20585 , \20580 , \20584 );
and \U$11454 ( \20586 , \19245 , \19249 );
and \U$11455 ( \20587 , \19249 , \19254 );
and \U$11456 ( \20588 , \19245 , \19254 );
or \U$11457 ( \20589 , \20586 , \20587 , \20588 );
and \U$11458 ( \20590 , \19260 , \19264 );
and \U$11459 ( \20591 , \19264 , \19541 );
and \U$11460 ( \20592 , \19260 , \19541 );
or \U$11461 ( \20593 , \20590 , \20591 , \20592 );
xor \U$11462 ( \20594 , \20589 , \20593 );
and \U$11463 ( \20595 , \19561 , \19563 );
xor \U$11464 ( \20596 , \20594 , \20595 );
xor \U$11465 ( \20597 , \20585 , \20596 );
xor \U$11466 ( \20598 , \20576 , \20597 );
and \U$11467 ( \20599 , \19237 , \19543 );
and \U$11468 ( \20600 , \19543 , \19575 );
and \U$11469 ( \20601 , \19237 , \19575 );
or \U$11470 ( \20602 , \20599 , \20600 , \20601 );
xor \U$11471 ( \20603 , \20598 , \20602 );
and \U$11472 ( \20604 , \19576 , \19580 );
and \U$11473 ( \20605 , \19581 , \19584 );
or \U$11474 ( \20606 , \20604 , \20605 );
xor \U$11475 ( \20607 , \20603 , \20606 );
buf g9bde ( \20608_nG9bde , \20607 );
and \U$11476 ( \20609 , \10704 , \20608_nG9bde );
or \U$11477 ( \20610 , \20259 , \20609 );
xor \U$11478 ( \20611 , \10703 , \20610 );
buf \U$11479 ( \20612 , \20611 );
buf \U$11481 ( \20613 , \20612 );
xor \U$11482 ( \20614 , \20258 , \20613 );
buf \U$11483 ( \20615 , \20614 );
xor \U$11484 ( \20616 , \20231 , \20615 );
buf \U$11485 ( \20617 , \20616 );
xor \U$11486 ( \20618 , \20173 , \20617 );
and \U$11487 ( \20619 , \19603 , \20618 );
and \U$11488 ( \20620 , \20161 , \20618 );
or \U$11489 ( \20621 , \20162 , \20619 , \20620 );
and \U$11490 ( \20622 , \20167 , \20172 );
and \U$11491 ( \20623 , \20167 , \20617 );
and \U$11492 ( \20624 , \20172 , \20617 );
or \U$11493 ( \20625 , \20622 , \20623 , \20624 );
xor \U$11494 ( \20626 , \20621 , \20625 );
and \U$11495 ( \20627 , \20178 , \20230 );
and \U$11496 ( \20628 , \20178 , \20615 );
and \U$11497 ( \20629 , \20230 , \20615 );
or \U$11498 ( \20630 , \20627 , \20628 , \20629 );
xor \U$11499 ( \20631 , \20626 , \20630 );
and \U$11500 ( \20632 , \20251 , \20257 );
and \U$11501 ( \20633 , \20251 , \20613 );
and \U$11502 ( \20634 , \20257 , \20613 );
or \U$11503 ( \20635 , \20632 , \20633 , \20634 );
buf \U$11504 ( \20636 , \20635 );
and \U$11505 ( \20637 , \20236 , \20242 );
and \U$11506 ( \20638 , \20236 , \20249 );
and \U$11507 ( \20639 , \20242 , \20249 );
or \U$11508 ( \20640 , \20637 , \20638 , \20639 );
buf \U$11509 ( \20641 , \20640 );
and \U$11510 ( \20642 , \20151 , \20158 );
buf \U$11511 ( \20643 , \20642 );
buf \U$11513 ( \20644 , \20643 );
and \U$11514 ( \20645 , \18702 , \11283_nG9c08 );
and \U$11515 ( \20646 , \18699 , \11598_nG9c05 );
or \U$11516 ( \20647 , \20645 , \20646 );
xor \U$11517 ( \20648 , \18698 , \20647 );
buf \U$11518 ( \20649 , \20648 );
buf \U$11520 ( \20650 , \20649 );
xor \U$11521 ( \20651 , \20644 , \20650 );
buf \U$11522 ( \20652 , \20651 );
and \U$11523 ( \20653 , \20155 , \10694_nG9c0e );
and \U$11524 ( \20654 , \20152 , \10995_nG9c0b );
or \U$11525 ( \20655 , \20653 , \20654 );
xor \U$11526 ( \20656 , \20151 , \20655 );
buf \U$11527 ( \20657 , \20656 );
buf \U$11529 ( \20658 , \20657 );
xor \U$11530 ( \20659 , \20652 , \20658 );
and \U$11531 ( \20660 , \17297 , \12470_nG9c02 );
and \U$11532 ( \20661 , \17294 , \12801_nG9bff );
or \U$11533 ( \20662 , \20660 , \20661 );
xor \U$11534 ( \20663 , \17293 , \20662 );
buf \U$11535 ( \20664 , \20663 );
buf \U$11537 ( \20665 , \20664 );
xor \U$11538 ( \20666 , \20659 , \20665 );
buf \U$11539 ( \20667 , \20666 );
and \U$11540 ( \20668 , \20196 , \20202 );
buf \U$11541 ( \20669 , \20668 );
xor \U$11542 ( \20670 , \20667 , \20669 );
and \U$11543 ( \20671 , \15940 , \13705_nG9bfc );
and \U$11544 ( \20672 , \15937 , \14070_nG9bf9 );
or \U$11545 ( \20673 , \20671 , \20672 );
xor \U$11546 ( \20674 , \15936 , \20673 );
buf \U$11547 ( \20675 , \20674 );
buf \U$11549 ( \20676 , \20675 );
xor \U$11550 ( \20677 , \20670 , \20676 );
buf \U$11551 ( \20678 , \20677 );
xor \U$11552 ( \20679 , \20641 , \20678 );
and \U$11553 ( \20680 , \12157 , \17665_nG9bea );
and \U$11554 ( \20681 , \12154 , \18107_nG9be7 );
or \U$11555 ( \20682 , \20680 , \20681 );
xor \U$11556 ( \20683 , \12153 , \20682 );
buf \U$11557 ( \20684 , \20683 );
buf \U$11559 ( \20685 , \20684 );
xor \U$11560 ( \20686 , \20679 , \20685 );
buf \U$11561 ( \20687 , \20686 );
xor \U$11562 ( \20688 , \20636 , \20687 );
and \U$11563 ( \20689 , \20188 , \20213 );
and \U$11564 ( \20690 , \20188 , \20220 );
and \U$11565 ( \20691 , \20213 , \20220 );
or \U$11566 ( \20692 , \20689 , \20690 , \20691 );
buf \U$11567 ( \20693 , \20692 );
xor \U$11568 ( \20694 , \20688 , \20693 );
buf \U$11569 ( \20695 , \20694 );
and \U$11570 ( \20696 , \20190 , \20204 );
and \U$11571 ( \20697 , \20190 , \20211 );
and \U$11572 ( \20698 , \20204 , \20211 );
or \U$11573 ( \20699 , \20696 , \20697 , \20698 );
buf \U$11574 ( \20700 , \20699 );
and \U$11575 ( \20701 , \14631 , \14984_nG9bf6 );
and \U$11576 ( \20702 , \14628 , \15373_nG9bf3 );
or \U$11577 ( \20703 , \20701 , \20702 );
xor \U$11578 ( \20704 , \14627 , \20703 );
buf \U$11579 ( \20705 , \20704 );
buf \U$11581 ( \20706 , \20705 );
xor \U$11582 ( \20707 , \20700 , \20706 );
and \U$11583 ( \20708 , \13370 , \16315_nG9bf0 );
and \U$11584 ( \20709 , \13367 , \16680_nG9bed );
or \U$11585 ( \20710 , \20708 , \20709 );
xor \U$11586 ( \20711 , \13366 , \20710 );
buf \U$11587 ( \20712 , \20711 );
buf \U$11589 ( \20713 , \20712 );
xor \U$11590 ( \20714 , \20707 , \20713 );
buf \U$11591 ( \20715 , \20714 );
and \U$11592 ( \20716 , \10421 , \19091_nG9be4 );
and \U$11593 ( \20717 , \10418 , \19586_nG9be1 );
or \U$11594 ( \20718 , \20716 , \20717 );
xor \U$11595 ( \20719 , \10417 , \20718 );
buf \U$11596 ( \20720 , \20719 );
buf \U$11598 ( \20721 , \20720 );
xor \U$11599 ( \20722 , \20715 , \20721 );
and \U$11600 ( \20723 , \10707 , \20608_nG9bde );
and \U$11601 ( \20724 , \20580 , \20584 );
and \U$11602 ( \20725 , \20584 , \20596 );
and \U$11603 ( \20726 , \20580 , \20596 );
or \U$11604 ( \20727 , \20724 , \20725 , \20726 );
and \U$11605 ( \20728 , \16267 , \14054 );
and \U$11606 ( \20729 , \16655 , \13692 );
nor \U$11607 ( \20730 , \20728 , \20729 );
xnor \U$11608 ( \20731 , \20730 , \14035 );
and \U$11609 ( \20732 , \11270 , \19534 );
and \U$11610 ( \20733 , \11586 , \19045 );
nor \U$11611 ( \20734 , \20732 , \20733 );
xnor \U$11612 ( \20735 , \20734 , \19540 );
xor \U$11613 ( \20736 , \20731 , \20735 );
and \U$11614 ( \20737 , RIdec4cd0_703, \9333 );
and \U$11615 ( \20738 , RIdec1fd0_671, \9335 );
and \U$11616 ( \20739 , RIfc7b4b8_6425, \9337 );
and \U$11617 ( \20740 , RIdebf2d0_639, \9339 );
and \U$11618 ( \20741 , RIfc7b1e8_6423, \9341 );
and \U$11619 ( \20742 , RIdebc5d0_607, \9343 );
and \U$11620 ( \20743 , RIdeb98d0_575, \9345 );
and \U$11621 ( \20744 , RIdeb6bd0_543, \9347 );
and \U$11622 ( \20745 , RIfe83358_7837, \9349 );
and \U$11623 ( \20746 , RIdeb11d0_479, \9351 );
and \U$11624 ( \20747 , RIee1e5c8_4804, \9353 );
and \U$11625 ( \20748 , RIdeae4d0_447, \9355 );
and \U$11626 ( \20749 , RIfc437c0_5790, \9357 );
and \U$11627 ( \20750 , RIdea93b8_415, \9359 );
and \U$11628 ( \20751 , RIdea2ab8_383, \9361 );
and \U$11629 ( \20752 , RIde9c1b8_351, \9363 );
and \U$11630 ( \20753 , RIfc90ea8_6671, \9365 );
and \U$11631 ( \20754 , RIfc7af18_6421, \9367 );
and \U$11632 ( \20755 , RIfe83088_7835, \9369 );
and \U$11633 ( \20756 , RIee1a950_4761, \9371 );
and \U$11634 ( \20757 , RIde906b0_294, \9373 );
and \U$11635 ( \20758 , RIde8cba0_276, \9375 );
and \U$11636 ( \20759 , RIfe82f20_7834, \9377 );
and \U$11637 ( \20760 , RIfe82db8_7833, \9379 );
and \U$11638 ( \20761 , RIee1a248_4756, \9381 );
and \U$11639 ( \20762 , RIfe831f0_7836, \9383 );
and \U$11640 ( \20763 , RIfcc2390_7232, \9385 );
and \U$11641 ( \20764 , RIee195a0_4747, \9387 );
and \U$11642 ( \20765 , RIfcbe718_7189, \9389 );
and \U$11643 ( \20766 , RIfea9e18_8249, \9391 );
and \U$11644 ( \20767 , RIfc43220_5786, \9393 );
and \U$11645 ( \20768 , RIe167868_2555, \9395 );
and \U$11646 ( \20769 , RIe164cd0_2524, \9397 );
and \U$11647 ( \20770 , RIe161fd0_2492, \9399 );
and \U$11648 ( \20771 , RIee36f88_5084, \9401 );
and \U$11649 ( \20772 , RIe15f2d0_2460, \9403 );
and \U$11650 ( \20773 , RIee35ea8_5072, \9405 );
and \U$11651 ( \20774 , RIe15c5d0_2428, \9407 );
and \U$11652 ( \20775 , RIe156bd0_2364, \9409 );
and \U$11653 ( \20776 , RIe153ed0_2332, \9411 );
and \U$11654 ( \20777 , RIfe83628_7839, \9413 );
and \U$11655 ( \20778 , RIe1511d0_2300, \9415 );
and \U$11656 ( \20779 , RIfebfda8_8303, \9417 );
and \U$11657 ( \20780 , RIe14e4d0_2268, \9419 );
and \U$11658 ( \20781 , RIfebfc40_8302, \9421 );
and \U$11659 ( \20782 , RIe14b7d0_2236, \9423 );
and \U$11660 ( \20783 , RIe148ad0_2204, \9425 );
and \U$11661 ( \20784 , RIe145dd0_2172, \9427 );
and \U$11662 ( \20785 , RIee34120_5051, \9429 );
and \U$11663 ( \20786 , RIee32ed8_5038, \9431 );
and \U$11664 ( \20787 , RIee31df8_5026, \9433 );
and \U$11665 ( \20788 , RIfcc1f58_7229, \9435 );
and \U$11666 ( \20789 , RIe140ad8_2113, \9437 );
and \U$11667 ( \20790 , RIdf3e878_2088, \9439 );
and \U$11668 ( \20791 , RIfe834c0_7838, \9441 );
and \U$11669 ( \20792 , RIdf3a390_2039, \9443 );
and \U$11670 ( \20793 , RIfc5a6c8_6051, \9445 );
and \U$11671 ( \20794 , RIfc91e20_6682, \9447 );
and \U$11672 ( \20795 , RIee2e888_4988, \9449 );
and \U$11673 ( \20796 , RIfc96a10_6736, \9451 );
and \U$11674 ( \20797 , RIdf35098_1980, \9453 );
and \U$11675 ( \20798 , RIfeab600_8266, \9455 );
and \U$11676 ( \20799 , RIdf30bb0_1931, \9457 );
and \U$11677 ( \20800 , RIfeab768_8267, \9459 );
or \U$11678 ( \20801 , \20737 , \20738 , \20739 , \20740 , \20741 , \20742 , \20743 , \20744 , \20745 , \20746 , \20747 , \20748 , \20749 , \20750 , \20751 , \20752 , \20753 , \20754 , \20755 , \20756 , \20757 , \20758 , \20759 , \20760 , \20761 , \20762 , \20763 , \20764 , \20765 , \20766 , \20767 , \20768 , \20769 , \20770 , \20771 , \20772 , \20773 , \20774 , \20775 , \20776 , \20777 , \20778 , \20779 , \20780 , \20781 , \20782 , \20783 , \20784 , \20785 , \20786 , \20787 , \20788 , \20789 , \20790 , \20791 , \20792 , \20793 , \20794 , \20795 , \20796 , \20797 , \20798 , \20799 , \20800 );
and \U$11679 ( \20802 , RIfcbe9e8_7191, \9462 );
and \U$11680 ( \20803 , RIfc79fa0_6410, \9464 );
and \U$11681 ( \20804 , RIfc96740_6734, \9466 );
and \U$11682 ( \20805 , RIfc92258_6685, \9468 );
and \U$11683 ( \20806 , RIfea7118_8217, \9470 );
and \U$11684 ( \20807 , RIfea95a8_8243, \9472 );
and \U$11685 ( \20808 , RIdf26020_1809, \9474 );
and \U$11686 ( \20809 , RIdf24400_1789, \9476 );
and \U$11687 ( \20810 , RIfc79a00_6406, \9478 );
and \U$11688 ( \20811 , RIfc5add0_6056, \9480 );
and \U$11689 ( \20812 , RIfce5d18_7637, \9482 );
and \U$11690 ( \20813 , RIfc92690_6688, \9484 );
and \U$11691 ( \20814 , RIfce3018_7605, \9486 );
and \U$11692 ( \20815 , RIdf1f270_1731, \9488 );
and \U$11693 ( \20816 , RIfc79730_6404, \9490 );
and \U$11694 ( \20817 , RIdf19000_1661, \9492 );
and \U$11695 ( \20818 , RIdf168a0_1633, \9494 );
and \U$11696 ( \20819 , RIdf13ba0_1601, \9496 );
and \U$11697 ( \20820 , RIdf10ea0_1569, \9498 );
and \U$11698 ( \20821 , RIdf0e1a0_1537, \9500 );
and \U$11699 ( \20822 , RIdf0b4a0_1505, \9502 );
and \U$11700 ( \20823 , RIdf087a0_1473, \9504 );
and \U$11701 ( \20824 , RIdf05aa0_1441, \9506 );
and \U$11702 ( \20825 , RIdf02da0_1409, \9508 );
and \U$11703 ( \20826 , RIdefd3a0_1345, \9510 );
and \U$11704 ( \20827 , RIdefa6a0_1313, \9512 );
and \U$11705 ( \20828 , RIdef79a0_1281, \9514 );
and \U$11706 ( \20829 , RIdef4ca0_1249, \9516 );
and \U$11707 ( \20830 , RIdef1fa0_1217, \9518 );
and \U$11708 ( \20831 , RIdeef2a0_1185, \9520 );
and \U$11709 ( \20832 , RIdeec5a0_1153, \9522 );
and \U$11710 ( \20833 , RIdee98a0_1121, \9524 );
and \U$11711 ( \20834 , RIfc5b7a8_6063, \9526 );
and \U$11712 ( \20835 , RIfc5b640_6062, \9528 );
and \U$11713 ( \20836 , RIfc931d0_6696, \9530 );
and \U$11714 ( \20837 , RIfcecac8_7715, \9532 );
and \U$11715 ( \20838 , RIdee4710_1063, \9534 );
and \U$11716 ( \20839 , RIdee26b8_1040, \9536 );
and \U$11717 ( \20840 , RIdee07c8_1018, \9538 );
and \U$11718 ( \20841 , RIdede4a0_993, \9540 );
and \U$11719 ( \20842 , RIfcbf0f0_7196, \9542 );
and \U$11720 ( \20843 , RIfcbf528_7199, \9544 );
and \U$11721 ( \20844 , RIfc792f8_6401, \9546 );
and \U$11722 ( \20845 , RIfc93068_6695, \9548 );
and \U$11723 ( \20846 , RIded91a8_934, \9550 );
and \U$11724 ( \20847 , RIded6d18_908, \9552 );
and \U$11725 ( \20848 , RIded4e28_886, \9554 );
and \U$11726 ( \20849 , RIded2998_860, \9556 );
and \U$11727 ( \20850 , RIded00d0_831, \9558 );
and \U$11728 ( \20851 , RIdecd3d0_799, \9560 );
and \U$11729 ( \20852 , RIdeca6d0_767, \9562 );
and \U$11730 ( \20853 , RIdec79d0_735, \9564 );
and \U$11731 ( \20854 , RIdeb3ed0_511, \9566 );
and \U$11732 ( \20855 , RIde958b8_319, \9568 );
and \U$11733 ( \20856 , RIe16dad8_2625, \9570 );
and \U$11734 ( \20857 , RIe1598d0_2396, \9572 );
and \U$11735 ( \20858 , RIe1430d0_2140, \9574 );
and \U$11736 ( \20859 , RIdf37ac8_2010, \9576 );
and \U$11737 ( \20860 , RIdf2c128_1878, \9578 );
and \U$11738 ( \20861 , RIdf1c9a8_1702, \9580 );
and \U$11739 ( \20862 , RIdf000a0_1377, \9582 );
and \U$11740 ( \20863 , RIdee6ba0_1089, \9584 );
and \U$11741 ( \20864 , RIdedb908_962, \9586 );
and \U$11742 ( \20865 , RIde7b800_192, \9588 );
or \U$11743 ( \20866 , \20802 , \20803 , \20804 , \20805 , \20806 , \20807 , \20808 , \20809 , \20810 , \20811 , \20812 , \20813 , \20814 , \20815 , \20816 , \20817 , \20818 , \20819 , \20820 , \20821 , \20822 , \20823 , \20824 , \20825 , \20826 , \20827 , \20828 , \20829 , \20830 , \20831 , \20832 , \20833 , \20834 , \20835 , \20836 , \20837 , \20838 , \20839 , \20840 , \20841 , \20842 , \20843 , \20844 , \20845 , \20846 , \20847 , \20848 , \20849 , \20850 , \20851 , \20852 , \20853 , \20854 , \20855 , \20856 , \20857 , \20858 , \20859 , \20860 , \20861 , \20862 , \20863 , \20864 , \20865 );
or \U$11744 ( \20867 , \20801 , \20866 );
_DC g5673 ( \20868_nG5673 , \20867 , \9597 );
and \U$11745 ( \20869 , RIe19cf68_3163, \9059 );
and \U$11746 ( \20870 , RIe19a268_3131, \9061 );
and \U$11747 ( \20871 , RIfc8d7d0_6632, \9063 );
and \U$11748 ( \20872 , RIe197568_3099, \9065 );
and \U$11749 ( \20873 , RIfc561e0_6002, \9067 );
and \U$11750 ( \20874 , RIe194868_3067, \9069 );
and \U$11751 ( \20875 , RIe191b68_3035, \9071 );
and \U$11752 ( \20876 , RIe18ee68_3003, \9073 );
and \U$11753 ( \20877 , RIe189468_2939, \9075 );
and \U$11754 ( \20878 , RIe186768_2907, \9077 );
and \U$11755 ( \20879 , RIf143330_5224, \9079 );
and \U$11756 ( \20880 , RIe183a68_2875, \9081 );
and \U$11757 ( \20881 , RIfc7d948_6451, \9083 );
and \U$11758 ( \20882 , RIe180d68_2843, \9085 );
and \U$11759 ( \20883 , RIe17e068_2811, \9087 );
and \U$11760 ( \20884 , RIe17b368_2779, \9089 );
and \U$11761 ( \20885 , RIfc564b0_6004, \9091 );
and \U$11762 ( \20886 , RIfcd6700_7462, \9093 );
and \U$11763 ( \20887 , RIfc461f0_5820, \9095 );
and \U$11764 ( \20888 , RIe175698_2713, \9097 );
and \U$11765 ( \20889 , RIfc46088_5819, \9099 );
and \U$11766 ( \20890 , RIfc45f20_5818, \9101 );
and \U$11767 ( \20891 , RIfc7dc18_6453, \9103 );
and \U$11768 ( \20892 , RIfcd69d0_7464, \9105 );
and \U$11769 ( \20893 , RIfc98630_6756, \9107 );
and \U$11770 ( \20894 , RIfcc2a98_7237, \9109 );
and \U$11771 ( \20895 , RIfc7d510_6448, \9111 );
and \U$11772 ( \20896 , RIe173208_2687, \9113 );
and \U$11773 ( \20897 , RIfc8e478_6641, \9115 );
and \U$11774 ( \20898 , RIfc45ae8_5815, \9117 );
and \U$11775 ( \20899 , RIfc8e8b0_6644, \9119 );
and \U$11776 ( \20900 , RIfc45980_5814, \9121 );
and \U$11777 ( \20901 , RIfe82ae8_7831, \9123 );
and \U$11778 ( \20902 , RIe2232c0_4690, \9125 );
and \U$11779 ( \20903 , RIf16ba10_5684, \9127 );
and \U$11780 ( \20904 , RIe2205c0_4658, \9129 );
and \U$11781 ( \20905 , RIfcd24e8_7415, \9131 );
and \U$11782 ( \20906 , RIe21d8c0_4626, \9133 );
and \U$11783 ( \20907 , RIe217ec0_4562, \9135 );
and \U$11784 ( \20908 , RIe2151c0_4530, \9137 );
and \U$11785 ( \20909 , RIfebf268_8295, \9139 );
and \U$11786 ( \20910 , RIe2124c0_4498, \9141 );
and \U$11787 ( \20911 , RIf168d10_5652, \9143 );
and \U$11788 ( \20912 , RIe20f7c0_4466, \9145 );
and \U$11789 ( \20913 , RIfc7d240_6446, \9147 );
and \U$11790 ( \20914 , RIe20cac0_4434, \9149 );
and \U$11791 ( \20915 , RIe209dc0_4402, \9151 );
and \U$11792 ( \20916 , RIe2070c0_4370, \9153 );
and \U$11793 ( \20917 , RIf166e20_5630, \9155 );
and \U$11794 ( \20918 , RIfebf6a0_8298, \9157 );
and \U$11795 ( \20919 , RIfebf808_8299, \9159 );
and \U$11796 ( \20920 , RIfebf538_8297, \9161 );
and \U$11797 ( \20921 , RIfc8eb80_6646, \9163 );
and \U$11798 ( \20922 , RIf164120_5598, \9165 );
and \U$11799 ( \20923 , RIfc453e0_5810, \9167 );
and \U$11800 ( \20924 , RIf161b28_5571, \9169 );
and \U$11801 ( \20925 , RIf15fc38_5549, \9171 );
and \U$11802 ( \20926 , RIf15dd48_5527, \9173 );
and \U$11803 ( \20927 , RIe1fc968_4251, \9175 );
and \U$11804 ( \20928 , RIe1fb888_4239, \9177 );
and \U$11805 ( \20929 , RIfebf3d0_8296, \9179 );
and \U$11806 ( \20930 , RIf15b318_5497, \9181 );
and \U$11807 ( \20931 , RIfca2518_6869, \9183 );
and \U$11808 ( \20932 , RIfc8f120_6650, \9185 );
or \U$11809 ( \20933 , \20869 , \20870 , \20871 , \20872 , \20873 , \20874 , \20875 , \20876 , \20877 , \20878 , \20879 , \20880 , \20881 , \20882 , \20883 , \20884 , \20885 , \20886 , \20887 , \20888 , \20889 , \20890 , \20891 , \20892 , \20893 , \20894 , \20895 , \20896 , \20897 , \20898 , \20899 , \20900 , \20901 , \20902 , \20903 , \20904 , \20905 , \20906 , \20907 , \20908 , \20909 , \20910 , \20911 , \20912 , \20913 , \20914 , \20915 , \20916 , \20917 , \20918 , \20919 , \20920 , \20921 , \20922 , \20923 , \20924 , \20925 , \20926 , \20927 , \20928 , \20929 , \20930 , \20931 , \20932 );
and \U$11810 ( \20934 , RIfebfad8_8301, \9188 );
and \U$11811 ( \20935 , RIfebf970_8300, \9190 );
and \U$11812 ( \20936 , RIfc7cca0_6442, \9192 );
and \U$11813 ( \20937 , RIe1f9dd0_4220, \9194 );
and \U$11814 ( \20938 , RIfe82c50_7832, \9196 );
and \U$11815 ( \20939 , RIf155648_5431, \9198 );
and \U$11816 ( \20940 , RIfc8f288_6651, \9200 );
and \U$11817 ( \20941 , RIe1f4f10_4164, \9202 );
and \U$11818 ( \20942 , RIf152d80_5402, \9204 );
and \U$11819 ( \20943 , RIfc8f828_6655, \9206 );
and \U$11820 ( \20944 , RIfcb3b88_7067, \9208 );
and \U$11821 ( \20945 , RIe1f2d50_4140, \9210 );
and \U$11822 ( \20946 , RIfc445d0_5800, \9212 );
and \U$11823 ( \20947 , RIfc8faf8_6657, \9214 );
and \U$11824 ( \20948 , RIf14da88_5343, \9216 );
and \U$11825 ( \20949 , RIe1eda58_4081, \9218 );
and \U$11826 ( \20950 , RIe1eb028_4051, \9220 );
and \U$11827 ( \20951 , RIe1e8328_4019, \9222 );
and \U$11828 ( \20952 , RIe1e5628_3987, \9224 );
and \U$11829 ( \20953 , RIe1e2928_3955, \9226 );
and \U$11830 ( \20954 , RIe1dfc28_3923, \9228 );
and \U$11831 ( \20955 , RIe1dcf28_3891, \9230 );
and \U$11832 ( \20956 , RIe1da228_3859, \9232 );
and \U$11833 ( \20957 , RIe1d7528_3827, \9234 );
and \U$11834 ( \20958 , RIe1d1b28_3763, \9236 );
and \U$11835 ( \20959 , RIe1cee28_3731, \9238 );
and \U$11836 ( \20960 , RIe1cc128_3699, \9240 );
and \U$11837 ( \20961 , RIe1c9428_3667, \9242 );
and \U$11838 ( \20962 , RIe1c6728_3635, \9244 );
and \U$11839 ( \20963 , RIe1c3a28_3603, \9246 );
and \U$11840 ( \20964 , RIe1c0d28_3571, \9248 );
and \U$11841 ( \20965 , RIe1be028_3539, \9250 );
and \U$11842 ( \20966 , RIfc7bff8_6433, \9252 );
and \U$11843 ( \20967 , RIfc44030_5796, \9254 );
and \U$11844 ( \20968 , RIe1b9000_3482, \9256 );
and \U$11845 ( \20969 , RIe1b6fa8_3459, \9258 );
and \U$11846 ( \20970 , RIfcbdd40_7182, \9260 );
and \U$11847 ( \20971 , RIfc8ff30_6660, \9262 );
and \U$11848 ( \20972 , RIe1b50b8_3437, \9264 );
and \U$11849 ( \20973 , RIe1b3d08_3423, \9266 );
and \U$11850 ( \20974 , RIfcbe178_7185, \9268 );
and \U$11851 ( \20975 , RIfc43d60_5794, \9270 );
and \U$11852 ( \20976 , RIe1b2520_3406, \9272 );
and \U$11853 ( \20977 , RIe1b0798_3385, \9274 );
and \U$11854 ( \20978 , RIfcdb5c0_7518, \9276 );
and \U$11855 ( \20979 , RIfc7ba58_6429, \9278 );
and \U$11856 ( \20980 , RIe1ac148_3335, \9280 );
and \U$11857 ( \20981 , RIe1aa960_3318, \9282 );
and \U$11858 ( \20982 , RIe1a8368_3291, \9284 );
and \U$11859 ( \20983 , RIe1a5668_3259, \9286 );
and \U$11860 ( \20984 , RIe1a2968_3227, \9288 );
and \U$11861 ( \20985 , RIe19fc68_3195, \9290 );
and \U$11862 ( \20986 , RIe18c168_2971, \9292 );
and \U$11863 ( \20987 , RIe178668_2747, \9294 );
and \U$11864 ( \20988 , RIe225fc0_4722, \9296 );
and \U$11865 ( \20989 , RIe21abc0_4594, \9298 );
and \U$11866 ( \20990 , RIe2043c0_4338, \9300 );
and \U$11867 ( \20991 , RIe1fe420_4270, \9302 );
and \U$11868 ( \20992 , RIe1f77d8_4193, \9304 );
and \U$11869 ( \20993 , RIe1f0320_4110, \9306 );
and \U$11870 ( \20994 , RIe1d4828_3795, \9308 );
and \U$11871 ( \20995 , RIe1bb328_3507, \9310 );
and \U$11872 ( \20996 , RIe1ae1a0_3358, \9312 );
and \U$11873 ( \20997 , RIe1707d8_2657, \9314 );
or \U$11874 ( \20998 , \20934 , \20935 , \20936 , \20937 , \20938 , \20939 , \20940 , \20941 , \20942 , \20943 , \20944 , \20945 , \20946 , \20947 , \20948 , \20949 , \20950 , \20951 , \20952 , \20953 , \20954 , \20955 , \20956 , \20957 , \20958 , \20959 , \20960 , \20961 , \20962 , \20963 , \20964 , \20965 , \20966 , \20967 , \20968 , \20969 , \20970 , \20971 , \20972 , \20973 , \20974 , \20975 , \20976 , \20977 , \20978 , \20979 , \20980 , \20981 , \20982 , \20983 , \20984 , \20985 , \20986 , \20987 , \20988 , \20989 , \20990 , \20991 , \20992 , \20993 , \20994 , \20995 , \20996 , \20997 );
or \U$11875 ( \20999 , \20933 , \20998 );
_DC g56f7 ( \21000_nG56f7 , \20999 , \9323 );
xor g56f8 ( \21001_nG56f8 , \20868_nG5673 , \21000_nG56f7 );
buf \U$11876 ( \21002 , \21001_nG56f8 );
xor \U$11877 ( \21003 , \21002 , \20556 );
not \U$11878 ( \21004 , \20557 );
and \U$11879 ( \21005 , \21003 , \21004 );
and \U$11880 ( \21006 , \10687 , \21005 );
and \U$11881 ( \21007 , \10988 , \20557 );
nor \U$11882 ( \21008 , \21006 , \21007 );
and \U$11883 ( \21009 , \20556 , \19531 );
not \U$11884 ( \21010 , \21009 );
and \U$11885 ( \21011 , \21002 , \21010 );
xnor \U$11886 ( \21012 , \21008 , \21011 );
xor \U$11887 ( \21013 , \20736 , \21012 );
and \U$11888 ( \21014 , \19032 , \11574 );
and \U$11889 ( \21015 , \19558 , \11278 );
nor \U$11890 ( \21016 , \21014 , \21015 );
xnor \U$11891 ( \21017 , \21016 , \11580 );
and \U$11892 ( \21018 , \17627 , \12790 );
and \U$11893 ( \21019 , \18035 , \12461 );
nor \U$11894 ( \21020 , \21018 , \21019 );
xnor \U$11895 ( \21021 , \21020 , \12780 );
xor \U$11896 ( \21022 , \21017 , \21021 );
and \U$11897 ( \21023 , \14950 , \15336 );
and \U$11898 ( \21024 , \15321 , \14963 );
nor \U$11899 ( \21025 , \21023 , \21024 );
xnor \U$11900 ( \21026 , \21025 , \15342 );
xor \U$11901 ( \21027 , \21022 , \21026 );
xor \U$11902 ( \21028 , \21013 , \21027 );
and \U$11903 ( \21029 , \20544 , \10983 );
_DC g65aa ( \21030_nG65aa , \20867 , \9597 );
_DC g65ab ( \21031_nG65ab , \20999 , \9323 );
and g65ac ( \21032_nG65ac , \21030_nG65aa , \21031_nG65ab );
buf \U$11904 ( \21033 , \21032_nG65ac );
and \U$11905 ( \21034 , \21033 , \10691 );
nor \U$11906 ( \21035 , \21029 , \21034 );
xnor \U$11907 ( \21036 , \21035 , \10980 );
not \U$11908 ( \21037 , \20558 );
and \U$11909 ( \21038 , \21037 , \21011 );
xor \U$11910 ( \21039 , \21036 , \21038 );
and \U$11911 ( \21040 , \13679 , \16635 );
and \U$11912 ( \21041 , \14024 , \16301 );
nor \U$11913 ( \21042 , \21040 , \21041 );
xnor \U$11914 ( \21043 , \21042 , \16625 );
xor \U$11915 ( \21044 , \21039 , \21043 );
and \U$11916 ( \21045 , \12448 , \18090 );
and \U$11917 ( \21046 , \12769 , \17655 );
nor \U$11918 ( \21047 , \21045 , \21046 );
xnor \U$11919 ( \21048 , \21047 , \18046 );
xor \U$11920 ( \21049 , \21044 , \21048 );
xor \U$11921 ( \21050 , \21028 , \21049 );
xor \U$11922 ( \21051 , \20727 , \21050 );
and \U$11923 ( \21052 , \20589 , \20593 );
and \U$11924 ( \21053 , \20593 , \20595 );
and \U$11925 ( \21054 , \20589 , \20595 );
or \U$11926 ( \21055 , \21052 , \21053 , \21054 );
and \U$11927 ( \21056 , \20277 , \20559 );
and \U$11928 ( \21057 , \20559 , \20574 );
and \U$11929 ( \21058 , \20277 , \20574 );
or \U$11930 ( \21059 , \21056 , \21057 , \21058 );
xor \U$11931 ( \21060 , \21055 , \21059 );
and \U$11932 ( \21061 , \20267 , \20271 );
and \U$11933 ( \21062 , \20271 , \20276 );
and \U$11934 ( \21063 , \20267 , \20276 );
or \U$11935 ( \21064 , \21061 , \21062 , \21063 );
and \U$11936 ( \21065 , \20547 , \20551 );
and \U$11937 ( \21066 , \20551 , \20558 );
and \U$11938 ( \21067 , \20547 , \20558 );
or \U$11939 ( \21068 , \21065 , \21066 , \21067 );
xor \U$11940 ( \21069 , \21064 , \21068 );
and \U$11941 ( \21070 , \20564 , \20568 );
and \U$11942 ( \21071 , \20568 , \20573 );
and \U$11943 ( \21072 , \20564 , \20573 );
or \U$11944 ( \21073 , \21070 , \21071 , \21072 );
xor \U$11945 ( \21074 , \21069 , \21073 );
xor \U$11946 ( \21075 , \21060 , \21074 );
xor \U$11947 ( \21076 , \21051 , \21075 );
and \U$11948 ( \21077 , \20263 , \20575 );
and \U$11949 ( \21078 , \20575 , \20597 );
and \U$11950 ( \21079 , \20263 , \20597 );
or \U$11951 ( \21080 , \21077 , \21078 , \21079 );
xor \U$11952 ( \21081 , \21076 , \21080 );
and \U$11953 ( \21082 , \20598 , \20602 );
and \U$11954 ( \21083 , \20603 , \20606 );
or \U$11955 ( \21084 , \21082 , \21083 );
xor \U$11956 ( \21085 , \21081 , \21084 );
buf g9bdb ( \21086_nG9bdb , \21085 );
and \U$11957 ( \21087 , \10704 , \21086_nG9bdb );
or \U$11958 ( \21088 , \20723 , \21087 );
xor \U$11959 ( \21089 , \10703 , \21088 );
buf \U$11960 ( \21090 , \21089 );
buf \U$11962 ( \21091 , \21090 );
xor \U$11963 ( \21092 , \20722 , \21091 );
buf \U$11964 ( \21093 , \21092 );
xor \U$11965 ( \21094 , \20695 , \21093 );
and \U$11966 ( \21095 , \20183 , \20222 );
and \U$11967 ( \21096 , \20183 , \20228 );
and \U$11968 ( \21097 , \20222 , \20228 );
or \U$11969 ( \21098 , \21095 , \21096 , \21097 );
buf \U$11970 ( \21099 , \21098 );
xor \U$11971 ( \21100 , \21094 , \21099 );
and \U$11972 ( \21101 , \20631 , \21100 );
and \U$11973 ( \21102 , \20621 , \20625 );
and \U$11974 ( \21103 , \20621 , \20630 );
and \U$11975 ( \21104 , \20625 , \20630 );
or \U$11976 ( \21105 , \21102 , \21103 , \21104 );
xor \U$11977 ( \21106 , \21101 , \21105 );
and \U$11978 ( \21107 , RIdec4fa0_705, \9059 );
and \U$11979 ( \21108 , RIdec22a0_673, \9061 );
and \U$11980 ( \21109 , RIee1fdb0_4821, \9063 );
and \U$11981 ( \21110 , RIdebf5a0_641, \9065 );
and \U$11982 ( \21111 , RIee1f270_4813, \9067 );
and \U$11983 ( \21112 , RIdebc8a0_609, \9069 );
and \U$11984 ( \21113 , RIdeb9ba0_577, \9071 );
and \U$11985 ( \21114 , RIdeb6ea0_545, \9073 );
and \U$11986 ( \21115 , RIee1ecd0_4809, \9075 );
and \U$11987 ( \21116 , RIdeb14a0_481, \9077 );
and \U$11988 ( \21117 , RIee1e730_4805, \9079 );
and \U$11989 ( \21118 , RIdeae7a0_449, \9081 );
and \U$11990 ( \21119 , RIee1d920_4795, \9083 );
and \U$11991 ( \21120 , RIdea9a48_417, \9085 );
and \U$11992 ( \21121 , RIdea3148_385, \9087 );
and \U$11993 ( \21122 , RIde9c848_353, \9089 );
and \U$11994 ( \21123 , RIee1cb10_4785, \9091 );
and \U$11995 ( \21124 , RIee1ba30_4773, \9093 );
and \U$11996 ( \21125 , RIee1b1c0_4767, \9095 );
and \U$11997 ( \21126 , RIfec04b0_8308, \9097 );
and \U$11998 ( \21127 , RIfe850e0_7858, \9099 );
and \U$11999 ( \21128 , RIde8d230_278, \9101 );
and \U$12000 ( \21129 , RIfea9cb0_8248, \9103 );
and \U$12001 ( \21130 , RIfe84f78_7857, \9105 );
and \U$12002 ( \21131 , RIee1a3b0_4757, \9107 );
and \U$12003 ( \21132 , RIfe853b0_7860, \9109 );
and \U$12004 ( \21133 , RIee199d8_4750, \9111 );
and \U$12005 ( \21134 , RIfe85248_7859, \9113 );
and \U$12006 ( \21135 , RIee39148_5108, \9115 );
and \U$12007 ( \21136 , RIe16b378_2597, \9117 );
and \U$12008 ( \21137 , RIee38608_5100, \9119 );
and \U$12009 ( \21138 , RIe167b38_2557, \9121 );
and \U$12010 ( \21139 , RIe164fa0_2526, \9123 );
and \U$12011 ( \21140 , RIe1622a0_2494, \9125 );
and \U$12012 ( \21141 , RIfe85950_7864, \9127 );
and \U$12013 ( \21142 , RIe15f5a0_2462, \9129 );
and \U$12014 ( \21143 , RIee36010_5073, \9131 );
and \U$12015 ( \21144 , RIe15c8a0_2430, \9133 );
and \U$12016 ( \21145 , RIe156ea0_2366, \9135 );
and \U$12017 ( \21146 , RIe1541a0_2334, \9137 );
and \U$12018 ( \21147 , RIfe85c20_7866, \9139 );
and \U$12019 ( \21148 , RIe1514a0_2302, \9141 );
and \U$12020 ( \21149 , RIee34dc8_5060, \9143 );
and \U$12021 ( \21150 , RIe14e7a0_2270, \9145 );
and \U$12022 ( \21151 , RIfc861b0_6548, \9147 );
and \U$12023 ( \21152 , RIe14baa0_2238, \9149 );
and \U$12024 ( \21153 , RIe148da0_2206, \9151 );
and \U$12025 ( \21154 , RIe1460a0_2174, \9153 );
and \U$12026 ( \21155 , RIee343f0_5053, \9155 );
and \U$12027 ( \21156 , RIfe85518_7861, \9157 );
and \U$12028 ( \21157 , RIfe857e8_7863, \9159 );
and \U$12029 ( \21158 , RIfe85680_7862, \9161 );
and \U$12030 ( \21159 , RIe140c40_2114, \9163 );
and \U$12031 ( \21160 , RIdf3eb48_2090, \9165 );
and \U$12032 ( \21161 , RIdf3c820_2065, \9167 );
and \U$12033 ( \21162 , RIdf3a660_2041, \9169 );
and \U$12034 ( \21163 , RIfc9d4f0_6812, \9171 );
and \U$12035 ( \21164 , RIee2f698_4998, \9173 );
and \U$12036 ( \21165 , RIfc52298_5957, \9175 );
and \U$12037 ( \21166 , RIee2d4d8_4974, \9177 );
and \U$12038 ( \21167 , RIdf35368_1982, \9179 );
and \U$12039 ( \21168 , RIdf32ed8_1956, \9181 );
and \U$12040 ( \21169 , RIdf30e80_1933, \9183 );
and \U$12041 ( \21170 , RIfe85ab8_7865, \9185 );
or \U$12042 ( \21171 , \21107 , \21108 , \21109 , \21110 , \21111 , \21112 , \21113 , \21114 , \21115 , \21116 , \21117 , \21118 , \21119 , \21120 , \21121 , \21122 , \21123 , \21124 , \21125 , \21126 , \21127 , \21128 , \21129 , \21130 , \21131 , \21132 , \21133 , \21134 , \21135 , \21136 , \21137 , \21138 , \21139 , \21140 , \21141 , \21142 , \21143 , \21144 , \21145 , \21146 , \21147 , \21148 , \21149 , \21150 , \21151 , \21152 , \21153 , \21154 , \21155 , \21156 , \21157 , \21158 , \21159 , \21160 , \21161 , \21162 , \21163 , \21164 , \21165 , \21166 , \21167 , \21168 , \21169 , \21170 );
and \U$12043 ( \21172 , RIee2b8b8_4954, \9188 );
and \U$12044 ( \21173 , RIee29f68_4936, \9190 );
and \U$12045 ( \21174 , RIee28bb8_4922, \9192 );
and \U$12046 ( \21175 , RIee27970_4909, \9194 );
and \U$12047 ( \21176 , RIdf2a0d0_1855, \9196 );
and \U$12048 ( \21177 , RIfe84e10_7856, \9198 );
and \U$12049 ( \21178 , RIdf262f0_1811, \9200 );
and \U$12050 ( \21179 , RIfe84ca8_7855, \9202 );
and \U$12051 ( \21180 , RIee27100_4903, \9204 );
and \U$12052 ( \21181 , RIee26b60_4899, \9206 );
and \U$12053 ( \21182 , RIfcd32f8_7425, \9208 );
and \U$12054 ( \21183 , RIee265c0_4895, \9210 );
and \U$12055 ( \21184 , RIfc9e300_6822, \9212 );
and \U$12056 ( \21185 , RIdf1f540_1733, \9214 );
and \U$12057 ( \21186 , RIee25eb8_4890, \9216 );
and \U$12058 ( \21187 , RIfe84b40_7854, \9218 );
and \U$12059 ( \21188 , RIdf16b70_1635, \9220 );
and \U$12060 ( \21189 , RIdf13e70_1603, \9222 );
and \U$12061 ( \21190 , RIdf11170_1571, \9224 );
and \U$12062 ( \21191 , RIdf0e470_1539, \9226 );
and \U$12063 ( \21192 , RIdf0b770_1507, \9228 );
and \U$12064 ( \21193 , RIdf08a70_1475, \9230 );
and \U$12065 ( \21194 , RIdf05d70_1443, \9232 );
and \U$12066 ( \21195 , RIdf03070_1411, \9234 );
and \U$12067 ( \21196 , RIdefd670_1347, \9236 );
and \U$12068 ( \21197 , RIdefa970_1315, \9238 );
and \U$12069 ( \21198 , RIdef7c70_1283, \9240 );
and \U$12070 ( \21199 , RIdef4f70_1251, \9242 );
and \U$12071 ( \21200 , RIdef2270_1219, \9244 );
and \U$12072 ( \21201 , RIdeef570_1187, \9246 );
and \U$12073 ( \21202 , RIdeec870_1155, \9248 );
and \U$12074 ( \21203 , RIdee9b70_1123, \9250 );
and \U$12075 ( \21204 , RIfec0348_8307, \9252 );
and \U$12076 ( \21205 , RIfcb54d8_7085, \9254 );
and \U$12077 ( \21206 , RIee23cf8_4866, \9256 );
and \U$12078 ( \21207 , RIfc54e30_5988, \9258 );
and \U$12079 ( \21208 , RIfec0078_8305, \9260 );
and \U$12080 ( \21209 , RIdee2988_1042, \9262 );
and \U$12081 ( \21210 , RIfec01e0_8306, \9264 );
and \U$12082 ( \21211 , RIdede770_995, \9266 );
and \U$12083 ( \21212 , RIfcd7ee8_7479, \9268 );
and \U$12084 ( \21213 , RIfcd43d8_7437, \9270 );
and \U$12085 ( \21214 , RIfc88eb0_6580, \9272 );
and \U$12086 ( \21215 , RIfc9e5d0_6824, \9274 );
and \U$12087 ( \21216 , RIded9478_936, \9276 );
and \U$12088 ( \21217 , RIded6fe8_910, \9278 );
and \U$12089 ( \21218 , RIded50f8_888, \9280 );
and \U$12090 ( \21219 , RIfeab330_8264, \9282 );
and \U$12091 ( \21220 , RIded03a0_833, \9284 );
and \U$12092 ( \21221 , RIdecd6a0_801, \9286 );
and \U$12093 ( \21222 , RIdeca9a0_769, \9288 );
and \U$12094 ( \21223 , RIdec7ca0_737, \9290 );
and \U$12095 ( \21224 , RIdeb41a0_513, \9292 );
and \U$12096 ( \21225 , RIde95f48_321, \9294 );
and \U$12097 ( \21226 , RIe16dda8_2627, \9296 );
and \U$12098 ( \21227 , RIe159ba0_2398, \9298 );
and \U$12099 ( \21228 , RIe1433a0_2142, \9300 );
and \U$12100 ( \21229 , RIdf37d98_2012, \9302 );
and \U$12101 ( \21230 , RIdf2c3f8_1880, \9304 );
and \U$12102 ( \21231 , RIdf1cc78_1704, \9306 );
and \U$12103 ( \21232 , RIdf00370_1379, \9308 );
and \U$12104 ( \21233 , RIdee6e70_1091, \9310 );
and \U$12105 ( \21234 , RIdedbbd8_964, \9312 );
and \U$12106 ( \21235 , RIde7be90_194, \9314 );
or \U$12107 ( \21236 , \21172 , \21173 , \21174 , \21175 , \21176 , \21177 , \21178 , \21179 , \21180 , \21181 , \21182 , \21183 , \21184 , \21185 , \21186 , \21187 , \21188 , \21189 , \21190 , \21191 , \21192 , \21193 , \21194 , \21195 , \21196 , \21197 , \21198 , \21199 , \21200 , \21201 , \21202 , \21203 , \21204 , \21205 , \21206 , \21207 , \21208 , \21209 , \21210 , \21211 , \21212 , \21213 , \21214 , \21215 , \21216 , \21217 , \21218 , \21219 , \21220 , \21221 , \21222 , \21223 , \21224 , \21225 , \21226 , \21227 , \21228 , \21229 , \21230 , \21231 , \21232 , \21233 , \21234 , \21235 );
or \U$12108 ( \21237 , \21171 , \21236 );
_DC g2871 ( \21238_nG2871 , \21237 , \9323 );
buf \U$12109 ( \21239 , \21238_nG2871 );
and \U$12110 ( \21240 , RIe19d238_3165, \9333 );
and \U$12111 ( \21241 , RIe19a538_3133, \9335 );
and \U$12112 ( \21242 , RIf145658_5249, \9337 );
and \U$12113 ( \21243 , RIe197838_3101, \9339 );
and \U$12114 ( \21244 , RIf1446e0_5238, \9341 );
and \U$12115 ( \21245 , RIe194b38_3069, \9343 );
and \U$12116 ( \21246 , RIe191e38_3037, \9345 );
and \U$12117 ( \21247 , RIe18f138_3005, \9347 );
and \U$12118 ( \21248 , RIe189738_2941, \9349 );
and \U$12119 ( \21249 , RIe186a38_2909, \9351 );
and \U$12120 ( \21250 , RIf143600_5226, \9353 );
and \U$12121 ( \21251 , RIe183d38_2877, \9355 );
and \U$12122 ( \21252 , RIf142c28_5219, \9357 );
and \U$12123 ( \21253 , RIe181038_2845, \9359 );
and \U$12124 ( \21254 , RIe17e338_2813, \9361 );
and \U$12125 ( \21255 , RIe17b638_2781, \9363 );
and \U$12126 ( \21256 , RIf1420e8_5211, \9365 );
and \U$12127 ( \21257 , RIf140a68_5195, \9367 );
and \U$12128 ( \21258 , RIf1401f8_5189, \9369 );
and \U$12129 ( \21259 , RIfebff10_8304, \9371 );
and \U$12130 ( \21260 , RIf13faf0_5184, \9373 );
and \U$12131 ( \21261 , RIf13ee48_5175, \9375 );
and \U$12132 ( \21262 , RIee3e2d8_5166, \9377 );
and \U$12133 ( \21263 , RIee3d1f8_5154, \9379 );
and \U$12134 ( \21264 , RIee3c118_5142, \9381 );
and \U$12135 ( \21265 , RIee3b038_5130, \9383 );
and \U$12136 ( \21266 , RIee39c88_5116, \9385 );
and \U$12137 ( \21267 , RIfe838f8_7841, \9387 );
and \U$12138 ( \21268 , RIf1701c8_5735, \9389 );
and \U$12139 ( \21269 , RIfc5ab00_6054, \9391 );
and \U$12140 ( \21270 , RIf16e008_5711, \9393 );
and \U$12141 ( \21271 , RIfcb0e88_7035, \9395 );
and \U$12142 ( \21272 , RIf16caf0_5696, \9397 );
and \U$12143 ( \21273 , RIe223590_4692, \9399 );
and \U$12144 ( \21274 , RIf16bce0_5686, \9401 );
and \U$12145 ( \21275 , RIe220890_4660, \9403 );
and \U$12146 ( \21276 , RIf16ac00_5674, \9405 );
and \U$12147 ( \21277 , RIe21db90_4628, \9407 );
and \U$12148 ( \21278 , RIe218190_4564, \9409 );
and \U$12149 ( \21279 , RIe215490_4532, \9411 );
and \U$12150 ( \21280 , RIf16a228_5667, \9413 );
and \U$12151 ( \21281 , RIe212790_4500, \9415 );
and \U$12152 ( \21282 , RIf168fe0_5654, \9417 );
and \U$12153 ( \21283 , RIe20fa90_4468, \9419 );
and \U$12154 ( \21284 , RIf167d98_5641, \9421 );
and \U$12155 ( \21285 , RIe20cd90_4436, \9423 );
and \U$12156 ( \21286 , RIe20a090_4404, \9425 );
and \U$12157 ( \21287 , RIe207390_4372, \9427 );
and \U$12158 ( \21288 , RIf1670f0_5632, \9429 );
and \U$12159 ( \21289 , RIf165ea8_5619, \9431 );
and \U$12160 ( \21290 , RIe202200_4314, \9433 );
and \U$12161 ( \21291 , RIfe83e98_7845, \9435 );
and \U$12162 ( \21292 , RIf164f30_5608, \9437 );
and \U$12163 ( \21293 , RIf1643f0_5600, \9439 );
and \U$12164 ( \21294 , RIfce8310_7664, \9441 );
and \U$12165 ( \21295 , RIf161df8_5573, \9443 );
and \U$12166 ( \21296 , RIf15ff08_5551, \9445 );
and \U$12167 ( \21297 , RIf15e018_5529, \9447 );
and \U$12168 ( \21298 , RIfe83d30_7844, \9449 );
and \U$12169 ( \21299 , RIfe84000_7846, \9451 );
and \U$12170 ( \21300 , RIf15cb00_5514, \9453 );
and \U$12171 ( \21301 , RIf15b5e8_5499, \9455 );
and \U$12172 ( \21302 , RIf15a508_5487, \9457 );
and \U$12173 ( \21303 , RIfc887a8_6575, \9459 );
or \U$12174 ( \21304 , \21240 , \21241 , \21242 , \21243 , \21244 , \21245 , \21246 , \21247 , \21248 , \21249 , \21250 , \21251 , \21252 , \21253 , \21254 , \21255 , \21256 , \21257 , \21258 , \21259 , \21260 , \21261 , \21262 , \21263 , \21264 , \21265 , \21266 , \21267 , \21268 , \21269 , \21270 , \21271 , \21272 , \21273 , \21274 , \21275 , \21276 , \21277 , \21278 , \21279 , \21280 , \21281 , \21282 , \21283 , \21284 , \21285 , \21286 , \21287 , \21288 , \21289 , \21290 , \21291 , \21292 , \21293 , \21294 , \21295 , \21296 , \21297 , \21298 , \21299 , \21300 , \21301 , \21302 , \21303 );
and \U$12175 ( \21305 , RIf158d20_5470, \9462 );
and \U$12176 ( \21306 , RIf157970_5456, \9464 );
and \U$12177 ( \21307 , RIf156cc8_5447, \9466 );
and \U$12178 ( \21308 , RIfe84438_7849, \9468 );
and \U$12179 ( \21309 , RIf156020_5438, \9470 );
and \U$12180 ( \21310 , RIfc51fc8_5955, \9472 );
and \U$12181 ( \21311 , RIf154568_5419, \9474 );
and \U$12182 ( \21312 , RIe1f51e0_4166, \9476 );
and \U$12183 ( \21313 , RIf153050_5404, \9478 );
and \U$12184 ( \21314 , RIf1519d0_5388, \9480 );
and \U$12185 ( \21315 , RIf150788_5375, \9482 );
and \U$12186 ( \21316 , RIfe842d0_7848, \9484 );
and \U$12187 ( \21317 , RIf14f810_5364, \9486 );
and \U$12188 ( \21318 , RIf14eb68_5355, \9488 );
and \U$12189 ( \21319 , RIf14dd58_5345, \9490 );
and \U$12190 ( \21320 , RIfe84168_7847, \9492 );
and \U$12191 ( \21321 , RIe1eb2f8_4053, \9494 );
and \U$12192 ( \21322 , RIe1e85f8_4021, \9496 );
and \U$12193 ( \21323 , RIe1e58f8_3989, \9498 );
and \U$12194 ( \21324 , RIe1e2bf8_3957, \9500 );
and \U$12195 ( \21325 , RIe1dfef8_3925, \9502 );
and \U$12196 ( \21326 , RIe1dd1f8_3893, \9504 );
and \U$12197 ( \21327 , RIe1da4f8_3861, \9506 );
and \U$12198 ( \21328 , RIe1d77f8_3829, \9508 );
and \U$12199 ( \21329 , RIe1d1df8_3765, \9510 );
and \U$12200 ( \21330 , RIe1cf0f8_3733, \9512 );
and \U$12201 ( \21331 , RIe1cc3f8_3701, \9514 );
and \U$12202 ( \21332 , RIe1c96f8_3669, \9516 );
and \U$12203 ( \21333 , RIe1c69f8_3637, \9518 );
and \U$12204 ( \21334 , RIe1c3cf8_3605, \9520 );
and \U$12205 ( \21335 , RIe1c0ff8_3573, \9522 );
and \U$12206 ( \21336 , RIe1be2f8_3541, \9524 );
and \U$12207 ( \21337 , RIf14c840_5330, \9526 );
and \U$12208 ( \21338 , RIf14b5f8_5317, \9528 );
and \U$12209 ( \21339 , RIfe83a60_7842, \9530 );
and \U$12210 ( \21340 , RIfe849d8_7853, \9532 );
and \U$12211 ( \21341 , RIfc74168_6343, \9534 );
and \U$12212 ( \21342 , RIf149b40_5298, \9536 );
and \U$12213 ( \21343 , RIfe83bc8_7843, \9538 );
and \U$12214 ( \21344 , RIfe84708_7851, \9540 );
and \U$12215 ( \21345 , RIf148d30_5288, \9542 );
and \U$12216 ( \21346 , RIf147ae8_5275, \9544 );
and \U$12217 ( \21347 , RIfe84870_7852, \9546 );
and \U$12218 ( \21348 , RIe1b0900_3386, \9548 );
and \U$12219 ( \21349 , RIf146fa8_5267, \9550 );
and \U$12220 ( \21350 , RIf146300_5258, \9552 );
and \U$12221 ( \21351 , RIfe845a0_7850, \9554 );
and \U$12222 ( \21352 , RIfe83790_7840, \9556 );
and \U$12223 ( \21353 , RIe1a8638_3293, \9558 );
and \U$12224 ( \21354 , RIe1a5938_3261, \9560 );
and \U$12225 ( \21355 , RIe1a2c38_3229, \9562 );
and \U$12226 ( \21356 , RIe19ff38_3197, \9564 );
and \U$12227 ( \21357 , RIe18c438_2973, \9566 );
and \U$12228 ( \21358 , RIe178938_2749, \9568 );
and \U$12229 ( \21359 , RIe226290_4724, \9570 );
and \U$12230 ( \21360 , RIe21ae90_4596, \9572 );
and \U$12231 ( \21361 , RIe204690_4340, \9574 );
and \U$12232 ( \21362 , RIe1fe6f0_4272, \9576 );
and \U$12233 ( \21363 , RIe1f7aa8_4195, \9578 );
and \U$12234 ( \21364 , RIe1f05f0_4112, \9580 );
and \U$12235 ( \21365 , RIe1d4af8_3797, \9582 );
and \U$12236 ( \21366 , RIe1bb5f8_3509, \9584 );
and \U$12237 ( \21367 , RIe1ae470_3360, \9586 );
and \U$12238 ( \21368 , RIe170aa8_2659, \9588 );
or \U$12239 ( \21369 , \21305 , \21306 , \21307 , \21308 , \21309 , \21310 , \21311 , \21312 , \21313 , \21314 , \21315 , \21316 , \21317 , \21318 , \21319 , \21320 , \21321 , \21322 , \21323 , \21324 , \21325 , \21326 , \21327 , \21328 , \21329 , \21330 , \21331 , \21332 , \21333 , \21334 , \21335 , \21336 , \21337 , \21338 , \21339 , \21340 , \21341 , \21342 , \21343 , \21344 , \21345 , \21346 , \21347 , \21348 , \21349 , \21350 , \21351 , \21352 , \21353 , \21354 , \21355 , \21356 , \21357 , \21358 , \21359 , \21360 , \21361 , \21362 , \21363 , \21364 , \21365 , \21366 , \21367 , \21368 );
or \U$12240 ( \21370 , \21304 , \21369 );
_DC g399e ( \21371_nG399e , \21370 , \9597 );
buf \U$12241 ( \21372 , \21371_nG399e );
xor \U$12242 ( \21373 , \21239 , \21372 );
and \U$12243 ( \21374 , RIdec4e38_704, \9059 );
and \U$12244 ( \21375 , RIdec2138_672, \9061 );
and \U$12245 ( \21376 , RIee1fc48_4820, \9063 );
and \U$12246 ( \21377 , RIdebf438_640, \9065 );
and \U$12247 ( \21378 , RIfc49490_5856, \9067 );
and \U$12248 ( \21379 , RIdebc738_608, \9069 );
and \U$12249 ( \21380 , RIdeb9a38_576, \9071 );
and \U$12250 ( \21381 , RIdeb6d38_544, \9073 );
and \U$12251 ( \21382 , RIfc48ef0_5852, \9075 );
and \U$12252 ( \21383 , RIdeb1338_480, \9077 );
and \U$12253 ( \21384 , RIfcd9b08_7499, \9079 );
and \U$12254 ( \21385 , RIdeae638_448, \9081 );
and \U$12255 ( \21386 , RIfc8b610_6608, \9083 );
and \U$12256 ( \21387 , RIdea9700_416, \9085 );
and \U$12257 ( \21388 , RIdea2e00_384, \9087 );
and \U$12258 ( \21389 , RIde9c500_352, \9089 );
and \U$12259 ( \21390 , RIee1c9a8_4784, \9091 );
and \U$12260 ( \21391 , RIee1b8c8_4772, \9093 );
and \U$12261 ( \21392 , RIfc80918_6485, \9095 );
and \U$12262 ( \21393 , RIfcdad50_7512, \9097 );
and \U$12263 ( \21394 , RIfe86e68_7879, \9099 );
and \U$12264 ( \21395 , RIde8cee8_277, \9101 );
and \U$12265 ( \21396 , RIfe86d00_7878, \9103 );
and \U$12266 ( \21397 , RIfec0d20_8314, \9105 );
and \U$12267 ( \21398 , RIde81098_219, \9107 );
and \U$12268 ( \21399 , RIfc8b8e0_6610, \9109 );
and \U$12269 ( \21400 , RIfcd2d58_7421, \9111 );
and \U$12270 ( \21401 , RIfce4530_7620, \9113 );
and \U$12271 ( \21402 , RIfc8ba48_6611, \9115 );
and \U$12272 ( \21403 , RIe16b210_2596, \9117 );
and \U$12273 ( \21404 , RIe1698c0_2578, \9119 );
and \U$12274 ( \21405 , RIe1679d0_2556, \9121 );
and \U$12275 ( \21406 , RIe164e38_2525, \9123 );
and \U$12276 ( \21407 , RIe162138_2493, \9125 );
and \U$12277 ( \21408 , RIee370f0_5085, \9127 );
and \U$12278 ( \21409 , RIe15f438_2461, \9129 );
and \U$12279 ( \21410 , RIfc999e0_6770, \9131 );
and \U$12280 ( \21411 , RIe15c738_2429, \9133 );
and \U$12281 ( \21412 , RIe156d38_2365, \9135 );
and \U$12282 ( \21413 , RIe154038_2333, \9137 );
and \U$12283 ( \21414 , RIfc3f260_5744, \9139 );
and \U$12284 ( \21415 , RIe151338_2301, \9141 );
and \U$12285 ( \21416 , RIfc48518_5845, \9143 );
and \U$12286 ( \21417 , RIe14e638_2269, \9145 );
and \U$12287 ( \21418 , RIfc99e18_6773, \9147 );
and \U$12288 ( \21419 , RIe14b938_2237, \9149 );
and \U$12289 ( \21420 , RIe148c38_2205, \9151 );
and \U$12290 ( \21421 , RIe145f38_2173, \9153 );
and \U$12291 ( \21422 , RIee34288_5052, \9155 );
and \U$12292 ( \21423 , RIee33040_5039, \9157 );
and \U$12293 ( \21424 , RIee31f60_5027, \9159 );
and \U$12294 ( \21425 , RIfcd99a0_7498, \9161 );
and \U$12295 ( \21426 , RIfe86b98_7877, \9163 );
and \U$12296 ( \21427 , RIdf3e9e0_2089, \9165 );
and \U$12297 ( \21428 , RIfe86a30_7876, \9167 );
and \U$12298 ( \21429 , RIdf3a4f8_2040, \9169 );
and \U$12299 ( \21430 , RIfcc3470_7244, \9171 );
and \U$12300 ( \21431 , RIee2f530_4997, \9173 );
and \U$12301 ( \21432 , RIfc7fdd8_6477, \9175 );
and \U$12302 ( \21433 , RIee2d370_4973, \9177 );
and \U$12303 ( \21434 , RIdf35200_1981, \9179 );
and \U$12304 ( \21435 , RIfec0ff0_8316, \9181 );
and \U$12305 ( \21436 , RIdf30d18_1932, \9183 );
and \U$12306 ( \21437 , RIfec0e88_8315, \9185 );
or \U$12307 ( \21438 , \21374 , \21375 , \21376 , \21377 , \21378 , \21379 , \21380 , \21381 , \21382 , \21383 , \21384 , \21385 , \21386 , \21387 , \21388 , \21389 , \21390 , \21391 , \21392 , \21393 , \21394 , \21395 , \21396 , \21397 , \21398 , \21399 , \21400 , \21401 , \21402 , \21403 , \21404 , \21405 , \21406 , \21407 , \21408 , \21409 , \21410 , \21411 , \21412 , \21413 , \21414 , \21415 , \21416 , \21417 , \21418 , \21419 , \21420 , \21421 , \21422 , \21423 , \21424 , \21425 , \21426 , \21427 , \21428 , \21429 , \21430 , \21431 , \21432 , \21433 , \21434 , \21435 , \21436 , \21437 );
and \U$12308 ( \21439 , RIfcd2a88_7419, \9188 );
and \U$12309 ( \21440 , RIfc8c858_6621, \9190 );
and \U$12310 ( \21441 , RIfc47ca8_5839, \9192 );
and \U$12311 ( \21442 , RIfcd6430_7460, \9194 );
and \U$12312 ( \21443 , RIdf29f68_1854, \9196 );
and \U$12313 ( \21444 , RIdf27da8_1830, \9198 );
and \U$12314 ( \21445 , RIdf26188_1810, \9200 );
and \U$12315 ( \21446 , RIdf24568_1790, \9202 );
and \U$12316 ( \21447 , RIfc8cb28_6623, \9204 );
and \U$12317 ( \21448 , RIfcdb188_7515, \9206 );
and \U$12318 ( \21449 , RIdf22948_1770, \9208 );
and \U$12319 ( \21450 , RIfc475a0_5834, \9210 );
and \U$12320 ( \21451 , RIdf21430_1755, \9212 );
and \U$12321 ( \21452 , RIdf1f3d8_1732, \9214 );
and \U$12322 ( \21453 , RIfec0bb8_8313, \9216 );
and \U$12323 ( \21454 , RIfe868c8_7875, \9218 );
and \U$12324 ( \21455 , RIdf16a08_1634, \9220 );
and \U$12325 ( \21456 , RIdf13d08_1602, \9222 );
and \U$12326 ( \21457 , RIdf11008_1570, \9224 );
and \U$12327 ( \21458 , RIdf0e308_1538, \9226 );
and \U$12328 ( \21459 , RIdf0b608_1506, \9228 );
and \U$12329 ( \21460 , RIdf08908_1474, \9230 );
and \U$12330 ( \21461 , RIdf05c08_1442, \9232 );
and \U$12331 ( \21462 , RIdf02f08_1410, \9234 );
and \U$12332 ( \21463 , RIdefd508_1346, \9236 );
and \U$12333 ( \21464 , RIdefa808_1314, \9238 );
and \U$12334 ( \21465 , RIdef7b08_1282, \9240 );
and \U$12335 ( \21466 , RIdef4e08_1250, \9242 );
and \U$12336 ( \21467 , RIdef2108_1218, \9244 );
and \U$12337 ( \21468 , RIdeef408_1186, \9246 );
and \U$12338 ( \21469 , RIdeec708_1154, \9248 );
and \U$12339 ( \21470 , RIdee9a08_1122, \9250 );
and \U$12340 ( \21471 , RIee254e0_4883, \9252 );
and \U$12341 ( \21472 , RIee246d0_4873, \9254 );
and \U$12342 ( \21473 , RIee23b90_4865, \9256 );
and \U$12343 ( \21474 , RIee231b8_4858, \9258 );
and \U$12344 ( \21475 , RIfe86fd0_7880, \9260 );
and \U$12345 ( \21476 , RIdee2820_1041, \9262 );
and \U$12346 ( \21477 , RIdee0930_1019, \9264 );
and \U$12347 ( \21478 , RIdede608_994, \9266 );
and \U$12348 ( \21479 , RIfc55da8_5999, \9268 );
and \U$12349 ( \21480 , RIfc98a68_6759, \9270 );
and \U$12350 ( \21481 , RIfcc3038_7241, \9272 );
and \U$12351 ( \21482 , RIfc464c0_5822, \9274 );
and \U$12352 ( \21483 , RIded9310_935, \9276 );
and \U$12353 ( \21484 , RIded6e80_909, \9278 );
and \U$12354 ( \21485 , RIded4f90_887, \9280 );
and \U$12355 ( \21486 , RIded2b00_861, \9282 );
and \U$12356 ( \21487 , RIded0238_832, \9284 );
and \U$12357 ( \21488 , RIdecd538_800, \9286 );
and \U$12358 ( \21489 , RIdeca838_768, \9288 );
and \U$12359 ( \21490 , RIdec7b38_736, \9290 );
and \U$12360 ( \21491 , RIdeb4038_512, \9292 );
and \U$12361 ( \21492 , RIde95c00_320, \9294 );
and \U$12362 ( \21493 , RIe16dc40_2626, \9296 );
and \U$12363 ( \21494 , RIe159a38_2397, \9298 );
and \U$12364 ( \21495 , RIe143238_2141, \9300 );
and \U$12365 ( \21496 , RIdf37c30_2011, \9302 );
and \U$12366 ( \21497 , RIdf2c290_1879, \9304 );
and \U$12367 ( \21498 , RIdf1cb10_1703, \9306 );
and \U$12368 ( \21499 , RIdf00208_1378, \9308 );
and \U$12369 ( \21500 , RIdee6d08_1090, \9310 );
and \U$12370 ( \21501 , RIdedba70_963, \9312 );
and \U$12371 ( \21502 , RIde7bb48_193, \9314 );
or \U$12372 ( \21503 , \21439 , \21440 , \21441 , \21442 , \21443 , \21444 , \21445 , \21446 , \21447 , \21448 , \21449 , \21450 , \21451 , \21452 , \21453 , \21454 , \21455 , \21456 , \21457 , \21458 , \21459 , \21460 , \21461 , \21462 , \21463 , \21464 , \21465 , \21466 , \21467 , \21468 , \21469 , \21470 , \21471 , \21472 , \21473 , \21474 , \21475 , \21476 , \21477 , \21478 , \21479 , \21480 , \21481 , \21482 , \21483 , \21484 , \21485 , \21486 , \21487 , \21488 , \21489 , \21490 , \21491 , \21492 , \21493 , \21494 , \21495 , \21496 , \21497 , \21498 , \21499 , \21500 , \21501 , \21502 );
or \U$12373 ( \21504 , \21438 , \21503 );
_DC g28f6 ( \21505_nG28f6 , \21504 , \9323 );
buf \U$12374 ( \21506 , \21505_nG28f6 );
and \U$12375 ( \21507 , RIe19d0d0_3164, \9333 );
and \U$12376 ( \21508 , RIe19a3d0_3132, \9335 );
and \U$12377 ( \21509 , RIf1454f0_5248, \9337 );
and \U$12378 ( \21510 , RIe1976d0_3100, \9339 );
and \U$12379 ( \21511 , RIf144578_5237, \9341 );
and \U$12380 ( \21512 , RIe1949d0_3068, \9343 );
and \U$12381 ( \21513 , RIe191cd0_3036, \9345 );
and \U$12382 ( \21514 , RIe18efd0_3004, \9347 );
and \U$12383 ( \21515 , RIe1895d0_2940, \9349 );
and \U$12384 ( \21516 , RIe1868d0_2908, \9351 );
and \U$12385 ( \21517 , RIf143498_5225, \9353 );
and \U$12386 ( \21518 , RIe183bd0_2876, \9355 );
and \U$12387 ( \21519 , RIfc51758_5949, \9357 );
and \U$12388 ( \21520 , RIe180ed0_2844, \9359 );
and \U$12389 ( \21521 , RIe17e1d0_2812, \9361 );
and \U$12390 ( \21522 , RIe17b4d0_2780, \9363 );
and \U$12391 ( \21523 , RIfc9b060_6786, \9365 );
and \U$12392 ( \21524 , RIfc9ee40_6830, \9367 );
and \U$12393 ( \21525 , RIe176e80_2730, \9369 );
and \U$12394 ( \21526 , RIe175800_2714, \9371 );
and \U$12395 ( \21527 , RIfcb70f8_7105, \9373 );
and \U$12396 ( \21528 , RIfce0cf0_7580, \9375 );
and \U$12397 ( \21529 , RIfcc4280_7254, \9377 );
and \U$12398 ( \21530 , RIfcba7d0_7144, \9379 );
and \U$12399 ( \21531 , RIee3bfb0_5141, \9381 );
and \U$12400 ( \21532 , RIee3aed0_5129, \9383 );
and \U$12401 ( \21533 , RIee39b20_5115, \9385 );
and \U$12402 ( \21534 , RIe173370_2688, \9387 );
and \U$12403 ( \21535 , RIf170060_5734, \9389 );
and \U$12404 ( \21536 , RIf16f3b8_5725, \9391 );
and \U$12405 ( \21537 , RIf16dea0_5710, \9393 );
and \U$12406 ( \21538 , RIf16d4c8_5703, \9395 );
and \U$12407 ( \21539 , RIf16c988_5695, \9397 );
and \U$12408 ( \21540 , RIe223428_4691, \9399 );
and \U$12409 ( \21541 , RIf16bb78_5685, \9401 );
and \U$12410 ( \21542 , RIe220728_4659, \9403 );
and \U$12411 ( \21543 , RIf16aa98_5673, \9405 );
and \U$12412 ( \21544 , RIe21da28_4627, \9407 );
and \U$12413 ( \21545 , RIe218028_4563, \9409 );
and \U$12414 ( \21546 , RIe215328_4531, \9411 );
and \U$12415 ( \21547 , RIf16a0c0_5666, \9413 );
and \U$12416 ( \21548 , RIe212628_4499, \9415 );
and \U$12417 ( \21549 , RIf168e78_5653, \9417 );
and \U$12418 ( \21550 , RIe20f928_4467, \9419 );
and \U$12419 ( \21551 , RIf167c30_5640, \9421 );
and \U$12420 ( \21552 , RIe20cc28_4435, \9423 );
and \U$12421 ( \21553 , RIe209f28_4403, \9425 );
and \U$12422 ( \21554 , RIe207228_4371, \9427 );
and \U$12423 ( \21555 , RIf166f88_5631, \9429 );
and \U$12424 ( \21556 , RIf165d40_5618, \9431 );
and \U$12425 ( \21557 , RIfec0618_8309, \9433 );
and \U$12426 ( \21558 , RIfe86760_7874, \9435 );
and \U$12427 ( \21559 , RIfc52b08_5963, \9437 );
and \U$12428 ( \21560 , RIf164288_5599, \9439 );
and \U$12429 ( \21561 , RIf163310_5588, \9441 );
and \U$12430 ( \21562 , RIf161c90_5572, \9443 );
and \U$12431 ( \21563 , RIf15fda0_5550, \9445 );
and \U$12432 ( \21564 , RIf15deb0_5528, \9447 );
and \U$12433 ( \21565 , RIfe865f8_7873, \9449 );
and \U$12434 ( \21566 , RIfe85d88_7867, \9451 );
and \U$12435 ( \21567 , RIf15c998_5513, \9453 );
and \U$12436 ( \21568 , RIf15b480_5498, \9455 );
and \U$12437 ( \21569 , RIf15a3a0_5486, \9457 );
and \U$12438 ( \21570 , RIf159b30_5480, \9459 );
or \U$12439 ( \21571 , \21507 , \21508 , \21509 , \21510 , \21511 , \21512 , \21513 , \21514 , \21515 , \21516 , \21517 , \21518 , \21519 , \21520 , \21521 , \21522 , \21523 , \21524 , \21525 , \21526 , \21527 , \21528 , \21529 , \21530 , \21531 , \21532 , \21533 , \21534 , \21535 , \21536 , \21537 , \21538 , \21539 , \21540 , \21541 , \21542 , \21543 , \21544 , \21545 , \21546 , \21547 , \21548 , \21549 , \21550 , \21551 , \21552 , \21553 , \21554 , \21555 , \21556 , \21557 , \21558 , \21559 , \21560 , \21561 , \21562 , \21563 , \21564 , \21565 , \21566 , \21567 , \21568 , \21569 , \21570 );
and \U$12440 ( \21572 , RIfc83348_6515, \9462 );
and \U$12441 ( \21573 , RIfc4ade0_5874, \9464 );
and \U$12442 ( \21574 , RIfc89720_6586, \9466 );
and \U$12443 ( \21575 , RIe1f9f38_4221, \9468 );
and \U$12444 ( \21576 , RIfc4ac78_5873, \9470 );
and \U$12445 ( \21577 , RIfc9f110_6832, \9472 );
and \U$12446 ( \21578 , RIfc4ab10_5872, \9474 );
and \U$12447 ( \21579 , RIe1f5078_4165, \9476 );
and \U$12448 ( \21580 , RIf152ee8_5403, \9478 );
and \U$12449 ( \21581 , RIfc899f0_6588, \9480 );
and \U$12450 ( \21582 , RIf150620_5374, \9482 );
and \U$12451 ( \21583 , RIe1f2eb8_4141, \9484 );
and \U$12452 ( \21584 , RIf14f6a8_5363, \9486 );
and \U$12453 ( \21585 , RIf14ea00_5354, \9488 );
and \U$12454 ( \21586 , RIf14dbf0_5344, \9490 );
and \U$12455 ( \21587 , RIe1edbc0_4082, \9492 );
and \U$12456 ( \21588 , RIe1eb190_4052, \9494 );
and \U$12457 ( \21589 , RIe1e8490_4020, \9496 );
and \U$12458 ( \21590 , RIe1e5790_3988, \9498 );
and \U$12459 ( \21591 , RIe1e2a90_3956, \9500 );
and \U$12460 ( \21592 , RIe1dfd90_3924, \9502 );
and \U$12461 ( \21593 , RIe1dd090_3892, \9504 );
and \U$12462 ( \21594 , RIe1da390_3860, \9506 );
and \U$12463 ( \21595 , RIe1d7690_3828, \9508 );
and \U$12464 ( \21596 , RIe1d1c90_3764, \9510 );
and \U$12465 ( \21597 , RIe1cef90_3732, \9512 );
and \U$12466 ( \21598 , RIe1cc290_3700, \9514 );
and \U$12467 ( \21599 , RIe1c9590_3668, \9516 );
and \U$12468 ( \21600 , RIe1c6890_3636, \9518 );
and \U$12469 ( \21601 , RIe1c3b90_3604, \9520 );
and \U$12470 ( \21602 , RIe1c0e90_3572, \9522 );
and \U$12471 ( \21603 , RIe1be190_3540, \9524 );
and \U$12472 ( \21604 , RIf14c6d8_5329, \9526 );
and \U$12473 ( \21605 , RIf14b490_5316, \9528 );
and \U$12474 ( \21606 , RIfe85ef0_7868, \9530 );
and \U$12475 ( \21607 , RIfe86490_7872, \9532 );
and \U$12476 ( \21608 , RIf14a248_5303, \9534 );
and \U$12477 ( \21609 , RIfc819f8_6497, \9536 );
and \U$12478 ( \21610 , RIfec0a50_8312, \9538 );
and \U$12479 ( \21611 , RIfe861c0_7870, \9540 );
and \U$12480 ( \21612 , RIf148bc8_5287, \9542 );
and \U$12481 ( \21613 , RIf147980_5274, \9544 );
and \U$12482 ( \21614 , RIfe86328_7871, \9546 );
and \U$12483 ( \21615 , RIfec0780_8310, \9548 );
and \U$12484 ( \21616 , RIfcbb478_7153, \9550 );
and \U$12485 ( \21617 , RIf146198_5257, \9552 );
and \U$12486 ( \21618 , RIfe86058_7869, \9554 );
and \U$12487 ( \21619 , RIfec08e8_8311, \9556 );
and \U$12488 ( \21620 , RIe1a84d0_3292, \9558 );
and \U$12489 ( \21621 , RIe1a57d0_3260, \9560 );
and \U$12490 ( \21622 , RIe1a2ad0_3228, \9562 );
and \U$12491 ( \21623 , RIe19fdd0_3196, \9564 );
and \U$12492 ( \21624 , RIe18c2d0_2972, \9566 );
and \U$12493 ( \21625 , RIe1787d0_2748, \9568 );
and \U$12494 ( \21626 , RIe226128_4723, \9570 );
and \U$12495 ( \21627 , RIe21ad28_4595, \9572 );
and \U$12496 ( \21628 , RIe204528_4339, \9574 );
and \U$12497 ( \21629 , RIe1fe588_4271, \9576 );
and \U$12498 ( \21630 , RIe1f7940_4194, \9578 );
and \U$12499 ( \21631 , RIe1f0488_4111, \9580 );
and \U$12500 ( \21632 , RIe1d4990_3796, \9582 );
and \U$12501 ( \21633 , RIe1bb490_3508, \9584 );
and \U$12502 ( \21634 , RIe1ae308_3359, \9586 );
and \U$12503 ( \21635 , RIe170940_2658, \9588 );
or \U$12504 ( \21636 , \21572 , \21573 , \21574 , \21575 , \21576 , \21577 , \21578 , \21579 , \21580 , \21581 , \21582 , \21583 , \21584 , \21585 , \21586 , \21587 , \21588 , \21589 , \21590 , \21591 , \21592 , \21593 , \21594 , \21595 , \21596 , \21597 , \21598 , \21599 , \21600 , \21601 , \21602 , \21603 , \21604 , \21605 , \21606 , \21607 , \21608 , \21609 , \21610 , \21611 , \21612 , \21613 , \21614 , \21615 , \21616 , \21617 , \21618 , \21619 , \21620 , \21621 , \21622 , \21623 , \21624 , \21625 , \21626 , \21627 , \21628 , \21629 , \21630 , \21631 , \21632 , \21633 , \21634 , \21635 );
or \U$12505 ( \21637 , \21571 , \21636 );
_DC g3a23 ( \21638_nG3a23 , \21637 , \9597 );
buf \U$12506 ( \21639 , \21638_nG3a23 );
and \U$12507 ( \21640 , \21506 , \21639 );
and \U$12508 ( \21641 , \19736 , \19869 );
and \U$12509 ( \21642 , \19869 , \20144 );
and \U$12510 ( \21643 , \19736 , \20144 );
or \U$12511 ( \21644 , \21641 , \21642 , \21643 );
and \U$12512 ( \21645 , \21639 , \21644 );
and \U$12513 ( \21646 , \21506 , \21644 );
or \U$12514 ( \21647 , \21640 , \21645 , \21646 );
xor \U$12515 ( \21648 , \21373 , \21647 );
buf g441e ( \21649_nG441e , \21648 );
xor \U$12516 ( \21650 , \21506 , \21639 );
xor \U$12517 ( \21651 , \21650 , \21644 );
buf g4421 ( \21652_nG4421 , \21651 );
nand \U$12518 ( \21653 , \21652_nG4421 , \20146_nG4424 );
and \U$12519 ( \21654 , \21649_nG441e , \21653 );
xor \U$12520 ( \21655 , \21652_nG4421 , \20146_nG4424 );
not \U$12521 ( \21656 , \21655 );
xor \U$12522 ( \21657 , \21649_nG441e , \21652_nG4421 );
and \U$12523 ( \21658 , \21656 , \21657 );
and \U$12525 ( \21659 , \21655 , \10694_nG9c0e );
or \U$12526 ( \21660 , 1'b0 , \21659 );
xor \U$12527 ( \21661 , \21654 , \21660 );
xor \U$12528 ( \21662 , \21654 , \21661 );
buf \U$12529 ( \21663 , \21662 );
buf \U$12530 ( \21664 , \21663 );
xor \U$12531 ( \21665 , \21106 , \21664 );
and \U$12532 ( \21666 , \20695 , \21093 );
and \U$12533 ( \21667 , \20695 , \21099 );
and \U$12534 ( \21668 , \21093 , \21099 );
or \U$12535 ( \21669 , \21666 , \21667 , \21668 );
and \U$12536 ( \21670 , \21665 , \21669 );
and \U$12537 ( \21671 , \20715 , \20721 );
and \U$12538 ( \21672 , \20715 , \21091 );
and \U$12539 ( \21673 , \20721 , \21091 );
or \U$12540 ( \21674 , \21671 , \21672 , \21673 );
buf \U$12541 ( \21675 , \21674 );
and \U$12542 ( \21676 , \20652 , \20658 );
and \U$12543 ( \21677 , \20652 , \20665 );
and \U$12544 ( \21678 , \20658 , \20665 );
or \U$12545 ( \21679 , \21676 , \21677 , \21678 );
buf \U$12546 ( \21680 , \21679 );
and \U$12547 ( \21681 , \15940 , \14070_nG9bf9 );
and \U$12548 ( \21682 , \15937 , \14984_nG9bf6 );
or \U$12549 ( \21683 , \21681 , \21682 );
xor \U$12550 ( \21684 , \15936 , \21683 );
buf \U$12551 ( \21685 , \21684 );
buf \U$12553 ( \21686 , \21685 );
xor \U$12554 ( \21687 , \21680 , \21686 );
and \U$12555 ( \21688 , \14631 , \15373_nG9bf3 );
and \U$12556 ( \21689 , \14628 , \16315_nG9bf0 );
or \U$12557 ( \21690 , \21688 , \21689 );
xor \U$12558 ( \21691 , \14627 , \21690 );
buf \U$12559 ( \21692 , \21691 );
buf \U$12561 ( \21693 , \21692 );
xor \U$12562 ( \21694 , \21687 , \21693 );
buf \U$12563 ( \21695 , \21694 );
and \U$12564 ( \21696 , \20667 , \20669 );
and \U$12565 ( \21697 , \20667 , \20676 );
and \U$12566 ( \21698 , \20669 , \20676 );
or \U$12567 ( \21699 , \21696 , \21697 , \21698 );
buf \U$12568 ( \21700 , \21699 );
xor \U$12569 ( \21701 , \21695 , \21700 );
and \U$12570 ( \21702 , \10421 , \19586_nG9be1 );
and \U$12571 ( \21703 , \10418 , \20608_nG9bde );
or \U$12572 ( \21704 , \21702 , \21703 );
xor \U$12573 ( \21705 , \10417 , \21704 );
buf \U$12574 ( \21706 , \21705 );
buf \U$12576 ( \21707 , \21706 );
xor \U$12577 ( \21708 , \21701 , \21707 );
buf \U$12578 ( \21709 , \21708 );
xor \U$12579 ( \21710 , \21675 , \21709 );
and \U$12580 ( \21711 , \20155 , \10995_nG9c0b );
and \U$12581 ( \21712 , \20152 , \11283_nG9c08 );
or \U$12582 ( \21713 , \21711 , \21712 );
xor \U$12583 ( \21714 , \20151 , \21713 );
buf \U$12584 ( \21715 , \21714 );
buf \U$12586 ( \21716 , \21715 );
and \U$12587 ( \21717 , \18702 , \11598_nG9c05 );
and \U$12588 ( \21718 , \18699 , \12470_nG9c02 );
or \U$12589 ( \21719 , \21717 , \21718 );
xor \U$12590 ( \21720 , \18698 , \21719 );
buf \U$12591 ( \21721 , \21720 );
buf \U$12593 ( \21722 , \21721 );
xor \U$12594 ( \21723 , \21716 , \21722 );
buf \U$12595 ( \21724 , \21723 );
and \U$12596 ( \21725 , \20644 , \20650 );
buf \U$12597 ( \21726 , \21725 );
xor \U$12598 ( \21727 , \21724 , \21726 );
and \U$12599 ( \21728 , \17297 , \12801_nG9bff );
and \U$12600 ( \21729 , \17294 , \13705_nG9bfc );
or \U$12601 ( \21730 , \21728 , \21729 );
xor \U$12602 ( \21731 , \17293 , \21730 );
buf \U$12603 ( \21732 , \21731 );
buf \U$12605 ( \21733 , \21732 );
xor \U$12606 ( \21734 , \21727 , \21733 );
buf \U$12607 ( \21735 , \21734 );
and \U$12608 ( \21736 , \13370 , \16680_nG9bed );
and \U$12609 ( \21737 , \13367 , \17665_nG9bea );
or \U$12610 ( \21738 , \21736 , \21737 );
xor \U$12611 ( \21739 , \13366 , \21738 );
buf \U$12612 ( \21740 , \21739 );
buf \U$12614 ( \21741 , \21740 );
xor \U$12615 ( \21742 , \21735 , \21741 );
and \U$12616 ( \21743 , \12157 , \18107_nG9be7 );
and \U$12617 ( \21744 , \12154 , \19091_nG9be4 );
or \U$12618 ( \21745 , \21743 , \21744 );
xor \U$12619 ( \21746 , \12153 , \21745 );
buf \U$12620 ( \21747 , \21746 );
buf \U$12622 ( \21748 , \21747 );
xor \U$12623 ( \21749 , \21742 , \21748 );
buf \U$12624 ( \21750 , \21749 );
xor \U$12625 ( \21751 , \21710 , \21750 );
buf \U$12626 ( \21752 , \21751 );
and \U$12627 ( \21753 , \20636 , \20687 );
and \U$12628 ( \21754 , \20636 , \20693 );
and \U$12629 ( \21755 , \20687 , \20693 );
or \U$12630 ( \21756 , \21753 , \21754 , \21755 );
buf \U$12631 ( \21757 , \21756 );
xor \U$12632 ( \21758 , \21752 , \21757 );
and \U$12633 ( \21759 , \20641 , \20678 );
and \U$12634 ( \21760 , \20641 , \20685 );
and \U$12635 ( \21761 , \20678 , \20685 );
or \U$12636 ( \21762 , \21759 , \21760 , \21761 );
buf \U$12637 ( \21763 , \21762 );
and \U$12638 ( \21764 , \20700 , \20706 );
and \U$12639 ( \21765 , \20700 , \20713 );
and \U$12640 ( \21766 , \20706 , \20713 );
or \U$12641 ( \21767 , \21764 , \21765 , \21766 );
buf \U$12642 ( \21768 , \21767 );
xor \U$12643 ( \21769 , \21763 , \21768 );
and \U$12644 ( \21770 , \10707 , \21086_nG9bdb );
and \U$12645 ( \21771 , \20727 , \21050 );
and \U$12646 ( \21772 , \21050 , \21075 );
and \U$12647 ( \21773 , \20727 , \21075 );
or \U$12648 ( \21774 , \21771 , \21772 , \21773 );
and \U$12649 ( \21775 , \21055 , \21059 );
and \U$12650 ( \21776 , \21059 , \21074 );
and \U$12651 ( \21777 , \21055 , \21074 );
or \U$12652 ( \21778 , \21775 , \21776 , \21777 );
and \U$12653 ( \21779 , \21039 , \21043 );
and \U$12654 ( \21780 , \21043 , \21048 );
and \U$12655 ( \21781 , \21039 , \21048 );
or \U$12656 ( \21782 , \21779 , \21780 , \21781 );
and \U$12657 ( \21783 , \19558 , \11574 );
and \U$12658 ( \21784 , \20544 , \11278 );
nor \U$12659 ( \21785 , \21783 , \21784 );
xnor \U$12660 ( \21786 , \21785 , \11580 );
and \U$12661 ( \21787 , \11586 , \19534 );
and \U$12662 ( \21788 , \12448 , \19045 );
nor \U$12663 ( \21789 , \21787 , \21788 );
xnor \U$12664 ( \21790 , \21789 , \19540 );
xor \U$12665 ( \21791 , \21786 , \21790 );
and \U$12666 ( \21792 , \10988 , \21005 );
and \U$12667 ( \21793 , \11270 , \20557 );
nor \U$12668 ( \21794 , \21792 , \21793 );
xnor \U$12669 ( \21795 , \21794 , \21011 );
xor \U$12670 ( \21796 , \21791 , \21795 );
xor \U$12671 ( \21797 , \21782 , \21796 );
and \U$12672 ( \21798 , \20731 , \20735 );
and \U$12673 ( \21799 , \20735 , \21012 );
and \U$12674 ( \21800 , \20731 , \21012 );
or \U$12675 ( \21801 , \21798 , \21799 , \21800 );
and \U$12676 ( \21802 , \21036 , \21038 );
xor \U$12677 ( \21803 , \21801 , \21802 );
and \U$12678 ( \21804 , \12769 , \18090 );
and \U$12679 ( \21805 , \13679 , \17655 );
nor \U$12680 ( \21806 , \21804 , \21805 );
xnor \U$12681 ( \21807 , \21806 , \18046 );
xor \U$12682 ( \21808 , \21803 , \21807 );
xor \U$12683 ( \21809 , \21797 , \21808 );
xor \U$12684 ( \21810 , \21778 , \21809 );
and \U$12685 ( \21811 , \21064 , \21068 );
and \U$12686 ( \21812 , \21068 , \21073 );
and \U$12687 ( \21813 , \21064 , \21073 );
or \U$12688 ( \21814 , \21811 , \21812 , \21813 );
and \U$12689 ( \21815 , \21013 , \21027 );
and \U$12690 ( \21816 , \21027 , \21049 );
and \U$12691 ( \21817 , \21013 , \21049 );
or \U$12692 ( \21818 , \21815 , \21816 , \21817 );
xor \U$12693 ( \21819 , \21814 , \21818 );
and \U$12694 ( \21820 , \21017 , \21021 );
and \U$12695 ( \21821 , \21021 , \21026 );
and \U$12696 ( \21822 , \21017 , \21026 );
or \U$12697 ( \21823 , \21820 , \21821 , \21822 );
and \U$12698 ( \21824 , \21033 , \10983 );
and \U$12699 ( \21825 , RIdec4e38_704, \9333 );
and \U$12700 ( \21826 , RIdec2138_672, \9335 );
and \U$12701 ( \21827 , RIee1fc48_4820, \9337 );
and \U$12702 ( \21828 , RIdebf438_640, \9339 );
and \U$12703 ( \21829 , RIfc49490_5856, \9341 );
and \U$12704 ( \21830 , RIdebc738_608, \9343 );
and \U$12705 ( \21831 , RIdeb9a38_576, \9345 );
and \U$12706 ( \21832 , RIdeb6d38_544, \9347 );
and \U$12707 ( \21833 , RIfc48ef0_5852, \9349 );
and \U$12708 ( \21834 , RIdeb1338_480, \9351 );
and \U$12709 ( \21835 , RIfcd9b08_7499, \9353 );
and \U$12710 ( \21836 , RIdeae638_448, \9355 );
and \U$12711 ( \21837 , RIfc8b610_6608, \9357 );
and \U$12712 ( \21838 , RIdea9700_416, \9359 );
and \U$12713 ( \21839 , RIdea2e00_384, \9361 );
and \U$12714 ( \21840 , RIde9c500_352, \9363 );
and \U$12715 ( \21841 , RIee1c9a8_4784, \9365 );
and \U$12716 ( \21842 , RIee1b8c8_4772, \9367 );
and \U$12717 ( \21843 , RIfc80918_6485, \9369 );
and \U$12718 ( \21844 , RIfcdad50_7512, \9371 );
and \U$12719 ( \21845 , RIfe86e68_7879, \9373 );
and \U$12720 ( \21846 , RIde8cee8_277, \9375 );
and \U$12721 ( \21847 , RIfe86d00_7878, \9377 );
and \U$12722 ( \21848 , RIfec0d20_8314, \9379 );
and \U$12723 ( \21849 , RIde81098_219, \9381 );
and \U$12724 ( \21850 , RIfc8b8e0_6610, \9383 );
and \U$12725 ( \21851 , RIfcd2d58_7421, \9385 );
and \U$12726 ( \21852 , RIfce4530_7620, \9387 );
and \U$12727 ( \21853 , RIfc8ba48_6611, \9389 );
and \U$12728 ( \21854 , RIe16b210_2596, \9391 );
and \U$12729 ( \21855 , RIe1698c0_2578, \9393 );
and \U$12730 ( \21856 , RIe1679d0_2556, \9395 );
and \U$12731 ( \21857 , RIe164e38_2525, \9397 );
and \U$12732 ( \21858 , RIe162138_2493, \9399 );
and \U$12733 ( \21859 , RIee370f0_5085, \9401 );
and \U$12734 ( \21860 , RIe15f438_2461, \9403 );
and \U$12735 ( \21861 , RIfc999e0_6770, \9405 );
and \U$12736 ( \21862 , RIe15c738_2429, \9407 );
and \U$12737 ( \21863 , RIe156d38_2365, \9409 );
and \U$12738 ( \21864 , RIe154038_2333, \9411 );
and \U$12739 ( \21865 , RIfc3f260_5744, \9413 );
and \U$12740 ( \21866 , RIe151338_2301, \9415 );
and \U$12741 ( \21867 , RIfc48518_5845, \9417 );
and \U$12742 ( \21868 , RIe14e638_2269, \9419 );
and \U$12743 ( \21869 , RIfc99e18_6773, \9421 );
and \U$12744 ( \21870 , RIe14b938_2237, \9423 );
and \U$12745 ( \21871 , RIe148c38_2205, \9425 );
and \U$12746 ( \21872 , RIe145f38_2173, \9427 );
and \U$12747 ( \21873 , RIee34288_5052, \9429 );
and \U$12748 ( \21874 , RIee33040_5039, \9431 );
and \U$12749 ( \21875 , RIee31f60_5027, \9433 );
and \U$12750 ( \21876 , RIfcd99a0_7498, \9435 );
and \U$12751 ( \21877 , RIfe86b98_7877, \9437 );
and \U$12752 ( \21878 , RIdf3e9e0_2089, \9439 );
and \U$12753 ( \21879 , RIfe86a30_7876, \9441 );
and \U$12754 ( \21880 , RIdf3a4f8_2040, \9443 );
and \U$12755 ( \21881 , RIfcc3470_7244, \9445 );
and \U$12756 ( \21882 , RIee2f530_4997, \9447 );
and \U$12757 ( \21883 , RIfc7fdd8_6477, \9449 );
and \U$12758 ( \21884 , RIee2d370_4973, \9451 );
and \U$12759 ( \21885 , RIdf35200_1981, \9453 );
and \U$12760 ( \21886 , RIfec0ff0_8316, \9455 );
and \U$12761 ( \21887 , RIdf30d18_1932, \9457 );
and \U$12762 ( \21888 , RIfec0e88_8315, \9459 );
or \U$12763 ( \21889 , \21825 , \21826 , \21827 , \21828 , \21829 , \21830 , \21831 , \21832 , \21833 , \21834 , \21835 , \21836 , \21837 , \21838 , \21839 , \21840 , \21841 , \21842 , \21843 , \21844 , \21845 , \21846 , \21847 , \21848 , \21849 , \21850 , \21851 , \21852 , \21853 , \21854 , \21855 , \21856 , \21857 , \21858 , \21859 , \21860 , \21861 , \21862 , \21863 , \21864 , \21865 , \21866 , \21867 , \21868 , \21869 , \21870 , \21871 , \21872 , \21873 , \21874 , \21875 , \21876 , \21877 , \21878 , \21879 , \21880 , \21881 , \21882 , \21883 , \21884 , \21885 , \21886 , \21887 , \21888 );
and \U$12764 ( \21890 , RIfcd2a88_7419, \9462 );
and \U$12765 ( \21891 , RIfc8c858_6621, \9464 );
and \U$12766 ( \21892 , RIfc47ca8_5839, \9466 );
and \U$12767 ( \21893 , RIfcd6430_7460, \9468 );
and \U$12768 ( \21894 , RIdf29f68_1854, \9470 );
and \U$12769 ( \21895 , RIdf27da8_1830, \9472 );
and \U$12770 ( \21896 , RIdf26188_1810, \9474 );
and \U$12771 ( \21897 , RIdf24568_1790, \9476 );
and \U$12772 ( \21898 , RIfc8cb28_6623, \9478 );
and \U$12773 ( \21899 , RIfcdb188_7515, \9480 );
and \U$12774 ( \21900 , RIdf22948_1770, \9482 );
and \U$12775 ( \21901 , RIfc475a0_5834, \9484 );
and \U$12776 ( \21902 , RIdf21430_1755, \9486 );
and \U$12777 ( \21903 , RIdf1f3d8_1732, \9488 );
and \U$12778 ( \21904 , RIfec0bb8_8313, \9490 );
and \U$12779 ( \21905 , RIfe868c8_7875, \9492 );
and \U$12780 ( \21906 , RIdf16a08_1634, \9494 );
and \U$12781 ( \21907 , RIdf13d08_1602, \9496 );
and \U$12782 ( \21908 , RIdf11008_1570, \9498 );
and \U$12783 ( \21909 , RIdf0e308_1538, \9500 );
and \U$12784 ( \21910 , RIdf0b608_1506, \9502 );
and \U$12785 ( \21911 , RIdf08908_1474, \9504 );
and \U$12786 ( \21912 , RIdf05c08_1442, \9506 );
and \U$12787 ( \21913 , RIdf02f08_1410, \9508 );
and \U$12788 ( \21914 , RIdefd508_1346, \9510 );
and \U$12789 ( \21915 , RIdefa808_1314, \9512 );
and \U$12790 ( \21916 , RIdef7b08_1282, \9514 );
and \U$12791 ( \21917 , RIdef4e08_1250, \9516 );
and \U$12792 ( \21918 , RIdef2108_1218, \9518 );
and \U$12793 ( \21919 , RIdeef408_1186, \9520 );
and \U$12794 ( \21920 , RIdeec708_1154, \9522 );
and \U$12795 ( \21921 , RIdee9a08_1122, \9524 );
and \U$12796 ( \21922 , RIee254e0_4883, \9526 );
and \U$12797 ( \21923 , RIee246d0_4873, \9528 );
and \U$12798 ( \21924 , RIee23b90_4865, \9530 );
and \U$12799 ( \21925 , RIee231b8_4858, \9532 );
and \U$12800 ( \21926 , RIfe86fd0_7880, \9534 );
and \U$12801 ( \21927 , RIdee2820_1041, \9536 );
and \U$12802 ( \21928 , RIdee0930_1019, \9538 );
and \U$12803 ( \21929 , RIdede608_994, \9540 );
and \U$12804 ( \21930 , RIfc55da8_5999, \9542 );
and \U$12805 ( \21931 , RIfc98a68_6759, \9544 );
and \U$12806 ( \21932 , RIfcc3038_7241, \9546 );
and \U$12807 ( \21933 , RIfc464c0_5822, \9548 );
and \U$12808 ( \21934 , RIded9310_935, \9550 );
and \U$12809 ( \21935 , RIded6e80_909, \9552 );
and \U$12810 ( \21936 , RIded4f90_887, \9554 );
and \U$12811 ( \21937 , RIded2b00_861, \9556 );
and \U$12812 ( \21938 , RIded0238_832, \9558 );
and \U$12813 ( \21939 , RIdecd538_800, \9560 );
and \U$12814 ( \21940 , RIdeca838_768, \9562 );
and \U$12815 ( \21941 , RIdec7b38_736, \9564 );
and \U$12816 ( \21942 , RIdeb4038_512, \9566 );
and \U$12817 ( \21943 , RIde95c00_320, \9568 );
and \U$12818 ( \21944 , RIe16dc40_2626, \9570 );
and \U$12819 ( \21945 , RIe159a38_2397, \9572 );
and \U$12820 ( \21946 , RIe143238_2141, \9574 );
and \U$12821 ( \21947 , RIdf37c30_2011, \9576 );
and \U$12822 ( \21948 , RIdf2c290_1879, \9578 );
and \U$12823 ( \21949 , RIdf1cb10_1703, \9580 );
and \U$12824 ( \21950 , RIdf00208_1378, \9582 );
and \U$12825 ( \21951 , RIdee6d08_1090, \9584 );
and \U$12826 ( \21952 , RIdedba70_963, \9586 );
and \U$12827 ( \21953 , RIde7bb48_193, \9588 );
or \U$12828 ( \21954 , \21890 , \21891 , \21892 , \21893 , \21894 , \21895 , \21896 , \21897 , \21898 , \21899 , \21900 , \21901 , \21902 , \21903 , \21904 , \21905 , \21906 , \21907 , \21908 , \21909 , \21910 , \21911 , \21912 , \21913 , \21914 , \21915 , \21916 , \21917 , \21918 , \21919 , \21920 , \21921 , \21922 , \21923 , \21924 , \21925 , \21926 , \21927 , \21928 , \21929 , \21930 , \21931 , \21932 , \21933 , \21934 , \21935 , \21936 , \21937 , \21938 , \21939 , \21940 , \21941 , \21942 , \21943 , \21944 , \21945 , \21946 , \21947 , \21948 , \21949 , \21950 , \21951 , \21952 , \21953 );
or \U$12829 ( \21955 , \21889 , \21954 );
_DC g65ad ( \21956_nG65ad , \21955 , \9597 );
and \U$12830 ( \21957 , RIe19d0d0_3164, \9059 );
and \U$12831 ( \21958 , RIe19a3d0_3132, \9061 );
and \U$12832 ( \21959 , RIf1454f0_5248, \9063 );
and \U$12833 ( \21960 , RIe1976d0_3100, \9065 );
and \U$12834 ( \21961 , RIf144578_5237, \9067 );
and \U$12835 ( \21962 , RIe1949d0_3068, \9069 );
and \U$12836 ( \21963 , RIe191cd0_3036, \9071 );
and \U$12837 ( \21964 , RIe18efd0_3004, \9073 );
and \U$12838 ( \21965 , RIe1895d0_2940, \9075 );
and \U$12839 ( \21966 , RIe1868d0_2908, \9077 );
and \U$12840 ( \21967 , RIf143498_5225, \9079 );
and \U$12841 ( \21968 , RIe183bd0_2876, \9081 );
and \U$12842 ( \21969 , RIfc51758_5949, \9083 );
and \U$12843 ( \21970 , RIe180ed0_2844, \9085 );
and \U$12844 ( \21971 , RIe17e1d0_2812, \9087 );
and \U$12845 ( \21972 , RIe17b4d0_2780, \9089 );
and \U$12846 ( \21973 , RIfc9b060_6786, \9091 );
and \U$12847 ( \21974 , RIfc9ee40_6830, \9093 );
and \U$12848 ( \21975 , RIe176e80_2730, \9095 );
and \U$12849 ( \21976 , RIe175800_2714, \9097 );
and \U$12850 ( \21977 , RIfcb70f8_7105, \9099 );
and \U$12851 ( \21978 , RIfce0cf0_7580, \9101 );
and \U$12852 ( \21979 , RIfcc4280_7254, \9103 );
and \U$12853 ( \21980 , RIfcba7d0_7144, \9105 );
and \U$12854 ( \21981 , RIee3bfb0_5141, \9107 );
and \U$12855 ( \21982 , RIee3aed0_5129, \9109 );
and \U$12856 ( \21983 , RIee39b20_5115, \9111 );
and \U$12857 ( \21984 , RIe173370_2688, \9113 );
and \U$12858 ( \21985 , RIf170060_5734, \9115 );
and \U$12859 ( \21986 , RIf16f3b8_5725, \9117 );
and \U$12860 ( \21987 , RIf16dea0_5710, \9119 );
and \U$12861 ( \21988 , RIf16d4c8_5703, \9121 );
and \U$12862 ( \21989 , RIf16c988_5695, \9123 );
and \U$12863 ( \21990 , RIe223428_4691, \9125 );
and \U$12864 ( \21991 , RIf16bb78_5685, \9127 );
and \U$12865 ( \21992 , RIe220728_4659, \9129 );
and \U$12866 ( \21993 , RIf16aa98_5673, \9131 );
and \U$12867 ( \21994 , RIe21da28_4627, \9133 );
and \U$12868 ( \21995 , RIe218028_4563, \9135 );
and \U$12869 ( \21996 , RIe215328_4531, \9137 );
and \U$12870 ( \21997 , RIf16a0c0_5666, \9139 );
and \U$12871 ( \21998 , RIe212628_4499, \9141 );
and \U$12872 ( \21999 , RIf168e78_5653, \9143 );
and \U$12873 ( \22000 , RIe20f928_4467, \9145 );
and \U$12874 ( \22001 , RIf167c30_5640, \9147 );
and \U$12875 ( \22002 , RIe20cc28_4435, \9149 );
and \U$12876 ( \22003 , RIe209f28_4403, \9151 );
and \U$12877 ( \22004 , RIe207228_4371, \9153 );
and \U$12878 ( \22005 , RIf166f88_5631, \9155 );
and \U$12879 ( \22006 , RIf165d40_5618, \9157 );
and \U$12880 ( \22007 , RIfec0618_8309, \9159 );
and \U$12881 ( \22008 , RIfe86760_7874, \9161 );
and \U$12882 ( \22009 , RIfc52b08_5963, \9163 );
and \U$12883 ( \22010 , RIf164288_5599, \9165 );
and \U$12884 ( \22011 , RIf163310_5588, \9167 );
and \U$12885 ( \22012 , RIf161c90_5572, \9169 );
and \U$12886 ( \22013 , RIf15fda0_5550, \9171 );
and \U$12887 ( \22014 , RIf15deb0_5528, \9173 );
and \U$12888 ( \22015 , RIfe865f8_7873, \9175 );
and \U$12889 ( \22016 , RIfe85d88_7867, \9177 );
and \U$12890 ( \22017 , RIf15c998_5513, \9179 );
and \U$12891 ( \22018 , RIf15b480_5498, \9181 );
and \U$12892 ( \22019 , RIf15a3a0_5486, \9183 );
and \U$12893 ( \22020 , RIf159b30_5480, \9185 );
or \U$12894 ( \22021 , \21957 , \21958 , \21959 , \21960 , \21961 , \21962 , \21963 , \21964 , \21965 , \21966 , \21967 , \21968 , \21969 , \21970 , \21971 , \21972 , \21973 , \21974 , \21975 , \21976 , \21977 , \21978 , \21979 , \21980 , \21981 , \21982 , \21983 , \21984 , \21985 , \21986 , \21987 , \21988 , \21989 , \21990 , \21991 , \21992 , \21993 , \21994 , \21995 , \21996 , \21997 , \21998 , \21999 , \22000 , \22001 , \22002 , \22003 , \22004 , \22005 , \22006 , \22007 , \22008 , \22009 , \22010 , \22011 , \22012 , \22013 , \22014 , \22015 , \22016 , \22017 , \22018 , \22019 , \22020 );
and \U$12895 ( \22022 , RIfc83348_6515, \9188 );
and \U$12896 ( \22023 , RIfc4ade0_5874, \9190 );
and \U$12897 ( \22024 , RIfc89720_6586, \9192 );
and \U$12898 ( \22025 , RIe1f9f38_4221, \9194 );
and \U$12899 ( \22026 , RIfc4ac78_5873, \9196 );
and \U$12900 ( \22027 , RIfc9f110_6832, \9198 );
and \U$12901 ( \22028 , RIfc4ab10_5872, \9200 );
and \U$12902 ( \22029 , RIe1f5078_4165, \9202 );
and \U$12903 ( \22030 , RIf152ee8_5403, \9204 );
and \U$12904 ( \22031 , RIfc899f0_6588, \9206 );
and \U$12905 ( \22032 , RIf150620_5374, \9208 );
and \U$12906 ( \22033 , RIe1f2eb8_4141, \9210 );
and \U$12907 ( \22034 , RIf14f6a8_5363, \9212 );
and \U$12908 ( \22035 , RIf14ea00_5354, \9214 );
and \U$12909 ( \22036 , RIf14dbf0_5344, \9216 );
and \U$12910 ( \22037 , RIe1edbc0_4082, \9218 );
and \U$12911 ( \22038 , RIe1eb190_4052, \9220 );
and \U$12912 ( \22039 , RIe1e8490_4020, \9222 );
and \U$12913 ( \22040 , RIe1e5790_3988, \9224 );
and \U$12914 ( \22041 , RIe1e2a90_3956, \9226 );
and \U$12915 ( \22042 , RIe1dfd90_3924, \9228 );
and \U$12916 ( \22043 , RIe1dd090_3892, \9230 );
and \U$12917 ( \22044 , RIe1da390_3860, \9232 );
and \U$12918 ( \22045 , RIe1d7690_3828, \9234 );
and \U$12919 ( \22046 , RIe1d1c90_3764, \9236 );
and \U$12920 ( \22047 , RIe1cef90_3732, \9238 );
and \U$12921 ( \22048 , RIe1cc290_3700, \9240 );
and \U$12922 ( \22049 , RIe1c9590_3668, \9242 );
and \U$12923 ( \22050 , RIe1c6890_3636, \9244 );
and \U$12924 ( \22051 , RIe1c3b90_3604, \9246 );
and \U$12925 ( \22052 , RIe1c0e90_3572, \9248 );
and \U$12926 ( \22053 , RIe1be190_3540, \9250 );
and \U$12927 ( \22054 , RIf14c6d8_5329, \9252 );
and \U$12928 ( \22055 , RIf14b490_5316, \9254 );
and \U$12929 ( \22056 , RIfe85ef0_7868, \9256 );
and \U$12930 ( \22057 , RIfe86490_7872, \9258 );
and \U$12931 ( \22058 , RIf14a248_5303, \9260 );
and \U$12932 ( \22059 , RIfc819f8_6497, \9262 );
and \U$12933 ( \22060 , RIfec0a50_8312, \9264 );
and \U$12934 ( \22061 , RIfe861c0_7870, \9266 );
and \U$12935 ( \22062 , RIf148bc8_5287, \9268 );
and \U$12936 ( \22063 , RIf147980_5274, \9270 );
and \U$12937 ( \22064 , RIfe86328_7871, \9272 );
and \U$12938 ( \22065 , RIfec0780_8310, \9274 );
and \U$12939 ( \22066 , RIfcbb478_7153, \9276 );
and \U$12940 ( \22067 , RIf146198_5257, \9278 );
and \U$12941 ( \22068 , RIfe86058_7869, \9280 );
and \U$12942 ( \22069 , RIfec08e8_8311, \9282 );
and \U$12943 ( \22070 , RIe1a84d0_3292, \9284 );
and \U$12944 ( \22071 , RIe1a57d0_3260, \9286 );
and \U$12945 ( \22072 , RIe1a2ad0_3228, \9288 );
and \U$12946 ( \22073 , RIe19fdd0_3196, \9290 );
and \U$12947 ( \22074 , RIe18c2d0_2972, \9292 );
and \U$12948 ( \22075 , RIe1787d0_2748, \9294 );
and \U$12949 ( \22076 , RIe226128_4723, \9296 );
and \U$12950 ( \22077 , RIe21ad28_4595, \9298 );
and \U$12951 ( \22078 , RIe204528_4339, \9300 );
and \U$12952 ( \22079 , RIe1fe588_4271, \9302 );
and \U$12953 ( \22080 , RIe1f7940_4194, \9304 );
and \U$12954 ( \22081 , RIe1f0488_4111, \9306 );
and \U$12955 ( \22082 , RIe1d4990_3796, \9308 );
and \U$12956 ( \22083 , RIe1bb490_3508, \9310 );
and \U$12957 ( \22084 , RIe1ae308_3359, \9312 );
and \U$12958 ( \22085 , RIe170940_2658, \9314 );
or \U$12959 ( \22086 , \22022 , \22023 , \22024 , \22025 , \22026 , \22027 , \22028 , \22029 , \22030 , \22031 , \22032 , \22033 , \22034 , \22035 , \22036 , \22037 , \22038 , \22039 , \22040 , \22041 , \22042 , \22043 , \22044 , \22045 , \22046 , \22047 , \22048 , \22049 , \22050 , \22051 , \22052 , \22053 , \22054 , \22055 , \22056 , \22057 , \22058 , \22059 , \22060 , \22061 , \22062 , \22063 , \22064 , \22065 , \22066 , \22067 , \22068 , \22069 , \22070 , \22071 , \22072 , \22073 , \22074 , \22075 , \22076 , \22077 , \22078 , \22079 , \22080 , \22081 , \22082 , \22083 , \22084 , \22085 );
or \U$12960 ( \22087 , \22021 , \22086 );
_DC g65ae ( \22088_nG65ae , \22087 , \9323 );
and g65af ( \22089_nG65af , \21956_nG65ad , \22088_nG65ae );
buf \U$12961 ( \22090 , \22089_nG65af );
and \U$12962 ( \22091 , \22090 , \10691 );
nor \U$12963 ( \22092 , \21824 , \22091 );
xnor \U$12964 ( \22093 , \22092 , \10980 );
and \U$12965 ( \22094 , \16655 , \14054 );
and \U$12966 ( \22095 , \17627 , \13692 );
nor \U$12967 ( \22096 , \22094 , \22095 );
xnor \U$12968 ( \22097 , \22096 , \14035 );
xor \U$12969 ( \22098 , \22093 , \22097 );
_DC g577c ( \22099_nG577c , \21955 , \9597 );
_DC g5800 ( \22100_nG5800 , \22087 , \9323 );
xor g5801 ( \22101_nG5801 , \22099_nG577c , \22100_nG5800 );
buf \U$12970 ( \22102 , \22101_nG5801 );
xor \U$12971 ( \22103 , \22102 , \21002 );
and \U$12972 ( \22104 , \10687 , \22103 );
xor \U$12973 ( \22105 , \22098 , \22104 );
xor \U$12974 ( \22106 , \21823 , \22105 );
and \U$12975 ( \22107 , \18035 , \12790 );
and \U$12976 ( \22108 , \19032 , \12461 );
nor \U$12977 ( \22109 , \22107 , \22108 );
xnor \U$12978 ( \22110 , \22109 , \12780 );
and \U$12979 ( \22111 , \15321 , \15336 );
and \U$12980 ( \22112 , \16267 , \14963 );
nor \U$12981 ( \22113 , \22111 , \22112 );
xnor \U$12982 ( \22114 , \22113 , \15342 );
xor \U$12983 ( \22115 , \22110 , \22114 );
and \U$12984 ( \22116 , \14024 , \16635 );
and \U$12985 ( \22117 , \14950 , \16301 );
nor \U$12986 ( \22118 , \22116 , \22117 );
xnor \U$12987 ( \22119 , \22118 , \16625 );
xor \U$12988 ( \22120 , \22115 , \22119 );
xor \U$12989 ( \22121 , \22106 , \22120 );
xor \U$12990 ( \22122 , \21819 , \22121 );
xor \U$12991 ( \22123 , \21810 , \22122 );
xor \U$12992 ( \22124 , \21774 , \22123 );
and \U$12993 ( \22125 , \21076 , \21080 );
and \U$12994 ( \22126 , \21081 , \21084 );
or \U$12995 ( \22127 , \22125 , \22126 );
xor \U$12996 ( \22128 , \22124 , \22127 );
buf g9bd8 ( \22129_nG9bd8 , \22128 );
and \U$12997 ( \22130 , \10704 , \22129_nG9bd8 );
or \U$12998 ( \22131 , \21770 , \22130 );
xor \U$12999 ( \22132 , \10703 , \22131 );
buf \U$13000 ( \22133 , \22132 );
buf \U$13002 ( \22134 , \22133 );
xor \U$13003 ( \22135 , \21769 , \22134 );
buf \U$13004 ( \22136 , \22135 );
xor \U$13005 ( \22137 , \21758 , \22136 );
and \U$13006 ( \22138 , \21665 , \22137 );
and \U$13007 ( \22139 , \21669 , \22137 );
or \U$13008 ( \22140 , \21670 , \22138 , \22139 );
and \U$13009 ( \22141 , \21101 , \21105 );
and \U$13010 ( \22142 , \21101 , \21664 );
and \U$13011 ( \22143 , \21105 , \21664 );
or \U$13012 ( \22144 , \22141 , \22142 , \22143 );
xor \U$13013 ( \22145 , \22140 , \22144 );
and \U$13014 ( \22146 , \21752 , \21757 );
and \U$13015 ( \22147 , \21752 , \22136 );
and \U$13016 ( \22148 , \21757 , \22136 );
or \U$13017 ( \22149 , \22146 , \22147 , \22148 );
xor \U$13018 ( \22150 , \22145 , \22149 );
and \U$13019 ( \22151 , \21763 , \21768 );
and \U$13020 ( \22152 , \21763 , \22134 );
and \U$13021 ( \22153 , \21768 , \22134 );
or \U$13022 ( \22154 , \22151 , \22152 , \22153 );
buf \U$13023 ( \22155 , \22154 );
and \U$13024 ( \22156 , \21724 , \21726 );
and \U$13025 ( \22157 , \21724 , \21733 );
and \U$13026 ( \22158 , \21726 , \21733 );
or \U$13027 ( \22159 , \22156 , \22157 , \22158 );
buf \U$13028 ( \22160 , \22159 );
and \U$13029 ( \22161 , \15940 , \14984_nG9bf6 );
and \U$13030 ( \22162 , \15937 , \15373_nG9bf3 );
or \U$13031 ( \22163 , \22161 , \22162 );
xor \U$13032 ( \22164 , \15936 , \22163 );
buf \U$13033 ( \22165 , \22164 );
buf \U$13035 ( \22166 , \22165 );
xor \U$13036 ( \22167 , \22160 , \22166 );
and \U$13037 ( \22168 , \14631 , \16315_nG9bf0 );
and \U$13038 ( \22169 , \14628 , \16680_nG9bed );
or \U$13039 ( \22170 , \22168 , \22169 );
xor \U$13040 ( \22171 , \14627 , \22170 );
buf \U$13041 ( \22172 , \22171 );
buf \U$13043 ( \22173 , \22172 );
xor \U$13044 ( \22174 , \22167 , \22173 );
buf \U$13045 ( \22175 , \22174 );
and \U$13046 ( \22176 , \12157 , \19091_nG9be4 );
and \U$13047 ( \22177 , \12154 , \19586_nG9be1 );
or \U$13048 ( \22178 , \22176 , \22177 );
xor \U$13049 ( \22179 , \12153 , \22178 );
buf \U$13050 ( \22180 , \22179 );
buf \U$13052 ( \22181 , \22180 );
xor \U$13053 ( \22182 , \22175 , \22181 );
and \U$13054 ( \22183 , \10421 , \20608_nG9bde );
and \U$13055 ( \22184 , \10418 , \21086_nG9bdb );
or \U$13056 ( \22185 , \22183 , \22184 );
xor \U$13057 ( \22186 , \10417 , \22185 );
buf \U$13058 ( \22187 , \22186 );
buf \U$13060 ( \22188 , \22187 );
xor \U$13061 ( \22189 , \22182 , \22188 );
buf \U$13062 ( \22190 , \22189 );
xor \U$13063 ( \22191 , \22155 , \22190 );
and \U$13064 ( \22192 , \21680 , \21686 );
and \U$13065 ( \22193 , \21680 , \21693 );
and \U$13066 ( \22194 , \21686 , \21693 );
or \U$13067 ( \22195 , \22192 , \22193 , \22194 );
buf \U$13068 ( \22196 , \22195 );
and \U$13069 ( \22197 , \21654 , \21661 );
buf \U$13070 ( \22198 , \22197 );
buf \U$13072 ( \22199 , \22198 );
and \U$13073 ( \22200 , \20155 , \11283_nG9c08 );
and \U$13074 ( \22201 , \20152 , \11598_nG9c05 );
or \U$13075 ( \22202 , \22200 , \22201 );
xor \U$13076 ( \22203 , \20151 , \22202 );
buf \U$13077 ( \22204 , \22203 );
buf \U$13079 ( \22205 , \22204 );
xor \U$13080 ( \22206 , \22199 , \22205 );
buf \U$13081 ( \22207 , \22206 );
and \U$13082 ( \22208 , \21658 , \10694_nG9c0e );
and \U$13083 ( \22209 , \21655 , \10995_nG9c0b );
or \U$13084 ( \22210 , \22208 , \22209 );
xor \U$13085 ( \22211 , \21654 , \22210 );
buf \U$13086 ( \22212 , \22211 );
buf \U$13088 ( \22213 , \22212 );
xor \U$13089 ( \22214 , \22207 , \22213 );
and \U$13090 ( \22215 , \18702 , \12470_nG9c02 );
and \U$13091 ( \22216 , \18699 , \12801_nG9bff );
or \U$13092 ( \22217 , \22215 , \22216 );
xor \U$13093 ( \22218 , \18698 , \22217 );
buf \U$13094 ( \22219 , \22218 );
buf \U$13096 ( \22220 , \22219 );
xor \U$13097 ( \22221 , \22214 , \22220 );
buf \U$13098 ( \22222 , \22221 );
and \U$13099 ( \22223 , \21716 , \21722 );
buf \U$13100 ( \22224 , \22223 );
xor \U$13101 ( \22225 , \22222 , \22224 );
and \U$13102 ( \22226 , \17297 , \13705_nG9bfc );
and \U$13103 ( \22227 , \17294 , \14070_nG9bf9 );
or \U$13104 ( \22228 , \22226 , \22227 );
xor \U$13105 ( \22229 , \17293 , \22228 );
buf \U$13106 ( \22230 , \22229 );
buf \U$13108 ( \22231 , \22230 );
xor \U$13109 ( \22232 , \22225 , \22231 );
buf \U$13110 ( \22233 , \22232 );
xor \U$13111 ( \22234 , \22196 , \22233 );
and \U$13112 ( \22235 , \13370 , \17665_nG9bea );
and \U$13113 ( \22236 , \13367 , \18107_nG9be7 );
or \U$13114 ( \22237 , \22235 , \22236 );
xor \U$13115 ( \22238 , \13366 , \22237 );
buf \U$13116 ( \22239 , \22238 );
buf \U$13118 ( \22240 , \22239 );
xor \U$13119 ( \22241 , \22234 , \22240 );
buf \U$13120 ( \22242 , \22241 );
xor \U$13121 ( \22243 , \22191 , \22242 );
buf \U$13122 ( \22244 , \22243 );
and \U$13123 ( \22245 , \21695 , \21700 );
and \U$13124 ( \22246 , \21695 , \21707 );
and \U$13125 ( \22247 , \21700 , \21707 );
or \U$13126 ( \22248 , \22245 , \22246 , \22247 );
buf \U$13127 ( \22249 , \22248 );
and \U$13128 ( \22250 , \21735 , \21741 );
and \U$13129 ( \22251 , \21735 , \21748 );
and \U$13130 ( \22252 , \21741 , \21748 );
or \U$13131 ( \22253 , \22250 , \22251 , \22252 );
buf \U$13132 ( \22254 , \22253 );
xor \U$13133 ( \22255 , \22249 , \22254 );
and \U$13134 ( \22256 , \10707 , \22129_nG9bd8 );
and \U$13135 ( \22257 , \21814 , \21818 );
and \U$13136 ( \22258 , \21818 , \22121 );
and \U$13137 ( \22259 , \21814 , \22121 );
or \U$13138 ( \22260 , \22257 , \22258 , \22259 );
and \U$13139 ( \22261 , \21801 , \21802 );
and \U$13140 ( \22262 , \21802 , \21807 );
and \U$13141 ( \22263 , \21801 , \21807 );
or \U$13142 ( \22264 , \22261 , \22262 , \22263 );
and \U$13143 ( \22265 , \20544 , \11574 );
and \U$13144 ( \22266 , \21033 , \11278 );
nor \U$13145 ( \22267 , \22265 , \22266 );
xnor \U$13146 ( \22268 , \22267 , \11580 );
and \U$13147 ( \22269 , \16267 , \15336 );
and \U$13148 ( \22270 , \16655 , \14963 );
nor \U$13149 ( \22271 , \22269 , \22270 );
xnor \U$13150 ( \22272 , \22271 , \15342 );
xor \U$13151 ( \22273 , \22268 , \22272 );
and \U$13152 ( \22274 , RIdec4fa0_705, \9333 );
and \U$13153 ( \22275 , RIdec22a0_673, \9335 );
and \U$13154 ( \22276 , RIee1fdb0_4821, \9337 );
and \U$13155 ( \22277 , RIdebf5a0_641, \9339 );
and \U$13156 ( \22278 , RIee1f270_4813, \9341 );
and \U$13157 ( \22279 , RIdebc8a0_609, \9343 );
and \U$13158 ( \22280 , RIdeb9ba0_577, \9345 );
and \U$13159 ( \22281 , RIdeb6ea0_545, \9347 );
and \U$13160 ( \22282 , RIee1ecd0_4809, \9349 );
and \U$13161 ( \22283 , RIdeb14a0_481, \9351 );
and \U$13162 ( \22284 , RIee1e730_4805, \9353 );
and \U$13163 ( \22285 , RIdeae7a0_449, \9355 );
and \U$13164 ( \22286 , RIee1d920_4795, \9357 );
and \U$13165 ( \22287 , RIdea9a48_417, \9359 );
and \U$13166 ( \22288 , RIdea3148_385, \9361 );
and \U$13167 ( \22289 , RIde9c848_353, \9363 );
and \U$13168 ( \22290 , RIee1cb10_4785, \9365 );
and \U$13169 ( \22291 , RIee1ba30_4773, \9367 );
and \U$13170 ( \22292 , RIee1b1c0_4767, \9369 );
and \U$13171 ( \22293 , RIfec04b0_8308, \9371 );
and \U$13172 ( \22294 , RIfe850e0_7858, \9373 );
and \U$13173 ( \22295 , RIde8d230_278, \9375 );
and \U$13174 ( \22296 , RIfea9cb0_8248, \9377 );
and \U$13175 ( \22297 , RIfe84f78_7857, \9379 );
and \U$13176 ( \22298 , RIee1a3b0_4757, \9381 );
and \U$13177 ( \22299 , RIfe853b0_7860, \9383 );
and \U$13178 ( \22300 , RIee199d8_4750, \9385 );
and \U$13179 ( \22301 , RIfe85248_7859, \9387 );
and \U$13180 ( \22302 , RIee39148_5108, \9389 );
and \U$13181 ( \22303 , RIe16b378_2597, \9391 );
and \U$13182 ( \22304 , RIee38608_5100, \9393 );
and \U$13183 ( \22305 , RIe167b38_2557, \9395 );
and \U$13184 ( \22306 , RIe164fa0_2526, \9397 );
and \U$13185 ( \22307 , RIe1622a0_2494, \9399 );
and \U$13186 ( \22308 , RIfe85950_7864, \9401 );
and \U$13187 ( \22309 , RIe15f5a0_2462, \9403 );
and \U$13188 ( \22310 , RIee36010_5073, \9405 );
and \U$13189 ( \22311 , RIe15c8a0_2430, \9407 );
and \U$13190 ( \22312 , RIe156ea0_2366, \9409 );
and \U$13191 ( \22313 , RIe1541a0_2334, \9411 );
and \U$13192 ( \22314 , RIfe85c20_7866, \9413 );
and \U$13193 ( \22315 , RIe1514a0_2302, \9415 );
and \U$13194 ( \22316 , RIee34dc8_5060, \9417 );
and \U$13195 ( \22317 , RIe14e7a0_2270, \9419 );
and \U$13196 ( \22318 , RIfc861b0_6548, \9421 );
and \U$13197 ( \22319 , RIe14baa0_2238, \9423 );
and \U$13198 ( \22320 , RIe148da0_2206, \9425 );
and \U$13199 ( \22321 , RIe1460a0_2174, \9427 );
and \U$13200 ( \22322 , RIee343f0_5053, \9429 );
and \U$13201 ( \22323 , RIfe85518_7861, \9431 );
and \U$13202 ( \22324 , RIfe857e8_7863, \9433 );
and \U$13203 ( \22325 , RIfe85680_7862, \9435 );
and \U$13204 ( \22326 , RIe140c40_2114, \9437 );
and \U$13205 ( \22327 , RIdf3eb48_2090, \9439 );
and \U$13206 ( \22328 , RIdf3c820_2065, \9441 );
and \U$13207 ( \22329 , RIdf3a660_2041, \9443 );
and \U$13208 ( \22330 , RIfc9d4f0_6812, \9445 );
and \U$13209 ( \22331 , RIee2f698_4998, \9447 );
and \U$13210 ( \22332 , RIfc52298_5957, \9449 );
and \U$13211 ( \22333 , RIee2d4d8_4974, \9451 );
and \U$13212 ( \22334 , RIdf35368_1982, \9453 );
and \U$13213 ( \22335 , RIdf32ed8_1956, \9455 );
and \U$13214 ( \22336 , RIdf30e80_1933, \9457 );
and \U$13215 ( \22337 , RIfe85ab8_7865, \9459 );
or \U$13216 ( \22338 , \22274 , \22275 , \22276 , \22277 , \22278 , \22279 , \22280 , \22281 , \22282 , \22283 , \22284 , \22285 , \22286 , \22287 , \22288 , \22289 , \22290 , \22291 , \22292 , \22293 , \22294 , \22295 , \22296 , \22297 , \22298 , \22299 , \22300 , \22301 , \22302 , \22303 , \22304 , \22305 , \22306 , \22307 , \22308 , \22309 , \22310 , \22311 , \22312 , \22313 , \22314 , \22315 , \22316 , \22317 , \22318 , \22319 , \22320 , \22321 , \22322 , \22323 , \22324 , \22325 , \22326 , \22327 , \22328 , \22329 , \22330 , \22331 , \22332 , \22333 , \22334 , \22335 , \22336 , \22337 );
and \U$13217 ( \22339 , RIee2b8b8_4954, \9462 );
and \U$13218 ( \22340 , RIee29f68_4936, \9464 );
and \U$13219 ( \22341 , RIee28bb8_4922, \9466 );
and \U$13220 ( \22342 , RIee27970_4909, \9468 );
and \U$13221 ( \22343 , RIdf2a0d0_1855, \9470 );
and \U$13222 ( \22344 , RIfe84e10_7856, \9472 );
and \U$13223 ( \22345 , RIdf262f0_1811, \9474 );
and \U$13224 ( \22346 , RIfe84ca8_7855, \9476 );
and \U$13225 ( \22347 , RIee27100_4903, \9478 );
and \U$13226 ( \22348 , RIee26b60_4899, \9480 );
and \U$13227 ( \22349 , RIfcd32f8_7425, \9482 );
and \U$13228 ( \22350 , RIee265c0_4895, \9484 );
and \U$13229 ( \22351 , RIfc9e300_6822, \9486 );
and \U$13230 ( \22352 , RIdf1f540_1733, \9488 );
and \U$13231 ( \22353 , RIee25eb8_4890, \9490 );
and \U$13232 ( \22354 , RIfe84b40_7854, \9492 );
and \U$13233 ( \22355 , RIdf16b70_1635, \9494 );
and \U$13234 ( \22356 , RIdf13e70_1603, \9496 );
and \U$13235 ( \22357 , RIdf11170_1571, \9498 );
and \U$13236 ( \22358 , RIdf0e470_1539, \9500 );
and \U$13237 ( \22359 , RIdf0b770_1507, \9502 );
and \U$13238 ( \22360 , RIdf08a70_1475, \9504 );
and \U$13239 ( \22361 , RIdf05d70_1443, \9506 );
and \U$13240 ( \22362 , RIdf03070_1411, \9508 );
and \U$13241 ( \22363 , RIdefd670_1347, \9510 );
and \U$13242 ( \22364 , RIdefa970_1315, \9512 );
and \U$13243 ( \22365 , RIdef7c70_1283, \9514 );
and \U$13244 ( \22366 , RIdef4f70_1251, \9516 );
and \U$13245 ( \22367 , RIdef2270_1219, \9518 );
and \U$13246 ( \22368 , RIdeef570_1187, \9520 );
and \U$13247 ( \22369 , RIdeec870_1155, \9522 );
and \U$13248 ( \22370 , RIdee9b70_1123, \9524 );
and \U$13249 ( \22371 , RIfec0348_8307, \9526 );
and \U$13250 ( \22372 , RIfcb54d8_7085, \9528 );
and \U$13251 ( \22373 , RIee23cf8_4866, \9530 );
and \U$13252 ( \22374 , RIfc54e30_5988, \9532 );
and \U$13253 ( \22375 , RIfec0078_8305, \9534 );
and \U$13254 ( \22376 , RIdee2988_1042, \9536 );
and \U$13255 ( \22377 , RIfec01e0_8306, \9538 );
and \U$13256 ( \22378 , RIdede770_995, \9540 );
and \U$13257 ( \22379 , RIfcd7ee8_7479, \9542 );
and \U$13258 ( \22380 , RIfcd43d8_7437, \9544 );
and \U$13259 ( \22381 , RIfc88eb0_6580, \9546 );
and \U$13260 ( \22382 , RIfc9e5d0_6824, \9548 );
and \U$13261 ( \22383 , RIded9478_936, \9550 );
and \U$13262 ( \22384 , RIded6fe8_910, \9552 );
and \U$13263 ( \22385 , RIded50f8_888, \9554 );
and \U$13264 ( \22386 , RIfeab330_8264, \9556 );
and \U$13265 ( \22387 , RIded03a0_833, \9558 );
and \U$13266 ( \22388 , RIdecd6a0_801, \9560 );
and \U$13267 ( \22389 , RIdeca9a0_769, \9562 );
and \U$13268 ( \22390 , RIdec7ca0_737, \9564 );
and \U$13269 ( \22391 , RIdeb41a0_513, \9566 );
and \U$13270 ( \22392 , RIde95f48_321, \9568 );
and \U$13271 ( \22393 , RIe16dda8_2627, \9570 );
and \U$13272 ( \22394 , RIe159ba0_2398, \9572 );
and \U$13273 ( \22395 , RIe1433a0_2142, \9574 );
and \U$13274 ( \22396 , RIdf37d98_2012, \9576 );
and \U$13275 ( \22397 , RIdf2c3f8_1880, \9578 );
and \U$13276 ( \22398 , RIdf1cc78_1704, \9580 );
and \U$13277 ( \22399 , RIdf00370_1379, \9582 );
and \U$13278 ( \22400 , RIdee6e70_1091, \9584 );
and \U$13279 ( \22401 , RIdedbbd8_964, \9586 );
and \U$13280 ( \22402 , RIde7be90_194, \9588 );
or \U$13281 ( \22403 , \22339 , \22340 , \22341 , \22342 , \22343 , \22344 , \22345 , \22346 , \22347 , \22348 , \22349 , \22350 , \22351 , \22352 , \22353 , \22354 , \22355 , \22356 , \22357 , \22358 , \22359 , \22360 , \22361 , \22362 , \22363 , \22364 , \22365 , \22366 , \22367 , \22368 , \22369 , \22370 , \22371 , \22372 , \22373 , \22374 , \22375 , \22376 , \22377 , \22378 , \22379 , \22380 , \22381 , \22382 , \22383 , \22384 , \22385 , \22386 , \22387 , \22388 , \22389 , \22390 , \22391 , \22392 , \22393 , \22394 , \22395 , \22396 , \22397 , \22398 , \22399 , \22400 , \22401 , \22402 );
or \U$13282 ( \22404 , \22338 , \22403 );
_DC g5885 ( \22405_nG5885 , \22404 , \9597 );
and \U$13283 ( \22406 , RIe19d238_3165, \9059 );
and \U$13284 ( \22407 , RIe19a538_3133, \9061 );
and \U$13285 ( \22408 , RIf145658_5249, \9063 );
and \U$13286 ( \22409 , RIe197838_3101, \9065 );
and \U$13287 ( \22410 , RIf1446e0_5238, \9067 );
and \U$13288 ( \22411 , RIe194b38_3069, \9069 );
and \U$13289 ( \22412 , RIe191e38_3037, \9071 );
and \U$13290 ( \22413 , RIe18f138_3005, \9073 );
and \U$13291 ( \22414 , RIe189738_2941, \9075 );
and \U$13292 ( \22415 , RIe186a38_2909, \9077 );
and \U$13293 ( \22416 , RIf143600_5226, \9079 );
and \U$13294 ( \22417 , RIe183d38_2877, \9081 );
and \U$13295 ( \22418 , RIf142c28_5219, \9083 );
and \U$13296 ( \22419 , RIe181038_2845, \9085 );
and \U$13297 ( \22420 , RIe17e338_2813, \9087 );
and \U$13298 ( \22421 , RIe17b638_2781, \9089 );
and \U$13299 ( \22422 , RIf1420e8_5211, \9091 );
and \U$13300 ( \22423 , RIf140a68_5195, \9093 );
and \U$13301 ( \22424 , RIf1401f8_5189, \9095 );
and \U$13302 ( \22425 , RIfebff10_8304, \9097 );
and \U$13303 ( \22426 , RIf13faf0_5184, \9099 );
and \U$13304 ( \22427 , RIf13ee48_5175, \9101 );
and \U$13305 ( \22428 , RIee3e2d8_5166, \9103 );
and \U$13306 ( \22429 , RIee3d1f8_5154, \9105 );
and \U$13307 ( \22430 , RIee3c118_5142, \9107 );
and \U$13308 ( \22431 , RIee3b038_5130, \9109 );
and \U$13309 ( \22432 , RIee39c88_5116, \9111 );
and \U$13310 ( \22433 , RIfe838f8_7841, \9113 );
and \U$13311 ( \22434 , RIf1701c8_5735, \9115 );
and \U$13312 ( \22435 , RIfc5ab00_6054, \9117 );
and \U$13313 ( \22436 , RIf16e008_5711, \9119 );
and \U$13314 ( \22437 , RIfcb0e88_7035, \9121 );
and \U$13315 ( \22438 , RIf16caf0_5696, \9123 );
and \U$13316 ( \22439 , RIe223590_4692, \9125 );
and \U$13317 ( \22440 , RIf16bce0_5686, \9127 );
and \U$13318 ( \22441 , RIe220890_4660, \9129 );
and \U$13319 ( \22442 , RIf16ac00_5674, \9131 );
and \U$13320 ( \22443 , RIe21db90_4628, \9133 );
and \U$13321 ( \22444 , RIe218190_4564, \9135 );
and \U$13322 ( \22445 , RIe215490_4532, \9137 );
and \U$13323 ( \22446 , RIf16a228_5667, \9139 );
and \U$13324 ( \22447 , RIe212790_4500, \9141 );
and \U$13325 ( \22448 , RIf168fe0_5654, \9143 );
and \U$13326 ( \22449 , RIe20fa90_4468, \9145 );
and \U$13327 ( \22450 , RIf167d98_5641, \9147 );
and \U$13328 ( \22451 , RIe20cd90_4436, \9149 );
and \U$13329 ( \22452 , RIe20a090_4404, \9151 );
and \U$13330 ( \22453 , RIe207390_4372, \9153 );
and \U$13331 ( \22454 , RIf1670f0_5632, \9155 );
and \U$13332 ( \22455 , RIf165ea8_5619, \9157 );
and \U$13333 ( \22456 , RIe202200_4314, \9159 );
and \U$13334 ( \22457 , RIfe83e98_7845, \9161 );
and \U$13335 ( \22458 , RIf164f30_5608, \9163 );
and \U$13336 ( \22459 , RIf1643f0_5600, \9165 );
and \U$13337 ( \22460 , RIfce8310_7664, \9167 );
and \U$13338 ( \22461 , RIf161df8_5573, \9169 );
and \U$13339 ( \22462 , RIf15ff08_5551, \9171 );
and \U$13340 ( \22463 , RIf15e018_5529, \9173 );
and \U$13341 ( \22464 , RIfe83d30_7844, \9175 );
and \U$13342 ( \22465 , RIfe84000_7846, \9177 );
and \U$13343 ( \22466 , RIf15cb00_5514, \9179 );
and \U$13344 ( \22467 , RIf15b5e8_5499, \9181 );
and \U$13345 ( \22468 , RIf15a508_5487, \9183 );
and \U$13346 ( \22469 , RIfc887a8_6575, \9185 );
or \U$13347 ( \22470 , \22406 , \22407 , \22408 , \22409 , \22410 , \22411 , \22412 , \22413 , \22414 , \22415 , \22416 , \22417 , \22418 , \22419 , \22420 , \22421 , \22422 , \22423 , \22424 , \22425 , \22426 , \22427 , \22428 , \22429 , \22430 , \22431 , \22432 , \22433 , \22434 , \22435 , \22436 , \22437 , \22438 , \22439 , \22440 , \22441 , \22442 , \22443 , \22444 , \22445 , \22446 , \22447 , \22448 , \22449 , \22450 , \22451 , \22452 , \22453 , \22454 , \22455 , \22456 , \22457 , \22458 , \22459 , \22460 , \22461 , \22462 , \22463 , \22464 , \22465 , \22466 , \22467 , \22468 , \22469 );
and \U$13348 ( \22471 , RIf158d20_5470, \9188 );
and \U$13349 ( \22472 , RIf157970_5456, \9190 );
and \U$13350 ( \22473 , RIf156cc8_5447, \9192 );
and \U$13351 ( \22474 , RIfe84438_7849, \9194 );
and \U$13352 ( \22475 , RIf156020_5438, \9196 );
and \U$13353 ( \22476 , RIfc51fc8_5955, \9198 );
and \U$13354 ( \22477 , RIf154568_5419, \9200 );
and \U$13355 ( \22478 , RIe1f51e0_4166, \9202 );
and \U$13356 ( \22479 , RIf153050_5404, \9204 );
and \U$13357 ( \22480 , RIf1519d0_5388, \9206 );
and \U$13358 ( \22481 , RIf150788_5375, \9208 );
and \U$13359 ( \22482 , RIfe842d0_7848, \9210 );
and \U$13360 ( \22483 , RIf14f810_5364, \9212 );
and \U$13361 ( \22484 , RIf14eb68_5355, \9214 );
and \U$13362 ( \22485 , RIf14dd58_5345, \9216 );
and \U$13363 ( \22486 , RIfe84168_7847, \9218 );
and \U$13364 ( \22487 , RIe1eb2f8_4053, \9220 );
and \U$13365 ( \22488 , RIe1e85f8_4021, \9222 );
and \U$13366 ( \22489 , RIe1e58f8_3989, \9224 );
and \U$13367 ( \22490 , RIe1e2bf8_3957, \9226 );
and \U$13368 ( \22491 , RIe1dfef8_3925, \9228 );
and \U$13369 ( \22492 , RIe1dd1f8_3893, \9230 );
and \U$13370 ( \22493 , RIe1da4f8_3861, \9232 );
and \U$13371 ( \22494 , RIe1d77f8_3829, \9234 );
and \U$13372 ( \22495 , RIe1d1df8_3765, \9236 );
and \U$13373 ( \22496 , RIe1cf0f8_3733, \9238 );
and \U$13374 ( \22497 , RIe1cc3f8_3701, \9240 );
and \U$13375 ( \22498 , RIe1c96f8_3669, \9242 );
and \U$13376 ( \22499 , RIe1c69f8_3637, \9244 );
and \U$13377 ( \22500 , RIe1c3cf8_3605, \9246 );
and \U$13378 ( \22501 , RIe1c0ff8_3573, \9248 );
and \U$13379 ( \22502 , RIe1be2f8_3541, \9250 );
and \U$13380 ( \22503 , RIf14c840_5330, \9252 );
and \U$13381 ( \22504 , RIf14b5f8_5317, \9254 );
and \U$13382 ( \22505 , RIfe83a60_7842, \9256 );
and \U$13383 ( \22506 , RIfe849d8_7853, \9258 );
and \U$13384 ( \22507 , RIfc74168_6343, \9260 );
and \U$13385 ( \22508 , RIf149b40_5298, \9262 );
and \U$13386 ( \22509 , RIfe83bc8_7843, \9264 );
and \U$13387 ( \22510 , RIfe84708_7851, \9266 );
and \U$13388 ( \22511 , RIf148d30_5288, \9268 );
and \U$13389 ( \22512 , RIf147ae8_5275, \9270 );
and \U$13390 ( \22513 , RIfe84870_7852, \9272 );
and \U$13391 ( \22514 , RIe1b0900_3386, \9274 );
and \U$13392 ( \22515 , RIf146fa8_5267, \9276 );
and \U$13393 ( \22516 , RIf146300_5258, \9278 );
and \U$13394 ( \22517 , RIfe845a0_7850, \9280 );
and \U$13395 ( \22518 , RIfe83790_7840, \9282 );
and \U$13396 ( \22519 , RIe1a8638_3293, \9284 );
and \U$13397 ( \22520 , RIe1a5938_3261, \9286 );
and \U$13398 ( \22521 , RIe1a2c38_3229, \9288 );
and \U$13399 ( \22522 , RIe19ff38_3197, \9290 );
and \U$13400 ( \22523 , RIe18c438_2973, \9292 );
and \U$13401 ( \22524 , RIe178938_2749, \9294 );
and \U$13402 ( \22525 , RIe226290_4724, \9296 );
and \U$13403 ( \22526 , RIe21ae90_4596, \9298 );
and \U$13404 ( \22527 , RIe204690_4340, \9300 );
and \U$13405 ( \22528 , RIe1fe6f0_4272, \9302 );
and \U$13406 ( \22529 , RIe1f7aa8_4195, \9304 );
and \U$13407 ( \22530 , RIe1f05f0_4112, \9306 );
and \U$13408 ( \22531 , RIe1d4af8_3797, \9308 );
and \U$13409 ( \22532 , RIe1bb5f8_3509, \9310 );
and \U$13410 ( \22533 , RIe1ae470_3360, \9312 );
and \U$13411 ( \22534 , RIe170aa8_2659, \9314 );
or \U$13412 ( \22535 , \22471 , \22472 , \22473 , \22474 , \22475 , \22476 , \22477 , \22478 , \22479 , \22480 , \22481 , \22482 , \22483 , \22484 , \22485 , \22486 , \22487 , \22488 , \22489 , \22490 , \22491 , \22492 , \22493 , \22494 , \22495 , \22496 , \22497 , \22498 , \22499 , \22500 , \22501 , \22502 , \22503 , \22504 , \22505 , \22506 , \22507 , \22508 , \22509 , \22510 , \22511 , \22512 , \22513 , \22514 , \22515 , \22516 , \22517 , \22518 , \22519 , \22520 , \22521 , \22522 , \22523 , \22524 , \22525 , \22526 , \22527 , \22528 , \22529 , \22530 , \22531 , \22532 , \22533 , \22534 );
or \U$13413 ( \22536 , \22470 , \22535 );
_DC g5909 ( \22537_nG5909 , \22536 , \9323 );
xor g590a ( \22538_nG590a , \22405_nG5885 , \22537_nG5909 );
buf \U$13414 ( \22539 , \22538_nG590a );
xor \U$13415 ( \22540 , \22539 , \22102 );
not \U$13416 ( \22541 , \22103 );
and \U$13417 ( \22542 , \22540 , \22541 );
and \U$13418 ( \22543 , \10687 , \22542 );
and \U$13419 ( \22544 , \10988 , \22103 );
nor \U$13420 ( \22545 , \22543 , \22544 );
and \U$13421 ( \22546 , \22102 , \21002 );
not \U$13422 ( \22547 , \22546 );
and \U$13423 ( \22548 , \22539 , \22547 );
xnor \U$13424 ( \22549 , \22545 , \22548 );
xor \U$13425 ( \22550 , \22273 , \22549 );
xor \U$13426 ( \22551 , \22264 , \22550 );
and \U$13427 ( \22552 , \22090 , \10983 );
_DC g65b0 ( \22553_nG65b0 , \22404 , \9597 );
_DC g65b1 ( \22554_nG65b1 , \22536 , \9323 );
and g65b2 ( \22555_nG65b2 , \22553_nG65b0 , \22554_nG65b1 );
buf \U$13428 ( \22556 , \22555_nG65b2 );
and \U$13429 ( \22557 , \22556 , \10691 );
nor \U$13430 ( \22558 , \22552 , \22557 );
xnor \U$13431 ( \22559 , \22558 , \10980 );
not \U$13432 ( \22560 , \22104 );
and \U$13433 ( \22561 , \22560 , \22548 );
xor \U$13434 ( \22562 , \22559 , \22561 );
and \U$13435 ( \22563 , \22093 , \22097 );
and \U$13436 ( \22564 , \22097 , \22104 );
and \U$13437 ( \22565 , \22093 , \22104 );
or \U$13438 ( \22566 , \22563 , \22564 , \22565 );
xor \U$13439 ( \22567 , \22562 , \22566 );
and \U$13440 ( \22568 , \21786 , \21790 );
and \U$13441 ( \22569 , \21790 , \21795 );
and \U$13442 ( \22570 , \21786 , \21795 );
or \U$13443 ( \22571 , \22568 , \22569 , \22570 );
xor \U$13444 ( \22572 , \22567 , \22571 );
xor \U$13445 ( \22573 , \22551 , \22572 );
xor \U$13446 ( \22574 , \22260 , \22573 );
and \U$13447 ( \22575 , \21823 , \22105 );
and \U$13448 ( \22576 , \22105 , \22120 );
and \U$13449 ( \22577 , \21823 , \22120 );
or \U$13450 ( \22578 , \22575 , \22576 , \22577 );
and \U$13451 ( \22579 , \21782 , \21796 );
and \U$13452 ( \22580 , \21796 , \21808 );
and \U$13453 ( \22581 , \21782 , \21808 );
or \U$13454 ( \22582 , \22579 , \22580 , \22581 );
xor \U$13455 ( \22583 , \22578 , \22582 );
and \U$13456 ( \22584 , \22110 , \22114 );
and \U$13457 ( \22585 , \22114 , \22119 );
and \U$13458 ( \22586 , \22110 , \22119 );
or \U$13459 ( \22587 , \22584 , \22585 , \22586 );
and \U$13460 ( \22588 , \19032 , \12790 );
and \U$13461 ( \22589 , \19558 , \12461 );
nor \U$13462 ( \22590 , \22588 , \22589 );
xnor \U$13463 ( \22591 , \22590 , \12780 );
and \U$13464 ( \22592 , \14950 , \16635 );
and \U$13465 ( \22593 , \15321 , \16301 );
nor \U$13466 ( \22594 , \22592 , \22593 );
xnor \U$13467 ( \22595 , \22594 , \16625 );
xor \U$13468 ( \22596 , \22591 , \22595 );
and \U$13469 ( \22597 , \13679 , \18090 );
and \U$13470 ( \22598 , \14024 , \17655 );
nor \U$13471 ( \22599 , \22597 , \22598 );
xnor \U$13472 ( \22600 , \22599 , \18046 );
xor \U$13473 ( \22601 , \22596 , \22600 );
xor \U$13474 ( \22602 , \22587 , \22601 );
and \U$13475 ( \22603 , \17627 , \14054 );
and \U$13476 ( \22604 , \18035 , \13692 );
nor \U$13477 ( \22605 , \22603 , \22604 );
xnor \U$13478 ( \22606 , \22605 , \14035 );
and \U$13479 ( \22607 , \12448 , \19534 );
and \U$13480 ( \22608 , \12769 , \19045 );
nor \U$13481 ( \22609 , \22607 , \22608 );
xnor \U$13482 ( \22610 , \22609 , \19540 );
xor \U$13483 ( \22611 , \22606 , \22610 );
and \U$13484 ( \22612 , \11270 , \21005 );
and \U$13485 ( \22613 , \11586 , \20557 );
nor \U$13486 ( \22614 , \22612 , \22613 );
xnor \U$13487 ( \22615 , \22614 , \21011 );
xor \U$13488 ( \22616 , \22611 , \22615 );
xor \U$13489 ( \22617 , \22602 , \22616 );
xor \U$13490 ( \22618 , \22583 , \22617 );
xor \U$13491 ( \22619 , \22574 , \22618 );
and \U$13492 ( \22620 , \21778 , \21809 );
and \U$13493 ( \22621 , \21809 , \22122 );
and \U$13494 ( \22622 , \21778 , \22122 );
or \U$13495 ( \22623 , \22620 , \22621 , \22622 );
xor \U$13496 ( \22624 , \22619 , \22623 );
and \U$13497 ( \22625 , \21774 , \22123 );
and \U$13498 ( \22626 , \22124 , \22127 );
or \U$13499 ( \22627 , \22625 , \22626 );
xor \U$13500 ( \22628 , \22624 , \22627 );
buf g9bd5 ( \22629_nG9bd5 , \22628 );
and \U$13501 ( \22630 , \10704 , \22629_nG9bd5 );
or \U$13502 ( \22631 , \22256 , \22630 );
xor \U$13503 ( \22632 , \10703 , \22631 );
buf \U$13504 ( \22633 , \22632 );
buf \U$13506 ( \22634 , \22633 );
xor \U$13507 ( \22635 , \22255 , \22634 );
buf \U$13508 ( \22636 , \22635 );
xor \U$13509 ( \22637 , \22244 , \22636 );
and \U$13510 ( \22638 , \21675 , \21709 );
and \U$13511 ( \22639 , \21675 , \21750 );
and \U$13512 ( \22640 , \21709 , \21750 );
or \U$13513 ( \22641 , \22638 , \22639 , \22640 );
buf \U$13514 ( \22642 , \22641 );
xor \U$13515 ( \22643 , \22637 , \22642 );
and \U$13516 ( \22644 , \22150 , \22643 );
and \U$13517 ( \22645 , \22140 , \22144 );
and \U$13518 ( \22646 , \22140 , \22149 );
and \U$13519 ( \22647 , \22144 , \22149 );
or \U$13520 ( \22648 , \22645 , \22646 , \22647 );
xor \U$13521 ( \22649 , \22644 , \22648 );
and \U$13522 ( \22650 , RIdec53d8_708, \9059 );
and \U$13523 ( \22651 , RIdec26d8_676, \9061 );
and \U$13524 ( \22652 , RIee20080_4823, \9063 );
and \U$13525 ( \22653 , RIdebf9d8_644, \9065 );
and \U$13526 ( \22654 , RIee1f3d8_4814, \9067 );
and \U$13527 ( \22655 , RIdebccd8_612, \9069 );
and \U$13528 ( \22656 , RIdeb9fd8_580, \9071 );
and \U$13529 ( \22657 , RIdeb72d8_548, \9073 );
and \U$13530 ( \22658 , RIee1ee38_4810, \9075 );
and \U$13531 ( \22659 , RIdeb18d8_484, \9077 );
and \U$13532 ( \22660 , RIee1e898_4806, \9079 );
and \U$13533 ( \22661 , RIdeaebd8_452, \9081 );
and \U$13534 ( \22662 , RIee1da88_4796, \9083 );
and \U$13535 ( \22663 , RIdeaa420_420, \9085 );
and \U$13536 ( \22664 , RIdea3b20_388, \9087 );
and \U$13537 ( \22665 , RIde9d220_356, \9089 );
and \U$13538 ( \22666 , RIee1cde0_4787, \9091 );
and \U$13539 ( \22667 , RIee1bd00_4775, \9093 );
and \U$13540 ( \22668 , RIee1b490_4769, \9095 );
and \U$13541 ( \22669 , RIfcd8a28_7487, \9097 );
and \U$13542 ( \22670 , RIde91088_297, \9099 );
and \U$13543 ( \22671 , RIde8d8c0_280, \9101 );
and \U$13544 ( \22672 , RIfe7dac0_7774, \9103 );
and \U$13545 ( \22673 , RIfe7d958_7773, \9105 );
and \U$13546 ( \22674 , RIee1a518_4758, \9107 );
and \U$13547 ( \22675 , RIee19e10_4753, \9109 );
and \U$13548 ( \22676 , RIee19b40_4751, \9111 );
and \U$13549 ( \22677 , RIfc768c8_6371, \9113 );
and \U$13550 ( \22678 , RIfcd05f8_7393, \9115 );
and \U$13551 ( \22679 , RIfe7dd90_7776, \9117 );
and \U$13552 ( \22680 , RIee38770_5101, \9119 );
and \U$13553 ( \22681 , RIfe7dc28_7775, \9121 );
and \U$13554 ( \22682 , RIe1653d8_2529, \9123 );
and \U$13555 ( \22683 , RIe1626d8_2497, \9125 );
and \U$13556 ( \22684 , RIee373c0_5087, \9127 );
and \U$13557 ( \22685 , RIe15f9d8_2465, \9129 );
and \U$13558 ( \22686 , RIee362e0_5075, \9131 );
and \U$13559 ( \22687 , RIe15ccd8_2433, \9133 );
and \U$13560 ( \22688 , RIe1572d8_2369, \9135 );
and \U$13561 ( \22689 , RIe1545d8_2337, \9137 );
and \U$13562 ( \22690 , RIfe7def8_7777, \9139 );
and \U$13563 ( \22691 , RIe1518d8_2305, \9141 );
and \U$13564 ( \22692 , RIfebdeb8_8281, \9143 );
and \U$13565 ( \22693 , RIe14ebd8_2273, \9145 );
and \U$13566 ( \22694 , RIfc649e8_6167, \9147 );
and \U$13567 ( \22695 , RIe14bed8_2241, \9149 );
and \U$13568 ( \22696 , RIe1491d8_2209, \9151 );
and \U$13569 ( \22697 , RIe1464d8_2177, \9153 );
and \U$13570 ( \22698 , RIfe7d7f0_7772, \9155 );
and \U$13571 ( \22699 , RIfe7d688_7771, \9157 );
and \U$13572 ( \22700 , RIee32230_5029, \9159 );
and \U$13573 ( \22701 , RIfceb9e8_7703, \9161 );
and \U$13574 ( \22702 , RIfebdd50_8280, \9163 );
and \U$13575 ( \22703 , RIfe7d520_7770, \9165 );
and \U$13576 ( \22704 , RIfebdbe8_8279, \9167 );
and \U$13577 ( \22705 , RIfe7d3b8_7769, \9169 );
and \U$13578 ( \22706 , RIfc734c0_6334, \9171 );
and \U$13579 ( \22707 , RIee2f968_5000, \9173 );
and \U$13580 ( \22708 , RIfccfab8_7385, \9175 );
and \U$13581 ( \22709 , RIee2d7a8_4976, \9177 );
and \U$13582 ( \22710 , RIdf357a0_1985, \9179 );
and \U$13583 ( \22711 , RIdf33310_1959, \9181 );
and \U$13584 ( \22712 , RIdf312b8_1936, \9183 );
and \U$13585 ( \22713 , RIdf2f0f8_1912, \9185 );
or \U$13586 ( \22714 , \22650 , \22651 , \22652 , \22653 , \22654 , \22655 , \22656 , \22657 , \22658 , \22659 , \22660 , \22661 , \22662 , \22663 , \22664 , \22665 , \22666 , \22667 , \22668 , \22669 , \22670 , \22671 , \22672 , \22673 , \22674 , \22675 , \22676 , \22677 , \22678 , \22679 , \22680 , \22681 , \22682 , \22683 , \22684 , \22685 , \22686 , \22687 , \22688 , \22689 , \22690 , \22691 , \22692 , \22693 , \22694 , \22695 , \22696 , \22697 , \22698 , \22699 , \22700 , \22701 , \22702 , \22703 , \22704 , \22705 , \22706 , \22707 , \22708 , \22709 , \22710 , \22711 , \22712 , \22713 );
and \U$13587 ( \22715 , RIee2bcf0_4957, \9188 );
and \U$13588 ( \22716 , RIee2a238_4938, \9190 );
and \U$13589 ( \22717 , RIee28e88_4924, \9192 );
and \U$13590 ( \22718 , RIee27c40_4911, \9194 );
and \U$13591 ( \22719 , RIfe7ce18_7765, \9196 );
and \U$13592 ( \22720 , RIfe7ccb0_7764, \9198 );
and \U$13593 ( \22721 , RIfe7cf80_7766, \9200 );
and \U$13594 ( \22722 , RIfe7cb48_7763, \9202 );
and \U$13595 ( \22723 , RIee27268_4904, \9204 );
and \U$13596 ( \22724 , RIee26e30_4901, \9206 );
and \U$13597 ( \22725 , RIee26890_4897, \9208 );
and \U$13598 ( \22726 , RIfcaa0d8_6957, \9210 );
and \U$13599 ( \22727 , RIee262f0_4893, \9212 );
and \U$13600 ( \22728 , RIfe7d250_7768, \9214 );
and \U$13601 ( \22729 , RIee26020_4891, \9216 );
and \U$13602 ( \22730 , RIfe7d0e8_7767, \9218 );
and \U$13603 ( \22731 , RIdf16fa8_1638, \9220 );
and \U$13604 ( \22732 , RIdf142a8_1606, \9222 );
and \U$13605 ( \22733 , RIdf115a8_1574, \9224 );
and \U$13606 ( \22734 , RIdf0e8a8_1542, \9226 );
and \U$13607 ( \22735 , RIdf0bba8_1510, \9228 );
and \U$13608 ( \22736 , RIdf08ea8_1478, \9230 );
and \U$13609 ( \22737 , RIdf061a8_1446, \9232 );
and \U$13610 ( \22738 , RIdf034a8_1414, \9234 );
and \U$13611 ( \22739 , RIdefdaa8_1350, \9236 );
and \U$13612 ( \22740 , RIdefada8_1318, \9238 );
and \U$13613 ( \22741 , RIdef80a8_1286, \9240 );
and \U$13614 ( \22742 , RIdef53a8_1254, \9242 );
and \U$13615 ( \22743 , RIdef26a8_1222, \9244 );
and \U$13616 ( \22744 , RIdeef9a8_1190, \9246 );
and \U$13617 ( \22745 , RIdeecca8_1158, \9248 );
and \U$13618 ( \22746 , RIdee9fa8_1126, \9250 );
and \U$13619 ( \22747 , RIee25648_4884, \9252 );
and \U$13620 ( \22748 , RIee249a0_4875, \9254 );
and \U$13621 ( \22749 , RIfebe020_8282, \9256 );
and \U$13622 ( \22750 , RIee23488_4860, \9258 );
and \U$13623 ( \22751 , RIfebe2f0_8284, \9260 );
and \U$13624 ( \22752 , RIfebe188_8283, \9262 );
and \U$13625 ( \22753 , RIfe7e1c8_7779, \9264 );
and \U$13626 ( \22754 , RIfe7e060_7778, \9266 );
and \U$13627 ( \22755 , RIfcbf7f8_7201, \9268 );
and \U$13628 ( \22756 , RIfc7aae0_6418, \9270 );
and \U$13629 ( \22757 , RIfc787b8_6393, \9272 );
and \U$13630 ( \22758 , RIfc618b0_6132, \9274 );
and \U$13631 ( \22759 , RIded98b0_939, \9276 );
and \U$13632 ( \22760 , RIded72b8_912, \9278 );
and \U$13633 ( \22761 , RIded5530_891, \9280 );
and \U$13634 ( \22762 , RIded2dd0_863, \9282 );
and \U$13635 ( \22763 , RIded07d8_836, \9284 );
and \U$13636 ( \22764 , RIdecdad8_804, \9286 );
and \U$13637 ( \22765 , RIdecadd8_772, \9288 );
and \U$13638 ( \22766 , RIdec80d8_740, \9290 );
and \U$13639 ( \22767 , RIdeb45d8_516, \9292 );
and \U$13640 ( \22768 , RIde96920_324, \9294 );
and \U$13641 ( \22769 , RIe16e1e0_2630, \9296 );
and \U$13642 ( \22770 , RIe159fd8_2401, \9298 );
and \U$13643 ( \22771 , RIe1437d8_2145, \9300 );
and \U$13644 ( \22772 , RIdf381d0_2015, \9302 );
and \U$13645 ( \22773 , RIdf2c830_1883, \9304 );
and \U$13646 ( \22774 , RIdf1d0b0_1707, \9306 );
and \U$13647 ( \22775 , RIdf007a8_1382, \9308 );
and \U$13648 ( \22776 , RIdee72a8_1094, \9310 );
and \U$13649 ( \22777 , RIdedc010_967, \9312 );
and \U$13650 ( \22778 , RIde7c868_197, \9314 );
or \U$13651 ( \22779 , \22715 , \22716 , \22717 , \22718 , \22719 , \22720 , \22721 , \22722 , \22723 , \22724 , \22725 , \22726 , \22727 , \22728 , \22729 , \22730 , \22731 , \22732 , \22733 , \22734 , \22735 , \22736 , \22737 , \22738 , \22739 , \22740 , \22741 , \22742 , \22743 , \22744 , \22745 , \22746 , \22747 , \22748 , \22749 , \22750 , \22751 , \22752 , \22753 , \22754 , \22755 , \22756 , \22757 , \22758 , \22759 , \22760 , \22761 , \22762 , \22763 , \22764 , \22765 , \22766 , \22767 , \22768 , \22769 , \22770 , \22771 , \22772 , \22773 , \22774 , \22775 , \22776 , \22777 , \22778 );
or \U$13652 ( \22780 , \22714 , \22779 );
_DC g2767 ( \22781_nG2767 , \22780 , \9323 );
buf \U$13653 ( \22782 , \22781_nG2767 );
and \U$13654 ( \22783 , RIe19d670_3168, \9333 );
and \U$13655 ( \22784 , RIe19a970_3136, \9335 );
and \U$13656 ( \22785 , RIfe7b630_7748, \9337 );
and \U$13657 ( \22786 , RIe197c70_3104, \9339 );
and \U$13658 ( \22787 , RIfe7b4c8_7747, \9341 );
and \U$13659 ( \22788 , RIe194f70_3072, \9343 );
and \U$13660 ( \22789 , RIe192270_3040, \9345 );
and \U$13661 ( \22790 , RIe18f570_3008, \9347 );
and \U$13662 ( \22791 , RIe189b70_2944, \9349 );
and \U$13663 ( \22792 , RIe186e70_2912, \9351 );
and \U$13664 ( \22793 , RIfe7b360_7746, \9353 );
and \U$13665 ( \22794 , RIe184170_2880, \9355 );
and \U$13666 ( \22795 , RIfe7b1f8_7745, \9357 );
and \U$13667 ( \22796 , RIe181470_2848, \9359 );
and \U$13668 ( \22797 , RIe17e770_2816, \9361 );
and \U$13669 ( \22798 , RIe17ba70_2784, \9363 );
and \U$13670 ( \22799 , RIf1423b8_5213, \9365 );
and \U$13671 ( \22800 , RIf140ea0_5198, \9367 );
and \U$13672 ( \22801 , RIf140360_5190, \9369 );
and \U$13673 ( \22802 , RIfe7b798_7749, \9371 );
and \U$13674 ( \22803 , RIf13fc58_5185, \9373 );
and \U$13675 ( \22804 , RIf13f280_5178, \9375 );
and \U$13676 ( \22805 , RIfc79460_6402, \9377 );
and \U$13677 ( \22806 , RIee3d4c8_5156, \9379 );
and \U$13678 ( \22807 , RIfe7b090_7744, \9381 );
and \U$13679 ( \22808 , RIfe7af28_7743, \9383 );
and \U$13680 ( \22809 , RIee39df0_5117, \9385 );
and \U$13681 ( \22810 , RIe1737a8_2691, \9387 );
and \U$13682 ( \22811 , RIfe7adc0_7742, \9389 );
and \U$13683 ( \22812 , RIfe7ac58_7741, \9391 );
and \U$13684 ( \22813 , RIf16e440_5714, \9393 );
and \U$13685 ( \22814 , RIfcb20d0_7048, \9395 );
and \U$13686 ( \22815 , RIfe7bd38_7753, \9397 );
and \U$13687 ( \22816 , RIe2239c8_4695, \9399 );
and \U$13688 ( \22817 , RIf16be48_5687, \9401 );
and \U$13689 ( \22818 , RIe220cc8_4663, \9403 );
and \U$13690 ( \22819 , RIf16aed0_5676, \9405 );
and \U$13691 ( \22820 , RIe21dfc8_4631, \9407 );
and \U$13692 ( \22821 , RIe2185c8_4567, \9409 );
and \U$13693 ( \22822 , RIe2158c8_4535, \9411 );
and \U$13694 ( \22823 , RIfebd7b0_8276, \9413 );
and \U$13695 ( \22824 , RIe212bc8_4503, \9415 );
and \U$13696 ( \22825 , RIfebd648_8275, \9417 );
and \U$13697 ( \22826 , RIe20fec8_4471, \9419 );
and \U$13698 ( \22827 , RIfe7b900_7750, \9421 );
and \U$13699 ( \22828 , RIe20d1c8_4439, \9423 );
and \U$13700 ( \22829 , RIe20a4c8_4407, \9425 );
and \U$13701 ( \22830 , RIe2077c8_4375, \9427 );
and \U$13702 ( \22831 , RIf167258_5633, \9429 );
and \U$13703 ( \22832 , RIf166178_5621, \9431 );
and \U$13704 ( \22833 , RIe2024d0_4316, \9433 );
and \U$13705 ( \22834 , RIfe7bbd0_7752, \9435 );
and \U$13706 ( \22835 , RIf165368_5611, \9437 );
and \U$13707 ( \22836 , RIf1646c0_5602, \9439 );
and \U$13708 ( \22837 , RIfcd0a30_7396, \9441 );
and \U$13709 ( \22838 , RIf1620c8_5575, \9443 );
and \U$13710 ( \22839 , RIf1601d8_5553, \9445 );
and \U$13711 ( \22840 , RIf15e2e8_5531, \9447 );
and \U$13712 ( \22841 , RIfe7ba68_7751, \9449 );
and \U$13713 ( \22842 , RIfe7bea0_7754, \9451 );
and \U$13714 ( \22843 , RIf15cdd0_5516, \9453 );
and \U$13715 ( \22844 , RIf15b8b8_5501, \9455 );
and \U$13716 ( \22845 , RIf15a7d8_5489, \9457 );
and \U$13717 ( \22846 , RIfca4840_6894, \9459 );
or \U$13718 ( \22847 , \22783 , \22784 , \22785 , \22786 , \22787 , \22788 , \22789 , \22790 , \22791 , \22792 , \22793 , \22794 , \22795 , \22796 , \22797 , \22798 , \22799 , \22800 , \22801 , \22802 , \22803 , \22804 , \22805 , \22806 , \22807 , \22808 , \22809 , \22810 , \22811 , \22812 , \22813 , \22814 , \22815 , \22816 , \22817 , \22818 , \22819 , \22820 , \22821 , \22822 , \22823 , \22824 , \22825 , \22826 , \22827 , \22828 , \22829 , \22830 , \22831 , \22832 , \22833 , \22834 , \22835 , \22836 , \22837 , \22838 , \22839 , \22840 , \22841 , \22842 , \22843 , \22844 , \22845 , \22846 );
and \U$13719 ( \22848 , RIf158ff0_5472, \9462 );
and \U$13720 ( \22849 , RIf157c40_5458, \9464 );
and \U$13721 ( \22850 , RIf156f98_5449, \9466 );
and \U$13722 ( \22851 , RIfe7c170_7756, \9468 );
and \U$13723 ( \22852 , RIf156458_5441, \9470 );
and \U$13724 ( \22853 , RIf155918_5433, \9472 );
and \U$13725 ( \22854 , RIf1549a0_5422, \9474 );
and \U$13726 ( \22855 , RIe1f54b0_4168, \9476 );
and \U$13727 ( \22856 , RIfe7c008_7755, \9478 );
and \U$13728 ( \22857 , RIf151b38_5389, \9480 );
and \U$13729 ( \22858 , RIf150bc0_5378, \9482 );
and \U$13730 ( \22859 , RIe1f32f0_4144, \9484 );
and \U$13731 ( \22860 , RIf14fae0_5366, \9486 );
and \U$13732 ( \22861 , RIf14ee38_5357, \9488 );
and \U$13733 ( \22862 , RIf14e028_5347, \9490 );
and \U$13734 ( \22863 , RIe1edff8_4085, \9492 );
and \U$13735 ( \22864 , RIe1eb730_4056, \9494 );
and \U$13736 ( \22865 , RIe1e8a30_4024, \9496 );
and \U$13737 ( \22866 , RIe1e5d30_3992, \9498 );
and \U$13738 ( \22867 , RIe1e3030_3960, \9500 );
and \U$13739 ( \22868 , RIe1e0330_3928, \9502 );
and \U$13740 ( \22869 , RIe1dd630_3896, \9504 );
and \U$13741 ( \22870 , RIe1da930_3864, \9506 );
and \U$13742 ( \22871 , RIe1d7c30_3832, \9508 );
and \U$13743 ( \22872 , RIe1d2230_3768, \9510 );
and \U$13744 ( \22873 , RIe1cf530_3736, \9512 );
and \U$13745 ( \22874 , RIe1cc830_3704, \9514 );
and \U$13746 ( \22875 , RIe1c9b30_3672, \9516 );
and \U$13747 ( \22876 , RIe1c6e30_3640, \9518 );
and \U$13748 ( \22877 , RIe1c4130_3608, \9520 );
and \U$13749 ( \22878 , RIe1c1430_3576, \9522 );
and \U$13750 ( \22879 , RIe1be730_3544, \9524 );
and \U$13751 ( \22880 , RIf14cb10_5332, \9526 );
and \U$13752 ( \22881 , RIf14b8c8_5319, \9528 );
and \U$13753 ( \22882 , RIfebda80_8278, \9530 );
and \U$13754 ( \22883 , RIfe7c878_7761, \9532 );
and \U$13755 ( \22884 , RIf14a680_5306, \9534 );
and \U$13756 ( \22885 , RIfe7c2d8_7757, \9536 );
and \U$13757 ( \22886 , RIfe7c9e0_7762, \9538 );
and \U$13758 ( \22887 , RIfe7c440_7758, \9540 );
and \U$13759 ( \22888 , RIf149000_5290, \9542 );
and \U$13760 ( \22889 , RIf147db8_5277, \9544 );
and \U$13761 ( \22890 , RIe1b2688_3407, \9546 );
and \U$13762 ( \22891 , RIfebd918_8277, \9548 );
and \U$13763 ( \22892 , RIfe7c5a8_7759, \9550 );
and \U$13764 ( \22893 , RIf146738_5261, \9552 );
and \U$13765 ( \22894 , RIfe7c710_7760, \9554 );
and \U$13766 ( \22895 , RIe1aad98_3321, \9556 );
and \U$13767 ( \22896 , RIe1a8a70_3296, \9558 );
and \U$13768 ( \22897 , RIe1a5d70_3264, \9560 );
and \U$13769 ( \22898 , RIe1a3070_3232, \9562 );
and \U$13770 ( \22899 , RIe1a0370_3200, \9564 );
and \U$13771 ( \22900 , RIe18c870_2976, \9566 );
and \U$13772 ( \22901 , RIe178d70_2752, \9568 );
and \U$13773 ( \22902 , RIe2266c8_4727, \9570 );
and \U$13774 ( \22903 , RIe21b2c8_4599, \9572 );
and \U$13775 ( \22904 , RIe204ac8_4343, \9574 );
and \U$13776 ( \22905 , RIe1feb28_4275, \9576 );
and \U$13777 ( \22906 , RIe1f7ee0_4198, \9578 );
and \U$13778 ( \22907 , RIe1f0a28_4115, \9580 );
and \U$13779 ( \22908 , RIe1d4f30_3800, \9582 );
and \U$13780 ( \22909 , RIe1bba30_3512, \9584 );
and \U$13781 ( \22910 , RIe1ae8a8_3363, \9586 );
and \U$13782 ( \22911 , RIe170ee0_2662, \9588 );
or \U$13783 ( \22912 , \22848 , \22849 , \22850 , \22851 , \22852 , \22853 , \22854 , \22855 , \22856 , \22857 , \22858 , \22859 , \22860 , \22861 , \22862 , \22863 , \22864 , \22865 , \22866 , \22867 , \22868 , \22869 , \22870 , \22871 , \22872 , \22873 , \22874 , \22875 , \22876 , \22877 , \22878 , \22879 , \22880 , \22881 , \22882 , \22883 , \22884 , \22885 , \22886 , \22887 , \22888 , \22889 , \22890 , \22891 , \22892 , \22893 , \22894 , \22895 , \22896 , \22897 , \22898 , \22899 , \22900 , \22901 , \22902 , \22903 , \22904 , \22905 , \22906 , \22907 , \22908 , \22909 , \22910 , \22911 );
or \U$13784 ( \22913 , \22847 , \22912 );
_DC g3894 ( \22914_nG3894 , \22913 , \9597 );
buf \U$13785 ( \22915 , \22914_nG3894 );
xor \U$13786 ( \22916 , \22782 , \22915 );
and \U$13787 ( \22917 , RIdec5270_707, \9059 );
and \U$13788 ( \22918 , RIdec2570_675, \9061 );
and \U$13789 ( \22919 , RIee1ff18_4822, \9063 );
and \U$13790 ( \22920 , RIdebf870_643, \9065 );
and \U$13791 ( \22921 , RIfe7f848_7795, \9067 );
and \U$13792 ( \22922 , RIdebcb70_611, \9069 );
and \U$13793 ( \22923 , RIdeb9e70_579, \9071 );
and \U$13794 ( \22924 , RIdeb7170_547, \9073 );
and \U$13795 ( \22925 , RIfe7fc80_7798, \9075 );
and \U$13796 ( \22926 , RIdeb1770_483, \9077 );
and \U$13797 ( \22927 , RIfca5d58_6909, \9079 );
and \U$13798 ( \22928 , RIdeaea70_451, \9081 );
and \U$13799 ( \22929 , RIfcaf808_7019, \9083 );
and \U$13800 ( \22930 , RIdeaa0d8_419, \9085 );
and \U$13801 ( \22931 , RIdea37d8_387, \9087 );
and \U$13802 ( \22932 , RIde9ced8_355, \9089 );
and \U$13803 ( \22933 , RIfcdc3d0_7528, \9091 );
and \U$13804 ( \22934 , RIfcce438_7369, \9093 );
and \U$13805 ( \22935 , RIfcb0a50_7032, \9095 );
and \U$13806 ( \22936 , RIfc75680_6358, \9097 );
and \U$13807 ( \22937 , RIde90d40_296, \9099 );
and \U$13808 ( \22938 , RIfe7f9b0_7796, \9101 );
and \U$13809 ( \22939 , RIde89720_260, \9103 );
and \U$13810 ( \22940 , RIde85580_240, \9105 );
and \U$13811 ( \22941 , RIde81728_221, \9107 );
and \U$13812 ( \22942 , RIfc52f40_5966, \9109 );
and \U$13813 ( \22943 , RIfc82100_6502, \9111 );
and \U$13814 ( \22944 , RIfca7108_6923, \9113 );
and \U$13815 ( \22945 , RIfe7fb18_7797, \9115 );
and \U$13816 ( \22946 , RIe16b648_2599, \9117 );
and \U$13817 ( \22947 , RIe169a28_2579, \9119 );
and \U$13818 ( \22948 , RIe167ca0_2558, \9121 );
and \U$13819 ( \22949 , RIe165270_2528, \9123 );
and \U$13820 ( \22950 , RIe162570_2496, \9125 );
and \U$13821 ( \22951 , RIee37258_5086, \9127 );
and \U$13822 ( \22952 , RIe15f870_2464, \9129 );
and \U$13823 ( \22953 , RIee36178_5074, \9131 );
and \U$13824 ( \22954 , RIe15cb70_2432, \9133 );
and \U$13825 ( \22955 , RIe157170_2368, \9135 );
and \U$13826 ( \22956 , RIe154470_2336, \9137 );
and \U$13827 ( \22957 , RIfc86fc0_6558, \9139 );
and \U$13828 ( \22958 , RIe151770_2304, \9141 );
and \U$13829 ( \22959 , RIfc4eff8_5921, \9143 );
and \U$13830 ( \22960 , RIe14ea70_2272, \9145 );
and \U$13831 ( \22961 , RIfce1290_7584, \9147 );
and \U$13832 ( \22962 , RIe14bd70_2240, \9149 );
and \U$13833 ( \22963 , RIe149070_2208, \9151 );
and \U$13834 ( \22964 , RIe146370_2176, \9153 );
and \U$13835 ( \22965 , RIee34558_5054, \9155 );
and \U$13836 ( \22966 , RIee331a8_5040, \9157 );
and \U$13837 ( \22967 , RIee320c8_5028, \9159 );
and \U$13838 ( \22968 , RIee31150_5017, \9161 );
and \U$13839 ( \22969 , RIfe800b8_7801, \9163 );
and \U$13840 ( \22970 , RIfe7ff50_7800, \9165 );
and \U$13841 ( \22971 , RIdf3caf0_2067, \9167 );
and \U$13842 ( \22972 , RIfe7fde8_7799, \9169 );
and \U$13843 ( \22973 , RIfcc8330_7300, \9171 );
and \U$13844 ( \22974 , RIee2f800_4999, \9173 );
and \U$13845 ( \22975 , RIfca0d30_6852, \9175 );
and \U$13846 ( \22976 , RIee2d640_4975, \9177 );
and \U$13847 ( \22977 , RIdf35638_1984, \9179 );
and \U$13848 ( \22978 , RIdf331a8_1958, \9181 );
and \U$13849 ( \22979 , RIdf31150_1935, \9183 );
and \U$13850 ( \22980 , RIdf2ef90_1911, \9185 );
or \U$13851 ( \22981 , \22917 , \22918 , \22919 , \22920 , \22921 , \22922 , \22923 , \22924 , \22925 , \22926 , \22927 , \22928 , \22929 , \22930 , \22931 , \22932 , \22933 , \22934 , \22935 , \22936 , \22937 , \22938 , \22939 , \22940 , \22941 , \22942 , \22943 , \22944 , \22945 , \22946 , \22947 , \22948 , \22949 , \22950 , \22951 , \22952 , \22953 , \22954 , \22955 , \22956 , \22957 , \22958 , \22959 , \22960 , \22961 , \22962 , \22963 , \22964 , \22965 , \22966 , \22967 , \22968 , \22969 , \22970 , \22971 , \22972 , \22973 , \22974 , \22975 , \22976 , \22977 , \22978 , \22979 , \22980 );
and \U$13852 ( \22982 , RIee2bb88_4956, \9188 );
and \U$13853 ( \22983 , RIee2a0d0_4937, \9190 );
and \U$13854 ( \22984 , RIee28d20_4923, \9192 );
and \U$13855 ( \22985 , RIfe7f578_7793, \9194 );
and \U$13856 ( \22986 , RIdf2a238_1856, \9196 );
and \U$13857 ( \22987 , RIdf27f10_1831, \9198 );
and \U$13858 ( \22988 , RIfe7f6e0_7794, \9200 );
and \U$13859 ( \22989 , RIdf246d0_1791, \9202 );
and \U$13860 ( \22990 , RIfcce9d8_7373, \9204 );
and \U$13861 ( \22991 , RIfc63638_6153, \9206 );
and \U$13862 ( \22992 , RIdf22c18_1772, \9208 );
and \U$13863 ( \22993 , RIfc62990_6144, \9210 );
and \U$13864 ( \22994 , RIdf21700_1757, \9212 );
and \U$13865 ( \22995 , RIdf1f810_1735, \9214 );
and \U$13866 ( \22996 , RIfeaa958_8257, \9216 );
and \U$13867 ( \22997 , RIdf19168_1662, \9218 );
and \U$13868 ( \22998 , RIdf16e40_1637, \9220 );
and \U$13869 ( \22999 , RIdf14140_1605, \9222 );
and \U$13870 ( \23000 , RIdf11440_1573, \9224 );
and \U$13871 ( \23001 , RIdf0e740_1541, \9226 );
and \U$13872 ( \23002 , RIdf0ba40_1509, \9228 );
and \U$13873 ( \23003 , RIdf08d40_1477, \9230 );
and \U$13874 ( \23004 , RIdf06040_1445, \9232 );
and \U$13875 ( \23005 , RIdf03340_1413, \9234 );
and \U$13876 ( \23006 , RIdefd940_1349, \9236 );
and \U$13877 ( \23007 , RIdefac40_1317, \9238 );
and \U$13878 ( \23008 , RIdef7f40_1285, \9240 );
and \U$13879 ( \23009 , RIdef5240_1253, \9242 );
and \U$13880 ( \23010 , RIdef2540_1221, \9244 );
and \U$13881 ( \23011 , RIdeef840_1189, \9246 );
and \U$13882 ( \23012 , RIdeecb40_1157, \9248 );
and \U$13883 ( \23013 , RIdee9e40_1125, \9250 );
and \U$13884 ( \23014 , RIfcb7800_7110, \9252 );
and \U$13885 ( \23015 , RIee24838_4874, \9254 );
and \U$13886 ( \23016 , RIfc4cb68_5895, \9256 );
and \U$13887 ( \23017 , RIee23320_4859, \9258 );
and \U$13888 ( \23018 , RIfe80388_7803, \9260 );
and \U$13889 ( \23019 , RIdee2c58_1044, \9262 );
and \U$13890 ( \23020 , RIfe80220_7802, \9264 );
and \U$13891 ( \23021 , RIdedea40_997, \9266 );
and \U$13892 ( \23022 , RIfc98900_6758, \9268 );
and \U$13893 ( \23023 , RIee223a8_4848, \9270 );
and \U$13894 ( \23024 , RIfcc8600_7302, \9272 );
and \U$13895 ( \23025 , RIee212c8_4836, \9274 );
and \U$13896 ( \23026 , RIded9748_938, \9276 );
and \U$13897 ( \23027 , RIfe804f0_7804, \9278 );
and \U$13898 ( \23028 , RIded53c8_890, \9280 );
and \U$13899 ( \23029 , RIded2c68_862, \9282 );
and \U$13900 ( \23030 , RIded0670_835, \9284 );
and \U$13901 ( \23031 , RIdecd970_803, \9286 );
and \U$13902 ( \23032 , RIdecac70_771, \9288 );
and \U$13903 ( \23033 , RIdec7f70_739, \9290 );
and \U$13904 ( \23034 , RIdeb4470_515, \9292 );
and \U$13905 ( \23035 , RIde965d8_323, \9294 );
and \U$13906 ( \23036 , RIe16e078_2629, \9296 );
and \U$13907 ( \23037 , RIe159e70_2400, \9298 );
and \U$13908 ( \23038 , RIe143670_2144, \9300 );
and \U$13909 ( \23039 , RIdf38068_2014, \9302 );
and \U$13910 ( \23040 , RIdf2c6c8_1882, \9304 );
and \U$13911 ( \23041 , RIdf1cf48_1706, \9306 );
and \U$13912 ( \23042 , RIdf00640_1381, \9308 );
and \U$13913 ( \23043 , RIdee7140_1093, \9310 );
and \U$13914 ( \23044 , RIdedbea8_966, \9312 );
and \U$13915 ( \23045 , RIde7c520_196, \9314 );
or \U$13916 ( \23046 , \22982 , \22983 , \22984 , \22985 , \22986 , \22987 , \22988 , \22989 , \22990 , \22991 , \22992 , \22993 , \22994 , \22995 , \22996 , \22997 , \22998 , \22999 , \23000 , \23001 , \23002 , \23003 , \23004 , \23005 , \23006 , \23007 , \23008 , \23009 , \23010 , \23011 , \23012 , \23013 , \23014 , \23015 , \23016 , \23017 , \23018 , \23019 , \23020 , \23021 , \23022 , \23023 , \23024 , \23025 , \23026 , \23027 , \23028 , \23029 , \23030 , \23031 , \23032 , \23033 , \23034 , \23035 , \23036 , \23037 , \23038 , \23039 , \23040 , \23041 , \23042 , \23043 , \23044 , \23045 );
or \U$13917 ( \23047 , \22981 , \23046 );
_DC g27ec ( \23048_nG27ec , \23047 , \9323 );
buf \U$13918 ( \23049 , \23048_nG27ec );
and \U$13919 ( \23050 , RIe19d508_3167, \9333 );
and \U$13920 ( \23051 , RIe19a808_3135, \9335 );
and \U$13921 ( \23052 , RIfe7ee70_7788, \9337 );
and \U$13922 ( \23053 , RIe197b08_3103, \9339 );
and \U$13923 ( \23054 , RIfe7efd8_7789, \9341 );
and \U$13924 ( \23055 , RIe194e08_3071, \9343 );
and \U$13925 ( \23056 , RIe192108_3039, \9345 );
and \U$13926 ( \23057 , RIe18f408_3007, \9347 );
and \U$13927 ( \23058 , RIe189a08_2943, \9349 );
and \U$13928 ( \23059 , RIe186d08_2911, \9351 );
and \U$13929 ( \23060 , RIf143768_5227, \9353 );
and \U$13930 ( \23061 , RIe184008_2879, \9355 );
and \U$13931 ( \23062 , RIfc4bbf0_5884, \9357 );
and \U$13932 ( \23063 , RIe181308_2847, \9359 );
and \U$13933 ( \23064 , RIe17e608_2815, \9361 );
and \U$13934 ( \23065 , RIe17b908_2783, \9363 );
and \U$13935 ( \23066 , RIfe7f410_7792, \9365 );
and \U$13936 ( \23067 , RIf140d38_5197, \9367 );
and \U$13937 ( \23068 , RIe176fe8_2731, \9369 );
and \U$13938 ( \23069 , RIe175ad0_2716, \9371 );
and \U$13939 ( \23070 , RIfe7f2a8_7791, \9373 );
and \U$13940 ( \23071 , RIf13f118_5177, \9375 );
and \U$13941 ( \23072 , RIee3e440_5167, \9377 );
and \U$13942 ( \23073 , RIee3d360_5155, \9379 );
and \U$13943 ( \23074 , RIee3c280_5143, \9381 );
and \U$13944 ( \23075 , RIee3b1a0_5131, \9383 );
and \U$13945 ( \23076 , RIfe7f140_7790, \9385 );
and \U$13946 ( \23077 , RIe173640_2690, \9387 );
and \U$13947 ( \23078 , RIf170330_5736, \9389 );
and \U$13948 ( \23079 , RIf16f520_5726, \9391 );
and \U$13949 ( \23080 , RIf16e2d8_5713, \9393 );
and \U$13950 ( \23081 , RIf16d630_5704, \9395 );
and \U$13951 ( \23082 , RIfe7ea38_7785, \9397 );
and \U$13952 ( \23083 , RIe223860_4694, \9399 );
and \U$13953 ( \23084 , RIfc9c410_6800, \9401 );
and \U$13954 ( \23085 , RIe220b60_4662, \9403 );
and \U$13955 ( \23086 , RIfcb8340_7118, \9405 );
and \U$13956 ( \23087 , RIe21de60_4630, \9407 );
and \U$13957 ( \23088 , RIe218460_4566, \9409 );
and \U$13958 ( \23089 , RIe215760_4534, \9411 );
and \U$13959 ( \23090 , RIfc9cc80_6806, \9413 );
and \U$13960 ( \23091 , RIe212a60_4502, \9415 );
and \U$13961 ( \23092 , RIfc4ddb0_5908, \9417 );
and \U$13962 ( \23093 , RIe20fd60_4470, \9419 );
and \U$13963 ( \23094 , RIfc873f8_6561, \9421 );
and \U$13964 ( \23095 , RIe20d060_4438, \9423 );
and \U$13965 ( \23096 , RIe20a360_4406, \9425 );
and \U$13966 ( \23097 , RIe207660_4374, \9427 );
and \U$13967 ( \23098 , RIfc86750_6552, \9429 );
and \U$13968 ( \23099 , RIfc4e4b8_5913, \9431 );
and \U$13969 ( \23100 , RIe202368_4315, \9433 );
and \U$13970 ( \23101 , RIe200a18_4297, \9435 );
and \U$13971 ( \23102 , RIf165200_5610, \9437 );
and \U$13972 ( \23103 , RIf164558_5601, \9439 );
and \U$13973 ( \23104 , RIf163478_5589, \9441 );
and \U$13974 ( \23105 , RIf161f60_5574, \9443 );
and \U$13975 ( \23106 , RIf160070_5552, \9445 );
and \U$13976 ( \23107 , RIf15e180_5530, \9447 );
and \U$13977 ( \23108 , RIe1fcc38_4253, \9449 );
and \U$13978 ( \23109 , RIe1fb9f0_4240, \9451 );
and \U$13979 ( \23110 , RIf15cc68_5515, \9453 );
and \U$13980 ( \23111 , RIf15b750_5500, \9455 );
and \U$13981 ( \23112 , RIf15a670_5488, \9457 );
and \U$13982 ( \23113 , RIf159c98_5481, \9459 );
or \U$13983 ( \23114 , \23050 , \23051 , \23052 , \23053 , \23054 , \23055 , \23056 , \23057 , \23058 , \23059 , \23060 , \23061 , \23062 , \23063 , \23064 , \23065 , \23066 , \23067 , \23068 , \23069 , \23070 , \23071 , \23072 , \23073 , \23074 , \23075 , \23076 , \23077 , \23078 , \23079 , \23080 , \23081 , \23082 , \23083 , \23084 , \23085 , \23086 , \23087 , \23088 , \23089 , \23090 , \23091 , \23092 , \23093 , \23094 , \23095 , \23096 , \23097 , \23098 , \23099 , \23100 , \23101 , \23102 , \23103 , \23104 , \23105 , \23106 , \23107 , \23108 , \23109 , \23110 , \23111 , \23112 , \23113 );
and \U$13984 ( \23115 , RIf158e88_5471, \9462 );
and \U$13985 ( \23116 , RIf157ad8_5457, \9464 );
and \U$13986 ( \23117 , RIf156e30_5448, \9466 );
and \U$13987 ( \23118 , RIfe7e768_7783, \9468 );
and \U$13988 ( \23119 , RIf1562f0_5440, \9470 );
and \U$13989 ( \23120 , RIf1557b0_5432, \9472 );
and \U$13990 ( \23121 , RIf154838_5421, \9474 );
and \U$13991 ( \23122 , RIfe7e8d0_7784, \9476 );
and \U$13992 ( \23123 , RIf1531b8_5405, \9478 );
and \U$13993 ( \23124 , RIfc52400_5958, \9480 );
and \U$13994 ( \23125 , RIf150a58_5377, \9482 );
and \U$13995 ( \23126 , RIe1f3188_4143, \9484 );
and \U$13996 ( \23127 , RIf14f978_5365, \9486 );
and \U$13997 ( \23128 , RIf14ecd0_5356, \9488 );
and \U$13998 ( \23129 , RIf14dec0_5346, \9490 );
and \U$13999 ( \23130 , RIe1ede90_4084, \9492 );
and \U$14000 ( \23131 , RIe1eb5c8_4055, \9494 );
and \U$14001 ( \23132 , RIe1e88c8_4023, \9496 );
and \U$14002 ( \23133 , RIe1e5bc8_3991, \9498 );
and \U$14003 ( \23134 , RIe1e2ec8_3959, \9500 );
and \U$14004 ( \23135 , RIe1e01c8_3927, \9502 );
and \U$14005 ( \23136 , RIe1dd4c8_3895, \9504 );
and \U$14006 ( \23137 , RIe1da7c8_3863, \9506 );
and \U$14007 ( \23138 , RIe1d7ac8_3831, \9508 );
and \U$14008 ( \23139 , RIe1d20c8_3767, \9510 );
and \U$14009 ( \23140 , RIe1cf3c8_3735, \9512 );
and \U$14010 ( \23141 , RIe1cc6c8_3703, \9514 );
and \U$14011 ( \23142 , RIe1c99c8_3671, \9516 );
and \U$14012 ( \23143 , RIe1c6cc8_3639, \9518 );
and \U$14013 ( \23144 , RIe1c3fc8_3607, \9520 );
and \U$14014 ( \23145 , RIe1c12c8_3575, \9522 );
and \U$14015 ( \23146 , RIe1be5c8_3543, \9524 );
and \U$14016 ( \23147 , RIf14c9a8_5331, \9526 );
and \U$14017 ( \23148 , RIf14b760_5318, \9528 );
and \U$14018 ( \23149 , RIfe7ed08_7787, \9530 );
and \U$14019 ( \23150 , RIfe7e600_7782, \9532 );
and \U$14020 ( \23151 , RIf14a518_5305, \9534 );
and \U$14021 ( \23152 , RIfca1f78_6865, \9536 );
and \U$14022 ( \23153 , RIfe7eba0_7786, \9538 );
and \U$14023 ( \23154 , RIfe7e498_7781, \9540 );
and \U$14024 ( \23155 , RIf148e98_5289, \9542 );
and \U$14025 ( \23156 , RIf147c50_5276, \9544 );
and \U$14026 ( \23157 , RIfe7e330_7780, \9546 );
and \U$14027 ( \23158 , RIe1b0a68_3387, \9548 );
and \U$14028 ( \23159 , RIf147278_5269, \9550 );
and \U$14029 ( \23160 , RIf1465d0_5260, \9552 );
and \U$14030 ( \23161 , RIe1ac418_3337, \9554 );
and \U$14031 ( \23162 , RIe1aac30_3320, \9556 );
and \U$14032 ( \23163 , RIe1a8908_3295, \9558 );
and \U$14033 ( \23164 , RIe1a5c08_3263, \9560 );
and \U$14034 ( \23165 , RIe1a2f08_3231, \9562 );
and \U$14035 ( \23166 , RIe1a0208_3199, \9564 );
and \U$14036 ( \23167 , RIe18c708_2975, \9566 );
and \U$14037 ( \23168 , RIe178c08_2751, \9568 );
and \U$14038 ( \23169 , RIe226560_4726, \9570 );
and \U$14039 ( \23170 , RIe21b160_4598, \9572 );
and \U$14040 ( \23171 , RIe204960_4342, \9574 );
and \U$14041 ( \23172 , RIe1fe9c0_4274, \9576 );
and \U$14042 ( \23173 , RIe1f7d78_4197, \9578 );
and \U$14043 ( \23174 , RIe1f08c0_4114, \9580 );
and \U$14044 ( \23175 , RIe1d4dc8_3799, \9582 );
and \U$14045 ( \23176 , RIe1bb8c8_3511, \9584 );
and \U$14046 ( \23177 , RIe1ae740_3362, \9586 );
and \U$14047 ( \23178 , RIe170d78_2661, \9588 );
or \U$14048 ( \23179 , \23115 , \23116 , \23117 , \23118 , \23119 , \23120 , \23121 , \23122 , \23123 , \23124 , \23125 , \23126 , \23127 , \23128 , \23129 , \23130 , \23131 , \23132 , \23133 , \23134 , \23135 , \23136 , \23137 , \23138 , \23139 , \23140 , \23141 , \23142 , \23143 , \23144 , \23145 , \23146 , \23147 , \23148 , \23149 , \23150 , \23151 , \23152 , \23153 , \23154 , \23155 , \23156 , \23157 , \23158 , \23159 , \23160 , \23161 , \23162 , \23163 , \23164 , \23165 , \23166 , \23167 , \23168 , \23169 , \23170 , \23171 , \23172 , \23173 , \23174 , \23175 , \23176 , \23177 , \23178 );
or \U$14049 ( \23180 , \23114 , \23179 );
_DC g3919 ( \23181_nG3919 , \23180 , \9597 );
buf \U$14050 ( \23182 , \23181_nG3919 );
and \U$14051 ( \23183 , \23049 , \23182 );
and \U$14052 ( \23184 , \21239 , \21372 );
and \U$14053 ( \23185 , \21372 , \21647 );
and \U$14054 ( \23186 , \21239 , \21647 );
or \U$14055 ( \23187 , \23184 , \23185 , \23186 );
and \U$14056 ( \23188 , \23182 , \23187 );
and \U$14057 ( \23189 , \23049 , \23187 );
or \U$14058 ( \23190 , \23183 , \23188 , \23189 );
xor \U$14059 ( \23191 , \22916 , \23190 );
buf g4418 ( \23192_nG4418 , \23191 );
xor \U$14060 ( \23193 , \23049 , \23182 );
xor \U$14061 ( \23194 , \23193 , \23187 );
buf g441b ( \23195_nG441b , \23194 );
nand \U$14062 ( \23196 , \23195_nG441b , \21649_nG441e );
and \U$14063 ( \23197 , \23192_nG4418 , \23196 );
xor \U$14064 ( \23198 , \23195_nG441b , \21649_nG441e );
not \U$14065 ( \23199 , \23198 );
xor \U$14066 ( \23200 , \23192_nG4418 , \23195_nG441b );
and \U$14067 ( \23201 , \23199 , \23200 );
and \U$14069 ( \23202 , \23198 , \10694_nG9c0e );
or \U$14070 ( \23203 , 1'b0 , \23202 );
xor \U$14071 ( \23204 , \23197 , \23203 );
xor \U$14072 ( \23205 , \23197 , \23204 );
buf \U$14073 ( \23206 , \23205 );
buf \U$14074 ( \23207 , \23206 );
xor \U$14075 ( \23208 , \22649 , \23207 );
and \U$14076 ( \23209 , \22244 , \22636 );
and \U$14077 ( \23210 , \22244 , \22642 );
and \U$14078 ( \23211 , \22636 , \22642 );
or \U$14079 ( \23212 , \23209 , \23210 , \23211 );
and \U$14080 ( \23213 , \23208 , \23212 );
and \U$14081 ( \23214 , \22175 , \22181 );
and \U$14082 ( \23215 , \22175 , \22188 );
and \U$14083 ( \23216 , \22181 , \22188 );
or \U$14084 ( \23217 , \23214 , \23215 , \23216 );
buf \U$14085 ( \23218 , \23217 );
and \U$14086 ( \23219 , \22196 , \22233 );
and \U$14087 ( \23220 , \22196 , \22240 );
and \U$14088 ( \23221 , \22233 , \22240 );
or \U$14089 ( \23222 , \23219 , \23220 , \23221 );
buf \U$14090 ( \23223 , \23222 );
and \U$14091 ( \23224 , \12157 , \19586_nG9be1 );
and \U$14092 ( \23225 , \12154 , \20608_nG9bde );
or \U$14093 ( \23226 , \23224 , \23225 );
xor \U$14094 ( \23227 , \12153 , \23226 );
buf \U$14095 ( \23228 , \23227 );
buf \U$14097 ( \23229 , \23228 );
xor \U$14098 ( \23230 , \23223 , \23229 );
and \U$14099 ( \23231 , \10421 , \21086_nG9bdb );
and \U$14100 ( \23232 , \10418 , \22129_nG9bd8 );
or \U$14101 ( \23233 , \23231 , \23232 );
xor \U$14102 ( \23234 , \10417 , \23233 );
buf \U$14103 ( \23235 , \23234 );
buf \U$14105 ( \23236 , \23235 );
xor \U$14106 ( \23237 , \23230 , \23236 );
buf \U$14107 ( \23238 , \23237 );
xor \U$14108 ( \23239 , \23218 , \23238 );
and \U$14109 ( \23240 , \22249 , \22254 );
and \U$14110 ( \23241 , \22249 , \22634 );
and \U$14111 ( \23242 , \22254 , \22634 );
or \U$14112 ( \23243 , \23240 , \23241 , \23242 );
buf \U$14113 ( \23244 , \23243 );
xor \U$14114 ( \23245 , \23239 , \23244 );
buf \U$14115 ( \23246 , \23245 );
and \U$14116 ( \23247 , \22155 , \22190 );
and \U$14117 ( \23248 , \22155 , \22242 );
and \U$14118 ( \23249 , \22190 , \22242 );
or \U$14119 ( \23250 , \23247 , \23248 , \23249 );
buf \U$14120 ( \23251 , \23250 );
xor \U$14121 ( \23252 , \23246 , \23251 );
and \U$14122 ( \23253 , \22160 , \22166 );
and \U$14123 ( \23254 , \22160 , \22173 );
and \U$14124 ( \23255 , \22166 , \22173 );
or \U$14125 ( \23256 , \23253 , \23254 , \23255 );
buf \U$14126 ( \23257 , \23256 );
and \U$14127 ( \23258 , \22207 , \22213 );
and \U$14128 ( \23259 , \22207 , \22220 );
and \U$14129 ( \23260 , \22213 , \22220 );
or \U$14130 ( \23261 , \23258 , \23259 , \23260 );
buf \U$14131 ( \23262 , \23261 );
and \U$14132 ( \23263 , \21658 , \10995_nG9c0b );
and \U$14133 ( \23264 , \21655 , \11283_nG9c08 );
or \U$14134 ( \23265 , \23263 , \23264 );
xor \U$14135 ( \23266 , \21654 , \23265 );
buf \U$14136 ( \23267 , \23266 );
buf \U$14138 ( \23268 , \23267 );
and \U$14139 ( \23269 , \20155 , \11598_nG9c05 );
and \U$14140 ( \23270 , \20152 , \12470_nG9c02 );
or \U$14141 ( \23271 , \23269 , \23270 );
xor \U$14142 ( \23272 , \20151 , \23271 );
buf \U$14143 ( \23273 , \23272 );
buf \U$14145 ( \23274 , \23273 );
xor \U$14146 ( \23275 , \23268 , \23274 );
buf \U$14147 ( \23276 , \23275 );
xor \U$14148 ( \23277 , \23262 , \23276 );
and \U$14149 ( \23278 , \15940 , \15373_nG9bf3 );
and \U$14150 ( \23279 , \15937 , \16315_nG9bf0 );
or \U$14151 ( \23280 , \23278 , \23279 );
xor \U$14152 ( \23281 , \15936 , \23280 );
buf \U$14153 ( \23282 , \23281 );
buf \U$14155 ( \23283 , \23282 );
xor \U$14156 ( \23284 , \23277 , \23283 );
buf \U$14157 ( \23285 , \23284 );
xor \U$14158 ( \23286 , \23257 , \23285 );
and \U$14159 ( \23287 , \22222 , \22224 );
and \U$14160 ( \23288 , \22222 , \22231 );
and \U$14161 ( \23289 , \22224 , \22231 );
or \U$14162 ( \23290 , \23287 , \23288 , \23289 );
buf \U$14163 ( \23291 , \23290 );
xor \U$14164 ( \23292 , \23286 , \23291 );
buf \U$14165 ( \23293 , \23292 );
and \U$14166 ( \23294 , \22199 , \22205 );
buf \U$14167 ( \23295 , \23294 );
and \U$14168 ( \23296 , \18702 , \12801_nG9bff );
and \U$14169 ( \23297 , \18699 , \13705_nG9bfc );
or \U$14170 ( \23298 , \23296 , \23297 );
xor \U$14171 ( \23299 , \18698 , \23298 );
buf \U$14172 ( \23300 , \23299 );
buf \U$14174 ( \23301 , \23300 );
xor \U$14175 ( \23302 , \23295 , \23301 );
and \U$14176 ( \23303 , \17297 , \14070_nG9bf9 );
and \U$14177 ( \23304 , \17294 , \14984_nG9bf6 );
or \U$14178 ( \23305 , \23303 , \23304 );
xor \U$14179 ( \23306 , \17293 , \23305 );
buf \U$14180 ( \23307 , \23306 );
buf \U$14182 ( \23308 , \23307 );
xor \U$14183 ( \23309 , \23302 , \23308 );
buf \U$14184 ( \23310 , \23309 );
and \U$14185 ( \23311 , \14631 , \16680_nG9bed );
and \U$14186 ( \23312 , \14628 , \17665_nG9bea );
or \U$14187 ( \23313 , \23311 , \23312 );
xor \U$14188 ( \23314 , \14627 , \23313 );
buf \U$14189 ( \23315 , \23314 );
buf \U$14191 ( \23316 , \23315 );
xor \U$14192 ( \23317 , \23310 , \23316 );
and \U$14193 ( \23318 , \13370 , \18107_nG9be7 );
and \U$14194 ( \23319 , \13367 , \19091_nG9be4 );
or \U$14195 ( \23320 , \23318 , \23319 );
xor \U$14196 ( \23321 , \13366 , \23320 );
buf \U$14197 ( \23322 , \23321 );
buf \U$14199 ( \23323 , \23322 );
xor \U$14200 ( \23324 , \23317 , \23323 );
buf \U$14201 ( \23325 , \23324 );
xor \U$14202 ( \23326 , \23293 , \23325 );
and \U$14203 ( \23327 , \10707 , \22629_nG9bd5 );
and \U$14204 ( \23328 , \22264 , \22550 );
and \U$14205 ( \23329 , \22550 , \22572 );
and \U$14206 ( \23330 , \22264 , \22572 );
or \U$14207 ( \23331 , \23328 , \23329 , \23330 );
and \U$14208 ( \23332 , \22578 , \22582 );
and \U$14209 ( \23333 , \22582 , \22617 );
and \U$14210 ( \23334 , \22578 , \22617 );
or \U$14211 ( \23335 , \23332 , \23333 , \23334 );
xor \U$14212 ( \23336 , \23331 , \23335 );
and \U$14213 ( \23337 , \22268 , \22272 );
and \U$14214 ( \23338 , \22272 , \22549 );
and \U$14215 ( \23339 , \22268 , \22549 );
or \U$14216 ( \23340 , \23337 , \23338 , \23339 );
and \U$14217 ( \23341 , \22591 , \22595 );
and \U$14218 ( \23342 , \22595 , \22600 );
and \U$14219 ( \23343 , \22591 , \22600 );
or \U$14220 ( \23344 , \23341 , \23342 , \23343 );
xor \U$14221 ( \23345 , \23340 , \23344 );
and \U$14222 ( \23346 , \22606 , \22610 );
and \U$14223 ( \23347 , \22610 , \22615 );
and \U$14224 ( \23348 , \22606 , \22615 );
or \U$14225 ( \23349 , \23346 , \23347 , \23348 );
xor \U$14226 ( \23350 , \23345 , \23349 );
and \U$14227 ( \23351 , \22556 , \10983 );
and \U$14228 ( \23352 , RIdec5270_707, \9333 );
and \U$14229 ( \23353 , RIdec2570_675, \9335 );
and \U$14230 ( \23354 , RIee1ff18_4822, \9337 );
and \U$14231 ( \23355 , RIdebf870_643, \9339 );
and \U$14232 ( \23356 , RIfe7f848_7795, \9341 );
and \U$14233 ( \23357 , RIdebcb70_611, \9343 );
and \U$14234 ( \23358 , RIdeb9e70_579, \9345 );
and \U$14235 ( \23359 , RIdeb7170_547, \9347 );
and \U$14236 ( \23360 , RIfe7fc80_7798, \9349 );
and \U$14237 ( \23361 , RIdeb1770_483, \9351 );
and \U$14238 ( \23362 , RIfca5d58_6909, \9353 );
and \U$14239 ( \23363 , RIdeaea70_451, \9355 );
and \U$14240 ( \23364 , RIfcaf808_7019, \9357 );
and \U$14241 ( \23365 , RIdeaa0d8_419, \9359 );
and \U$14242 ( \23366 , RIdea37d8_387, \9361 );
and \U$14243 ( \23367 , RIde9ced8_355, \9363 );
and \U$14244 ( \23368 , RIfcdc3d0_7528, \9365 );
and \U$14245 ( \23369 , RIfcce438_7369, \9367 );
and \U$14246 ( \23370 , RIfcb0a50_7032, \9369 );
and \U$14247 ( \23371 , RIfc75680_6358, \9371 );
and \U$14248 ( \23372 , RIde90d40_296, \9373 );
and \U$14249 ( \23373 , RIfe7f9b0_7796, \9375 );
and \U$14250 ( \23374 , RIde89720_260, \9377 );
and \U$14251 ( \23375 , RIde85580_240, \9379 );
and \U$14252 ( \23376 , RIde81728_221, \9381 );
and \U$14253 ( \23377 , RIfc52f40_5966, \9383 );
and \U$14254 ( \23378 , RIfc82100_6502, \9385 );
and \U$14255 ( \23379 , RIfca7108_6923, \9387 );
and \U$14256 ( \23380 , RIfe7fb18_7797, \9389 );
and \U$14257 ( \23381 , RIe16b648_2599, \9391 );
and \U$14258 ( \23382 , RIe169a28_2579, \9393 );
and \U$14259 ( \23383 , RIe167ca0_2558, \9395 );
and \U$14260 ( \23384 , RIe165270_2528, \9397 );
and \U$14261 ( \23385 , RIe162570_2496, \9399 );
and \U$14262 ( \23386 , RIee37258_5086, \9401 );
and \U$14263 ( \23387 , RIe15f870_2464, \9403 );
and \U$14264 ( \23388 , RIee36178_5074, \9405 );
and \U$14265 ( \23389 , RIe15cb70_2432, \9407 );
and \U$14266 ( \23390 , RIe157170_2368, \9409 );
and \U$14267 ( \23391 , RIe154470_2336, \9411 );
and \U$14268 ( \23392 , RIfc86fc0_6558, \9413 );
and \U$14269 ( \23393 , RIe151770_2304, \9415 );
and \U$14270 ( \23394 , RIfc4eff8_5921, \9417 );
and \U$14271 ( \23395 , RIe14ea70_2272, \9419 );
and \U$14272 ( \23396 , RIfce1290_7584, \9421 );
and \U$14273 ( \23397 , RIe14bd70_2240, \9423 );
and \U$14274 ( \23398 , RIe149070_2208, \9425 );
and \U$14275 ( \23399 , RIe146370_2176, \9427 );
and \U$14276 ( \23400 , RIee34558_5054, \9429 );
and \U$14277 ( \23401 , RIee331a8_5040, \9431 );
and \U$14278 ( \23402 , RIee320c8_5028, \9433 );
and \U$14279 ( \23403 , RIee31150_5017, \9435 );
and \U$14280 ( \23404 , RIfe800b8_7801, \9437 );
and \U$14281 ( \23405 , RIfe7ff50_7800, \9439 );
and \U$14282 ( \23406 , RIdf3caf0_2067, \9441 );
and \U$14283 ( \23407 , RIfe7fde8_7799, \9443 );
and \U$14284 ( \23408 , RIfcc8330_7300, \9445 );
and \U$14285 ( \23409 , RIee2f800_4999, \9447 );
and \U$14286 ( \23410 , RIfca0d30_6852, \9449 );
and \U$14287 ( \23411 , RIee2d640_4975, \9451 );
and \U$14288 ( \23412 , RIdf35638_1984, \9453 );
and \U$14289 ( \23413 , RIdf331a8_1958, \9455 );
and \U$14290 ( \23414 , RIdf31150_1935, \9457 );
and \U$14291 ( \23415 , RIdf2ef90_1911, \9459 );
or \U$14292 ( \23416 , \23352 , \23353 , \23354 , \23355 , \23356 , \23357 , \23358 , \23359 , \23360 , \23361 , \23362 , \23363 , \23364 , \23365 , \23366 , \23367 , \23368 , \23369 , \23370 , \23371 , \23372 , \23373 , \23374 , \23375 , \23376 , \23377 , \23378 , \23379 , \23380 , \23381 , \23382 , \23383 , \23384 , \23385 , \23386 , \23387 , \23388 , \23389 , \23390 , \23391 , \23392 , \23393 , \23394 , \23395 , \23396 , \23397 , \23398 , \23399 , \23400 , \23401 , \23402 , \23403 , \23404 , \23405 , \23406 , \23407 , \23408 , \23409 , \23410 , \23411 , \23412 , \23413 , \23414 , \23415 );
and \U$14293 ( \23417 , RIee2bb88_4956, \9462 );
and \U$14294 ( \23418 , RIee2a0d0_4937, \9464 );
and \U$14295 ( \23419 , RIee28d20_4923, \9466 );
and \U$14296 ( \23420 , RIfe7f578_7793, \9468 );
and \U$14297 ( \23421 , RIdf2a238_1856, \9470 );
and \U$14298 ( \23422 , RIdf27f10_1831, \9472 );
and \U$14299 ( \23423 , RIfe7f6e0_7794, \9474 );
and \U$14300 ( \23424 , RIdf246d0_1791, \9476 );
and \U$14301 ( \23425 , RIfcce9d8_7373, \9478 );
and \U$14302 ( \23426 , RIfc63638_6153, \9480 );
and \U$14303 ( \23427 , RIdf22c18_1772, \9482 );
and \U$14304 ( \23428 , RIfc62990_6144, \9484 );
and \U$14305 ( \23429 , RIdf21700_1757, \9486 );
and \U$14306 ( \23430 , RIdf1f810_1735, \9488 );
and \U$14307 ( \23431 , RIfeaa958_8257, \9490 );
and \U$14308 ( \23432 , RIdf19168_1662, \9492 );
and \U$14309 ( \23433 , RIdf16e40_1637, \9494 );
and \U$14310 ( \23434 , RIdf14140_1605, \9496 );
and \U$14311 ( \23435 , RIdf11440_1573, \9498 );
and \U$14312 ( \23436 , RIdf0e740_1541, \9500 );
and \U$14313 ( \23437 , RIdf0ba40_1509, \9502 );
and \U$14314 ( \23438 , RIdf08d40_1477, \9504 );
and \U$14315 ( \23439 , RIdf06040_1445, \9506 );
and \U$14316 ( \23440 , RIdf03340_1413, \9508 );
and \U$14317 ( \23441 , RIdefd940_1349, \9510 );
and \U$14318 ( \23442 , RIdefac40_1317, \9512 );
and \U$14319 ( \23443 , RIdef7f40_1285, \9514 );
and \U$14320 ( \23444 , RIdef5240_1253, \9516 );
and \U$14321 ( \23445 , RIdef2540_1221, \9518 );
and \U$14322 ( \23446 , RIdeef840_1189, \9520 );
and \U$14323 ( \23447 , RIdeecb40_1157, \9522 );
and \U$14324 ( \23448 , RIdee9e40_1125, \9524 );
and \U$14325 ( \23449 , RIfcb7800_7110, \9526 );
and \U$14326 ( \23450 , RIee24838_4874, \9528 );
and \U$14327 ( \23451 , RIfc4cb68_5895, \9530 );
and \U$14328 ( \23452 , RIee23320_4859, \9532 );
and \U$14329 ( \23453 , RIfe80388_7803, \9534 );
and \U$14330 ( \23454 , RIdee2c58_1044, \9536 );
and \U$14331 ( \23455 , RIfe80220_7802, \9538 );
and \U$14332 ( \23456 , RIdedea40_997, \9540 );
and \U$14333 ( \23457 , RIfc98900_6758, \9542 );
and \U$14334 ( \23458 , RIee223a8_4848, \9544 );
and \U$14335 ( \23459 , RIfcc8600_7302, \9546 );
and \U$14336 ( \23460 , RIee212c8_4836, \9548 );
and \U$14337 ( \23461 , RIded9748_938, \9550 );
and \U$14338 ( \23462 , RIfe804f0_7804, \9552 );
and \U$14339 ( \23463 , RIded53c8_890, \9554 );
and \U$14340 ( \23464 , RIded2c68_862, \9556 );
and \U$14341 ( \23465 , RIded0670_835, \9558 );
and \U$14342 ( \23466 , RIdecd970_803, \9560 );
and \U$14343 ( \23467 , RIdecac70_771, \9562 );
and \U$14344 ( \23468 , RIdec7f70_739, \9564 );
and \U$14345 ( \23469 , RIdeb4470_515, \9566 );
and \U$14346 ( \23470 , RIde965d8_323, \9568 );
and \U$14347 ( \23471 , RIe16e078_2629, \9570 );
and \U$14348 ( \23472 , RIe159e70_2400, \9572 );
and \U$14349 ( \23473 , RIe143670_2144, \9574 );
and \U$14350 ( \23474 , RIdf38068_2014, \9576 );
and \U$14351 ( \23475 , RIdf2c6c8_1882, \9578 );
and \U$14352 ( \23476 , RIdf1cf48_1706, \9580 );
and \U$14353 ( \23477 , RIdf00640_1381, \9582 );
and \U$14354 ( \23478 , RIdee7140_1093, \9584 );
and \U$14355 ( \23479 , RIdedbea8_966, \9586 );
and \U$14356 ( \23480 , RIde7c520_196, \9588 );
or \U$14357 ( \23481 , \23417 , \23418 , \23419 , \23420 , \23421 , \23422 , \23423 , \23424 , \23425 , \23426 , \23427 , \23428 , \23429 , \23430 , \23431 , \23432 , \23433 , \23434 , \23435 , \23436 , \23437 , \23438 , \23439 , \23440 , \23441 , \23442 , \23443 , \23444 , \23445 , \23446 , \23447 , \23448 , \23449 , \23450 , \23451 , \23452 , \23453 , \23454 , \23455 , \23456 , \23457 , \23458 , \23459 , \23460 , \23461 , \23462 , \23463 , \23464 , \23465 , \23466 , \23467 , \23468 , \23469 , \23470 , \23471 , \23472 , \23473 , \23474 , \23475 , \23476 , \23477 , \23478 , \23479 , \23480 );
or \U$14358 ( \23482 , \23416 , \23481 );
_DC g65b3 ( \23483_nG65b3 , \23482 , \9597 );
and \U$14359 ( \23484 , RIe19d508_3167, \9059 );
and \U$14360 ( \23485 , RIe19a808_3135, \9061 );
and \U$14361 ( \23486 , RIfe7ee70_7788, \9063 );
and \U$14362 ( \23487 , RIe197b08_3103, \9065 );
and \U$14363 ( \23488 , RIfe7efd8_7789, \9067 );
and \U$14364 ( \23489 , RIe194e08_3071, \9069 );
and \U$14365 ( \23490 , RIe192108_3039, \9071 );
and \U$14366 ( \23491 , RIe18f408_3007, \9073 );
and \U$14367 ( \23492 , RIe189a08_2943, \9075 );
and \U$14368 ( \23493 , RIe186d08_2911, \9077 );
and \U$14369 ( \23494 , RIf143768_5227, \9079 );
and \U$14370 ( \23495 , RIe184008_2879, \9081 );
and \U$14371 ( \23496 , RIfc4bbf0_5884, \9083 );
and \U$14372 ( \23497 , RIe181308_2847, \9085 );
and \U$14373 ( \23498 , RIe17e608_2815, \9087 );
and \U$14374 ( \23499 , RIe17b908_2783, \9089 );
and \U$14375 ( \23500 , RIfe7f410_7792, \9091 );
and \U$14376 ( \23501 , RIf140d38_5197, \9093 );
and \U$14377 ( \23502 , RIe176fe8_2731, \9095 );
and \U$14378 ( \23503 , RIe175ad0_2716, \9097 );
and \U$14379 ( \23504 , RIfe7f2a8_7791, \9099 );
and \U$14380 ( \23505 , RIf13f118_5177, \9101 );
and \U$14381 ( \23506 , RIee3e440_5167, \9103 );
and \U$14382 ( \23507 , RIee3d360_5155, \9105 );
and \U$14383 ( \23508 , RIee3c280_5143, \9107 );
and \U$14384 ( \23509 , RIee3b1a0_5131, \9109 );
and \U$14385 ( \23510 , RIfe7f140_7790, \9111 );
and \U$14386 ( \23511 , RIe173640_2690, \9113 );
and \U$14387 ( \23512 , RIf170330_5736, \9115 );
and \U$14388 ( \23513 , RIf16f520_5726, \9117 );
and \U$14389 ( \23514 , RIf16e2d8_5713, \9119 );
and \U$14390 ( \23515 , RIf16d630_5704, \9121 );
and \U$14391 ( \23516 , RIfe7ea38_7785, \9123 );
and \U$14392 ( \23517 , RIe223860_4694, \9125 );
and \U$14393 ( \23518 , RIfc9c410_6800, \9127 );
and \U$14394 ( \23519 , RIe220b60_4662, \9129 );
and \U$14395 ( \23520 , RIfcb8340_7118, \9131 );
and \U$14396 ( \23521 , RIe21de60_4630, \9133 );
and \U$14397 ( \23522 , RIe218460_4566, \9135 );
and \U$14398 ( \23523 , RIe215760_4534, \9137 );
and \U$14399 ( \23524 , RIfc9cc80_6806, \9139 );
and \U$14400 ( \23525 , RIe212a60_4502, \9141 );
and \U$14401 ( \23526 , RIfc4ddb0_5908, \9143 );
and \U$14402 ( \23527 , RIe20fd60_4470, \9145 );
and \U$14403 ( \23528 , RIfc873f8_6561, \9147 );
and \U$14404 ( \23529 , RIe20d060_4438, \9149 );
and \U$14405 ( \23530 , RIe20a360_4406, \9151 );
and \U$14406 ( \23531 , RIe207660_4374, \9153 );
and \U$14407 ( \23532 , RIfc86750_6552, \9155 );
and \U$14408 ( \23533 , RIfc4e4b8_5913, \9157 );
and \U$14409 ( \23534 , RIe202368_4315, \9159 );
and \U$14410 ( \23535 , RIe200a18_4297, \9161 );
and \U$14411 ( \23536 , RIf165200_5610, \9163 );
and \U$14412 ( \23537 , RIf164558_5601, \9165 );
and \U$14413 ( \23538 , RIf163478_5589, \9167 );
and \U$14414 ( \23539 , RIf161f60_5574, \9169 );
and \U$14415 ( \23540 , RIf160070_5552, \9171 );
and \U$14416 ( \23541 , RIf15e180_5530, \9173 );
and \U$14417 ( \23542 , RIe1fcc38_4253, \9175 );
and \U$14418 ( \23543 , RIe1fb9f0_4240, \9177 );
and \U$14419 ( \23544 , RIf15cc68_5515, \9179 );
and \U$14420 ( \23545 , RIf15b750_5500, \9181 );
and \U$14421 ( \23546 , RIf15a670_5488, \9183 );
and \U$14422 ( \23547 , RIf159c98_5481, \9185 );
or \U$14423 ( \23548 , \23484 , \23485 , \23486 , \23487 , \23488 , \23489 , \23490 , \23491 , \23492 , \23493 , \23494 , \23495 , \23496 , \23497 , \23498 , \23499 , \23500 , \23501 , \23502 , \23503 , \23504 , \23505 , \23506 , \23507 , \23508 , \23509 , \23510 , \23511 , \23512 , \23513 , \23514 , \23515 , \23516 , \23517 , \23518 , \23519 , \23520 , \23521 , \23522 , \23523 , \23524 , \23525 , \23526 , \23527 , \23528 , \23529 , \23530 , \23531 , \23532 , \23533 , \23534 , \23535 , \23536 , \23537 , \23538 , \23539 , \23540 , \23541 , \23542 , \23543 , \23544 , \23545 , \23546 , \23547 );
and \U$14424 ( \23549 , RIf158e88_5471, \9188 );
and \U$14425 ( \23550 , RIf157ad8_5457, \9190 );
and \U$14426 ( \23551 , RIf156e30_5448, \9192 );
and \U$14427 ( \23552 , RIfe7e768_7783, \9194 );
and \U$14428 ( \23553 , RIf1562f0_5440, \9196 );
and \U$14429 ( \23554 , RIf1557b0_5432, \9198 );
and \U$14430 ( \23555 , RIf154838_5421, \9200 );
and \U$14431 ( \23556 , RIfe7e8d0_7784, \9202 );
and \U$14432 ( \23557 , RIf1531b8_5405, \9204 );
and \U$14433 ( \23558 , RIfc52400_5958, \9206 );
and \U$14434 ( \23559 , RIf150a58_5377, \9208 );
and \U$14435 ( \23560 , RIe1f3188_4143, \9210 );
and \U$14436 ( \23561 , RIf14f978_5365, \9212 );
and \U$14437 ( \23562 , RIf14ecd0_5356, \9214 );
and \U$14438 ( \23563 , RIf14dec0_5346, \9216 );
and \U$14439 ( \23564 , RIe1ede90_4084, \9218 );
and \U$14440 ( \23565 , RIe1eb5c8_4055, \9220 );
and \U$14441 ( \23566 , RIe1e88c8_4023, \9222 );
and \U$14442 ( \23567 , RIe1e5bc8_3991, \9224 );
and \U$14443 ( \23568 , RIe1e2ec8_3959, \9226 );
and \U$14444 ( \23569 , RIe1e01c8_3927, \9228 );
and \U$14445 ( \23570 , RIe1dd4c8_3895, \9230 );
and \U$14446 ( \23571 , RIe1da7c8_3863, \9232 );
and \U$14447 ( \23572 , RIe1d7ac8_3831, \9234 );
and \U$14448 ( \23573 , RIe1d20c8_3767, \9236 );
and \U$14449 ( \23574 , RIe1cf3c8_3735, \9238 );
and \U$14450 ( \23575 , RIe1cc6c8_3703, \9240 );
and \U$14451 ( \23576 , RIe1c99c8_3671, \9242 );
and \U$14452 ( \23577 , RIe1c6cc8_3639, \9244 );
and \U$14453 ( \23578 , RIe1c3fc8_3607, \9246 );
and \U$14454 ( \23579 , RIe1c12c8_3575, \9248 );
and \U$14455 ( \23580 , RIe1be5c8_3543, \9250 );
and \U$14456 ( \23581 , RIf14c9a8_5331, \9252 );
and \U$14457 ( \23582 , RIf14b760_5318, \9254 );
and \U$14458 ( \23583 , RIfe7ed08_7787, \9256 );
and \U$14459 ( \23584 , RIfe7e600_7782, \9258 );
and \U$14460 ( \23585 , RIf14a518_5305, \9260 );
and \U$14461 ( \23586 , RIfca1f78_6865, \9262 );
and \U$14462 ( \23587 , RIfe7eba0_7786, \9264 );
and \U$14463 ( \23588 , RIfe7e498_7781, \9266 );
and \U$14464 ( \23589 , RIf148e98_5289, \9268 );
and \U$14465 ( \23590 , RIf147c50_5276, \9270 );
and \U$14466 ( \23591 , RIfe7e330_7780, \9272 );
and \U$14467 ( \23592 , RIe1b0a68_3387, \9274 );
and \U$14468 ( \23593 , RIf147278_5269, \9276 );
and \U$14469 ( \23594 , RIf1465d0_5260, \9278 );
and \U$14470 ( \23595 , RIe1ac418_3337, \9280 );
and \U$14471 ( \23596 , RIe1aac30_3320, \9282 );
and \U$14472 ( \23597 , RIe1a8908_3295, \9284 );
and \U$14473 ( \23598 , RIe1a5c08_3263, \9286 );
and \U$14474 ( \23599 , RIe1a2f08_3231, \9288 );
and \U$14475 ( \23600 , RIe1a0208_3199, \9290 );
and \U$14476 ( \23601 , RIe18c708_2975, \9292 );
and \U$14477 ( \23602 , RIe178c08_2751, \9294 );
and \U$14478 ( \23603 , RIe226560_4726, \9296 );
and \U$14479 ( \23604 , RIe21b160_4598, \9298 );
and \U$14480 ( \23605 , RIe204960_4342, \9300 );
and \U$14481 ( \23606 , RIe1fe9c0_4274, \9302 );
and \U$14482 ( \23607 , RIe1f7d78_4197, \9304 );
and \U$14483 ( \23608 , RIe1f08c0_4114, \9306 );
and \U$14484 ( \23609 , RIe1d4dc8_3799, \9308 );
and \U$14485 ( \23610 , RIe1bb8c8_3511, \9310 );
and \U$14486 ( \23611 , RIe1ae740_3362, \9312 );
and \U$14487 ( \23612 , RIe170d78_2661, \9314 );
or \U$14488 ( \23613 , \23549 , \23550 , \23551 , \23552 , \23553 , \23554 , \23555 , \23556 , \23557 , \23558 , \23559 , \23560 , \23561 , \23562 , \23563 , \23564 , \23565 , \23566 , \23567 , \23568 , \23569 , \23570 , \23571 , \23572 , \23573 , \23574 , \23575 , \23576 , \23577 , \23578 , \23579 , \23580 , \23581 , \23582 , \23583 , \23584 , \23585 , \23586 , \23587 , \23588 , \23589 , \23590 , \23591 , \23592 , \23593 , \23594 , \23595 , \23596 , \23597 , \23598 , \23599 , \23600 , \23601 , \23602 , \23603 , \23604 , \23605 , \23606 , \23607 , \23608 , \23609 , \23610 , \23611 , \23612 );
or \U$14489 ( \23614 , \23548 , \23613 );
_DC g65b4 ( \23615_nG65b4 , \23614 , \9323 );
and g65b5 ( \23616_nG65b5 , \23483_nG65b3 , \23615_nG65b4 );
buf \U$14490 ( \23617 , \23616_nG65b5 );
and \U$14491 ( \23618 , \23617 , \10691 );
nor \U$14492 ( \23619 , \23351 , \23618 );
xnor \U$14493 ( \23620 , \23619 , \10980 );
and \U$14494 ( \23621 , \18035 , \14054 );
and \U$14495 ( \23622 , \19032 , \13692 );
nor \U$14496 ( \23623 , \23621 , \23622 );
xnor \U$14497 ( \23624 , \23623 , \14035 );
xor \U$14498 ( \23625 , \23620 , \23624 );
_DC g598e ( \23626_nG598e , \23482 , \9597 );
_DC g5a12 ( \23627_nG5a12 , \23614 , \9323 );
xor g5a13 ( \23628_nG5a13 , \23626_nG598e , \23627_nG5a12 );
buf \U$14499 ( \23629 , \23628_nG5a13 );
xor \U$14500 ( \23630 , \23629 , \22539 );
and \U$14501 ( \23631 , \10687 , \23630 );
xor \U$14502 ( \23632 , \23625 , \23631 );
and \U$14503 ( \23633 , \19558 , \12790 );
and \U$14504 ( \23634 , \20544 , \12461 );
nor \U$14505 ( \23635 , \23633 , \23634 );
xnor \U$14506 ( \23636 , \23635 , \12780 );
and \U$14507 ( \23637 , \16655 , \15336 );
and \U$14508 ( \23638 , \17627 , \14963 );
nor \U$14509 ( \23639 , \23637 , \23638 );
xnor \U$14510 ( \23640 , \23639 , \15342 );
xor \U$14511 ( \23641 , \23636 , \23640 );
and \U$14512 ( \23642 , \10988 , \22542 );
and \U$14513 ( \23643 , \11270 , \22103 );
nor \U$14514 ( \23644 , \23642 , \23643 );
xnor \U$14515 ( \23645 , \23644 , \22548 );
xor \U$14516 ( \23646 , \23641 , \23645 );
xor \U$14517 ( \23647 , \23632 , \23646 );
and \U$14518 ( \23648 , \21033 , \11574 );
and \U$14519 ( \23649 , \22090 , \11278 );
nor \U$14520 ( \23650 , \23648 , \23649 );
xnor \U$14521 ( \23651 , \23650 , \11580 );
and \U$14522 ( \23652 , \12769 , \19534 );
and \U$14523 ( \23653 , \13679 , \19045 );
nor \U$14524 ( \23654 , \23652 , \23653 );
xnor \U$14525 ( \23655 , \23654 , \19540 );
xor \U$14526 ( \23656 , \23651 , \23655 );
and \U$14527 ( \23657 , \11586 , \21005 );
and \U$14528 ( \23658 , \12448 , \20557 );
nor \U$14529 ( \23659 , \23657 , \23658 );
xnor \U$14530 ( \23660 , \23659 , \21011 );
xor \U$14531 ( \23661 , \23656 , \23660 );
xor \U$14532 ( \23662 , \23647 , \23661 );
xor \U$14533 ( \23663 , \23350 , \23662 );
and \U$14534 ( \23664 , \22562 , \22566 );
and \U$14535 ( \23665 , \22566 , \22571 );
and \U$14536 ( \23666 , \22562 , \22571 );
or \U$14537 ( \23667 , \23664 , \23665 , \23666 );
and \U$14538 ( \23668 , \22587 , \22601 );
and \U$14539 ( \23669 , \22601 , \22616 );
and \U$14540 ( \23670 , \22587 , \22616 );
or \U$14541 ( \23671 , \23668 , \23669 , \23670 );
xor \U$14542 ( \23672 , \23667 , \23671 );
and \U$14543 ( \23673 , \22559 , \22561 );
and \U$14544 ( \23674 , \15321 , \16635 );
and \U$14545 ( \23675 , \16267 , \16301 );
nor \U$14546 ( \23676 , \23674 , \23675 );
xnor \U$14547 ( \23677 , \23676 , \16625 );
xor \U$14548 ( \23678 , \23673 , \23677 );
and \U$14549 ( \23679 , \14024 , \18090 );
and \U$14550 ( \23680 , \14950 , \17655 );
nor \U$14551 ( \23681 , \23679 , \23680 );
xnor \U$14552 ( \23682 , \23681 , \18046 );
xor \U$14553 ( \23683 , \23678 , \23682 );
xor \U$14554 ( \23684 , \23672 , \23683 );
xor \U$14555 ( \23685 , \23663 , \23684 );
xor \U$14556 ( \23686 , \23336 , \23685 );
and \U$14557 ( \23687 , \22260 , \22573 );
and \U$14558 ( \23688 , \22573 , \22618 );
and \U$14559 ( \23689 , \22260 , \22618 );
or \U$14560 ( \23690 , \23687 , \23688 , \23689 );
xor \U$14561 ( \23691 , \23686 , \23690 );
and \U$14562 ( \23692 , \22619 , \22623 );
and \U$14563 ( \23693 , \22624 , \22627 );
or \U$14564 ( \23694 , \23692 , \23693 );
xor \U$14565 ( \23695 , \23691 , \23694 );
buf g9bd2 ( \23696_nG9bd2 , \23695 );
and \U$14566 ( \23697 , \10704 , \23696_nG9bd2 );
or \U$14567 ( \23698 , \23327 , \23697 );
xor \U$14568 ( \23699 , \10703 , \23698 );
buf \U$14569 ( \23700 , \23699 );
buf \U$14571 ( \23701 , \23700 );
xor \U$14572 ( \23702 , \23326 , \23701 );
buf \U$14573 ( \23703 , \23702 );
xor \U$14574 ( \23704 , \23252 , \23703 );
and \U$14575 ( \23705 , \23208 , \23704 );
and \U$14576 ( \23706 , \23212 , \23704 );
or \U$14577 ( \23707 , \23213 , \23705 , \23706 );
and \U$14578 ( \23708 , \22644 , \22648 );
and \U$14579 ( \23709 , \22644 , \23207 );
and \U$14580 ( \23710 , \22648 , \23207 );
or \U$14581 ( \23711 , \23708 , \23709 , \23710 );
xor \U$14582 ( \23712 , \23707 , \23711 );
and \U$14583 ( \23713 , \23246 , \23251 );
and \U$14584 ( \23714 , \23246 , \23703 );
and \U$14585 ( \23715 , \23251 , \23703 );
or \U$14586 ( \23716 , \23713 , \23714 , \23715 );
xor \U$14587 ( \23717 , \23712 , \23716 );
and \U$14588 ( \23718 , \23310 , \23316 );
and \U$14589 ( \23719 , \23310 , \23323 );
and \U$14590 ( \23720 , \23316 , \23323 );
or \U$14591 ( \23721 , \23718 , \23719 , \23720 );
buf \U$14592 ( \23722 , \23721 );
and \U$14593 ( \23723 , \23257 , \23285 );
and \U$14594 ( \23724 , \23257 , \23291 );
and \U$14595 ( \23725 , \23285 , \23291 );
or \U$14596 ( \23726 , \23723 , \23724 , \23725 );
buf \U$14597 ( \23727 , \23726 );
xor \U$14598 ( \23728 , \23722 , \23727 );
and \U$14599 ( \23729 , \10421 , \22129_nG9bd8 );
and \U$14600 ( \23730 , \10418 , \22629_nG9bd5 );
or \U$14601 ( \23731 , \23729 , \23730 );
xor \U$14602 ( \23732 , \10417 , \23731 );
buf \U$14603 ( \23733 , \23732 );
buf \U$14605 ( \23734 , \23733 );
xor \U$14606 ( \23735 , \23728 , \23734 );
buf \U$14607 ( \23736 , \23735 );
and \U$14608 ( \23737 , \23293 , \23325 );
and \U$14609 ( \23738 , \23293 , \23701 );
and \U$14610 ( \23739 , \23325 , \23701 );
or \U$14611 ( \23740 , \23737 , \23738 , \23739 );
buf \U$14612 ( \23741 , \23740 );
xor \U$14613 ( \23742 , \23736 , \23741 );
and \U$14614 ( \23743 , \23223 , \23229 );
and \U$14615 ( \23744 , \23223 , \23236 );
and \U$14616 ( \23745 , \23229 , \23236 );
or \U$14617 ( \23746 , \23743 , \23744 , \23745 );
buf \U$14618 ( \23747 , \23746 );
xor \U$14619 ( \23748 , \23742 , \23747 );
buf \U$14620 ( \23749 , \23748 );
and \U$14621 ( \23750 , \23218 , \23238 );
and \U$14622 ( \23751 , \23218 , \23244 );
and \U$14623 ( \23752 , \23238 , \23244 );
or \U$14624 ( \23753 , \23750 , \23751 , \23752 );
buf \U$14625 ( \23754 , \23753 );
xor \U$14626 ( \23755 , \23749 , \23754 );
and \U$14627 ( \23756 , \23262 , \23276 );
and \U$14628 ( \23757 , \23262 , \23283 );
and \U$14629 ( \23758 , \23276 , \23283 );
or \U$14630 ( \23759 , \23756 , \23757 , \23758 );
buf \U$14631 ( \23760 , \23759 );
and \U$14632 ( \23761 , \23268 , \23274 );
buf \U$14633 ( \23762 , \23761 );
and \U$14634 ( \23763 , \18702 , \13705_nG9bfc );
and \U$14635 ( \23764 , \18699 , \14070_nG9bf9 );
or \U$14636 ( \23765 , \23763 , \23764 );
xor \U$14637 ( \23766 , \18698 , \23765 );
buf \U$14638 ( \23767 , \23766 );
buf \U$14640 ( \23768 , \23767 );
xor \U$14641 ( \23769 , \23762 , \23768 );
and \U$14642 ( \23770 , \17297 , \14984_nG9bf6 );
and \U$14643 ( \23771 , \17294 , \15373_nG9bf3 );
or \U$14644 ( \23772 , \23770 , \23771 );
xor \U$14645 ( \23773 , \17293 , \23772 );
buf \U$14646 ( \23774 , \23773 );
buf \U$14648 ( \23775 , \23774 );
xor \U$14649 ( \23776 , \23769 , \23775 );
buf \U$14650 ( \23777 , \23776 );
xor \U$14651 ( \23778 , \23760 , \23777 );
and \U$14652 ( \23779 , \14631 , \17665_nG9bea );
and \U$14653 ( \23780 , \14628 , \18107_nG9be7 );
or \U$14654 ( \23781 , \23779 , \23780 );
xor \U$14655 ( \23782 , \14627 , \23781 );
buf \U$14656 ( \23783 , \23782 );
buf \U$14658 ( \23784 , \23783 );
xor \U$14659 ( \23785 , \23778 , \23784 );
buf \U$14660 ( \23786 , \23785 );
and \U$14661 ( \23787 , \23295 , \23301 );
and \U$14662 ( \23788 , \23295 , \23308 );
and \U$14663 ( \23789 , \23301 , \23308 );
or \U$14664 ( \23790 , \23787 , \23788 , \23789 );
buf \U$14665 ( \23791 , \23790 );
and \U$14666 ( \23792 , \23197 , \23204 );
buf \U$14667 ( \23793 , \23792 );
buf \U$14669 ( \23794 , \23793 );
and \U$14670 ( \23795 , \23201 , \10694_nG9c0e );
and \U$14671 ( \23796 , \23198 , \10995_nG9c0b );
or \U$14672 ( \23797 , \23795 , \23796 );
xor \U$14673 ( \23798 , \23197 , \23797 );
buf \U$14674 ( \23799 , \23798 );
buf \U$14676 ( \23800 , \23799 );
xor \U$14677 ( \23801 , \23794 , \23800 );
buf \U$14678 ( \23802 , \23801 );
and \U$14679 ( \23803 , \21658 , \11283_nG9c08 );
and \U$14680 ( \23804 , \21655 , \11598_nG9c05 );
or \U$14681 ( \23805 , \23803 , \23804 );
xor \U$14682 ( \23806 , \21654 , \23805 );
buf \U$14683 ( \23807 , \23806 );
buf \U$14685 ( \23808 , \23807 );
xor \U$14686 ( \23809 , \23802 , \23808 );
and \U$14687 ( \23810 , \20155 , \12470_nG9c02 );
and \U$14688 ( \23811 , \20152 , \12801_nG9bff );
or \U$14689 ( \23812 , \23810 , \23811 );
xor \U$14690 ( \23813 , \20151 , \23812 );
buf \U$14691 ( \23814 , \23813 );
buf \U$14693 ( \23815 , \23814 );
xor \U$14694 ( \23816 , \23809 , \23815 );
buf \U$14695 ( \23817 , \23816 );
xor \U$14696 ( \23818 , \23791 , \23817 );
and \U$14697 ( \23819 , \15940 , \16315_nG9bf0 );
and \U$14698 ( \23820 , \15937 , \16680_nG9bed );
or \U$14699 ( \23821 , \23819 , \23820 );
xor \U$14700 ( \23822 , \15936 , \23821 );
buf \U$14701 ( \23823 , \23822 );
buf \U$14703 ( \23824 , \23823 );
xor \U$14704 ( \23825 , \23818 , \23824 );
buf \U$14705 ( \23826 , \23825 );
and \U$14706 ( \23827 , \13370 , \19091_nG9be4 );
and \U$14707 ( \23828 , \13367 , \19586_nG9be1 );
or \U$14708 ( \23829 , \23827 , \23828 );
xor \U$14709 ( \23830 , \13366 , \23829 );
buf \U$14710 ( \23831 , \23830 );
buf \U$14712 ( \23832 , \23831 );
xor \U$14713 ( \23833 , \23826 , \23832 );
and \U$14714 ( \23834 , \12157 , \20608_nG9bde );
and \U$14715 ( \23835 , \12154 , \21086_nG9bdb );
or \U$14716 ( \23836 , \23834 , \23835 );
xor \U$14717 ( \23837 , \12153 , \23836 );
buf \U$14718 ( \23838 , \23837 );
buf \U$14720 ( \23839 , \23838 );
xor \U$14721 ( \23840 , \23833 , \23839 );
buf \U$14722 ( \23841 , \23840 );
xor \U$14723 ( \23842 , \23786 , \23841 );
and \U$14724 ( \23843 , \10707 , \23696_nG9bd2 );
and \U$14725 ( \23844 , \23667 , \23671 );
and \U$14726 ( \23845 , \23671 , \23683 );
and \U$14727 ( \23846 , \23667 , \23683 );
or \U$14728 ( \23847 , \23844 , \23845 , \23846 );
and \U$14729 ( \23848 , \23350 , \23662 );
and \U$14730 ( \23849 , \23662 , \23684 );
and \U$14731 ( \23850 , \23350 , \23684 );
or \U$14732 ( \23851 , \23848 , \23849 , \23850 );
xor \U$14733 ( \23852 , \23847 , \23851 );
and \U$14734 ( \23853 , \23632 , \23646 );
and \U$14735 ( \23854 , \23646 , \23661 );
and \U$14736 ( \23855 , \23632 , \23661 );
or \U$14737 ( \23856 , \23853 , \23854 , \23855 );
and \U$14738 ( \23857 , \23673 , \23677 );
and \U$14739 ( \23858 , \23677 , \23682 );
and \U$14740 ( \23859 , \23673 , \23682 );
or \U$14741 ( \23860 , \23857 , \23858 , \23859 );
and \U$14742 ( \23861 , \17627 , \15336 );
and \U$14743 ( \23862 , \18035 , \14963 );
nor \U$14744 ( \23863 , \23861 , \23862 );
xnor \U$14745 ( \23864 , \23863 , \15342 );
and \U$14746 ( \23865 , \11270 , \22542 );
and \U$14747 ( \23866 , \11586 , \22103 );
nor \U$14748 ( \23867 , \23865 , \23866 );
xnor \U$14749 ( \23868 , \23867 , \22548 );
xor \U$14750 ( \23869 , \23864 , \23868 );
and \U$14751 ( \23870 , RIdec53d8_708, \9333 );
and \U$14752 ( \23871 , RIdec26d8_676, \9335 );
and \U$14753 ( \23872 , RIee20080_4823, \9337 );
and \U$14754 ( \23873 , RIdebf9d8_644, \9339 );
and \U$14755 ( \23874 , RIee1f3d8_4814, \9341 );
and \U$14756 ( \23875 , RIdebccd8_612, \9343 );
and \U$14757 ( \23876 , RIdeb9fd8_580, \9345 );
and \U$14758 ( \23877 , RIdeb72d8_548, \9347 );
and \U$14759 ( \23878 , RIee1ee38_4810, \9349 );
and \U$14760 ( \23879 , RIdeb18d8_484, \9351 );
and \U$14761 ( \23880 , RIee1e898_4806, \9353 );
and \U$14762 ( \23881 , RIdeaebd8_452, \9355 );
and \U$14763 ( \23882 , RIee1da88_4796, \9357 );
and \U$14764 ( \23883 , RIdeaa420_420, \9359 );
and \U$14765 ( \23884 , RIdea3b20_388, \9361 );
and \U$14766 ( \23885 , RIde9d220_356, \9363 );
and \U$14767 ( \23886 , RIee1cde0_4787, \9365 );
and \U$14768 ( \23887 , RIee1bd00_4775, \9367 );
and \U$14769 ( \23888 , RIee1b490_4769, \9369 );
and \U$14770 ( \23889 , RIfcd8a28_7487, \9371 );
and \U$14771 ( \23890 , RIde91088_297, \9373 );
and \U$14772 ( \23891 , RIde8d8c0_280, \9375 );
and \U$14773 ( \23892 , RIfe7dac0_7774, \9377 );
and \U$14774 ( \23893 , RIfe7d958_7773, \9379 );
and \U$14775 ( \23894 , RIee1a518_4758, \9381 );
and \U$14776 ( \23895 , RIee19e10_4753, \9383 );
and \U$14777 ( \23896 , RIee19b40_4751, \9385 );
and \U$14778 ( \23897 , RIfc768c8_6371, \9387 );
and \U$14779 ( \23898 , RIfcd05f8_7393, \9389 );
and \U$14780 ( \23899 , RIfe7dd90_7776, \9391 );
and \U$14781 ( \23900 , RIee38770_5101, \9393 );
and \U$14782 ( \23901 , RIfe7dc28_7775, \9395 );
and \U$14783 ( \23902 , RIe1653d8_2529, \9397 );
and \U$14784 ( \23903 , RIe1626d8_2497, \9399 );
and \U$14785 ( \23904 , RIee373c0_5087, \9401 );
and \U$14786 ( \23905 , RIe15f9d8_2465, \9403 );
and \U$14787 ( \23906 , RIee362e0_5075, \9405 );
and \U$14788 ( \23907 , RIe15ccd8_2433, \9407 );
and \U$14789 ( \23908 , RIe1572d8_2369, \9409 );
and \U$14790 ( \23909 , RIe1545d8_2337, \9411 );
and \U$14791 ( \23910 , RIfe7def8_7777, \9413 );
and \U$14792 ( \23911 , RIe1518d8_2305, \9415 );
and \U$14793 ( \23912 , RIfebdeb8_8281, \9417 );
and \U$14794 ( \23913 , RIe14ebd8_2273, \9419 );
and \U$14795 ( \23914 , RIfc649e8_6167, \9421 );
and \U$14796 ( \23915 , RIe14bed8_2241, \9423 );
and \U$14797 ( \23916 , RIe1491d8_2209, \9425 );
and \U$14798 ( \23917 , RIe1464d8_2177, \9427 );
and \U$14799 ( \23918 , RIfe7d7f0_7772, \9429 );
and \U$14800 ( \23919 , RIfe7d688_7771, \9431 );
and \U$14801 ( \23920 , RIee32230_5029, \9433 );
and \U$14802 ( \23921 , RIfceb9e8_7703, \9435 );
and \U$14803 ( \23922 , RIfebdd50_8280, \9437 );
and \U$14804 ( \23923 , RIfe7d520_7770, \9439 );
and \U$14805 ( \23924 , RIfebdbe8_8279, \9441 );
and \U$14806 ( \23925 , RIfe7d3b8_7769, \9443 );
and \U$14807 ( \23926 , RIfc734c0_6334, \9445 );
and \U$14808 ( \23927 , RIee2f968_5000, \9447 );
and \U$14809 ( \23928 , RIfccfab8_7385, \9449 );
and \U$14810 ( \23929 , RIee2d7a8_4976, \9451 );
and \U$14811 ( \23930 , RIdf357a0_1985, \9453 );
and \U$14812 ( \23931 , RIdf33310_1959, \9455 );
and \U$14813 ( \23932 , RIdf312b8_1936, \9457 );
and \U$14814 ( \23933 , RIdf2f0f8_1912, \9459 );
or \U$14815 ( \23934 , \23870 , \23871 , \23872 , \23873 , \23874 , \23875 , \23876 , \23877 , \23878 , \23879 , \23880 , \23881 , \23882 , \23883 , \23884 , \23885 , \23886 , \23887 , \23888 , \23889 , \23890 , \23891 , \23892 , \23893 , \23894 , \23895 , \23896 , \23897 , \23898 , \23899 , \23900 , \23901 , \23902 , \23903 , \23904 , \23905 , \23906 , \23907 , \23908 , \23909 , \23910 , \23911 , \23912 , \23913 , \23914 , \23915 , \23916 , \23917 , \23918 , \23919 , \23920 , \23921 , \23922 , \23923 , \23924 , \23925 , \23926 , \23927 , \23928 , \23929 , \23930 , \23931 , \23932 , \23933 );
and \U$14816 ( \23935 , RIee2bcf0_4957, \9462 );
and \U$14817 ( \23936 , RIee2a238_4938, \9464 );
and \U$14818 ( \23937 , RIee28e88_4924, \9466 );
and \U$14819 ( \23938 , RIee27c40_4911, \9468 );
and \U$14820 ( \23939 , RIfe7ce18_7765, \9470 );
and \U$14821 ( \23940 , RIfe7ccb0_7764, \9472 );
and \U$14822 ( \23941 , RIfe7cf80_7766, \9474 );
and \U$14823 ( \23942 , RIfe7cb48_7763, \9476 );
and \U$14824 ( \23943 , RIee27268_4904, \9478 );
and \U$14825 ( \23944 , RIee26e30_4901, \9480 );
and \U$14826 ( \23945 , RIee26890_4897, \9482 );
and \U$14827 ( \23946 , RIfcaa0d8_6957, \9484 );
and \U$14828 ( \23947 , RIee262f0_4893, \9486 );
and \U$14829 ( \23948 , RIfe7d250_7768, \9488 );
and \U$14830 ( \23949 , RIee26020_4891, \9490 );
and \U$14831 ( \23950 , RIfe7d0e8_7767, \9492 );
and \U$14832 ( \23951 , RIdf16fa8_1638, \9494 );
and \U$14833 ( \23952 , RIdf142a8_1606, \9496 );
and \U$14834 ( \23953 , RIdf115a8_1574, \9498 );
and \U$14835 ( \23954 , RIdf0e8a8_1542, \9500 );
and \U$14836 ( \23955 , RIdf0bba8_1510, \9502 );
and \U$14837 ( \23956 , RIdf08ea8_1478, \9504 );
and \U$14838 ( \23957 , RIdf061a8_1446, \9506 );
and \U$14839 ( \23958 , RIdf034a8_1414, \9508 );
and \U$14840 ( \23959 , RIdefdaa8_1350, \9510 );
and \U$14841 ( \23960 , RIdefada8_1318, \9512 );
and \U$14842 ( \23961 , RIdef80a8_1286, \9514 );
and \U$14843 ( \23962 , RIdef53a8_1254, \9516 );
and \U$14844 ( \23963 , RIdef26a8_1222, \9518 );
and \U$14845 ( \23964 , RIdeef9a8_1190, \9520 );
and \U$14846 ( \23965 , RIdeecca8_1158, \9522 );
and \U$14847 ( \23966 , RIdee9fa8_1126, \9524 );
and \U$14848 ( \23967 , RIee25648_4884, \9526 );
and \U$14849 ( \23968 , RIee249a0_4875, \9528 );
and \U$14850 ( \23969 , RIfebe020_8282, \9530 );
and \U$14851 ( \23970 , RIee23488_4860, \9532 );
and \U$14852 ( \23971 , RIfebe2f0_8284, \9534 );
and \U$14853 ( \23972 , RIfebe188_8283, \9536 );
and \U$14854 ( \23973 , RIfe7e1c8_7779, \9538 );
and \U$14855 ( \23974 , RIfe7e060_7778, \9540 );
and \U$14856 ( \23975 , RIfcbf7f8_7201, \9542 );
and \U$14857 ( \23976 , RIfc7aae0_6418, \9544 );
and \U$14858 ( \23977 , RIfc787b8_6393, \9546 );
and \U$14859 ( \23978 , RIfc618b0_6132, \9548 );
and \U$14860 ( \23979 , RIded98b0_939, \9550 );
and \U$14861 ( \23980 , RIded72b8_912, \9552 );
and \U$14862 ( \23981 , RIded5530_891, \9554 );
and \U$14863 ( \23982 , RIded2dd0_863, \9556 );
and \U$14864 ( \23983 , RIded07d8_836, \9558 );
and \U$14865 ( \23984 , RIdecdad8_804, \9560 );
and \U$14866 ( \23985 , RIdecadd8_772, \9562 );
and \U$14867 ( \23986 , RIdec80d8_740, \9564 );
and \U$14868 ( \23987 , RIdeb45d8_516, \9566 );
and \U$14869 ( \23988 , RIde96920_324, \9568 );
and \U$14870 ( \23989 , RIe16e1e0_2630, \9570 );
and \U$14871 ( \23990 , RIe159fd8_2401, \9572 );
and \U$14872 ( \23991 , RIe1437d8_2145, \9574 );
and \U$14873 ( \23992 , RIdf381d0_2015, \9576 );
and \U$14874 ( \23993 , RIdf2c830_1883, \9578 );
and \U$14875 ( \23994 , RIdf1d0b0_1707, \9580 );
and \U$14876 ( \23995 , RIdf007a8_1382, \9582 );
and \U$14877 ( \23996 , RIdee72a8_1094, \9584 );
and \U$14878 ( \23997 , RIdedc010_967, \9586 );
and \U$14879 ( \23998 , RIde7c868_197, \9588 );
or \U$14880 ( \23999 , \23935 , \23936 , \23937 , \23938 , \23939 , \23940 , \23941 , \23942 , \23943 , \23944 , \23945 , \23946 , \23947 , \23948 , \23949 , \23950 , \23951 , \23952 , \23953 , \23954 , \23955 , \23956 , \23957 , \23958 , \23959 , \23960 , \23961 , \23962 , \23963 , \23964 , \23965 , \23966 , \23967 , \23968 , \23969 , \23970 , \23971 , \23972 , \23973 , \23974 , \23975 , \23976 , \23977 , \23978 , \23979 , \23980 , \23981 , \23982 , \23983 , \23984 , \23985 , \23986 , \23987 , \23988 , \23989 , \23990 , \23991 , \23992 , \23993 , \23994 , \23995 , \23996 , \23997 , \23998 );
or \U$14881 ( \24000 , \23934 , \23999 );
_DC g5a97 ( \24001_nG5a97 , \24000 , \9597 );
and \U$14882 ( \24002 , RIe19d670_3168, \9059 );
and \U$14883 ( \24003 , RIe19a970_3136, \9061 );
and \U$14884 ( \24004 , RIfe7b630_7748, \9063 );
and \U$14885 ( \24005 , RIe197c70_3104, \9065 );
and \U$14886 ( \24006 , RIfe7b4c8_7747, \9067 );
and \U$14887 ( \24007 , RIe194f70_3072, \9069 );
and \U$14888 ( \24008 , RIe192270_3040, \9071 );
and \U$14889 ( \24009 , RIe18f570_3008, \9073 );
and \U$14890 ( \24010 , RIe189b70_2944, \9075 );
and \U$14891 ( \24011 , RIe186e70_2912, \9077 );
and \U$14892 ( \24012 , RIfe7b360_7746, \9079 );
and \U$14893 ( \24013 , RIe184170_2880, \9081 );
and \U$14894 ( \24014 , RIfe7b1f8_7745, \9083 );
and \U$14895 ( \24015 , RIe181470_2848, \9085 );
and \U$14896 ( \24016 , RIe17e770_2816, \9087 );
and \U$14897 ( \24017 , RIe17ba70_2784, \9089 );
and \U$14898 ( \24018 , RIf1423b8_5213, \9091 );
and \U$14899 ( \24019 , RIf140ea0_5198, \9093 );
and \U$14900 ( \24020 , RIf140360_5190, \9095 );
and \U$14901 ( \24021 , RIfe7b798_7749, \9097 );
and \U$14902 ( \24022 , RIf13fc58_5185, \9099 );
and \U$14903 ( \24023 , RIf13f280_5178, \9101 );
and \U$14904 ( \24024 , RIfc79460_6402, \9103 );
and \U$14905 ( \24025 , RIee3d4c8_5156, \9105 );
and \U$14906 ( \24026 , RIfe7b090_7744, \9107 );
and \U$14907 ( \24027 , RIfe7af28_7743, \9109 );
and \U$14908 ( \24028 , RIee39df0_5117, \9111 );
and \U$14909 ( \24029 , RIe1737a8_2691, \9113 );
and \U$14910 ( \24030 , RIfe7adc0_7742, \9115 );
and \U$14911 ( \24031 , RIfe7ac58_7741, \9117 );
and \U$14912 ( \24032 , RIf16e440_5714, \9119 );
and \U$14913 ( \24033 , RIfcb20d0_7048, \9121 );
and \U$14914 ( \24034 , RIfe7bd38_7753, \9123 );
and \U$14915 ( \24035 , RIe2239c8_4695, \9125 );
and \U$14916 ( \24036 , RIf16be48_5687, \9127 );
and \U$14917 ( \24037 , RIe220cc8_4663, \9129 );
and \U$14918 ( \24038 , RIf16aed0_5676, \9131 );
and \U$14919 ( \24039 , RIe21dfc8_4631, \9133 );
and \U$14920 ( \24040 , RIe2185c8_4567, \9135 );
and \U$14921 ( \24041 , RIe2158c8_4535, \9137 );
and \U$14922 ( \24042 , RIfebd7b0_8276, \9139 );
and \U$14923 ( \24043 , RIe212bc8_4503, \9141 );
and \U$14924 ( \24044 , RIfebd648_8275, \9143 );
and \U$14925 ( \24045 , RIe20fec8_4471, \9145 );
and \U$14926 ( \24046 , RIfe7b900_7750, \9147 );
and \U$14927 ( \24047 , RIe20d1c8_4439, \9149 );
and \U$14928 ( \24048 , RIe20a4c8_4407, \9151 );
and \U$14929 ( \24049 , RIe2077c8_4375, \9153 );
and \U$14930 ( \24050 , RIf167258_5633, \9155 );
and \U$14931 ( \24051 , RIf166178_5621, \9157 );
and \U$14932 ( \24052 , RIe2024d0_4316, \9159 );
and \U$14933 ( \24053 , RIfe7bbd0_7752, \9161 );
and \U$14934 ( \24054 , RIf165368_5611, \9163 );
and \U$14935 ( \24055 , RIf1646c0_5602, \9165 );
and \U$14936 ( \24056 , RIfcd0a30_7396, \9167 );
and \U$14937 ( \24057 , RIf1620c8_5575, \9169 );
and \U$14938 ( \24058 , RIf1601d8_5553, \9171 );
and \U$14939 ( \24059 , RIf15e2e8_5531, \9173 );
and \U$14940 ( \24060 , RIfe7ba68_7751, \9175 );
and \U$14941 ( \24061 , RIfe7bea0_7754, \9177 );
and \U$14942 ( \24062 , RIf15cdd0_5516, \9179 );
and \U$14943 ( \24063 , RIf15b8b8_5501, \9181 );
and \U$14944 ( \24064 , RIf15a7d8_5489, \9183 );
and \U$14945 ( \24065 , RIfca4840_6894, \9185 );
or \U$14946 ( \24066 , \24002 , \24003 , \24004 , \24005 , \24006 , \24007 , \24008 , \24009 , \24010 , \24011 , \24012 , \24013 , \24014 , \24015 , \24016 , \24017 , \24018 , \24019 , \24020 , \24021 , \24022 , \24023 , \24024 , \24025 , \24026 , \24027 , \24028 , \24029 , \24030 , \24031 , \24032 , \24033 , \24034 , \24035 , \24036 , \24037 , \24038 , \24039 , \24040 , \24041 , \24042 , \24043 , \24044 , \24045 , \24046 , \24047 , \24048 , \24049 , \24050 , \24051 , \24052 , \24053 , \24054 , \24055 , \24056 , \24057 , \24058 , \24059 , \24060 , \24061 , \24062 , \24063 , \24064 , \24065 );
and \U$14947 ( \24067 , RIf158ff0_5472, \9188 );
and \U$14948 ( \24068 , RIf157c40_5458, \9190 );
and \U$14949 ( \24069 , RIf156f98_5449, \9192 );
and \U$14950 ( \24070 , RIfe7c170_7756, \9194 );
and \U$14951 ( \24071 , RIf156458_5441, \9196 );
and \U$14952 ( \24072 , RIf155918_5433, \9198 );
and \U$14953 ( \24073 , RIf1549a0_5422, \9200 );
and \U$14954 ( \24074 , RIe1f54b0_4168, \9202 );
and \U$14955 ( \24075 , RIfe7c008_7755, \9204 );
and \U$14956 ( \24076 , RIf151b38_5389, \9206 );
and \U$14957 ( \24077 , RIf150bc0_5378, \9208 );
and \U$14958 ( \24078 , RIe1f32f0_4144, \9210 );
and \U$14959 ( \24079 , RIf14fae0_5366, \9212 );
and \U$14960 ( \24080 , RIf14ee38_5357, \9214 );
and \U$14961 ( \24081 , RIf14e028_5347, \9216 );
and \U$14962 ( \24082 , RIe1edff8_4085, \9218 );
and \U$14963 ( \24083 , RIe1eb730_4056, \9220 );
and \U$14964 ( \24084 , RIe1e8a30_4024, \9222 );
and \U$14965 ( \24085 , RIe1e5d30_3992, \9224 );
and \U$14966 ( \24086 , RIe1e3030_3960, \9226 );
and \U$14967 ( \24087 , RIe1e0330_3928, \9228 );
and \U$14968 ( \24088 , RIe1dd630_3896, \9230 );
and \U$14969 ( \24089 , RIe1da930_3864, \9232 );
and \U$14970 ( \24090 , RIe1d7c30_3832, \9234 );
and \U$14971 ( \24091 , RIe1d2230_3768, \9236 );
and \U$14972 ( \24092 , RIe1cf530_3736, \9238 );
and \U$14973 ( \24093 , RIe1cc830_3704, \9240 );
and \U$14974 ( \24094 , RIe1c9b30_3672, \9242 );
and \U$14975 ( \24095 , RIe1c6e30_3640, \9244 );
and \U$14976 ( \24096 , RIe1c4130_3608, \9246 );
and \U$14977 ( \24097 , RIe1c1430_3576, \9248 );
and \U$14978 ( \24098 , RIe1be730_3544, \9250 );
and \U$14979 ( \24099 , RIf14cb10_5332, \9252 );
and \U$14980 ( \24100 , RIf14b8c8_5319, \9254 );
and \U$14981 ( \24101 , RIfebda80_8278, \9256 );
and \U$14982 ( \24102 , RIfe7c878_7761, \9258 );
and \U$14983 ( \24103 , RIf14a680_5306, \9260 );
and \U$14984 ( \24104 , RIfe7c2d8_7757, \9262 );
and \U$14985 ( \24105 , RIfe7c9e0_7762, \9264 );
and \U$14986 ( \24106 , RIfe7c440_7758, \9266 );
and \U$14987 ( \24107 , RIf149000_5290, \9268 );
and \U$14988 ( \24108 , RIf147db8_5277, \9270 );
and \U$14989 ( \24109 , RIe1b2688_3407, \9272 );
and \U$14990 ( \24110 , RIfebd918_8277, \9274 );
and \U$14991 ( \24111 , RIfe7c5a8_7759, \9276 );
and \U$14992 ( \24112 , RIf146738_5261, \9278 );
and \U$14993 ( \24113 , RIfe7c710_7760, \9280 );
and \U$14994 ( \24114 , RIe1aad98_3321, \9282 );
and \U$14995 ( \24115 , RIe1a8a70_3296, \9284 );
and \U$14996 ( \24116 , RIe1a5d70_3264, \9286 );
and \U$14997 ( \24117 , RIe1a3070_3232, \9288 );
and \U$14998 ( \24118 , RIe1a0370_3200, \9290 );
and \U$14999 ( \24119 , RIe18c870_2976, \9292 );
and \U$15000 ( \24120 , RIe178d70_2752, \9294 );
and \U$15001 ( \24121 , RIe2266c8_4727, \9296 );
and \U$15002 ( \24122 , RIe21b2c8_4599, \9298 );
and \U$15003 ( \24123 , RIe204ac8_4343, \9300 );
and \U$15004 ( \24124 , RIe1feb28_4275, \9302 );
and \U$15005 ( \24125 , RIe1f7ee0_4198, \9304 );
and \U$15006 ( \24126 , RIe1f0a28_4115, \9306 );
and \U$15007 ( \24127 , RIe1d4f30_3800, \9308 );
and \U$15008 ( \24128 , RIe1bba30_3512, \9310 );
and \U$15009 ( \24129 , RIe1ae8a8_3363, \9312 );
and \U$15010 ( \24130 , RIe170ee0_2662, \9314 );
or \U$15011 ( \24131 , \24067 , \24068 , \24069 , \24070 , \24071 , \24072 , \24073 , \24074 , \24075 , \24076 , \24077 , \24078 , \24079 , \24080 , \24081 , \24082 , \24083 , \24084 , \24085 , \24086 , \24087 , \24088 , \24089 , \24090 , \24091 , \24092 , \24093 , \24094 , \24095 , \24096 , \24097 , \24098 , \24099 , \24100 , \24101 , \24102 , \24103 , \24104 , \24105 , \24106 , \24107 , \24108 , \24109 , \24110 , \24111 , \24112 , \24113 , \24114 , \24115 , \24116 , \24117 , \24118 , \24119 , \24120 , \24121 , \24122 , \24123 , \24124 , \24125 , \24126 , \24127 , \24128 , \24129 , \24130 );
or \U$15012 ( \24132 , \24066 , \24131 );
_DC g5b1b ( \24133_nG5b1b , \24132 , \9323 );
xor g5b1c ( \24134_nG5b1c , \24001_nG5a97 , \24133_nG5b1b );
buf \U$15013 ( \24135 , \24134_nG5b1c );
xor \U$15014 ( \24136 , \24135 , \23629 );
not \U$15015 ( \24137 , \23630 );
and \U$15016 ( \24138 , \24136 , \24137 );
and \U$15017 ( \24139 , \10687 , \24138 );
and \U$15018 ( \24140 , \10988 , \23630 );
nor \U$15019 ( \24141 , \24139 , \24140 );
and \U$15020 ( \24142 , \23629 , \22539 );
not \U$15021 ( \24143 , \24142 );
and \U$15022 ( \24144 , \24135 , \24143 );
xnor \U$15023 ( \24145 , \24141 , \24144 );
xor \U$15024 ( \24146 , \23869 , \24145 );
xor \U$15025 ( \24147 , \23860 , \24146 );
and \U$15026 ( \24148 , \19032 , \14054 );
and \U$15027 ( \24149 , \19558 , \13692 );
nor \U$15028 ( \24150 , \24148 , \24149 );
xnor \U$15029 ( \24151 , \24150 , \14035 );
and \U$15030 ( \24152 , \13679 , \19534 );
and \U$15031 ( \24153 , \14024 , \19045 );
nor \U$15032 ( \24154 , \24152 , \24153 );
xnor \U$15033 ( \24155 , \24154 , \19540 );
xor \U$15034 ( \24156 , \24151 , \24155 );
and \U$15035 ( \24157 , \12448 , \21005 );
and \U$15036 ( \24158 , \12769 , \20557 );
nor \U$15037 ( \24159 , \24157 , \24158 );
xnor \U$15038 ( \24160 , \24159 , \21011 );
xor \U$15039 ( \24161 , \24156 , \24160 );
xor \U$15040 ( \24162 , \24147 , \24161 );
xor \U$15041 ( \24163 , \23856 , \24162 );
and \U$15042 ( \24164 , \23340 , \23344 );
and \U$15043 ( \24165 , \23344 , \23349 );
and \U$15044 ( \24166 , \23340 , \23349 );
or \U$15045 ( \24167 , \24164 , \24165 , \24166 );
and \U$15046 ( \24168 , \22090 , \11574 );
and \U$15047 ( \24169 , \22556 , \11278 );
nor \U$15048 ( \24170 , \24168 , \24169 );
xnor \U$15049 ( \24171 , \24170 , \11580 );
not \U$15050 ( \24172 , \23631 );
and \U$15051 ( \24173 , \24172 , \24144 );
xor \U$15052 ( \24174 , \24171 , \24173 );
and \U$15053 ( \24175 , \23651 , \23655 );
and \U$15054 ( \24176 , \23655 , \23660 );
and \U$15055 ( \24177 , \23651 , \23660 );
or \U$15056 ( \24178 , \24175 , \24176 , \24177 );
xor \U$15057 ( \24179 , \24174 , \24178 );
and \U$15058 ( \24180 , \14950 , \18090 );
and \U$15059 ( \24181 , \15321 , \17655 );
nor \U$15060 ( \24182 , \24180 , \24181 );
xnor \U$15061 ( \24183 , \24182 , \18046 );
xor \U$15062 ( \24184 , \24179 , \24183 );
xor \U$15063 ( \24185 , \24167 , \24184 );
and \U$15064 ( \24186 , \23620 , \23624 );
and \U$15065 ( \24187 , \23624 , \23631 );
and \U$15066 ( \24188 , \23620 , \23631 );
or \U$15067 ( \24189 , \24186 , \24187 , \24188 );
and \U$15068 ( \24190 , \23636 , \23640 );
and \U$15069 ( \24191 , \23640 , \23645 );
and \U$15070 ( \24192 , \23636 , \23645 );
or \U$15071 ( \24193 , \24190 , \24191 , \24192 );
xor \U$15072 ( \24194 , \24189 , \24193 );
and \U$15073 ( \24195 , \23617 , \10983 );
_DC g65b6 ( \24196_nG65b6 , \24000 , \9597 );
_DC g65b7 ( \24197_nG65b7 , \24132 , \9323 );
and g65b8 ( \24198_nG65b8 , \24196_nG65b6 , \24197_nG65b7 );
buf \U$15074 ( \24199 , \24198_nG65b8 );
and \U$15075 ( \24200 , \24199 , \10691 );
nor \U$15076 ( \24201 , \24195 , \24200 );
xnor \U$15077 ( \24202 , \24201 , \10980 );
and \U$15078 ( \24203 , \20544 , \12790 );
and \U$15079 ( \24204 , \21033 , \12461 );
nor \U$15080 ( \24205 , \24203 , \24204 );
xnor \U$15081 ( \24206 , \24205 , \12780 );
xor \U$15082 ( \24207 , \24202 , \24206 );
and \U$15083 ( \24208 , \16267 , \16635 );
and \U$15084 ( \24209 , \16655 , \16301 );
nor \U$15085 ( \24210 , \24208 , \24209 );
xnor \U$15086 ( \24211 , \24210 , \16625 );
xor \U$15087 ( \24212 , \24207 , \24211 );
xor \U$15088 ( \24213 , \24194 , \24212 );
xor \U$15089 ( \24214 , \24185 , \24213 );
xor \U$15090 ( \24215 , \24163 , \24214 );
xor \U$15091 ( \24216 , \23852 , \24215 );
and \U$15092 ( \24217 , \23331 , \23335 );
and \U$15093 ( \24218 , \23335 , \23685 );
and \U$15094 ( \24219 , \23331 , \23685 );
or \U$15095 ( \24220 , \24217 , \24218 , \24219 );
xor \U$15096 ( \24221 , \24216 , \24220 );
and \U$15097 ( \24222 , \23686 , \23690 );
and \U$15098 ( \24223 , \23691 , \23694 );
or \U$15099 ( \24224 , \24222 , \24223 );
xor \U$15100 ( \24225 , \24221 , \24224 );
buf g9bcf ( \24226_nG9bcf , \24225 );
and \U$15101 ( \24227 , \10704 , \24226_nG9bcf );
or \U$15102 ( \24228 , \23843 , \24227 );
xor \U$15103 ( \24229 , \10703 , \24228 );
buf \U$15104 ( \24230 , \24229 );
buf \U$15106 ( \24231 , \24230 );
xor \U$15107 ( \24232 , \23842 , \24231 );
buf \U$15108 ( \24233 , \24232 );
xor \U$15109 ( \24234 , \23755 , \24233 );
and \U$15110 ( \24235 , \23717 , \24234 );
and \U$15111 ( \24236 , \23707 , \23711 );
and \U$15112 ( \24237 , \23707 , \23716 );
and \U$15113 ( \24238 , \23711 , \23716 );
or \U$15114 ( \24239 , \24236 , \24237 , \24238 );
xor \U$15115 ( \24240 , \24235 , \24239 );
and \U$15116 ( \24241 , RIdec56a8_710, \9059 );
and \U$15117 ( \24242 , RIdec29a8_678, \9061 );
and \U$15118 ( \24243 , RIfc54020_5978, \9063 );
and \U$15119 ( \24244 , RIdebfca8_646, \9065 );
and \U$15120 ( \24245 , RIee1f540_4815, \9067 );
and \U$15121 ( \24246 , RIdebcfa8_614, \9069 );
and \U$15122 ( \24247 , RIdeba2a8_582, \9071 );
and \U$15123 ( \24248 , RIdeb75a8_550, \9073 );
and \U$15124 ( \24249 , RIfc4fe08_5931, \9075 );
and \U$15125 ( \24250 , RIdeb1ba8_486, \9077 );
and \U$15126 ( \24251 , RIfc6b630_6244, \9079 );
and \U$15127 ( \24252 , RIdeaeea8_454, \9081 );
and \U$15128 ( \24253 , RIfc6a118_6229, \9083 );
and \U$15129 ( \24254 , RIdeaaab0_422, \9085 );
and \U$15130 ( \24255 , RIdea41b0_390, \9087 );
and \U$15131 ( \24256 , RIde9d8b0_358, \9089 );
and \U$15132 ( \24257 , RIfc69ce0_6226, \9091 );
and \U$15133 ( \24258 , RIee1be68_4776, \9093 );
and \U$15134 ( \24259 , RIfc653c0_6174, \9095 );
and \U$15135 ( \24260 , RIee1ac20_4763, \9097 );
and \U$15136 ( \24261 , RIde91718_299, \9099 );
and \U$15137 ( \24262 , RIde8df50_282, \9101 );
and \U$15138 ( \24263 , RIde89db0_262, \9103 );
and \U$15139 ( \24264 , RIde85c10_242, \9105 );
and \U$15140 ( \24265 , RIde81db8_223, \9107 );
and \U$15141 ( \24266 , RIfca76a8_6927, \9109 );
and \U$15142 ( \24267 , RIfcca4f0_7324, \9111 );
and \U$15143 ( \24268 , RIfc4ce38_5897, \9113 );
and \U$15144 ( \24269 , RIfc6b360_6242, \9115 );
and \U$15145 ( \24270 , RIe16b918_2601, \9117 );
and \U$15146 ( \24271 , RIe169cf8_2581, \9119 );
and \U$15147 ( \24272 , RIe167f70_2560, \9121 );
and \U$15148 ( \24273 , RIe1656a8_2531, \9123 );
and \U$15149 ( \24274 , RIe1629a8_2499, \9125 );
and \U$15150 ( \24275 , RIee37690_5089, \9127 );
and \U$15151 ( \24276 , RIe15fca8_2467, \9129 );
and \U$15152 ( \24277 , RIfce93f0_7676, \9131 );
and \U$15153 ( \24278 , RIe15cfa8_2435, \9133 );
and \U$15154 ( \24279 , RIe1575a8_2371, \9135 );
and \U$15155 ( \24280 , RIe1548a8_2339, \9137 );
and \U$15156 ( \24281 , RIee35908_5068, \9139 );
and \U$15157 ( \24282 , RIe151ba8_2307, \9141 );
and \U$15158 ( \24283 , RIee34f30_5061, \9143 );
and \U$15159 ( \24284 , RIe14eea8_2275, \9145 );
and \U$15160 ( \24285 , RIfce32e8_7607, \9147 );
and \U$15161 ( \24286 , RIe14c1a8_2243, \9149 );
and \U$15162 ( \24287 , RIe1494a8_2211, \9151 );
and \U$15163 ( \24288 , RIe1467a8_2179, \9153 );
and \U$15164 ( \24289 , RIfcde2c0_7550, \9155 );
and \U$15165 ( \24290 , RIfc687c8_6211, \9157 );
and \U$15166 ( \24291 , RIfca9160_6946, \9159 );
and \U$15167 ( \24292 , RIfcb1590_7040, \9161 );
and \U$15168 ( \24293 , RIe141078_2117, \9163 );
and \U$15169 ( \24294 , RIdf3ef80_2093, \9165 );
and \U$15170 ( \24295 , RIdf3cdc0_2069, \9167 );
and \U$15171 ( \24296 , RIfebeb60_8290, \9169 );
and \U$15172 ( \24297 , RIfc64448_6163, \9171 );
and \U$15173 ( \24298 , RIee2fad0_5001, \9173 );
and \U$15174 ( \24299 , RIfca7978_6929, \9175 );
and \U$15175 ( \24300 , RIfc676e8_6199, \9177 );
and \U$15176 ( \24301 , RIdf35a70_1987, \9179 );
and \U$15177 ( \24302 , RIdf335e0_1961, \9181 );
and \U$15178 ( \24303 , RIdf31420_1937, \9183 );
and \U$15179 ( \24304 , RIdf2f3c8_1914, \9185 );
or \U$15180 ( \24305 , \24241 , \24242 , \24243 , \24244 , \24245 , \24246 , \24247 , \24248 , \24249 , \24250 , \24251 , \24252 , \24253 , \24254 , \24255 , \24256 , \24257 , \24258 , \24259 , \24260 , \24261 , \24262 , \24263 , \24264 , \24265 , \24266 , \24267 , \24268 , \24269 , \24270 , \24271 , \24272 , \24273 , \24274 , \24275 , \24276 , \24277 , \24278 , \24279 , \24280 , \24281 , \24282 , \24283 , \24284 , \24285 , \24286 , \24287 , \24288 , \24289 , \24290 , \24291 , \24292 , \24293 , \24294 , \24295 , \24296 , \24297 , \24298 , \24299 , \24300 , \24301 , \24302 , \24303 , \24304 );
and \U$15181 ( \24306 , RIfccef78_7377, \9188 );
and \U$15182 ( \24307 , RIfca6fa0_6922, \9190 );
and \U$15183 ( \24308 , RIfc62558_6141, \9192 );
and \U$15184 ( \24309 , RIfc61fb8_6137, \9194 );
and \U$15185 ( \24310 , RIfe81b70_7820, \9196 );
and \U$15186 ( \24311 , RIdf281e0_1833, \9198 );
and \U$15187 ( \24312 , RIfe81cd8_7821, \9200 );
and \U$15188 ( \24313 , RIdf249a0_1793, \9202 );
and \U$15189 ( \24314 , RIfc44300_5798, \9204 );
and \U$15190 ( \24315 , RIfcafc40_7022, \9206 );
and \U$15191 ( \24316 , RIdf22ee8_1774, \9208 );
and \U$15192 ( \24317 , RIfcaac18_6965, \9210 );
and \U$15193 ( \24318 , RIdf219d0_1759, \9212 );
and \U$15194 ( \24319 , RIdf1fae0_1737, \9214 );
and \U$15195 ( \24320 , RIdf1b1c0_1685, \9216 );
and \U$15196 ( \24321 , RIdf19438_1664, \9218 );
and \U$15197 ( \24322 , RIdf17278_1640, \9220 );
and \U$15198 ( \24323 , RIdf14578_1608, \9222 );
and \U$15199 ( \24324 , RIdf11878_1576, \9224 );
and \U$15200 ( \24325 , RIdf0eb78_1544, \9226 );
and \U$15201 ( \24326 , RIdf0be78_1512, \9228 );
and \U$15202 ( \24327 , RIdf09178_1480, \9230 );
and \U$15203 ( \24328 , RIdf06478_1448, \9232 );
and \U$15204 ( \24329 , RIdf03778_1416, \9234 );
and \U$15205 ( \24330 , RIdefdd78_1352, \9236 );
and \U$15206 ( \24331 , RIdefb078_1320, \9238 );
and \U$15207 ( \24332 , RIdef8378_1288, \9240 );
and \U$15208 ( \24333 , RIdef5678_1256, \9242 );
and \U$15209 ( \24334 , RIdef2978_1224, \9244 );
and \U$15210 ( \24335 , RIdeefc78_1192, \9246 );
and \U$15211 ( \24336 , RIdeecf78_1160, \9248 );
and \U$15212 ( \24337 , RIdeea278_1128, \9250 );
and \U$15213 ( \24338 , RIfc611a8_6127, \9252 );
and \U$15214 ( \24339 , RIfc61a18_6133, \9254 );
and \U$15215 ( \24340 , RIfca65c8_6915, \9256 );
and \U$15216 ( \24341 , RIfca6b68_6919, \9258 );
and \U$15217 ( \24342 , RIdee4b48_1066, \9260 );
and \U$15218 ( \24343 , RIdee2dc0_1045, \9262 );
and \U$15219 ( \24344 , RIdee0c00_1021, \9264 );
and \U$15220 ( \24345 , RIdedeba8_998, \9266 );
and \U$15221 ( \24346 , RIfc626c0_6142, \9268 );
and \U$15222 ( \24347 , RIfc738f8_6337, \9270 );
and \U$15223 ( \24348 , RIfcb31b0_7060, \9272 );
and \U$15224 ( \24349 , RIee21430_4837, \9274 );
and \U$15225 ( \24350 , RIded9a18_940, \9276 );
and \U$15226 ( \24351 , RIded7588_914, \9278 );
and \U$15227 ( \24352 , RIded5698_892, \9280 );
and \U$15228 ( \24353 , RIded30a0_865, \9282 );
and \U$15229 ( \24354 , RIded0aa8_838, \9284 );
and \U$15230 ( \24355 , RIdecdda8_806, \9286 );
and \U$15231 ( \24356 , RIdecb0a8_774, \9288 );
and \U$15232 ( \24357 , RIdec83a8_742, \9290 );
and \U$15233 ( \24358 , RIdeb48a8_518, \9292 );
and \U$15234 ( \24359 , RIde96fb0_326, \9294 );
and \U$15235 ( \24360 , RIe16e4b0_2632, \9296 );
and \U$15236 ( \24361 , RIe15a2a8_2403, \9298 );
and \U$15237 ( \24362 , RIe143aa8_2147, \9300 );
and \U$15238 ( \24363 , RIdf384a0_2017, \9302 );
and \U$15239 ( \24364 , RIdf2cb00_1885, \9304 );
and \U$15240 ( \24365 , RIdf1d380_1709, \9306 );
and \U$15241 ( \24366 , RIdf00a78_1384, \9308 );
and \U$15242 ( \24367 , RIdee7578_1096, \9310 );
and \U$15243 ( \24368 , RIdedc2e0_969, \9312 );
and \U$15244 ( \24369 , RIde7cef8_199, \9314 );
or \U$15245 ( \24370 , \24306 , \24307 , \24308 , \24309 , \24310 , \24311 , \24312 , \24313 , \24314 , \24315 , \24316 , \24317 , \24318 , \24319 , \24320 , \24321 , \24322 , \24323 , \24324 , \24325 , \24326 , \24327 , \24328 , \24329 , \24330 , \24331 , \24332 , \24333 , \24334 , \24335 , \24336 , \24337 , \24338 , \24339 , \24340 , \24341 , \24342 , \24343 , \24344 , \24345 , \24346 , \24347 , \24348 , \24349 , \24350 , \24351 , \24352 , \24353 , \24354 , \24355 , \24356 , \24357 , \24358 , \24359 , \24360 , \24361 , \24362 , \24363 , \24364 , \24365 , \24366 , \24367 , \24368 , \24369 );
or \U$15246 ( \24371 , \24305 , \24370 );
_DC g265d ( \24372_nG265d , \24371 , \9323 );
buf \U$15247 ( \24373 , \24372_nG265d );
and \U$15248 ( \24374 , RIe19d940_3170, \9333 );
and \U$15249 ( \24375 , RIe19ac40_3138, \9335 );
and \U$15250 ( \24376 , RIfc64880_6166, \9337 );
and \U$15251 ( \24377 , RIe197f40_3106, \9339 );
and \U$15252 ( \24378 , RIf144848_5239, \9341 );
and \U$15253 ( \24379 , RIe195240_3074, \9343 );
and \U$15254 ( \24380 , RIe192540_3042, \9345 );
and \U$15255 ( \24381 , RIe18f840_3010, \9347 );
and \U$15256 ( \24382 , RIe189e40_2946, \9349 );
and \U$15257 ( \24383 , RIe187140_2914, \9351 );
and \U$15258 ( \24384 , RIf143a38_5229, \9353 );
and \U$15259 ( \24385 , RIe184440_2882, \9355 );
and \U$15260 ( \24386 , RIfc6f140_6286, \9357 );
and \U$15261 ( \24387 , RIe181740_2850, \9359 );
and \U$15262 ( \24388 , RIe17ea40_2818, \9361 );
and \U$15263 ( \24389 , RIe17bd40_2786, \9363 );
and \U$15264 ( \24390 , RIfc64f88_6171, \9365 );
and \U$15265 ( \24391 , RIf141008_5199, \9367 );
and \U$15266 ( \24392 , RIe177150_2732, \9369 );
and \U$15267 ( \24393 , RIfe81738_7817, \9371 );
and \U$15268 ( \24394 , RIfccabf8_7329, \9373 );
and \U$15269 ( \24395 , RIf13f3e8_5179, \9375 );
and \U$15270 ( \24396 , RIfca81e8_6935, \9377 );
and \U$15271 ( \24397 , RIee3d630_5157, \9379 );
and \U$15272 ( \24398 , RIfc66068_6183, \9381 );
and \U$15273 ( \24399 , RIfc6ed08_6283, \9383 );
and \U$15274 ( \24400 , RIfcdde88_7547, \9385 );
and \U$15275 ( \24401 , RIe173a78_2693, \9387 );
and \U$15276 ( \24402 , RIfc66338_6185, \9389 );
and \U$15277 ( \24403 , RIfc6eba0_6282, \9391 );
and \U$15278 ( \24404 , RIfc664a0_6186, \9393 );
and \U$15279 ( \24405 , RIfcacdd8_6989, \9395 );
and \U$15280 ( \24406 , RIfe81468_7815, \9397 );
and \U$15281 ( \24407 , RIe223c98_4697, \9399 );
and \U$15282 ( \24408 , RIfc66d10_6192, \9401 );
and \U$15283 ( \24409 , RIe220f98_4665, \9403 );
and \U$15284 ( \24410 , RIf16b038_5677, \9405 );
and \U$15285 ( \24411 , RIe21e298_4633, \9407 );
and \U$15286 ( \24412 , RIe218898_4569, \9409 );
and \U$15287 ( \24413 , RIe215b98_4537, \9411 );
and \U$15288 ( \24414 , RIfc3fc38_5751, \9413 );
and \U$15289 ( \24415 , RIe212e98_4505, \9415 );
and \U$15290 ( \24416 , RIfc67850_6200, \9417 );
and \U$15291 ( \24417 , RIe210198_4473, \9419 );
and \U$15292 ( \24418 , RIf167f00_5642, \9421 );
and \U$15293 ( \24419 , RIe20d498_4441, \9423 );
and \U$15294 ( \24420 , RIe20a798_4409, \9425 );
and \U$15295 ( \24421 , RIe207a98_4377, \9427 );
and \U$15296 ( \24422 , RIfcacb08_6987, \9429 );
and \U$15297 ( \24423 , RIfcac9a0_6986, \9431 );
and \U$15298 ( \24424 , RIfea8900_8234, \9433 );
and \U$15299 ( \24425 , RIfe818a0_7818, \9435 );
and \U$15300 ( \24426 , RIfca8a58_6941, \9437 );
and \U$15301 ( \24427 , RIfccad60_7330, \9439 );
and \U$15302 ( \24428 , RIfcac838_6985, \9441 );
and \U$15303 ( \24429 , RIfc67418_6197, \9443 );
and \U$15304 ( \24430 , RIf160340_5554, \9445 );
and \U$15305 ( \24431 , RIf15e450_5532, \9447 );
and \U$15306 ( \24432 , RIfe81a08_7819, \9449 );
and \U$15307 ( \24433 , RIfe81300_7814, \9451 );
and \U$15308 ( \24434 , RIfc6dac0_6270, \9453 );
and \U$15309 ( \24435 , RIf15ba20_5502, \9455 );
and \U$15310 ( \24436 , RIfc6d958_6269, \9457 );
and \U$15311 ( \24437 , RIfc6d7f0_6268, \9459 );
or \U$15312 ( \24438 , \24374 , \24375 , \24376 , \24377 , \24378 , \24379 , \24380 , \24381 , \24382 , \24383 , \24384 , \24385 , \24386 , \24387 , \24388 , \24389 , \24390 , \24391 , \24392 , \24393 , \24394 , \24395 , \24396 , \24397 , \24398 , \24399 , \24400 , \24401 , \24402 , \24403 , \24404 , \24405 , \24406 , \24407 , \24408 , \24409 , \24410 , \24411 , \24412 , \24413 , \24414 , \24415 , \24416 , \24417 , \24418 , \24419 , \24420 , \24421 , \24422 , \24423 , \24424 , \24425 , \24426 , \24427 , \24428 , \24429 , \24430 , \24431 , \24432 , \24433 , \24434 , \24435 , \24436 , \24437 );
and \U$15313 ( \24439 , RIfc587d8_6029, \9462 );
and \U$15314 ( \24440 , RIfc6cf80_6262, \9464 );
and \U$15315 ( \24441 , RIfc6d3b8_6265, \9466 );
and \U$15316 ( \24442 , RIfe815d0_7816, \9468 );
and \U$15317 ( \24443 , RIfc6d520_6266, \9470 );
and \U$15318 ( \24444 , RIfcabe60_6978, \9472 );
and \U$15319 ( \24445 , RIfc6d0e8_6263, \9474 );
and \U$15320 ( \24446 , RIe1f5780_4170, \9476 );
and \U$15321 ( \24447 , RIfc6c5a8_6255, \9478 );
and \U$15322 ( \24448 , RIfc68d68_6215, \9480 );
and \U$15323 ( \24449 , RIfc68c00_6214, \9482 );
and \U$15324 ( \24450 , RIe1f3458_4145, \9484 );
and \U$15325 ( \24451 , RIfc68a98_6213, \9486 );
and \U$15326 ( \24452 , RIfccb8a0_7338, \9488 );
and \U$15327 ( \24453 , RIfca9b38_6953, \9490 );
and \U$15328 ( \24454 , RIe1ee160_4086, \9492 );
and \U$15329 ( \24455 , RIe1eba00_4058, \9494 );
and \U$15330 ( \24456 , RIe1e8d00_4026, \9496 );
and \U$15331 ( \24457 , RIe1e6000_3994, \9498 );
and \U$15332 ( \24458 , RIe1e3300_3962, \9500 );
and \U$15333 ( \24459 , RIe1e0600_3930, \9502 );
and \U$15334 ( \24460 , RIe1dd900_3898, \9504 );
and \U$15335 ( \24461 , RIe1dac00_3866, \9506 );
and \U$15336 ( \24462 , RIe1d7f00_3834, \9508 );
and \U$15337 ( \24463 , RIe1d2500_3770, \9510 );
and \U$15338 ( \24464 , RIe1cf800_3738, \9512 );
and \U$15339 ( \24465 , RIe1ccb00_3706, \9514 );
and \U$15340 ( \24466 , RIe1c9e00_3674, \9516 );
and \U$15341 ( \24467 , RIe1c7100_3642, \9518 );
and \U$15342 ( \24468 , RIe1c4400_3610, \9520 );
and \U$15343 ( \24469 , RIe1c1700_3578, \9522 );
and \U$15344 ( \24470 , RIe1bea00_3546, \9524 );
and \U$15345 ( \24471 , RIfc6bbd0_6248, \9526 );
and \U$15346 ( \24472 , RIfcdd348_7539, \9528 );
and \U$15347 ( \24473 , RIe1b9438_3485, \9530 );
and \U$15348 ( \24474 , RIe1b73e0_3462, \9532 );
and \U$15349 ( \24475 , RIfcab5f0_6972, \9534 );
and \U$15350 ( \24476 , RIfccbb70_7340, \9536 );
and \U$15351 ( \24477 , RIe1b5220_3438, \9538 );
and \U$15352 ( \24478 , RIe1b3e70_3424, \9540 );
and \U$15353 ( \24479 , RIfc6c9e0_6258, \9542 );
and \U$15354 ( \24480 , RIfcab488_6971, \9544 );
and \U$15355 ( \24481 , RIfea7dc0_8226, \9546 );
and \U$15356 ( \24482 , RIe1b0bd0_3388, \9548 );
and \U$15357 ( \24483 , RIfc6ce18_6261, \9550 );
and \U$15358 ( \24484 , RIfcabfc8_6979, \9552 );
and \U$15359 ( \24485 , RIe1ac580_3338, \9554 );
and \U$15360 ( \24486 , RIe1aaf00_3322, \9556 );
and \U$15361 ( \24487 , RIe1a8d40_3298, \9558 );
and \U$15362 ( \24488 , RIe1a6040_3266, \9560 );
and \U$15363 ( \24489 , RIe1a3340_3234, \9562 );
and \U$15364 ( \24490 , RIe1a0640_3202, \9564 );
and \U$15365 ( \24491 , RIe18cb40_2978, \9566 );
and \U$15366 ( \24492 , RIe179040_2754, \9568 );
and \U$15367 ( \24493 , RIe226998_4729, \9570 );
and \U$15368 ( \24494 , RIe21b598_4601, \9572 );
and \U$15369 ( \24495 , RIe204d98_4345, \9574 );
and \U$15370 ( \24496 , RIe1fedf8_4277, \9576 );
and \U$15371 ( \24497 , RIe1f81b0_4200, \9578 );
and \U$15372 ( \24498 , RIe1f0cf8_4117, \9580 );
and \U$15373 ( \24499 , RIe1d5200_3802, \9582 );
and \U$15374 ( \24500 , RIe1bbd00_3514, \9584 );
and \U$15375 ( \24501 , RIe1aeb78_3365, \9586 );
and \U$15376 ( \24502 , RIe1711b0_2664, \9588 );
or \U$15377 ( \24503 , \24439 , \24440 , \24441 , \24442 , \24443 , \24444 , \24445 , \24446 , \24447 , \24448 , \24449 , \24450 , \24451 , \24452 , \24453 , \24454 , \24455 , \24456 , \24457 , \24458 , \24459 , \24460 , \24461 , \24462 , \24463 , \24464 , \24465 , \24466 , \24467 , \24468 , \24469 , \24470 , \24471 , \24472 , \24473 , \24474 , \24475 , \24476 , \24477 , \24478 , \24479 , \24480 , \24481 , \24482 , \24483 , \24484 , \24485 , \24486 , \24487 , \24488 , \24489 , \24490 , \24491 , \24492 , \24493 , \24494 , \24495 , \24496 , \24497 , \24498 , \24499 , \24500 , \24501 , \24502 );
or \U$15378 ( \24504 , \24438 , \24503 );
_DC g378a ( \24505_nG378a , \24504 , \9597 );
buf \U$15379 ( \24506 , \24505_nG378a );
xor \U$15380 ( \24507 , \24373 , \24506 );
and \U$15381 ( \24508 , RIdec5540_709, \9059 );
and \U$15382 ( \24509 , RIdec2840_677, \9061 );
and \U$15383 ( \24510 , RIfcc4dc0_7262, \9063 );
and \U$15384 ( \24511 , RIdebfb40_645, \9065 );
and \U$15385 ( \24512 , RIfc9d7c0_6814, \9067 );
and \U$15386 ( \24513 , RIdebce40_613, \9069 );
and \U$15387 ( \24514 , RIdeba140_581, \9071 );
and \U$15388 ( \24515 , RIdeb7440_549, \9073 );
and \U$15389 ( \24516 , RIfc4d978_5905, \9075 );
and \U$15390 ( \24517 , RIdeb1a40_485, \9077 );
and \U$15391 ( \24518 , RIfc9dbf8_6817, \9079 );
and \U$15392 ( \24519 , RIdeaed40_453, \9081 );
and \U$15393 ( \24520 , RIfcb8610_7120, \9083 );
and \U$15394 ( \24521 , RIdeaa768_421, \9085 );
and \U$15395 ( \24522 , RIdea3e68_389, \9087 );
and \U$15396 ( \24523 , RIde9d568_357, \9089 );
and \U$15397 ( \24524 , RIfc50678_5937, \9091 );
and \U$15398 ( \24525 , RIfc507e0_5938, \9093 );
and \U$15399 ( \24526 , RIfc9dec8_6819, \9095 );
and \U$15400 ( \24527 , RIfc853a0_6538, \9097 );
and \U$15401 ( \24528 , RIde913d0_298, \9099 );
and \U$15402 ( \24529 , RIde8dc08_281, \9101 );
and \U$15403 ( \24530 , RIde89a68_261, \9103 );
and \U$15404 ( \24531 , RIde858c8_241, \9105 );
and \U$15405 ( \24532 , RIde81a70_222, \9107 );
and \U$15406 ( \24533 , RIfc84860_6530, \9109 );
and \U$15407 ( \24534 , RIfc50948_5939, \9111 );
and \U$15408 ( \24535 , RIfc84c98_6533, \9113 );
and \U$15409 ( \24536 , RIfcb7da0_7114, \9115 );
and \U$15410 ( \24537 , RIe16b7b0_2600, \9117 );
and \U$15411 ( \24538 , RIe169b90_2580, \9119 );
and \U$15412 ( \24539 , RIe167e08_2559, \9121 );
and \U$15413 ( \24540 , RIe165540_2530, \9123 );
and \U$15414 ( \24541 , RIe162840_2498, \9125 );
and \U$15415 ( \24542 , RIee37528_5088, \9127 );
and \U$15416 ( \24543 , RIe15fb40_2466, \9129 );
and \U$15417 ( \24544 , RIfcb5be0_7090, \9131 );
and \U$15418 ( \24545 , RIe15ce40_2434, \9133 );
and \U$15419 ( \24546 , RIe157440_2370, \9135 );
and \U$15420 ( \24547 , RIe154740_2338, \9137 );
and \U$15421 ( \24548 , RIfcd35c8_7427, \9139 );
and \U$15422 ( \24549 , RIe151a40_2306, \9141 );
and \U$15423 ( \24550 , RIfc53a80_5974, \9143 );
and \U$15424 ( \24551 , RIe14ed40_2274, \9145 );
and \U$15425 ( \24552 , RIfcc6170_7276, \9147 );
and \U$15426 ( \24553 , RIe14c040_2242, \9149 );
and \U$15427 ( \24554 , RIe149340_2210, \9151 );
and \U$15428 ( \24555 , RIe146640_2178, \9153 );
and \U$15429 ( \24556 , RIfc7f130_6468, \9155 );
and \U$15430 ( \24557 , RIee33310_5041, \9157 );
and \U$15431 ( \24558 , RIfcb4f38_7081, \9159 );
and \U$15432 ( \24559 , RIfc47f78_5841, \9161 );
and \U$15433 ( \24560 , RIe140f10_2116, \9163 );
and \U$15434 ( \24561 , RIdf3ee18_2092, \9165 );
and \U$15435 ( \24562 , RIdf3cc58_2068, \9167 );
and \U$15436 ( \24563 , RIdf3a7c8_2042, \9169 );
and \U$15437 ( \24564 , RIfc7fc70_6476, \9171 );
and \U$15438 ( \24565 , RIfcd27b8_7417, \9173 );
and \U$15439 ( \24566 , RIfca1000_6854, \9175 );
and \U$15440 ( \24567 , RIfcc6b48_7283, \9177 );
and \U$15441 ( \24568 , RIdf35908_1986, \9179 );
and \U$15442 ( \24569 , RIdf33478_1960, \9181 );
and \U$15443 ( \24570 , RIfebe9f8_8289, \9183 );
and \U$15444 ( \24571 , RIdf2f260_1913, \9185 );
or \U$15445 ( \24572 , \24508 , \24509 , \24510 , \24511 , \24512 , \24513 , \24514 , \24515 , \24516 , \24517 , \24518 , \24519 , \24520 , \24521 , \24522 , \24523 , \24524 , \24525 , \24526 , \24527 , \24528 , \24529 , \24530 , \24531 , \24532 , \24533 , \24534 , \24535 , \24536 , \24537 , \24538 , \24539 , \24540 , \24541 , \24542 , \24543 , \24544 , \24545 , \24546 , \24547 , \24548 , \24549 , \24550 , \24551 , \24552 , \24553 , \24554 , \24555 , \24556 , \24557 , \24558 , \24559 , \24560 , \24561 , \24562 , \24563 , \24564 , \24565 , \24566 , \24567 , \24568 , \24569 , \24570 , \24571 );
and \U$15446 ( \24573 , RIfcb7968_7111, \9188 );
and \U$15447 ( \24574 , RIee2a3a0_4939, \9190 );
and \U$15448 ( \24575 , RIfc51050_5944, \9192 );
and \U$15449 ( \24576 , RIfcd3fa0_7434, \9194 );
and \U$15450 ( \24577 , RIdf2a3a0_1857, \9196 );
and \U$15451 ( \24578 , RIdf28078_1832, \9198 );
and \U$15452 ( \24579 , RIfe81198_7813, \9200 );
and \U$15453 ( \24580 , RIdf24838_1792, \9202 );
and \U$15454 ( \24581 , RIfc84428_6527, \9204 );
and \U$15455 ( \24582 , RIfce7ed8_7661, \9206 );
and \U$15456 ( \24583 , RIdf22d80_1773, \9208 );
and \U$15457 ( \24584 , RIfc515f0_5948, \9210 );
and \U$15458 ( \24585 , RIdf21868_1758, \9212 );
and \U$15459 ( \24586 , RIdf1f978_1736, \9214 );
and \U$15460 ( \24587 , RIdf1b058_1684, \9216 );
and \U$15461 ( \24588 , RIdf192d0_1663, \9218 );
and \U$15462 ( \24589 , RIdf17110_1639, \9220 );
and \U$15463 ( \24590 , RIdf14410_1607, \9222 );
and \U$15464 ( \24591 , RIdf11710_1575, \9224 );
and \U$15465 ( \24592 , RIdf0ea10_1543, \9226 );
and \U$15466 ( \24593 , RIdf0bd10_1511, \9228 );
and \U$15467 ( \24594 , RIdf09010_1479, \9230 );
and \U$15468 ( \24595 , RIdf06310_1447, \9232 );
and \U$15469 ( \24596 , RIdf03610_1415, \9234 );
and \U$15470 ( \24597 , RIdefdc10_1351, \9236 );
and \U$15471 ( \24598 , RIdefaf10_1319, \9238 );
and \U$15472 ( \24599 , RIdef8210_1287, \9240 );
and \U$15473 ( \24600 , RIdef5510_1255, \9242 );
and \U$15474 ( \24601 , RIdef2810_1223, \9244 );
and \U$15475 ( \24602 , RIdeefb10_1191, \9246 );
and \U$15476 ( \24603 , RIdeece10_1159, \9248 );
and \U$15477 ( \24604 , RIdeea110_1127, \9250 );
and \U$15478 ( \24605 , RIfc7e1b8_6457, \9252 );
and \U$15479 ( \24606 , RIfca19d8_6861, \9254 );
and \U$15480 ( \24607 , RIfc7dab0_6452, \9256 );
and \U$15481 ( \24608 , RIfc7e488_6459, \9258 );
and \U$15482 ( \24609 , RIdee49e0_1065, \9260 );
and \U$15483 ( \24610 , RIfe80d60_7810, \9262 );
and \U$15484 ( \24611 , RIfeabba0_8270, \9264 );
and \U$15485 ( \24612 , RIfe80bf8_7809, \9266 );
and \U$15486 ( \24613 , RIfcb3750_7064, \9268 );
and \U$15487 ( \24614 , RIfce9f30_7684, \9270 );
and \U$15488 ( \24615 , RIfc7e5f0_6460, \9272 );
and \U$15489 ( \24616 , RIfc56a50_6008, \9274 );
and \U$15490 ( \24617 , RIfe81030_7812, \9276 );
and \U$15491 ( \24618 , RIded7420_913, \9278 );
and \U$15492 ( \24619 , RIfe80ec8_7811, \9280 );
and \U$15493 ( \24620 , RIded2f38_864, \9282 );
and \U$15494 ( \24621 , RIded0940_837, \9284 );
and \U$15495 ( \24622 , RIdecdc40_805, \9286 );
and \U$15496 ( \24623 , RIdecaf40_773, \9288 );
and \U$15497 ( \24624 , RIdec8240_741, \9290 );
and \U$15498 ( \24625 , RIdeb4740_517, \9292 );
and \U$15499 ( \24626 , RIde96c68_325, \9294 );
and \U$15500 ( \24627 , RIe16e348_2631, \9296 );
and \U$15501 ( \24628 , RIe15a140_2402, \9298 );
and \U$15502 ( \24629 , RIe143940_2146, \9300 );
and \U$15503 ( \24630 , RIdf38338_2016, \9302 );
and \U$15504 ( \24631 , RIdf2c998_1884, \9304 );
and \U$15505 ( \24632 , RIdf1d218_1708, \9306 );
and \U$15506 ( \24633 , RIdf00910_1383, \9308 );
and \U$15507 ( \24634 , RIdee7410_1095, \9310 );
and \U$15508 ( \24635 , RIdedc178_968, \9312 );
and \U$15509 ( \24636 , RIde7cbb0_198, \9314 );
or \U$15510 ( \24637 , \24573 , \24574 , \24575 , \24576 , \24577 , \24578 , \24579 , \24580 , \24581 , \24582 , \24583 , \24584 , \24585 , \24586 , \24587 , \24588 , \24589 , \24590 , \24591 , \24592 , \24593 , \24594 , \24595 , \24596 , \24597 , \24598 , \24599 , \24600 , \24601 , \24602 , \24603 , \24604 , \24605 , \24606 , \24607 , \24608 , \24609 , \24610 , \24611 , \24612 , \24613 , \24614 , \24615 , \24616 , \24617 , \24618 , \24619 , \24620 , \24621 , \24622 , \24623 , \24624 , \24625 , \24626 , \24627 , \24628 , \24629 , \24630 , \24631 , \24632 , \24633 , \24634 , \24635 , \24636 );
or \U$15511 ( \24638 , \24572 , \24637 );
_DC g26e2 ( \24639_nG26e2 , \24638 , \9323 );
buf \U$15512 ( \24640 , \24639_nG26e2 );
and \U$15513 ( \24641 , RIe19d7d8_3169, \9333 );
and \U$15514 ( \24642 , RIe19aad8_3137, \9335 );
and \U$15515 ( \24643 , RIfcc2d68_7239, \9337 );
and \U$15516 ( \24644 , RIe197dd8_3105, \9339 );
and \U$15517 ( \24645 , RIfc5c5b8_6073, \9341 );
and \U$15518 ( \24646 , RIe1950d8_3073, \9343 );
and \U$15519 ( \24647 , RIe1923d8_3041, \9345 );
and \U$15520 ( \24648 , RIe18f6d8_3009, \9347 );
and \U$15521 ( \24649 , RIe189cd8_2945, \9349 );
and \U$15522 ( \24650 , RIe186fd8_2913, \9351 );
and \U$15523 ( \24651 , RIf1438d0_5228, \9353 );
and \U$15524 ( \24652 , RIe1842d8_2881, \9355 );
and \U$15525 ( \24653 , RIfc5b370_6060, \9357 );
and \U$15526 ( \24654 , RIe1815d8_2849, \9359 );
and \U$15527 ( \24655 , RIe17e8d8_2817, \9361 );
and \U$15528 ( \24656 , RIe17bbd8_2785, \9363 );
and \U$15529 ( \24657 , RIfcbb748_7155, \9365 );
and \U$15530 ( \24658 , RIfc59480_6038, \9367 );
and \U$15531 ( \24659 , RIfcbbce8_7159, \9369 );
and \U$15532 ( \24660 , RIe175c38_2717, \9371 );
and \U$15533 ( \24661 , RIfcdb890_7520, \9373 );
and \U$15534 ( \24662 , RIfc59b88_6043, \9375 );
and \U$15535 ( \24663 , RIfc8ada0_6602, \9377 );
and \U$15536 ( \24664 , RIfcb5eb0_7092, \9379 );
and \U$15537 ( \24665 , RIfc57c98_6021, \9381 );
and \U$15538 ( \24666 , RIfc57158_6013, \9383 );
and \U$15539 ( \24667 , RIfc58aa8_6031, \9385 );
and \U$15540 ( \24668 , RIe173910_2692, \9387 );
and \U$15541 ( \24669 , RIfcc62d8_7277, \9389 );
and \U$15542 ( \24670 , RIfc8a968_6599, \9391 );
and \U$15543 ( \24671 , RIfc57428_6015, \9393 );
and \U$15544 ( \24672 , RIfc56d20_6010, \9395 );
and \U$15545 ( \24673 , RIfc408e0_5760, \9397 );
and \U$15546 ( \24674 , RIe223b30_4696, \9399 );
and \U$15547 ( \24675 , RIfc82970_6508, \9401 );
and \U$15548 ( \24676 , RIe220e30_4664, \9403 );
and \U$15549 ( \24677 , RIfcecc30_7716, \9405 );
and \U$15550 ( \24678 , RIe21e130_4632, \9407 );
and \U$15551 ( \24679 , RIe218730_4568, \9409 );
and \U$15552 ( \24680 , RIe215a30_4536, \9411 );
and \U$15553 ( \24681 , RIfc3fad0_5750, \9413 );
and \U$15554 ( \24682 , RIe212d30_4504, \9415 );
and \U$15555 ( \24683 , RIf169148_5655, \9417 );
and \U$15556 ( \24684 , RIe210030_4472, \9419 );
and \U$15557 ( \24685 , RIfc545c0_5982, \9421 );
and \U$15558 ( \24686 , RIe20d330_4440, \9423 );
and \U$15559 ( \24687 , RIe20a630_4408, \9425 );
and \U$15560 ( \24688 , RIe207930_4376, \9427 );
and \U$15561 ( \24689 , RIfc88d48_6579, \9429 );
and \U$15562 ( \24690 , RIfc4bec0_5886, \9431 );
and \U$15563 ( \24691 , RIe202638_4317, \9433 );
and \U$15564 ( \24692 , RIe200b80_4298, \9435 );
and \U$15565 ( \24693 , RIfc88910_6576, \9437 );
and \U$15566 ( \24694 , RIfc4c190_5888, \9439 );
and \U$15567 ( \24695 , RIfc4c2f8_5889, \9441 );
and \U$15568 ( \24696 , RIfcba398_7141, \9443 );
and \U$15569 ( \24697 , RIfcd4270_7436, \9445 );
and \U$15570 ( \24698 , RIfcba0c8_7139, \9447 );
and \U$15571 ( \24699 , RIe1fcda0_4254, \9449 );
and \U$15572 ( \24700 , RIe1fbb58_4241, \9451 );
and \U$15573 ( \24701 , RIfc53d50_5976, \9453 );
and \U$15574 ( \24702 , RIfc9b768_6791, \9455 );
and \U$15575 ( \24703 , RIfc537b0_5972, \9457 );
and \U$15576 ( \24704 , RIfc4c5c8_5891, \9459 );
or \U$15577 ( \24705 , \24641 , \24642 , \24643 , \24644 , \24645 , \24646 , \24647 , \24648 , \24649 , \24650 , \24651 , \24652 , \24653 , \24654 , \24655 , \24656 , \24657 , \24658 , \24659 , \24660 , \24661 , \24662 , \24663 , \24664 , \24665 , \24666 , \24667 , \24668 , \24669 , \24670 , \24671 , \24672 , \24673 , \24674 , \24675 , \24676 , \24677 , \24678 , \24679 , \24680 , \24681 , \24682 , \24683 , \24684 , \24685 , \24686 , \24687 , \24688 , \24689 , \24690 , \24691 , \24692 , \24693 , \24694 , \24695 , \24696 , \24697 , \24698 , \24699 , \24700 , \24701 , \24702 , \24703 , \24704 );
and \U$15578 ( \24706 , RIfc9e468_6823, \9462 );
and \U$15579 ( \24707 , RIf157da8_5459, \9464 );
and \U$15580 ( \24708 , RIfcb9f60_7138, \9466 );
and \U$15581 ( \24709 , RIe1fa208_4223, \9468 );
and \U$15582 ( \24710 , RIfc849c8_6531, \9470 );
and \U$15583 ( \24711 , RIfc529a0_5962, \9472 );
and \U$15584 ( \24712 , RIfc9f6b0_6836, \9474 );
and \U$15585 ( \24713 , RIe1f5618_4169, \9476 );
and \U$15586 ( \24714 , RIf153320_5406, \9478 );
and \U$15587 ( \24715 , RIfcc4988_7259, \9480 );
and \U$15588 ( \24716 , RIf150d28_5379, \9482 );
and \U$15589 ( \24717 , RIfebe458_8285, \9484 );
and \U$15590 ( \24718 , RIfc87f38_6569, \9486 );
and \U$15591 ( \24719 , RIfcb7f08_7115, \9488 );
and \U$15592 ( \24720 , RIf14e190_5348, \9490 );
and \U$15593 ( \24721 , RIfe80658_7805, \9492 );
and \U$15594 ( \24722 , RIe1eb898_4057, \9494 );
and \U$15595 ( \24723 , RIe1e8b98_4025, \9496 );
and \U$15596 ( \24724 , RIe1e5e98_3993, \9498 );
and \U$15597 ( \24725 , RIe1e3198_3961, \9500 );
and \U$15598 ( \24726 , RIe1e0498_3929, \9502 );
and \U$15599 ( \24727 , RIe1dd798_3897, \9504 );
and \U$15600 ( \24728 , RIe1daa98_3865, \9506 );
and \U$15601 ( \24729 , RIe1d7d98_3833, \9508 );
and \U$15602 ( \24730 , RIe1d2398_3769, \9510 );
and \U$15603 ( \24731 , RIe1cf698_3737, \9512 );
and \U$15604 ( \24732 , RIe1cc998_3705, \9514 );
and \U$15605 ( \24733 , RIe1c9c98_3673, \9516 );
and \U$15606 ( \24734 , RIe1c6f98_3641, \9518 );
and \U$15607 ( \24735 , RIe1c4298_3609, \9520 );
and \U$15608 ( \24736 , RIe1c1598_3577, \9522 );
and \U$15609 ( \24737 , RIe1be898_3545, \9524 );
and \U$15610 ( \24738 , RIf14cc78_5333, \9526 );
and \U$15611 ( \24739 , RIf14ba30_5320, \9528 );
and \U$15612 ( \24740 , RIe1b92d0_3484, \9530 );
and \U$15613 ( \24741 , RIe1b7278_3461, \9532 );
and \U$15614 ( \24742 , RIf14a7e8_5307, \9534 );
and \U$15615 ( \24743 , RIf149ca8_5299, \9536 );
and \U$15616 ( \24744 , RIfebe5c0_8286, \9538 );
and \U$15617 ( \24745 , RIfe807c0_7806, \9540 );
and \U$15618 ( \24746 , RIfc50510_5936, \9542 );
and \U$15619 ( \24747 , RIfce4f08_7627, \9544 );
and \U$15620 ( \24748 , RIfe80a90_7808, \9546 );
and \U$15621 ( \24749 , RIfebe890_8288, \9548 );
and \U$15622 ( \24750 , RIfc9cde8_6807, \9550 );
and \U$15623 ( \24751 , RIfc87560_6562, \9552 );
and \U$15624 ( \24752 , RIfe80928_7807, \9554 );
and \U$15625 ( \24753 , RIfebe728_8287, \9556 );
and \U$15626 ( \24754 , RIe1a8bd8_3297, \9558 );
and \U$15627 ( \24755 , RIe1a5ed8_3265, \9560 );
and \U$15628 ( \24756 , RIe1a31d8_3233, \9562 );
and \U$15629 ( \24757 , RIe1a04d8_3201, \9564 );
and \U$15630 ( \24758 , RIe18c9d8_2977, \9566 );
and \U$15631 ( \24759 , RIe178ed8_2753, \9568 );
and \U$15632 ( \24760 , RIe226830_4728, \9570 );
and \U$15633 ( \24761 , RIe21b430_4600, \9572 );
and \U$15634 ( \24762 , RIe204c30_4344, \9574 );
and \U$15635 ( \24763 , RIe1fec90_4276, \9576 );
and \U$15636 ( \24764 , RIe1f8048_4199, \9578 );
and \U$15637 ( \24765 , RIe1f0b90_4116, \9580 );
and \U$15638 ( \24766 , RIe1d5098_3801, \9582 );
and \U$15639 ( \24767 , RIe1bbb98_3513, \9584 );
and \U$15640 ( \24768 , RIe1aea10_3364, \9586 );
and \U$15641 ( \24769 , RIe171048_2663, \9588 );
or \U$15642 ( \24770 , \24706 , \24707 , \24708 , \24709 , \24710 , \24711 , \24712 , \24713 , \24714 , \24715 , \24716 , \24717 , \24718 , \24719 , \24720 , \24721 , \24722 , \24723 , \24724 , \24725 , \24726 , \24727 , \24728 , \24729 , \24730 , \24731 , \24732 , \24733 , \24734 , \24735 , \24736 , \24737 , \24738 , \24739 , \24740 , \24741 , \24742 , \24743 , \24744 , \24745 , \24746 , \24747 , \24748 , \24749 , \24750 , \24751 , \24752 , \24753 , \24754 , \24755 , \24756 , \24757 , \24758 , \24759 , \24760 , \24761 , \24762 , \24763 , \24764 , \24765 , \24766 , \24767 , \24768 , \24769 );
or \U$15643 ( \24771 , \24705 , \24770 );
_DC g380f ( \24772_nG380f , \24771 , \9597 );
buf \U$15644 ( \24773 , \24772_nG380f );
and \U$15645 ( \24774 , \24640 , \24773 );
and \U$15646 ( \24775 , \22782 , \22915 );
and \U$15647 ( \24776 , \22915 , \23190 );
and \U$15648 ( \24777 , \22782 , \23190 );
or \U$15649 ( \24778 , \24775 , \24776 , \24777 );
and \U$15650 ( \24779 , \24773 , \24778 );
and \U$15651 ( \24780 , \24640 , \24778 );
or \U$15652 ( \24781 , \24774 , \24779 , \24780 );
xor \U$15653 ( \24782 , \24507 , \24781 );
buf g4412 ( \24783_nG4412 , \24782 );
xor \U$15654 ( \24784 , \24640 , \24773 );
xor \U$15655 ( \24785 , \24784 , \24778 );
buf g4415 ( \24786_nG4415 , \24785 );
nand \U$15656 ( \24787 , \24786_nG4415 , \23192_nG4418 );
and \U$15657 ( \24788 , \24783_nG4412 , \24787 );
xor \U$15658 ( \24789 , \24786_nG4415 , \23192_nG4418 );
not \U$15659 ( \24790 , \24789 );
xor \U$15660 ( \24791 , \24783_nG4412 , \24786_nG4415 );
and \U$15661 ( \24792 , \24790 , \24791 );
and \U$15663 ( \24793 , \24789 , \10694_nG9c0e );
or \U$15664 ( \24794 , 1'b0 , \24793 );
xor \U$15665 ( \24795 , \24788 , \24794 );
xor \U$15666 ( \24796 , \24788 , \24795 );
buf \U$15667 ( \24797 , \24796 );
buf \U$15668 ( \24798 , \24797 );
xor \U$15669 ( \24799 , \24240 , \24798 );
and \U$15670 ( \24800 , \23736 , \23741 );
and \U$15671 ( \24801 , \23736 , \23747 );
and \U$15672 ( \24802 , \23741 , \23747 );
or \U$15673 ( \24803 , \24800 , \24801 , \24802 );
buf \U$15674 ( \24804 , \24803 );
and \U$15675 ( \24805 , \23826 , \23832 );
and \U$15676 ( \24806 , \23826 , \23839 );
and \U$15677 ( \24807 , \23832 , \23839 );
or \U$15678 ( \24808 , \24805 , \24806 , \24807 );
buf \U$15679 ( \24809 , \24808 );
and \U$15680 ( \24810 , \23802 , \23808 );
and \U$15681 ( \24811 , \23802 , \23815 );
and \U$15682 ( \24812 , \23808 , \23815 );
or \U$15683 ( \24813 , \24810 , \24811 , \24812 );
buf \U$15684 ( \24814 , \24813 );
and \U$15685 ( \24815 , \23201 , \10995_nG9c0b );
and \U$15686 ( \24816 , \23198 , \11283_nG9c08 );
or \U$15687 ( \24817 , \24815 , \24816 );
xor \U$15688 ( \24818 , \23197 , \24817 );
buf \U$15689 ( \24819 , \24818 );
buf \U$15691 ( \24820 , \24819 );
and \U$15692 ( \24821 , \21658 , \11598_nG9c05 );
and \U$15693 ( \24822 , \21655 , \12470_nG9c02 );
or \U$15694 ( \24823 , \24821 , \24822 );
xor \U$15695 ( \24824 , \21654 , \24823 );
buf \U$15696 ( \24825 , \24824 );
buf \U$15698 ( \24826 , \24825 );
xor \U$15699 ( \24827 , \24820 , \24826 );
buf \U$15700 ( \24828 , \24827 );
xor \U$15701 ( \24829 , \24814 , \24828 );
and \U$15702 ( \24830 , \17297 , \15373_nG9bf3 );
and \U$15703 ( \24831 , \17294 , \16315_nG9bf0 );
or \U$15704 ( \24832 , \24830 , \24831 );
xor \U$15705 ( \24833 , \17293 , \24832 );
buf \U$15706 ( \24834 , \24833 );
buf \U$15708 ( \24835 , \24834 );
xor \U$15709 ( \24836 , \24829 , \24835 );
buf \U$15710 ( \24837 , \24836 );
and \U$15711 ( \24838 , \23762 , \23768 );
and \U$15712 ( \24839 , \23762 , \23775 );
and \U$15713 ( \24840 , \23768 , \23775 );
or \U$15714 ( \24841 , \24838 , \24839 , \24840 );
buf \U$15715 ( \24842 , \24841 );
xor \U$15716 ( \24843 , \24837 , \24842 );
and \U$15717 ( \24844 , \12157 , \21086_nG9bdb );
and \U$15718 ( \24845 , \12154 , \22129_nG9bd8 );
or \U$15719 ( \24846 , \24844 , \24845 );
xor \U$15720 ( \24847 , \12153 , \24846 );
buf \U$15721 ( \24848 , \24847 );
buf \U$15723 ( \24849 , \24848 );
xor \U$15724 ( \24850 , \24843 , \24849 );
buf \U$15725 ( \24851 , \24850 );
xor \U$15726 ( \24852 , \24809 , \24851 );
and \U$15727 ( \24853 , \23760 , \23777 );
and \U$15728 ( \24854 , \23760 , \23784 );
and \U$15729 ( \24855 , \23777 , \23784 );
or \U$15730 ( \24856 , \24853 , \24854 , \24855 );
buf \U$15731 ( \24857 , \24856 );
and \U$15732 ( \24858 , \23791 , \23817 );
and \U$15733 ( \24859 , \23791 , \23824 );
and \U$15734 ( \24860 , \23817 , \23824 );
or \U$15735 ( \24861 , \24858 , \24859 , \24860 );
buf \U$15736 ( \24862 , \24861 );
xor \U$15737 ( \24863 , \24857 , \24862 );
and \U$15738 ( \24864 , \13370 , \19586_nG9be1 );
and \U$15739 ( \24865 , \13367 , \20608_nG9bde );
or \U$15740 ( \24866 , \24864 , \24865 );
xor \U$15741 ( \24867 , \13366 , \24866 );
buf \U$15742 ( \24868 , \24867 );
buf \U$15744 ( \24869 , \24868 );
xor \U$15745 ( \24870 , \24863 , \24869 );
buf \U$15746 ( \24871 , \24870 );
xor \U$15747 ( \24872 , \24852 , \24871 );
buf \U$15748 ( \24873 , \24872 );
xor \U$15749 ( \24874 , \24804 , \24873 );
and \U$15750 ( \24875 , \23722 , \23727 );
and \U$15751 ( \24876 , \23722 , \23734 );
and \U$15752 ( \24877 , \23727 , \23734 );
or \U$15753 ( \24878 , \24875 , \24876 , \24877 );
buf \U$15754 ( \24879 , \24878 );
and \U$15755 ( \24880 , \23794 , \23800 );
buf \U$15756 ( \24881 , \24880 );
and \U$15757 ( \24882 , \20155 , \12801_nG9bff );
and \U$15758 ( \24883 , \20152 , \13705_nG9bfc );
or \U$15759 ( \24884 , \24882 , \24883 );
xor \U$15760 ( \24885 , \20151 , \24884 );
buf \U$15761 ( \24886 , \24885 );
buf \U$15763 ( \24887 , \24886 );
xor \U$15764 ( \24888 , \24881 , \24887 );
and \U$15765 ( \24889 , \18702 , \14070_nG9bf9 );
and \U$15766 ( \24890 , \18699 , \14984_nG9bf6 );
or \U$15767 ( \24891 , \24889 , \24890 );
xor \U$15768 ( \24892 , \18698 , \24891 );
buf \U$15769 ( \24893 , \24892 );
buf \U$15771 ( \24894 , \24893 );
xor \U$15772 ( \24895 , \24888 , \24894 );
buf \U$15773 ( \24896 , \24895 );
and \U$15774 ( \24897 , \15940 , \16680_nG9bed );
and \U$15775 ( \24898 , \15937 , \17665_nG9bea );
or \U$15776 ( \24899 , \24897 , \24898 );
xor \U$15777 ( \24900 , \15936 , \24899 );
buf \U$15778 ( \24901 , \24900 );
buf \U$15780 ( \24902 , \24901 );
xor \U$15781 ( \24903 , \24896 , \24902 );
and \U$15782 ( \24904 , \14631 , \18107_nG9be7 );
and \U$15783 ( \24905 , \14628 , \19091_nG9be4 );
or \U$15784 ( \24906 , \24904 , \24905 );
xor \U$15785 ( \24907 , \14627 , \24906 );
buf \U$15786 ( \24908 , \24907 );
buf \U$15788 ( \24909 , \24908 );
xor \U$15789 ( \24910 , \24903 , \24909 );
buf \U$15790 ( \24911 , \24910 );
and \U$15791 ( \24912 , \10421 , \22629_nG9bd5 );
and \U$15792 ( \24913 , \10418 , \23696_nG9bd2 );
or \U$15793 ( \24914 , \24912 , \24913 );
xor \U$15794 ( \24915 , \10417 , \24914 );
buf \U$15795 ( \24916 , \24915 );
buf \U$15797 ( \24917 , \24916 );
xor \U$15798 ( \24918 , \24911 , \24917 );
and \U$15799 ( \24919 , \10707 , \24226_nG9bcf );
and \U$15800 ( \24920 , \23856 , \24162 );
and \U$15801 ( \24921 , \24162 , \24214 );
and \U$15802 ( \24922 , \23856 , \24214 );
or \U$15803 ( \24923 , \24920 , \24921 , \24922 );
and \U$15804 ( \24924 , \24189 , \24193 );
and \U$15805 ( \24925 , \24193 , \24212 );
and \U$15806 ( \24926 , \24189 , \24212 );
or \U$15807 ( \24927 , \24924 , \24925 , \24926 );
and \U$15808 ( \24928 , \23860 , \24146 );
and \U$15809 ( \24929 , \24146 , \24161 );
and \U$15810 ( \24930 , \23860 , \24161 );
or \U$15811 ( \24931 , \24928 , \24929 , \24930 );
xor \U$15812 ( \24932 , \24927 , \24931 );
and \U$15813 ( \24933 , \24202 , \24206 );
and \U$15814 ( \24934 , \24206 , \24211 );
and \U$15815 ( \24935 , \24202 , \24211 );
or \U$15816 ( \24936 , \24933 , \24934 , \24935 );
and \U$15817 ( \24937 , \23864 , \23868 );
and \U$15818 ( \24938 , \23868 , \24145 );
and \U$15819 ( \24939 , \23864 , \24145 );
or \U$15820 ( \24940 , \24937 , \24938 , \24939 );
xor \U$15821 ( \24941 , \24936 , \24940 );
and \U$15822 ( \24942 , \24171 , \24173 );
xor \U$15823 ( \24943 , \24941 , \24942 );
xor \U$15824 ( \24944 , \24932 , \24943 );
xor \U$15825 ( \24945 , \24923 , \24944 );
and \U$15826 ( \24946 , \24167 , \24184 );
and \U$15827 ( \24947 , \24184 , \24213 );
and \U$15828 ( \24948 , \24167 , \24213 );
or \U$15829 ( \24949 , \24946 , \24947 , \24948 );
and \U$15830 ( \24950 , \24151 , \24155 );
and \U$15831 ( \24951 , \24155 , \24160 );
and \U$15832 ( \24952 , \24151 , \24160 );
or \U$15833 ( \24953 , \24950 , \24951 , \24952 );
and \U$15834 ( \24954 , \18035 , \15336 );
and \U$15835 ( \24955 , \19032 , \14963 );
nor \U$15836 ( \24956 , \24954 , \24955 );
xnor \U$15837 ( \24957 , \24956 , \15342 );
and \U$15838 ( \24958 , \14024 , \19534 );
and \U$15839 ( \24959 , \14950 , \19045 );
nor \U$15840 ( \24960 , \24958 , \24959 );
xnor \U$15841 ( \24961 , \24960 , \19540 );
xor \U$15842 ( \24962 , \24957 , \24961 );
and \U$15843 ( \24963 , \12769 , \21005 );
and \U$15844 ( \24964 , \13679 , \20557 );
nor \U$15845 ( \24965 , \24963 , \24964 );
xnor \U$15846 ( \24966 , \24965 , \21011 );
xor \U$15847 ( \24967 , \24962 , \24966 );
xor \U$15848 ( \24968 , \24953 , \24967 );
and \U$15849 ( \24969 , \21033 , \12790 );
and \U$15850 ( \24970 , \22090 , \12461 );
nor \U$15851 ( \24971 , \24969 , \24970 );
xnor \U$15852 ( \24972 , \24971 , \12780 );
and \U$15853 ( \24973 , \16655 , \16635 );
and \U$15854 ( \24974 , \17627 , \16301 );
nor \U$15855 ( \24975 , \24973 , \24974 );
xnor \U$15856 ( \24976 , \24975 , \16625 );
xor \U$15857 ( \24977 , \24972 , \24976 );
and \U$15858 ( \24978 , \15321 , \18090 );
and \U$15859 ( \24979 , \16267 , \17655 );
nor \U$15860 ( \24980 , \24978 , \24979 );
xnor \U$15861 ( \24981 , \24980 , \18046 );
xor \U$15862 ( \24982 , \24977 , \24981 );
xor \U$15863 ( \24983 , \24968 , \24982 );
xor \U$15864 ( \24984 , \24949 , \24983 );
and \U$15865 ( \24985 , \24174 , \24178 );
and \U$15866 ( \24986 , \24178 , \24183 );
and \U$15867 ( \24987 , \24174 , \24183 );
or \U$15868 ( \24988 , \24985 , \24986 , \24987 );
and \U$15869 ( \24989 , \22556 , \11574 );
and \U$15870 ( \24990 , \23617 , \11278 );
nor \U$15871 ( \24991 , \24989 , \24990 );
xnor \U$15872 ( \24992 , \24991 , \11580 );
and \U$15873 ( \24993 , \19558 , \14054 );
and \U$15874 ( \24994 , \20544 , \13692 );
nor \U$15875 ( \24995 , \24993 , \24994 );
xnor \U$15876 ( \24996 , \24995 , \14035 );
xor \U$15877 ( \24997 , \24992 , \24996 );
and \U$15878 ( \24998 , RIdec5540_709, \9333 );
and \U$15879 ( \24999 , RIdec2840_677, \9335 );
and \U$15880 ( \25000 , RIfcc4dc0_7262, \9337 );
and \U$15881 ( \25001 , RIdebfb40_645, \9339 );
and \U$15882 ( \25002 , RIfc9d7c0_6814, \9341 );
and \U$15883 ( \25003 , RIdebce40_613, \9343 );
and \U$15884 ( \25004 , RIdeba140_581, \9345 );
and \U$15885 ( \25005 , RIdeb7440_549, \9347 );
and \U$15886 ( \25006 , RIfc4d978_5905, \9349 );
and \U$15887 ( \25007 , RIdeb1a40_485, \9351 );
and \U$15888 ( \25008 , RIfc9dbf8_6817, \9353 );
and \U$15889 ( \25009 , RIdeaed40_453, \9355 );
and \U$15890 ( \25010 , RIfcb8610_7120, \9357 );
and \U$15891 ( \25011 , RIdeaa768_421, \9359 );
and \U$15892 ( \25012 , RIdea3e68_389, \9361 );
and \U$15893 ( \25013 , RIde9d568_357, \9363 );
and \U$15894 ( \25014 , RIfc50678_5937, \9365 );
and \U$15895 ( \25015 , RIfc507e0_5938, \9367 );
and \U$15896 ( \25016 , RIfc9dec8_6819, \9369 );
and \U$15897 ( \25017 , RIfc853a0_6538, \9371 );
and \U$15898 ( \25018 , RIde913d0_298, \9373 );
and \U$15899 ( \25019 , RIde8dc08_281, \9375 );
and \U$15900 ( \25020 , RIde89a68_261, \9377 );
and \U$15901 ( \25021 , RIde858c8_241, \9379 );
and \U$15902 ( \25022 , RIde81a70_222, \9381 );
and \U$15903 ( \25023 , RIfc84860_6530, \9383 );
and \U$15904 ( \25024 , RIfc50948_5939, \9385 );
and \U$15905 ( \25025 , RIfc84c98_6533, \9387 );
and \U$15906 ( \25026 , RIfcb7da0_7114, \9389 );
and \U$15907 ( \25027 , RIe16b7b0_2600, \9391 );
and \U$15908 ( \25028 , RIe169b90_2580, \9393 );
and \U$15909 ( \25029 , RIe167e08_2559, \9395 );
and \U$15910 ( \25030 , RIe165540_2530, \9397 );
and \U$15911 ( \25031 , RIe162840_2498, \9399 );
and \U$15912 ( \25032 , RIee37528_5088, \9401 );
and \U$15913 ( \25033 , RIe15fb40_2466, \9403 );
and \U$15914 ( \25034 , RIfcb5be0_7090, \9405 );
and \U$15915 ( \25035 , RIe15ce40_2434, \9407 );
and \U$15916 ( \25036 , RIe157440_2370, \9409 );
and \U$15917 ( \25037 , RIe154740_2338, \9411 );
and \U$15918 ( \25038 , RIfcd35c8_7427, \9413 );
and \U$15919 ( \25039 , RIe151a40_2306, \9415 );
and \U$15920 ( \25040 , RIfc53a80_5974, \9417 );
and \U$15921 ( \25041 , RIe14ed40_2274, \9419 );
and \U$15922 ( \25042 , RIfcc6170_7276, \9421 );
and \U$15923 ( \25043 , RIe14c040_2242, \9423 );
and \U$15924 ( \25044 , RIe149340_2210, \9425 );
and \U$15925 ( \25045 , RIe146640_2178, \9427 );
and \U$15926 ( \25046 , RIfc7f130_6468, \9429 );
and \U$15927 ( \25047 , RIee33310_5041, \9431 );
and \U$15928 ( \25048 , RIfcb4f38_7081, \9433 );
and \U$15929 ( \25049 , RIfc47f78_5841, \9435 );
and \U$15930 ( \25050 , RIe140f10_2116, \9437 );
and \U$15931 ( \25051 , RIdf3ee18_2092, \9439 );
and \U$15932 ( \25052 , RIdf3cc58_2068, \9441 );
and \U$15933 ( \25053 , RIdf3a7c8_2042, \9443 );
and \U$15934 ( \25054 , RIfc7fc70_6476, \9445 );
and \U$15935 ( \25055 , RIfcd27b8_7417, \9447 );
and \U$15936 ( \25056 , RIfca1000_6854, \9449 );
and \U$15937 ( \25057 , RIfcc6b48_7283, \9451 );
and \U$15938 ( \25058 , RIdf35908_1986, \9453 );
and \U$15939 ( \25059 , RIdf33478_1960, \9455 );
and \U$15940 ( \25060 , RIfebe9f8_8289, \9457 );
and \U$15941 ( \25061 , RIdf2f260_1913, \9459 );
or \U$15942 ( \25062 , \24998 , \24999 , \25000 , \25001 , \25002 , \25003 , \25004 , \25005 , \25006 , \25007 , \25008 , \25009 , \25010 , \25011 , \25012 , \25013 , \25014 , \25015 , \25016 , \25017 , \25018 , \25019 , \25020 , \25021 , \25022 , \25023 , \25024 , \25025 , \25026 , \25027 , \25028 , \25029 , \25030 , \25031 , \25032 , \25033 , \25034 , \25035 , \25036 , \25037 , \25038 , \25039 , \25040 , \25041 , \25042 , \25043 , \25044 , \25045 , \25046 , \25047 , \25048 , \25049 , \25050 , \25051 , \25052 , \25053 , \25054 , \25055 , \25056 , \25057 , \25058 , \25059 , \25060 , \25061 );
and \U$15943 ( \25063 , RIfcb7968_7111, \9462 );
and \U$15944 ( \25064 , RIee2a3a0_4939, \9464 );
and \U$15945 ( \25065 , RIfc51050_5944, \9466 );
and \U$15946 ( \25066 , RIfcd3fa0_7434, \9468 );
and \U$15947 ( \25067 , RIdf2a3a0_1857, \9470 );
and \U$15948 ( \25068 , RIdf28078_1832, \9472 );
and \U$15949 ( \25069 , RIfe81198_7813, \9474 );
and \U$15950 ( \25070 , RIdf24838_1792, \9476 );
and \U$15951 ( \25071 , RIfc84428_6527, \9478 );
and \U$15952 ( \25072 , RIfce7ed8_7661, \9480 );
and \U$15953 ( \25073 , RIdf22d80_1773, \9482 );
and \U$15954 ( \25074 , RIfc515f0_5948, \9484 );
and \U$15955 ( \25075 , RIdf21868_1758, \9486 );
and \U$15956 ( \25076 , RIdf1f978_1736, \9488 );
and \U$15957 ( \25077 , RIdf1b058_1684, \9490 );
and \U$15958 ( \25078 , RIdf192d0_1663, \9492 );
and \U$15959 ( \25079 , RIdf17110_1639, \9494 );
and \U$15960 ( \25080 , RIdf14410_1607, \9496 );
and \U$15961 ( \25081 , RIdf11710_1575, \9498 );
and \U$15962 ( \25082 , RIdf0ea10_1543, \9500 );
and \U$15963 ( \25083 , RIdf0bd10_1511, \9502 );
and \U$15964 ( \25084 , RIdf09010_1479, \9504 );
and \U$15965 ( \25085 , RIdf06310_1447, \9506 );
and \U$15966 ( \25086 , RIdf03610_1415, \9508 );
and \U$15967 ( \25087 , RIdefdc10_1351, \9510 );
and \U$15968 ( \25088 , RIdefaf10_1319, \9512 );
and \U$15969 ( \25089 , RIdef8210_1287, \9514 );
and \U$15970 ( \25090 , RIdef5510_1255, \9516 );
and \U$15971 ( \25091 , RIdef2810_1223, \9518 );
and \U$15972 ( \25092 , RIdeefb10_1191, \9520 );
and \U$15973 ( \25093 , RIdeece10_1159, \9522 );
and \U$15974 ( \25094 , RIdeea110_1127, \9524 );
and \U$15975 ( \25095 , RIfc7e1b8_6457, \9526 );
and \U$15976 ( \25096 , RIfca19d8_6861, \9528 );
and \U$15977 ( \25097 , RIfc7dab0_6452, \9530 );
and \U$15978 ( \25098 , RIfc7e488_6459, \9532 );
and \U$15979 ( \25099 , RIdee49e0_1065, \9534 );
and \U$15980 ( \25100 , RIfe80d60_7810, \9536 );
and \U$15981 ( \25101 , RIfeabba0_8270, \9538 );
and \U$15982 ( \25102 , RIfe80bf8_7809, \9540 );
and \U$15983 ( \25103 , RIfcb3750_7064, \9542 );
and \U$15984 ( \25104 , RIfce9f30_7684, \9544 );
and \U$15985 ( \25105 , RIfc7e5f0_6460, \9546 );
and \U$15986 ( \25106 , RIfc56a50_6008, \9548 );
and \U$15987 ( \25107 , RIfe81030_7812, \9550 );
and \U$15988 ( \25108 , RIded7420_913, \9552 );
and \U$15989 ( \25109 , RIfe80ec8_7811, \9554 );
and \U$15990 ( \25110 , RIded2f38_864, \9556 );
and \U$15991 ( \25111 , RIded0940_837, \9558 );
and \U$15992 ( \25112 , RIdecdc40_805, \9560 );
and \U$15993 ( \25113 , RIdecaf40_773, \9562 );
and \U$15994 ( \25114 , RIdec8240_741, \9564 );
and \U$15995 ( \25115 , RIdeb4740_517, \9566 );
and \U$15996 ( \25116 , RIde96c68_325, \9568 );
and \U$15997 ( \25117 , RIe16e348_2631, \9570 );
and \U$15998 ( \25118 , RIe15a140_2402, \9572 );
and \U$15999 ( \25119 , RIe143940_2146, \9574 );
and \U$16000 ( \25120 , RIdf38338_2016, \9576 );
and \U$16001 ( \25121 , RIdf2c998_1884, \9578 );
and \U$16002 ( \25122 , RIdf1d218_1708, \9580 );
and \U$16003 ( \25123 , RIdf00910_1383, \9582 );
and \U$16004 ( \25124 , RIdee7410_1095, \9584 );
and \U$16005 ( \25125 , RIdedc178_968, \9586 );
and \U$16006 ( \25126 , RIde7cbb0_198, \9588 );
or \U$16007 ( \25127 , \25063 , \25064 , \25065 , \25066 , \25067 , \25068 , \25069 , \25070 , \25071 , \25072 , \25073 , \25074 , \25075 , \25076 , \25077 , \25078 , \25079 , \25080 , \25081 , \25082 , \25083 , \25084 , \25085 , \25086 , \25087 , \25088 , \25089 , \25090 , \25091 , \25092 , \25093 , \25094 , \25095 , \25096 , \25097 , \25098 , \25099 , \25100 , \25101 , \25102 , \25103 , \25104 , \25105 , \25106 , \25107 , \25108 , \25109 , \25110 , \25111 , \25112 , \25113 , \25114 , \25115 , \25116 , \25117 , \25118 , \25119 , \25120 , \25121 , \25122 , \25123 , \25124 , \25125 , \25126 );
or \U$16008 ( \25128 , \25062 , \25127 );
_DC g5ba0 ( \25129_nG5ba0 , \25128 , \9597 );
and \U$16009 ( \25130 , RIe19d7d8_3169, \9059 );
and \U$16010 ( \25131 , RIe19aad8_3137, \9061 );
and \U$16011 ( \25132 , RIfcc2d68_7239, \9063 );
and \U$16012 ( \25133 , RIe197dd8_3105, \9065 );
and \U$16013 ( \25134 , RIfc5c5b8_6073, \9067 );
and \U$16014 ( \25135 , RIe1950d8_3073, \9069 );
and \U$16015 ( \25136 , RIe1923d8_3041, \9071 );
and \U$16016 ( \25137 , RIe18f6d8_3009, \9073 );
and \U$16017 ( \25138 , RIe189cd8_2945, \9075 );
and \U$16018 ( \25139 , RIe186fd8_2913, \9077 );
and \U$16019 ( \25140 , RIf1438d0_5228, \9079 );
and \U$16020 ( \25141 , RIe1842d8_2881, \9081 );
and \U$16021 ( \25142 , RIfc5b370_6060, \9083 );
and \U$16022 ( \25143 , RIe1815d8_2849, \9085 );
and \U$16023 ( \25144 , RIe17e8d8_2817, \9087 );
and \U$16024 ( \25145 , RIe17bbd8_2785, \9089 );
and \U$16025 ( \25146 , RIfcbb748_7155, \9091 );
and \U$16026 ( \25147 , RIfc59480_6038, \9093 );
and \U$16027 ( \25148 , RIfcbbce8_7159, \9095 );
and \U$16028 ( \25149 , RIe175c38_2717, \9097 );
and \U$16029 ( \25150 , RIfcdb890_7520, \9099 );
and \U$16030 ( \25151 , RIfc59b88_6043, \9101 );
and \U$16031 ( \25152 , RIfc8ada0_6602, \9103 );
and \U$16032 ( \25153 , RIfcb5eb0_7092, \9105 );
and \U$16033 ( \25154 , RIfc57c98_6021, \9107 );
and \U$16034 ( \25155 , RIfc57158_6013, \9109 );
and \U$16035 ( \25156 , RIfc58aa8_6031, \9111 );
and \U$16036 ( \25157 , RIe173910_2692, \9113 );
and \U$16037 ( \25158 , RIfcc62d8_7277, \9115 );
and \U$16038 ( \25159 , RIfc8a968_6599, \9117 );
and \U$16039 ( \25160 , RIfc57428_6015, \9119 );
and \U$16040 ( \25161 , RIfc56d20_6010, \9121 );
and \U$16041 ( \25162 , RIfc408e0_5760, \9123 );
and \U$16042 ( \25163 , RIe223b30_4696, \9125 );
and \U$16043 ( \25164 , RIfc82970_6508, \9127 );
and \U$16044 ( \25165 , RIe220e30_4664, \9129 );
and \U$16045 ( \25166 , RIfcecc30_7716, \9131 );
and \U$16046 ( \25167 , RIe21e130_4632, \9133 );
and \U$16047 ( \25168 , RIe218730_4568, \9135 );
and \U$16048 ( \25169 , RIe215a30_4536, \9137 );
and \U$16049 ( \25170 , RIfc3fad0_5750, \9139 );
and \U$16050 ( \25171 , RIe212d30_4504, \9141 );
and \U$16051 ( \25172 , RIf169148_5655, \9143 );
and \U$16052 ( \25173 , RIe210030_4472, \9145 );
and \U$16053 ( \25174 , RIfc545c0_5982, \9147 );
and \U$16054 ( \25175 , RIe20d330_4440, \9149 );
and \U$16055 ( \25176 , RIe20a630_4408, \9151 );
and \U$16056 ( \25177 , RIe207930_4376, \9153 );
and \U$16057 ( \25178 , RIfc88d48_6579, \9155 );
and \U$16058 ( \25179 , RIfc4bec0_5886, \9157 );
and \U$16059 ( \25180 , RIe202638_4317, \9159 );
and \U$16060 ( \25181 , RIe200b80_4298, \9161 );
and \U$16061 ( \25182 , RIfc88910_6576, \9163 );
and \U$16062 ( \25183 , RIfc4c190_5888, \9165 );
and \U$16063 ( \25184 , RIfc4c2f8_5889, \9167 );
and \U$16064 ( \25185 , RIfcba398_7141, \9169 );
and \U$16065 ( \25186 , RIfcd4270_7436, \9171 );
and \U$16066 ( \25187 , RIfcba0c8_7139, \9173 );
and \U$16067 ( \25188 , RIe1fcda0_4254, \9175 );
and \U$16068 ( \25189 , RIe1fbb58_4241, \9177 );
and \U$16069 ( \25190 , RIfc53d50_5976, \9179 );
and \U$16070 ( \25191 , RIfc9b768_6791, \9181 );
and \U$16071 ( \25192 , RIfc537b0_5972, \9183 );
and \U$16072 ( \25193 , RIfc4c5c8_5891, \9185 );
or \U$16073 ( \25194 , \25130 , \25131 , \25132 , \25133 , \25134 , \25135 , \25136 , \25137 , \25138 , \25139 , \25140 , \25141 , \25142 , \25143 , \25144 , \25145 , \25146 , \25147 , \25148 , \25149 , \25150 , \25151 , \25152 , \25153 , \25154 , \25155 , \25156 , \25157 , \25158 , \25159 , \25160 , \25161 , \25162 , \25163 , \25164 , \25165 , \25166 , \25167 , \25168 , \25169 , \25170 , \25171 , \25172 , \25173 , \25174 , \25175 , \25176 , \25177 , \25178 , \25179 , \25180 , \25181 , \25182 , \25183 , \25184 , \25185 , \25186 , \25187 , \25188 , \25189 , \25190 , \25191 , \25192 , \25193 );
and \U$16074 ( \25195 , RIfc9e468_6823, \9188 );
and \U$16075 ( \25196 , RIf157da8_5459, \9190 );
and \U$16076 ( \25197 , RIfcb9f60_7138, \9192 );
and \U$16077 ( \25198 , RIe1fa208_4223, \9194 );
and \U$16078 ( \25199 , RIfc849c8_6531, \9196 );
and \U$16079 ( \25200 , RIfc529a0_5962, \9198 );
and \U$16080 ( \25201 , RIfc9f6b0_6836, \9200 );
and \U$16081 ( \25202 , RIe1f5618_4169, \9202 );
and \U$16082 ( \25203 , RIf153320_5406, \9204 );
and \U$16083 ( \25204 , RIfcc4988_7259, \9206 );
and \U$16084 ( \25205 , RIf150d28_5379, \9208 );
and \U$16085 ( \25206 , RIfebe458_8285, \9210 );
and \U$16086 ( \25207 , RIfc87f38_6569, \9212 );
and \U$16087 ( \25208 , RIfcb7f08_7115, \9214 );
and \U$16088 ( \25209 , RIf14e190_5348, \9216 );
and \U$16089 ( \25210 , RIfe80658_7805, \9218 );
and \U$16090 ( \25211 , RIe1eb898_4057, \9220 );
and \U$16091 ( \25212 , RIe1e8b98_4025, \9222 );
and \U$16092 ( \25213 , RIe1e5e98_3993, \9224 );
and \U$16093 ( \25214 , RIe1e3198_3961, \9226 );
and \U$16094 ( \25215 , RIe1e0498_3929, \9228 );
and \U$16095 ( \25216 , RIe1dd798_3897, \9230 );
and \U$16096 ( \25217 , RIe1daa98_3865, \9232 );
and \U$16097 ( \25218 , RIe1d7d98_3833, \9234 );
and \U$16098 ( \25219 , RIe1d2398_3769, \9236 );
and \U$16099 ( \25220 , RIe1cf698_3737, \9238 );
and \U$16100 ( \25221 , RIe1cc998_3705, \9240 );
and \U$16101 ( \25222 , RIe1c9c98_3673, \9242 );
and \U$16102 ( \25223 , RIe1c6f98_3641, \9244 );
and \U$16103 ( \25224 , RIe1c4298_3609, \9246 );
and \U$16104 ( \25225 , RIe1c1598_3577, \9248 );
and \U$16105 ( \25226 , RIe1be898_3545, \9250 );
and \U$16106 ( \25227 , RIf14cc78_5333, \9252 );
and \U$16107 ( \25228 , RIf14ba30_5320, \9254 );
and \U$16108 ( \25229 , RIe1b92d0_3484, \9256 );
and \U$16109 ( \25230 , RIe1b7278_3461, \9258 );
and \U$16110 ( \25231 , RIf14a7e8_5307, \9260 );
and \U$16111 ( \25232 , RIf149ca8_5299, \9262 );
and \U$16112 ( \25233 , RIfebe5c0_8286, \9264 );
and \U$16113 ( \25234 , RIfe807c0_7806, \9266 );
and \U$16114 ( \25235 , RIfc50510_5936, \9268 );
and \U$16115 ( \25236 , RIfce4f08_7627, \9270 );
and \U$16116 ( \25237 , RIfe80a90_7808, \9272 );
and \U$16117 ( \25238 , RIfebe890_8288, \9274 );
and \U$16118 ( \25239 , RIfc9cde8_6807, \9276 );
and \U$16119 ( \25240 , RIfc87560_6562, \9278 );
and \U$16120 ( \25241 , RIfe80928_7807, \9280 );
and \U$16121 ( \25242 , RIfebe728_8287, \9282 );
and \U$16122 ( \25243 , RIe1a8bd8_3297, \9284 );
and \U$16123 ( \25244 , RIe1a5ed8_3265, \9286 );
and \U$16124 ( \25245 , RIe1a31d8_3233, \9288 );
and \U$16125 ( \25246 , RIe1a04d8_3201, \9290 );
and \U$16126 ( \25247 , RIe18c9d8_2977, \9292 );
and \U$16127 ( \25248 , RIe178ed8_2753, \9294 );
and \U$16128 ( \25249 , RIe226830_4728, \9296 );
and \U$16129 ( \25250 , RIe21b430_4600, \9298 );
and \U$16130 ( \25251 , RIe204c30_4344, \9300 );
and \U$16131 ( \25252 , RIe1fec90_4276, \9302 );
and \U$16132 ( \25253 , RIe1f8048_4199, \9304 );
and \U$16133 ( \25254 , RIe1f0b90_4116, \9306 );
and \U$16134 ( \25255 , RIe1d5098_3801, \9308 );
and \U$16135 ( \25256 , RIe1bbb98_3513, \9310 );
and \U$16136 ( \25257 , RIe1aea10_3364, \9312 );
and \U$16137 ( \25258 , RIe171048_2663, \9314 );
or \U$16138 ( \25259 , \25195 , \25196 , \25197 , \25198 , \25199 , \25200 , \25201 , \25202 , \25203 , \25204 , \25205 , \25206 , \25207 , \25208 , \25209 , \25210 , \25211 , \25212 , \25213 , \25214 , \25215 , \25216 , \25217 , \25218 , \25219 , \25220 , \25221 , \25222 , \25223 , \25224 , \25225 , \25226 , \25227 , \25228 , \25229 , \25230 , \25231 , \25232 , \25233 , \25234 , \25235 , \25236 , \25237 , \25238 , \25239 , \25240 , \25241 , \25242 , \25243 , \25244 , \25245 , \25246 , \25247 , \25248 , \25249 , \25250 , \25251 , \25252 , \25253 , \25254 , \25255 , \25256 , \25257 , \25258 );
or \U$16139 ( \25260 , \25194 , \25259 );
_DC g5c24 ( \25261_nG5c24 , \25260 , \9323 );
xor g5c25 ( \25262_nG5c25 , \25129_nG5ba0 , \25261_nG5c24 );
buf \U$16140 ( \25263 , \25262_nG5c25 );
xor \U$16141 ( \25264 , \25263 , \24135 );
and \U$16142 ( \25265 , \10687 , \25264 );
xor \U$16143 ( \25266 , \24997 , \25265 );
xor \U$16144 ( \25267 , \24988 , \25266 );
and \U$16145 ( \25268 , \24199 , \10983 );
_DC g65b9 ( \25269_nG65b9 , \25128 , \9597 );
_DC g65ba ( \25270_nG65ba , \25260 , \9323 );
and g65bb ( \25271_nG65bb , \25269_nG65b9 , \25270_nG65ba );
buf \U$16146 ( \25272 , \25271_nG65bb );
and \U$16147 ( \25273 , \25272 , \10691 );
nor \U$16148 ( \25274 , \25268 , \25273 );
xnor \U$16149 ( \25275 , \25274 , \10980 );
and \U$16150 ( \25276 , \11586 , \22542 );
and \U$16151 ( \25277 , \12448 , \22103 );
nor \U$16152 ( \25278 , \25276 , \25277 );
xnor \U$16153 ( \25279 , \25278 , \22548 );
xor \U$16154 ( \25280 , \25275 , \25279 );
and \U$16155 ( \25281 , \10988 , \24138 );
and \U$16156 ( \25282 , \11270 , \23630 );
nor \U$16157 ( \25283 , \25281 , \25282 );
xnor \U$16158 ( \25284 , \25283 , \24144 );
xor \U$16159 ( \25285 , \25280 , \25284 );
xor \U$16160 ( \25286 , \25267 , \25285 );
xor \U$16161 ( \25287 , \24984 , \25286 );
xor \U$16162 ( \25288 , \24945 , \25287 );
and \U$16163 ( \25289 , \23847 , \23851 );
and \U$16164 ( \25290 , \23851 , \24215 );
and \U$16165 ( \25291 , \23847 , \24215 );
or \U$16166 ( \25292 , \25289 , \25290 , \25291 );
xor \U$16167 ( \25293 , \25288 , \25292 );
and \U$16168 ( \25294 , \24216 , \24220 );
and \U$16169 ( \25295 , \24221 , \24224 );
or \U$16170 ( \25296 , \25294 , \25295 );
xor \U$16171 ( \25297 , \25293 , \25296 );
buf g9bcc ( \25298_nG9bcc , \25297 );
and \U$16172 ( \25299 , \10704 , \25298_nG9bcc );
or \U$16173 ( \25300 , \24919 , \25299 );
xor \U$16174 ( \25301 , \10703 , \25300 );
buf \U$16175 ( \25302 , \25301 );
buf \U$16177 ( \25303 , \25302 );
xor \U$16178 ( \25304 , \24918 , \25303 );
buf \U$16179 ( \25305 , \25304 );
xor \U$16180 ( \25306 , \24879 , \25305 );
and \U$16181 ( \25307 , \23786 , \23841 );
and \U$16182 ( \25308 , \23786 , \24231 );
and \U$16183 ( \25309 , \23841 , \24231 );
or \U$16184 ( \25310 , \25307 , \25308 , \25309 );
buf \U$16185 ( \25311 , \25310 );
xor \U$16186 ( \25312 , \25306 , \25311 );
buf \U$16187 ( \25313 , \25312 );
xor \U$16188 ( \25314 , \24874 , \25313 );
and \U$16189 ( \25315 , \24799 , \25314 );
and \U$16190 ( \25316 , \23749 , \23754 );
and \U$16191 ( \25317 , \23749 , \24233 );
and \U$16192 ( \25318 , \23754 , \24233 );
or \U$16193 ( \25319 , \25316 , \25317 , \25318 );
and \U$16194 ( \25320 , \24799 , \25319 );
and \U$16195 ( \25321 , \25314 , \25319 );
or \U$16196 ( \25322 , \25315 , \25320 , \25321 );
and \U$16197 ( \25323 , \24235 , \24239 );
and \U$16198 ( \25324 , \24235 , \24798 );
and \U$16199 ( \25325 , \24239 , \24798 );
or \U$16200 ( \25326 , \25323 , \25324 , \25325 );
xor \U$16201 ( \25327 , \25322 , \25326 );
and \U$16202 ( \25328 , \24881 , \24887 );
and \U$16203 ( \25329 , \24881 , \24894 );
and \U$16204 ( \25330 , \24887 , \24894 );
or \U$16205 ( \25331 , \25328 , \25329 , \25330 );
buf \U$16206 ( \25332 , \25331 );
and \U$16207 ( \25333 , \24788 , \24795 );
buf \U$16208 ( \25334 , \25333 );
buf \U$16210 ( \25335 , \25334 );
and \U$16211 ( \25336 , \23201 , \11283_nG9c08 );
and \U$16212 ( \25337 , \23198 , \11598_nG9c05 );
or \U$16213 ( \25338 , \25336 , \25337 );
xor \U$16214 ( \25339 , \23197 , \25338 );
buf \U$16215 ( \25340 , \25339 );
buf \U$16217 ( \25341 , \25340 );
xor \U$16218 ( \25342 , \25335 , \25341 );
buf \U$16219 ( \25343 , \25342 );
and \U$16220 ( \25344 , \24792 , \10694_nG9c0e );
and \U$16221 ( \25345 , \24789 , \10995_nG9c0b );
or \U$16222 ( \25346 , \25344 , \25345 );
xor \U$16223 ( \25347 , \24788 , \25346 );
buf \U$16224 ( \25348 , \25347 );
buf \U$16226 ( \25349 , \25348 );
xor \U$16227 ( \25350 , \25343 , \25349 );
and \U$16228 ( \25351 , \21658 , \12470_nG9c02 );
and \U$16229 ( \25352 , \21655 , \12801_nG9bff );
or \U$16230 ( \25353 , \25351 , \25352 );
xor \U$16231 ( \25354 , \21654 , \25353 );
buf \U$16232 ( \25355 , \25354 );
buf \U$16234 ( \25356 , \25355 );
xor \U$16235 ( \25357 , \25350 , \25356 );
buf \U$16236 ( \25358 , \25357 );
xor \U$16237 ( \25359 , \25332 , \25358 );
and \U$16238 ( \25360 , \17297 , \16315_nG9bf0 );
and \U$16239 ( \25361 , \17294 , \16680_nG9bed );
or \U$16240 ( \25362 , \25360 , \25361 );
xor \U$16241 ( \25363 , \17293 , \25362 );
buf \U$16242 ( \25364 , \25363 );
buf \U$16244 ( \25365 , \25364 );
xor \U$16245 ( \25366 , \25359 , \25365 );
buf \U$16246 ( \25367 , \25366 );
and \U$16247 ( \25368 , \14631 , \19091_nG9be4 );
and \U$16248 ( \25369 , \14628 , \19586_nG9be1 );
or \U$16249 ( \25370 , \25368 , \25369 );
xor \U$16250 ( \25371 , \14627 , \25370 );
buf \U$16251 ( \25372 , \25371 );
buf \U$16253 ( \25373 , \25372 );
xor \U$16254 ( \25374 , \25367 , \25373 );
and \U$16255 ( \25375 , \13370 , \20608_nG9bde );
and \U$16256 ( \25376 , \13367 , \21086_nG9bdb );
or \U$16257 ( \25377 , \25375 , \25376 );
xor \U$16258 ( \25378 , \13366 , \25377 );
buf \U$16259 ( \25379 , \25378 );
buf \U$16261 ( \25380 , \25379 );
xor \U$16262 ( \25381 , \25374 , \25380 );
buf \U$16263 ( \25382 , \25381 );
and \U$16264 ( \25383 , \24814 , \24828 );
and \U$16265 ( \25384 , \24814 , \24835 );
and \U$16266 ( \25385 , \24828 , \24835 );
or \U$16267 ( \25386 , \25383 , \25384 , \25385 );
buf \U$16268 ( \25387 , \25386 );
and \U$16269 ( \25388 , \24820 , \24826 );
buf \U$16270 ( \25389 , \25388 );
and \U$16271 ( \25390 , \20155 , \13705_nG9bfc );
and \U$16272 ( \25391 , \20152 , \14070_nG9bf9 );
or \U$16273 ( \25392 , \25390 , \25391 );
xor \U$16274 ( \25393 , \20151 , \25392 );
buf \U$16275 ( \25394 , \25393 );
buf \U$16277 ( \25395 , \25394 );
xor \U$16278 ( \25396 , \25389 , \25395 );
and \U$16279 ( \25397 , \18702 , \14984_nG9bf6 );
and \U$16280 ( \25398 , \18699 , \15373_nG9bf3 );
or \U$16281 ( \25399 , \25397 , \25398 );
xor \U$16282 ( \25400 , \18698 , \25399 );
buf \U$16283 ( \25401 , \25400 );
buf \U$16285 ( \25402 , \25401 );
xor \U$16286 ( \25403 , \25396 , \25402 );
buf \U$16287 ( \25404 , \25403 );
xor \U$16288 ( \25405 , \25387 , \25404 );
and \U$16289 ( \25406 , \15940 , \17665_nG9bea );
and \U$16290 ( \25407 , \15937 , \18107_nG9be7 );
or \U$16291 ( \25408 , \25406 , \25407 );
xor \U$16292 ( \25409 , \15936 , \25408 );
buf \U$16293 ( \25410 , \25409 );
buf \U$16295 ( \25411 , \25410 );
xor \U$16296 ( \25412 , \25405 , \25411 );
buf \U$16297 ( \25413 , \25412 );
xor \U$16298 ( \25414 , \25382 , \25413 );
and \U$16299 ( \25415 , \10421 , \23696_nG9bd2 );
and \U$16300 ( \25416 , \10418 , \24226_nG9bcf );
or \U$16301 ( \25417 , \25415 , \25416 );
xor \U$16302 ( \25418 , \10417 , \25417 );
buf \U$16303 ( \25419 , \25418 );
buf \U$16305 ( \25420 , \25419 );
xor \U$16306 ( \25421 , \25414 , \25420 );
buf \U$16307 ( \25422 , \25421 );
and \U$16308 ( \25423 , \24809 , \24851 );
and \U$16309 ( \25424 , \24809 , \24871 );
and \U$16310 ( \25425 , \24851 , \24871 );
or \U$16311 ( \25426 , \25423 , \25424 , \25425 );
buf \U$16312 ( \25427 , \25426 );
xor \U$16313 ( \25428 , \25422 , \25427 );
and \U$16314 ( \25429 , \24837 , \24842 );
and \U$16315 ( \25430 , \24837 , \24849 );
and \U$16316 ( \25431 , \24842 , \24849 );
or \U$16317 ( \25432 , \25429 , \25430 , \25431 );
buf \U$16318 ( \25433 , \25432 );
and \U$16319 ( \25434 , \24896 , \24902 );
and \U$16320 ( \25435 , \24896 , \24909 );
and \U$16321 ( \25436 , \24902 , \24909 );
or \U$16322 ( \25437 , \25434 , \25435 , \25436 );
buf \U$16323 ( \25438 , \25437 );
xor \U$16324 ( \25439 , \25433 , \25438 );
and \U$16325 ( \25440 , \12157 , \22129_nG9bd8 );
and \U$16326 ( \25441 , \12154 , \22629_nG9bd5 );
or \U$16327 ( \25442 , \25440 , \25441 );
xor \U$16328 ( \25443 , \12153 , \25442 );
buf \U$16329 ( \25444 , \25443 );
buf \U$16331 ( \25445 , \25444 );
xor \U$16332 ( \25446 , \25439 , \25445 );
buf \U$16333 ( \25447 , \25446 );
xor \U$16334 ( \25448 , \25428 , \25447 );
buf \U$16335 ( \25449 , \25448 );
and \U$16336 ( \25450 , \24879 , \25305 );
and \U$16337 ( \25451 , \24879 , \25311 );
and \U$16338 ( \25452 , \25305 , \25311 );
or \U$16339 ( \25453 , \25450 , \25451 , \25452 );
buf \U$16340 ( \25454 , \25453 );
xor \U$16341 ( \25455 , \25449 , \25454 );
and \U$16342 ( \25456 , \24911 , \24917 );
and \U$16343 ( \25457 , \24911 , \25303 );
and \U$16344 ( \25458 , \24917 , \25303 );
or \U$16345 ( \25459 , \25456 , \25457 , \25458 );
buf \U$16346 ( \25460 , \25459 );
and \U$16347 ( \25461 , \24857 , \24862 );
and \U$16348 ( \25462 , \24857 , \24869 );
and \U$16349 ( \25463 , \24862 , \24869 );
or \U$16350 ( \25464 , \25461 , \25462 , \25463 );
buf \U$16351 ( \25465 , \25464 );
xor \U$16352 ( \25466 , \25460 , \25465 );
and \U$16353 ( \25467 , \10707 , \25298_nG9bcc );
and \U$16354 ( \25468 , \24927 , \24931 );
and \U$16355 ( \25469 , \24931 , \24943 );
and \U$16356 ( \25470 , \24927 , \24943 );
or \U$16357 ( \25471 , \25468 , \25469 , \25470 );
and \U$16358 ( \25472 , \24949 , \24983 );
and \U$16359 ( \25473 , \24983 , \25286 );
and \U$16360 ( \25474 , \24949 , \25286 );
or \U$16361 ( \25475 , \25472 , \25473 , \25474 );
xor \U$16362 ( \25476 , \25471 , \25475 );
and \U$16363 ( \25477 , \24988 , \25266 );
and \U$16364 ( \25478 , \25266 , \25285 );
and \U$16365 ( \25479 , \24988 , \25285 );
or \U$16366 ( \25480 , \25477 , \25478 , \25479 );
and \U$16367 ( \25481 , \24936 , \24940 );
and \U$16368 ( \25482 , \24940 , \24942 );
and \U$16369 ( \25483 , \24936 , \24942 );
or \U$16370 ( \25484 , \25481 , \25482 , \25483 );
and \U$16371 ( \25485 , \20544 , \14054 );
and \U$16372 ( \25486 , \21033 , \13692 );
nor \U$16373 ( \25487 , \25485 , \25486 );
xnor \U$16374 ( \25488 , \25487 , \14035 );
and \U$16375 ( \25489 , \14950 , \19534 );
and \U$16376 ( \25490 , \15321 , \19045 );
nor \U$16377 ( \25491 , \25489 , \25490 );
xnor \U$16378 ( \25492 , \25491 , \19540 );
xor \U$16379 ( \25493 , \25488 , \25492 );
and \U$16380 ( \25494 , \13679 , \21005 );
and \U$16381 ( \25495 , \14024 , \20557 );
nor \U$16382 ( \25496 , \25494 , \25495 );
xnor \U$16383 ( \25497 , \25496 , \21011 );
xor \U$16384 ( \25498 , \25493 , \25497 );
xor \U$16385 ( \25499 , \25484 , \25498 );
and \U$16386 ( \25500 , \23617 , \11574 );
and \U$16387 ( \25501 , \24199 , \11278 );
nor \U$16388 ( \25502 , \25500 , \25501 );
xnor \U$16389 ( \25503 , \25502 , \11580 );
not \U$16390 ( \25504 , \25265 );
and \U$16391 ( \25505 , RIdec56a8_710, \9333 );
and \U$16392 ( \25506 , RIdec29a8_678, \9335 );
and \U$16393 ( \25507 , RIfc54020_5978, \9337 );
and \U$16394 ( \25508 , RIdebfca8_646, \9339 );
and \U$16395 ( \25509 , RIee1f540_4815, \9341 );
and \U$16396 ( \25510 , RIdebcfa8_614, \9343 );
and \U$16397 ( \25511 , RIdeba2a8_582, \9345 );
and \U$16398 ( \25512 , RIdeb75a8_550, \9347 );
and \U$16399 ( \25513 , RIfc4fe08_5931, \9349 );
and \U$16400 ( \25514 , RIdeb1ba8_486, \9351 );
and \U$16401 ( \25515 , RIfc6b630_6244, \9353 );
and \U$16402 ( \25516 , RIdeaeea8_454, \9355 );
and \U$16403 ( \25517 , RIfc6a118_6229, \9357 );
and \U$16404 ( \25518 , RIdeaaab0_422, \9359 );
and \U$16405 ( \25519 , RIdea41b0_390, \9361 );
and \U$16406 ( \25520 , RIde9d8b0_358, \9363 );
and \U$16407 ( \25521 , RIfc69ce0_6226, \9365 );
and \U$16408 ( \25522 , RIee1be68_4776, \9367 );
and \U$16409 ( \25523 , RIfc653c0_6174, \9369 );
and \U$16410 ( \25524 , RIee1ac20_4763, \9371 );
and \U$16411 ( \25525 , RIde91718_299, \9373 );
and \U$16412 ( \25526 , RIde8df50_282, \9375 );
and \U$16413 ( \25527 , RIde89db0_262, \9377 );
and \U$16414 ( \25528 , RIde85c10_242, \9379 );
and \U$16415 ( \25529 , RIde81db8_223, \9381 );
and \U$16416 ( \25530 , RIfca76a8_6927, \9383 );
and \U$16417 ( \25531 , RIfcca4f0_7324, \9385 );
and \U$16418 ( \25532 , RIfc4ce38_5897, \9387 );
and \U$16419 ( \25533 , RIfc6b360_6242, \9389 );
and \U$16420 ( \25534 , RIe16b918_2601, \9391 );
and \U$16421 ( \25535 , RIe169cf8_2581, \9393 );
and \U$16422 ( \25536 , RIe167f70_2560, \9395 );
and \U$16423 ( \25537 , RIe1656a8_2531, \9397 );
and \U$16424 ( \25538 , RIe1629a8_2499, \9399 );
and \U$16425 ( \25539 , RIee37690_5089, \9401 );
and \U$16426 ( \25540 , RIe15fca8_2467, \9403 );
and \U$16427 ( \25541 , RIfce93f0_7676, \9405 );
and \U$16428 ( \25542 , RIe15cfa8_2435, \9407 );
and \U$16429 ( \25543 , RIe1575a8_2371, \9409 );
and \U$16430 ( \25544 , RIe1548a8_2339, \9411 );
and \U$16431 ( \25545 , RIee35908_5068, \9413 );
and \U$16432 ( \25546 , RIe151ba8_2307, \9415 );
and \U$16433 ( \25547 , RIee34f30_5061, \9417 );
and \U$16434 ( \25548 , RIe14eea8_2275, \9419 );
and \U$16435 ( \25549 , RIfce32e8_7607, \9421 );
and \U$16436 ( \25550 , RIe14c1a8_2243, \9423 );
and \U$16437 ( \25551 , RIe1494a8_2211, \9425 );
and \U$16438 ( \25552 , RIe1467a8_2179, \9427 );
and \U$16439 ( \25553 , RIfcde2c0_7550, \9429 );
and \U$16440 ( \25554 , RIfc687c8_6211, \9431 );
and \U$16441 ( \25555 , RIfca9160_6946, \9433 );
and \U$16442 ( \25556 , RIfcb1590_7040, \9435 );
and \U$16443 ( \25557 , RIe141078_2117, \9437 );
and \U$16444 ( \25558 , RIdf3ef80_2093, \9439 );
and \U$16445 ( \25559 , RIdf3cdc0_2069, \9441 );
and \U$16446 ( \25560 , RIfebeb60_8290, \9443 );
and \U$16447 ( \25561 , RIfc64448_6163, \9445 );
and \U$16448 ( \25562 , RIee2fad0_5001, \9447 );
and \U$16449 ( \25563 , RIfca7978_6929, \9449 );
and \U$16450 ( \25564 , RIfc676e8_6199, \9451 );
and \U$16451 ( \25565 , RIdf35a70_1987, \9453 );
and \U$16452 ( \25566 , RIdf335e0_1961, \9455 );
and \U$16453 ( \25567 , RIdf31420_1937, \9457 );
and \U$16454 ( \25568 , RIdf2f3c8_1914, \9459 );
or \U$16455 ( \25569 , \25505 , \25506 , \25507 , \25508 , \25509 , \25510 , \25511 , \25512 , \25513 , \25514 , \25515 , \25516 , \25517 , \25518 , \25519 , \25520 , \25521 , \25522 , \25523 , \25524 , \25525 , \25526 , \25527 , \25528 , \25529 , \25530 , \25531 , \25532 , \25533 , \25534 , \25535 , \25536 , \25537 , \25538 , \25539 , \25540 , \25541 , \25542 , \25543 , \25544 , \25545 , \25546 , \25547 , \25548 , \25549 , \25550 , \25551 , \25552 , \25553 , \25554 , \25555 , \25556 , \25557 , \25558 , \25559 , \25560 , \25561 , \25562 , \25563 , \25564 , \25565 , \25566 , \25567 , \25568 );
and \U$16456 ( \25570 , RIfccef78_7377, \9462 );
and \U$16457 ( \25571 , RIfca6fa0_6922, \9464 );
and \U$16458 ( \25572 , RIfc62558_6141, \9466 );
and \U$16459 ( \25573 , RIfc61fb8_6137, \9468 );
and \U$16460 ( \25574 , RIfe81b70_7820, \9470 );
and \U$16461 ( \25575 , RIdf281e0_1833, \9472 );
and \U$16462 ( \25576 , RIfe81cd8_7821, \9474 );
and \U$16463 ( \25577 , RIdf249a0_1793, \9476 );
and \U$16464 ( \25578 , RIfc44300_5798, \9478 );
and \U$16465 ( \25579 , RIfcafc40_7022, \9480 );
and \U$16466 ( \25580 , RIdf22ee8_1774, \9482 );
and \U$16467 ( \25581 , RIfcaac18_6965, \9484 );
and \U$16468 ( \25582 , RIdf219d0_1759, \9486 );
and \U$16469 ( \25583 , RIdf1fae0_1737, \9488 );
and \U$16470 ( \25584 , RIdf1b1c0_1685, \9490 );
and \U$16471 ( \25585 , RIdf19438_1664, \9492 );
and \U$16472 ( \25586 , RIdf17278_1640, \9494 );
and \U$16473 ( \25587 , RIdf14578_1608, \9496 );
and \U$16474 ( \25588 , RIdf11878_1576, \9498 );
and \U$16475 ( \25589 , RIdf0eb78_1544, \9500 );
and \U$16476 ( \25590 , RIdf0be78_1512, \9502 );
and \U$16477 ( \25591 , RIdf09178_1480, \9504 );
and \U$16478 ( \25592 , RIdf06478_1448, \9506 );
and \U$16479 ( \25593 , RIdf03778_1416, \9508 );
and \U$16480 ( \25594 , RIdefdd78_1352, \9510 );
and \U$16481 ( \25595 , RIdefb078_1320, \9512 );
and \U$16482 ( \25596 , RIdef8378_1288, \9514 );
and \U$16483 ( \25597 , RIdef5678_1256, \9516 );
and \U$16484 ( \25598 , RIdef2978_1224, \9518 );
and \U$16485 ( \25599 , RIdeefc78_1192, \9520 );
and \U$16486 ( \25600 , RIdeecf78_1160, \9522 );
and \U$16487 ( \25601 , RIdeea278_1128, \9524 );
and \U$16488 ( \25602 , RIfc611a8_6127, \9526 );
and \U$16489 ( \25603 , RIfc61a18_6133, \9528 );
and \U$16490 ( \25604 , RIfca65c8_6915, \9530 );
and \U$16491 ( \25605 , RIfca6b68_6919, \9532 );
and \U$16492 ( \25606 , RIdee4b48_1066, \9534 );
and \U$16493 ( \25607 , RIdee2dc0_1045, \9536 );
and \U$16494 ( \25608 , RIdee0c00_1021, \9538 );
and \U$16495 ( \25609 , RIdedeba8_998, \9540 );
and \U$16496 ( \25610 , RIfc626c0_6142, \9542 );
and \U$16497 ( \25611 , RIfc738f8_6337, \9544 );
and \U$16498 ( \25612 , RIfcb31b0_7060, \9546 );
and \U$16499 ( \25613 , RIee21430_4837, \9548 );
and \U$16500 ( \25614 , RIded9a18_940, \9550 );
and \U$16501 ( \25615 , RIded7588_914, \9552 );
and \U$16502 ( \25616 , RIded5698_892, \9554 );
and \U$16503 ( \25617 , RIded30a0_865, \9556 );
and \U$16504 ( \25618 , RIded0aa8_838, \9558 );
and \U$16505 ( \25619 , RIdecdda8_806, \9560 );
and \U$16506 ( \25620 , RIdecb0a8_774, \9562 );
and \U$16507 ( \25621 , RIdec83a8_742, \9564 );
and \U$16508 ( \25622 , RIdeb48a8_518, \9566 );
and \U$16509 ( \25623 , RIde96fb0_326, \9568 );
and \U$16510 ( \25624 , RIe16e4b0_2632, \9570 );
and \U$16511 ( \25625 , RIe15a2a8_2403, \9572 );
and \U$16512 ( \25626 , RIe143aa8_2147, \9574 );
and \U$16513 ( \25627 , RIdf384a0_2017, \9576 );
and \U$16514 ( \25628 , RIdf2cb00_1885, \9578 );
and \U$16515 ( \25629 , RIdf1d380_1709, \9580 );
and \U$16516 ( \25630 , RIdf00a78_1384, \9582 );
and \U$16517 ( \25631 , RIdee7578_1096, \9584 );
and \U$16518 ( \25632 , RIdedc2e0_969, \9586 );
and \U$16519 ( \25633 , RIde7cef8_199, \9588 );
or \U$16520 ( \25634 , \25570 , \25571 , \25572 , \25573 , \25574 , \25575 , \25576 , \25577 , \25578 , \25579 , \25580 , \25581 , \25582 , \25583 , \25584 , \25585 , \25586 , \25587 , \25588 , \25589 , \25590 , \25591 , \25592 , \25593 , \25594 , \25595 , \25596 , \25597 , \25598 , \25599 , \25600 , \25601 , \25602 , \25603 , \25604 , \25605 , \25606 , \25607 , \25608 , \25609 , \25610 , \25611 , \25612 , \25613 , \25614 , \25615 , \25616 , \25617 , \25618 , \25619 , \25620 , \25621 , \25622 , \25623 , \25624 , \25625 , \25626 , \25627 , \25628 , \25629 , \25630 , \25631 , \25632 , \25633 );
or \U$16521 ( \25635 , \25569 , \25634 );
_DC g5ca9 ( \25636_nG5ca9 , \25635 , \9597 );
and \U$16522 ( \25637 , RIe19d940_3170, \9059 );
and \U$16523 ( \25638 , RIe19ac40_3138, \9061 );
and \U$16524 ( \25639 , RIfc64880_6166, \9063 );
and \U$16525 ( \25640 , RIe197f40_3106, \9065 );
and \U$16526 ( \25641 , RIf144848_5239, \9067 );
and \U$16527 ( \25642 , RIe195240_3074, \9069 );
and \U$16528 ( \25643 , RIe192540_3042, \9071 );
and \U$16529 ( \25644 , RIe18f840_3010, \9073 );
and \U$16530 ( \25645 , RIe189e40_2946, \9075 );
and \U$16531 ( \25646 , RIe187140_2914, \9077 );
and \U$16532 ( \25647 , RIf143a38_5229, \9079 );
and \U$16533 ( \25648 , RIe184440_2882, \9081 );
and \U$16534 ( \25649 , RIfc6f140_6286, \9083 );
and \U$16535 ( \25650 , RIe181740_2850, \9085 );
and \U$16536 ( \25651 , RIe17ea40_2818, \9087 );
and \U$16537 ( \25652 , RIe17bd40_2786, \9089 );
and \U$16538 ( \25653 , RIfc64f88_6171, \9091 );
and \U$16539 ( \25654 , RIf141008_5199, \9093 );
and \U$16540 ( \25655 , RIe177150_2732, \9095 );
and \U$16541 ( \25656 , RIfe81738_7817, \9097 );
and \U$16542 ( \25657 , RIfccabf8_7329, \9099 );
and \U$16543 ( \25658 , RIf13f3e8_5179, \9101 );
and \U$16544 ( \25659 , RIfca81e8_6935, \9103 );
and \U$16545 ( \25660 , RIee3d630_5157, \9105 );
and \U$16546 ( \25661 , RIfc66068_6183, \9107 );
and \U$16547 ( \25662 , RIfc6ed08_6283, \9109 );
and \U$16548 ( \25663 , RIfcdde88_7547, \9111 );
and \U$16549 ( \25664 , RIe173a78_2693, \9113 );
and \U$16550 ( \25665 , RIfc66338_6185, \9115 );
and \U$16551 ( \25666 , RIfc6eba0_6282, \9117 );
and \U$16552 ( \25667 , RIfc664a0_6186, \9119 );
and \U$16553 ( \25668 , RIfcacdd8_6989, \9121 );
and \U$16554 ( \25669 , RIfe81468_7815, \9123 );
and \U$16555 ( \25670 , RIe223c98_4697, \9125 );
and \U$16556 ( \25671 , RIfc66d10_6192, \9127 );
and \U$16557 ( \25672 , RIe220f98_4665, \9129 );
and \U$16558 ( \25673 , RIf16b038_5677, \9131 );
and \U$16559 ( \25674 , RIe21e298_4633, \9133 );
and \U$16560 ( \25675 , RIe218898_4569, \9135 );
and \U$16561 ( \25676 , RIe215b98_4537, \9137 );
and \U$16562 ( \25677 , RIfc3fc38_5751, \9139 );
and \U$16563 ( \25678 , RIe212e98_4505, \9141 );
and \U$16564 ( \25679 , RIfc67850_6200, \9143 );
and \U$16565 ( \25680 , RIe210198_4473, \9145 );
and \U$16566 ( \25681 , RIf167f00_5642, \9147 );
and \U$16567 ( \25682 , RIe20d498_4441, \9149 );
and \U$16568 ( \25683 , RIe20a798_4409, \9151 );
and \U$16569 ( \25684 , RIe207a98_4377, \9153 );
and \U$16570 ( \25685 , RIfcacb08_6987, \9155 );
and \U$16571 ( \25686 , RIfcac9a0_6986, \9157 );
and \U$16572 ( \25687 , RIfea8900_8234, \9159 );
and \U$16573 ( \25688 , RIfe818a0_7818, \9161 );
and \U$16574 ( \25689 , RIfca8a58_6941, \9163 );
and \U$16575 ( \25690 , RIfccad60_7330, \9165 );
and \U$16576 ( \25691 , RIfcac838_6985, \9167 );
and \U$16577 ( \25692 , RIfc67418_6197, \9169 );
and \U$16578 ( \25693 , RIf160340_5554, \9171 );
and \U$16579 ( \25694 , RIf15e450_5532, \9173 );
and \U$16580 ( \25695 , RIfe81a08_7819, \9175 );
and \U$16581 ( \25696 , RIfe81300_7814, \9177 );
and \U$16582 ( \25697 , RIfc6dac0_6270, \9179 );
and \U$16583 ( \25698 , RIf15ba20_5502, \9181 );
and \U$16584 ( \25699 , RIfc6d958_6269, \9183 );
and \U$16585 ( \25700 , RIfc6d7f0_6268, \9185 );
or \U$16586 ( \25701 , \25637 , \25638 , \25639 , \25640 , \25641 , \25642 , \25643 , \25644 , \25645 , \25646 , \25647 , \25648 , \25649 , \25650 , \25651 , \25652 , \25653 , \25654 , \25655 , \25656 , \25657 , \25658 , \25659 , \25660 , \25661 , \25662 , \25663 , \25664 , \25665 , \25666 , \25667 , \25668 , \25669 , \25670 , \25671 , \25672 , \25673 , \25674 , \25675 , \25676 , \25677 , \25678 , \25679 , \25680 , \25681 , \25682 , \25683 , \25684 , \25685 , \25686 , \25687 , \25688 , \25689 , \25690 , \25691 , \25692 , \25693 , \25694 , \25695 , \25696 , \25697 , \25698 , \25699 , \25700 );
and \U$16587 ( \25702 , RIfc587d8_6029, \9188 );
and \U$16588 ( \25703 , RIfc6cf80_6262, \9190 );
and \U$16589 ( \25704 , RIfc6d3b8_6265, \9192 );
and \U$16590 ( \25705 , RIfe815d0_7816, \9194 );
and \U$16591 ( \25706 , RIfc6d520_6266, \9196 );
and \U$16592 ( \25707 , RIfcabe60_6978, \9198 );
and \U$16593 ( \25708 , RIfc6d0e8_6263, \9200 );
and \U$16594 ( \25709 , RIe1f5780_4170, \9202 );
and \U$16595 ( \25710 , RIfc6c5a8_6255, \9204 );
and \U$16596 ( \25711 , RIfc68d68_6215, \9206 );
and \U$16597 ( \25712 , RIfc68c00_6214, \9208 );
and \U$16598 ( \25713 , RIe1f3458_4145, \9210 );
and \U$16599 ( \25714 , RIfc68a98_6213, \9212 );
and \U$16600 ( \25715 , RIfccb8a0_7338, \9214 );
and \U$16601 ( \25716 , RIfca9b38_6953, \9216 );
and \U$16602 ( \25717 , RIe1ee160_4086, \9218 );
and \U$16603 ( \25718 , RIe1eba00_4058, \9220 );
and \U$16604 ( \25719 , RIe1e8d00_4026, \9222 );
and \U$16605 ( \25720 , RIe1e6000_3994, \9224 );
and \U$16606 ( \25721 , RIe1e3300_3962, \9226 );
and \U$16607 ( \25722 , RIe1e0600_3930, \9228 );
and \U$16608 ( \25723 , RIe1dd900_3898, \9230 );
and \U$16609 ( \25724 , RIe1dac00_3866, \9232 );
and \U$16610 ( \25725 , RIe1d7f00_3834, \9234 );
and \U$16611 ( \25726 , RIe1d2500_3770, \9236 );
and \U$16612 ( \25727 , RIe1cf800_3738, \9238 );
and \U$16613 ( \25728 , RIe1ccb00_3706, \9240 );
and \U$16614 ( \25729 , RIe1c9e00_3674, \9242 );
and \U$16615 ( \25730 , RIe1c7100_3642, \9244 );
and \U$16616 ( \25731 , RIe1c4400_3610, \9246 );
and \U$16617 ( \25732 , RIe1c1700_3578, \9248 );
and \U$16618 ( \25733 , RIe1bea00_3546, \9250 );
and \U$16619 ( \25734 , RIfc6bbd0_6248, \9252 );
and \U$16620 ( \25735 , RIfcdd348_7539, \9254 );
and \U$16621 ( \25736 , RIe1b9438_3485, \9256 );
and \U$16622 ( \25737 , RIe1b73e0_3462, \9258 );
and \U$16623 ( \25738 , RIfcab5f0_6972, \9260 );
and \U$16624 ( \25739 , RIfccbb70_7340, \9262 );
and \U$16625 ( \25740 , RIe1b5220_3438, \9264 );
and \U$16626 ( \25741 , RIe1b3e70_3424, \9266 );
and \U$16627 ( \25742 , RIfc6c9e0_6258, \9268 );
and \U$16628 ( \25743 , RIfcab488_6971, \9270 );
and \U$16629 ( \25744 , RIfea7dc0_8226, \9272 );
and \U$16630 ( \25745 , RIe1b0bd0_3388, \9274 );
and \U$16631 ( \25746 , RIfc6ce18_6261, \9276 );
and \U$16632 ( \25747 , RIfcabfc8_6979, \9278 );
and \U$16633 ( \25748 , RIe1ac580_3338, \9280 );
and \U$16634 ( \25749 , RIe1aaf00_3322, \9282 );
and \U$16635 ( \25750 , RIe1a8d40_3298, \9284 );
and \U$16636 ( \25751 , RIe1a6040_3266, \9286 );
and \U$16637 ( \25752 , RIe1a3340_3234, \9288 );
and \U$16638 ( \25753 , RIe1a0640_3202, \9290 );
and \U$16639 ( \25754 , RIe18cb40_2978, \9292 );
and \U$16640 ( \25755 , RIe179040_2754, \9294 );
and \U$16641 ( \25756 , RIe226998_4729, \9296 );
and \U$16642 ( \25757 , RIe21b598_4601, \9298 );
and \U$16643 ( \25758 , RIe204d98_4345, \9300 );
and \U$16644 ( \25759 , RIe1fedf8_4277, \9302 );
and \U$16645 ( \25760 , RIe1f81b0_4200, \9304 );
and \U$16646 ( \25761 , RIe1f0cf8_4117, \9306 );
and \U$16647 ( \25762 , RIe1d5200_3802, \9308 );
and \U$16648 ( \25763 , RIe1bbd00_3514, \9310 );
and \U$16649 ( \25764 , RIe1aeb78_3365, \9312 );
and \U$16650 ( \25765 , RIe1711b0_2664, \9314 );
or \U$16651 ( \25766 , \25702 , \25703 , \25704 , \25705 , \25706 , \25707 , \25708 , \25709 , \25710 , \25711 , \25712 , \25713 , \25714 , \25715 , \25716 , \25717 , \25718 , \25719 , \25720 , \25721 , \25722 , \25723 , \25724 , \25725 , \25726 , \25727 , \25728 , \25729 , \25730 , \25731 , \25732 , \25733 , \25734 , \25735 , \25736 , \25737 , \25738 , \25739 , \25740 , \25741 , \25742 , \25743 , \25744 , \25745 , \25746 , \25747 , \25748 , \25749 , \25750 , \25751 , \25752 , \25753 , \25754 , \25755 , \25756 , \25757 , \25758 , \25759 , \25760 , \25761 , \25762 , \25763 , \25764 , \25765 );
or \U$16652 ( \25767 , \25701 , \25766 );
_DC g5d2d ( \25768_nG5d2d , \25767 , \9323 );
xor g5d2e ( \25769_nG5d2e , \25636_nG5ca9 , \25768_nG5d2d );
buf \U$16653 ( \25770 , \25769_nG5d2e );
and \U$16654 ( \25771 , \25263 , \24135 );
not \U$16655 ( \25772 , \25771 );
and \U$16656 ( \25773 , \25770 , \25772 );
and \U$16657 ( \25774 , \25504 , \25773 );
xor \U$16658 ( \25775 , \25503 , \25774 );
and \U$16659 ( \25776 , \17627 , \16635 );
and \U$16660 ( \25777 , \18035 , \16301 );
nor \U$16661 ( \25778 , \25776 , \25777 );
xnor \U$16662 ( \25779 , \25778 , \16625 );
xor \U$16663 ( \25780 , \25775 , \25779 );
and \U$16664 ( \25781 , \16267 , \18090 );
and \U$16665 ( \25782 , \16655 , \17655 );
nor \U$16666 ( \25783 , \25781 , \25782 );
xnor \U$16667 ( \25784 , \25783 , \18046 );
xor \U$16668 ( \25785 , \25780 , \25784 );
xor \U$16669 ( \25786 , \25499 , \25785 );
xor \U$16670 ( \25787 , \25480 , \25786 );
and \U$16671 ( \25788 , \24953 , \24967 );
and \U$16672 ( \25789 , \24967 , \24982 );
and \U$16673 ( \25790 , \24953 , \24982 );
or \U$16674 ( \25791 , \25788 , \25789 , \25790 );
and \U$16675 ( \25792 , \24992 , \24996 );
and \U$16676 ( \25793 , \24996 , \25265 );
and \U$16677 ( \25794 , \24992 , \25265 );
or \U$16678 ( \25795 , \25792 , \25793 , \25794 );
and \U$16679 ( \25796 , \25275 , \25279 );
and \U$16680 ( \25797 , \25279 , \25284 );
and \U$16681 ( \25798 , \25275 , \25284 );
or \U$16682 ( \25799 , \25796 , \25797 , \25798 );
xor \U$16683 ( \25800 , \25795 , \25799 );
and \U$16684 ( \25801 , \24972 , \24976 );
and \U$16685 ( \25802 , \24976 , \24981 );
and \U$16686 ( \25803 , \24972 , \24981 );
or \U$16687 ( \25804 , \25801 , \25802 , \25803 );
xor \U$16688 ( \25805 , \25800 , \25804 );
xor \U$16689 ( \25806 , \25791 , \25805 );
and \U$16690 ( \25807 , \24957 , \24961 );
and \U$16691 ( \25808 , \24961 , \24966 );
and \U$16692 ( \25809 , \24957 , \24966 );
or \U$16693 ( \25810 , \25807 , \25808 , \25809 );
and \U$16694 ( \25811 , \25272 , \10983 );
_DC g65bc ( \25812_nG65bc , \25635 , \9597 );
_DC g65bd ( \25813_nG65bd , \25767 , \9323 );
and g65be ( \25814_nG65be , \25812_nG65bc , \25813_nG65bd );
buf \U$16695 ( \25815 , \25814_nG65be );
and \U$16696 ( \25816 , \25815 , \10691 );
nor \U$16697 ( \25817 , \25811 , \25816 );
xnor \U$16698 ( \25818 , \25817 , \10980 );
and \U$16699 ( \25819 , \22090 , \12790 );
and \U$16700 ( \25820 , \22556 , \12461 );
nor \U$16701 ( \25821 , \25819 , \25820 );
xnor \U$16702 ( \25822 , \25821 , \12780 );
xor \U$16703 ( \25823 , \25818 , \25822 );
xor \U$16704 ( \25824 , \25770 , \25263 );
not \U$16705 ( \25825 , \25264 );
and \U$16706 ( \25826 , \25824 , \25825 );
and \U$16707 ( \25827 , \10687 , \25826 );
and \U$16708 ( \25828 , \10988 , \25264 );
nor \U$16709 ( \25829 , \25827 , \25828 );
xnor \U$16710 ( \25830 , \25829 , \25773 );
xor \U$16711 ( \25831 , \25823 , \25830 );
xor \U$16712 ( \25832 , \25810 , \25831 );
and \U$16713 ( \25833 , \19032 , \15336 );
and \U$16714 ( \25834 , \19558 , \14963 );
nor \U$16715 ( \25835 , \25833 , \25834 );
xnor \U$16716 ( \25836 , \25835 , \15342 );
and \U$16717 ( \25837 , \12448 , \22542 );
and \U$16718 ( \25838 , \12769 , \22103 );
nor \U$16719 ( \25839 , \25837 , \25838 );
xnor \U$16720 ( \25840 , \25839 , \22548 );
xor \U$16721 ( \25841 , \25836 , \25840 );
and \U$16722 ( \25842 , \11270 , \24138 );
and \U$16723 ( \25843 , \11586 , \23630 );
nor \U$16724 ( \25844 , \25842 , \25843 );
xnor \U$16725 ( \25845 , \25844 , \24144 );
xor \U$16726 ( \25846 , \25841 , \25845 );
xor \U$16727 ( \25847 , \25832 , \25846 );
xor \U$16728 ( \25848 , \25806 , \25847 );
xor \U$16729 ( \25849 , \25787 , \25848 );
xor \U$16730 ( \25850 , \25476 , \25849 );
and \U$16731 ( \25851 , \24923 , \24944 );
and \U$16732 ( \25852 , \24944 , \25287 );
and \U$16733 ( \25853 , \24923 , \25287 );
or \U$16734 ( \25854 , \25851 , \25852 , \25853 );
xor \U$16735 ( \25855 , \25850 , \25854 );
and \U$16736 ( \25856 , \25288 , \25292 );
and \U$16737 ( \25857 , \25293 , \25296 );
or \U$16738 ( \25858 , \25856 , \25857 );
xor \U$16739 ( \25859 , \25855 , \25858 );
buf g9bc9 ( \25860_nG9bc9 , \25859 );
and \U$16740 ( \25861 , \10704 , \25860_nG9bc9 );
or \U$16741 ( \25862 , \25467 , \25861 );
xor \U$16742 ( \25863 , \10703 , \25862 );
buf \U$16743 ( \25864 , \25863 );
buf \U$16745 ( \25865 , \25864 );
xor \U$16746 ( \25866 , \25466 , \25865 );
buf \U$16747 ( \25867 , \25866 );
xor \U$16748 ( \25868 , \25455 , \25867 );
xor \U$16749 ( \25869 , \25327 , \25868 );
and \U$16750 ( \25870 , \24804 , \24873 );
and \U$16751 ( \25871 , \24804 , \25313 );
and \U$16752 ( \25872 , \24873 , \25313 );
or \U$16753 ( \25873 , \25870 , \25871 , \25872 );
and \U$16754 ( \25874 , \25869 , \25873 );
and \U$16755 ( \25875 , \25322 , \25326 );
and \U$16756 ( \25876 , \25322 , \25868 );
and \U$16757 ( \25877 , \25326 , \25868 );
or \U$16758 ( \25878 , \25875 , \25876 , \25877 );
xor \U$16759 ( \25879 , \25874 , \25878 );
and \U$16760 ( \25880 , RIdec5978_712, \9059 );
and \U$16761 ( \25881 , RIdec2c78_680, \9061 );
and \U$16762 ( \25882 , RIfc8aad0_6600, \9063 );
and \U$16763 ( \25883 , RIdebff78_648, \9065 );
and \U$16764 ( \25884 , RIfc8ac38_6601, \9067 );
and \U$16765 ( \25885 , RIdebd278_616, \9069 );
and \U$16766 ( \25886 , RIdeba578_584, \9071 );
and \U$16767 ( \25887 , RIdeb7878_552, \9073 );
and \U$16768 ( \25888 , RIfc40e80_5764, \9075 );
and \U$16769 ( \25889 , RIdeb1e78_488, \9077 );
and \U$16770 ( \25890 , RIfcdaeb8_7513, \9079 );
and \U$16771 ( \25891 , RIdeaf178_456, \9081 );
and \U$16772 ( \25892 , RIee1dbf0_4797, \9083 );
and \U$16773 ( \25893 , RIdeab140_424, \9085 );
and \U$16774 ( \25894 , RIdea4840_392, \9087 );
and \U$16775 ( \25895 , RIde9df40_360, \9089 );
and \U$16776 ( \25896 , RIfc8b070_6604, \9091 );
and \U$16777 ( \25897 , RIfcc38a8_7247, \9093 );
and \U$16778 ( \25898 , RIfc807b0_6484, \9095 );
and \U$16779 ( \25899 , RIfcbb8b0_7156, \9097 );
and \U$16780 ( \25900 , RIde91a60_300, \9099 );
and \U$16781 ( \25901 , RIde8e298_283, \9101 );
and \U$16782 ( \25902 , RIde8a440_264, \9103 );
and \U$16783 ( \25903 , RIde862a0_244, \9105 );
and \U$16784 ( \25904 , RIde82100_224, \9107 );
and \U$16785 ( \25905 , RIfcbbb80_7158, \9109 );
and \U$16786 ( \25906 , RIfc8c150_6616, \9111 );
and \U$16787 ( \25907 , RIfcbbfb8_7161, \9113 );
and \U$16788 ( \25908 , RIfc54458_5981, \9115 );
and \U$16789 ( \25909 , RIe16bbe8_2603, \9117 );
and \U$16790 ( \25910 , RIfc8c2b8_6617, \9119 );
and \U$16791 ( \25911 , RIe168240_2562, \9121 );
and \U$16792 ( \25912 , RIe165978_2533, \9123 );
and \U$16793 ( \25913 , RIe162c78_2501, \9125 );
and \U$16794 ( \25914 , RIee37960_5091, \9127 );
and \U$16795 ( \25915 , RIe15ff78_2469, \9129 );
and \U$16796 ( \25916 , RIfcd6b38_7465, \9131 );
and \U$16797 ( \25917 , RIe15d278_2437, \9133 );
and \U$16798 ( \25918 , RIe157878_2373, \9135 );
and \U$16799 ( \25919 , RIe154b78_2341, \9137 );
and \U$16800 ( \25920 , RIfc8e5e0_6642, \9139 );
and \U$16801 ( \25921 , RIe151e78_2309, \9141 );
and \U$16802 ( \25922 , RIfcb4290_7072, \9143 );
and \U$16803 ( \25923 , RIe14f178_2277, \9145 );
and \U$16804 ( \25924 , RIfc56ff0_6012, \9147 );
and \U$16805 ( \25925 , RIe14c478_2245, \9149 );
and \U$16806 ( \25926 , RIe149778_2213, \9151 );
and \U$16807 ( \25927 , RIe146a78_2181, \9153 );
and \U$16808 ( \25928 , RIee346c0_5055, \9155 );
and \U$16809 ( \25929 , RIee335e0_5043, \9157 );
and \U$16810 ( \25930 , RIee32398_5030, \9159 );
and \U$16811 ( \25931 , RIee31420_5019, \9161 );
and \U$16812 ( \25932 , RIe141348_2119, \9163 );
and \U$16813 ( \25933 , RIe13f020_2094, \9165 );
and \U$16814 ( \25934 , RIfec16f8_8321, \9167 );
and \U$16815 ( \25935 , RIdf3a930_2043, \9169 );
and \U$16816 ( \25936 , RIfce3e28_7615, \9171 );
and \U$16817 ( \25937 , RIfc56780_6006, \9173 );
and \U$16818 ( \25938 , RIfcb4128_7071, \9175 );
and \U$16819 ( \25939 , RIfce2eb0_7604, \9177 );
and \U$16820 ( \25940 , RIdf35d40_1989, \9179 );
and \U$16821 ( \25941 , RIfe88218_7893, \9181 );
and \U$16822 ( \25942 , RIdf316f0_1939, \9183 );
and \U$16823 ( \25943 , RIdf2f698_1916, \9185 );
or \U$16824 ( \25944 , \25880 , \25881 , \25882 , \25883 , \25884 , \25885 , \25886 , \25887 , \25888 , \25889 , \25890 , \25891 , \25892 , \25893 , \25894 , \25895 , \25896 , \25897 , \25898 , \25899 , \25900 , \25901 , \25902 , \25903 , \25904 , \25905 , \25906 , \25907 , \25908 , \25909 , \25910 , \25911 , \25912 , \25913 , \25914 , \25915 , \25916 , \25917 , \25918 , \25919 , \25920 , \25921 , \25922 , \25923 , \25924 , \25925 , \25926 , \25927 , \25928 , \25929 , \25930 , \25931 , \25932 , \25933 , \25934 , \25935 , \25936 , \25937 , \25938 , \25939 , \25940 , \25941 , \25942 , \25943 );
and \U$16825 ( \25945 , RIfc7f9a0_6474, \9188 );
and \U$16826 ( \25946 , RIfce4260_7618, \9190 );
and \U$16827 ( \25947 , RIfcd62c8_7459, \9192 );
and \U$16828 ( \25948 , RIfce9990_7680, \9194 );
and \U$16829 ( \25949 , RIdf2a670_1859, \9196 );
and \U$16830 ( \25950 , RIdf284b0_1835, \9198 );
and \U$16831 ( \25951 , RIdf26728_1814, \9200 );
and \U$16832 ( \25952 , RIdf24c70_1795, \9202 );
and \U$16833 ( \25953 , RIfc7ecf8_6465, \9204 );
and \U$16834 ( \25954 , RIfcc31a0_7242, \9206 );
and \U$16835 ( \25955 , RIfc99008_6763, \9208 );
and \U$16836 ( \25956 , RIfc46e98_5829, \9210 );
and \U$16837 ( \25957 , RIfce2a78_7601, \9212 );
and \U$16838 ( \25958 , RIdf1fdb0_1739, \9214 );
and \U$16839 ( \25959 , RIfcc6e18_7285, \9216 );
and \U$16840 ( \25960 , RIdf19708_1666, \9218 );
and \U$16841 ( \25961 , RIdf17548_1642, \9220 );
and \U$16842 ( \25962 , RIdf14848_1610, \9222 );
and \U$16843 ( \25963 , RIdf11b48_1578, \9224 );
and \U$16844 ( \25964 , RIdf0ee48_1546, \9226 );
and \U$16845 ( \25965 , RIdf0c148_1514, \9228 );
and \U$16846 ( \25966 , RIdf09448_1482, \9230 );
and \U$16847 ( \25967 , RIdf06748_1450, \9232 );
and \U$16848 ( \25968 , RIdf03a48_1418, \9234 );
and \U$16849 ( \25969 , RIdefe048_1354, \9236 );
and \U$16850 ( \25970 , RIdefb348_1322, \9238 );
and \U$16851 ( \25971 , RIdef8648_1290, \9240 );
and \U$16852 ( \25972 , RIdef5948_1258, \9242 );
and \U$16853 ( \25973 , RIdef2c48_1226, \9244 );
and \U$16854 ( \25974 , RIdeeff48_1194, \9246 );
and \U$16855 ( \25975 , RIdeed248_1162, \9248 );
and \U$16856 ( \25976 , RIdeea548_1130, \9250 );
and \U$16857 ( \25977 , RIfcd9130_7492, \9252 );
and \U$16858 ( \25978 , RIfc7cb38_6441, \9254 );
and \U$16859 ( \25979 , RIfc97af0_6748, \9256 );
and \U$16860 ( \25980 , RIfcb3e58_7069, \9258 );
and \U$16861 ( \25981 , RIdee4e18_1068, \9260 );
and \U$16862 ( \25982 , RIdee3090_1047, \9262 );
and \U$16863 ( \25983 , RIdee0ed0_1023, \9264 );
and \U$16864 ( \25984 , RIfe88380_7894, \9266 );
and \U$16865 ( \25985 , RIfc97dc0_6750, \9268 );
and \U$16866 ( \25986 , RIfcc2930_7236, \9270 );
and \U$16867 ( \25987 , RIfcd9298_7493, \9272 );
and \U$16868 ( \25988 , RIfc7c868_6439, \9274 );
and \U$16869 ( \25989 , RIded9ce8_942, \9276 );
and \U$16870 ( \25990 , RIded76f0_915, \9278 );
and \U$16871 ( \25991 , RIded5968_894, \9280 );
and \U$16872 ( \25992 , RIded3370_867, \9282 );
and \U$16873 ( \25993 , RIded0d78_840, \9284 );
and \U$16874 ( \25994 , RIdece078_808, \9286 );
and \U$16875 ( \25995 , RIdecb378_776, \9288 );
and \U$16876 ( \25996 , RIdec8678_744, \9290 );
and \U$16877 ( \25997 , RIdeb4b78_520, \9292 );
and \U$16878 ( \25998 , RIde97640_328, \9294 );
and \U$16879 ( \25999 , RIe16e780_2634, \9296 );
and \U$16880 ( \26000 , RIe15a578_2405, \9298 );
and \U$16881 ( \26001 , RIe143d78_2149, \9300 );
and \U$16882 ( \26002 , RIdf38770_2019, \9302 );
and \U$16883 ( \26003 , RIdf2cdd0_1887, \9304 );
and \U$16884 ( \26004 , RIdf1d650_1711, \9306 );
and \U$16885 ( \26005 , RIdf00d48_1386, \9308 );
and \U$16886 ( \26006 , RIdee7848_1098, \9310 );
and \U$16887 ( \26007 , RIdedc5b0_971, \9312 );
and \U$16888 ( \26008 , RIde7d588_201, \9314 );
or \U$16889 ( \26009 , \25945 , \25946 , \25947 , \25948 , \25949 , \25950 , \25951 , \25952 , \25953 , \25954 , \25955 , \25956 , \25957 , \25958 , \25959 , \25960 , \25961 , \25962 , \25963 , \25964 , \25965 , \25966 , \25967 , \25968 , \25969 , \25970 , \25971 , \25972 , \25973 , \25974 , \25975 , \25976 , \25977 , \25978 , \25979 , \25980 , \25981 , \25982 , \25983 , \25984 , \25985 , \25986 , \25987 , \25988 , \25989 , \25990 , \25991 , \25992 , \25993 , \25994 , \25995 , \25996 , \25997 , \25998 , \25999 , \26000 , \26001 , \26002 , \26003 , \26004 , \26005 , \26006 , \26007 , \26008 );
or \U$16890 ( \26010 , \25944 , \26009 );
_DC g2553 ( \26011_nG2553 , \26010 , \9323 );
buf \U$16891 ( \26012 , \26011_nG2553 );
and \U$16892 ( \26013 , RIe19dc10_3172, \9333 );
and \U$16893 ( \26014 , RIe19af10_3140, \9335 );
and \U$16894 ( \26015 , RIfec1590_8320, \9337 );
and \U$16895 ( \26016 , RIe198210_3108, \9339 );
and \U$16896 ( \26017 , RIfec1428_8319, \9341 );
and \U$16897 ( \26018 , RIe195510_3076, \9343 );
and \U$16898 ( \26019 , RIe192810_3044, \9345 );
and \U$16899 ( \26020 , RIe18fb10_3012, \9347 );
and \U$16900 ( \26021 , RIe18a110_2948, \9349 );
and \U$16901 ( \26022 , RIe187410_2916, \9351 );
and \U$16902 ( \26023 , RIfec12c0_8318, \9353 );
and \U$16903 ( \26024 , RIe184710_2884, \9355 );
and \U$16904 ( \26025 , RIfc88370_6572, \9357 );
and \U$16905 ( \26026 , RIe181a10_2852, \9359 );
and \U$16906 ( \26027 , RIe17ed10_2820, \9361 );
and \U$16907 ( \26028 , RIe17c010_2788, \9363 );
and \U$16908 ( \26029 , RIfc6ccb0_6260, \9365 );
and \U$16909 ( \26030 , RIfc5f858_6109, \9367 );
and \U$16910 ( \26031 , RIfca88f0_6940, \9369 );
and \U$16911 ( \26032 , RIe175f08_2719, \9371 );
and \U$16912 ( \26033 , RIfc81020_6490, \9373 );
and \U$16913 ( \26034 , RIfcc6008_7275, \9375 );
and \U$16914 ( \26035 , RIfc4ea58_5917, \9377 );
and \U$16915 ( \26036 , RIfc42140_5774, \9379 );
and \U$16916 ( \26037 , RIfca3b98_6885, \9381 );
and \U$16917 ( \26038 , RIfc5ac68_6055, \9383 );
and \U$16918 ( \26039 , RIfc984c8_6755, \9385 );
and \U$16919 ( \26040 , RIe173d48_2695, \9387 );
and \U$16920 ( \26041 , RIfc9b330_6788, \9389 );
and \U$16921 ( \26042 , RIf16f688_5727, \9391 );
and \U$16922 ( \26043 , RIfc42410_5776, \9393 );
and \U$16923 ( \26044 , RIfc5f588_6107, \9395 );
and \U$16924 ( \26045 , RIfe880b0_7892, \9397 );
and \U$16925 ( \26046 , RIe223f68_4699, \9399 );
and \U$16926 ( \26047 , RIf16bfb0_5688, \9401 );
and \U$16927 ( \26048 , RIe221268_4667, \9403 );
and \U$16928 ( \26049 , RIfc86cf0_6556, \9405 );
and \U$16929 ( \26050 , RIe21e568_4635, \9407 );
and \U$16930 ( \26051 , RIe218b68_4571, \9409 );
and \U$16931 ( \26052 , RIe215e68_4539, \9411 );
and \U$16932 ( \26053 , RIfe87de0_7890, \9413 );
and \U$16933 ( \26054 , RIe213168_4507, \9415 );
and \U$16934 ( \26055 , RIf1692b0_5656, \9417 );
and \U$16935 ( \26056 , RIe210468_4475, \9419 );
and \U$16936 ( \26057 , RIfcdf670_7564, \9421 );
and \U$16937 ( \26058 , RIe20d768_4443, \9423 );
and \U$16938 ( \26059 , RIe20aa68_4411, \9425 );
and \U$16939 ( \26060 , RIe207d68_4379, \9427 );
and \U$16940 ( \26061 , RIfca6460_6914, \9429 );
and \U$16941 ( \26062 , RIf1662e0_5622, \9431 );
and \U$16942 ( \26063 , RIe202908_4319, \9433 );
and \U$16943 ( \26064 , RIfe87b10_7888, \9435 );
and \U$16944 ( \26065 , RIfc58c10_6032, \9437 );
and \U$16945 ( \26066 , RIfc50ab0_5940, \9439 );
and \U$16946 ( \26067 , RIfccd790_7360, \9441 );
and \U$16947 ( \26068 , RIfccd1f0_7356, \9443 );
and \U$16948 ( \26069 , RIf160610_5556, \9445 );
and \U$16949 ( \26070 , RIf15e720_5534, \9447 );
and \U$16950 ( \26071 , RIfe87c78_7889, \9449 );
and \U$16951 ( \26072 , RIfe87f48_7891, \9451 );
and \U$16952 ( \26073 , RIfce7668_7655, \9453 );
and \U$16953 ( \26074 , RIfc86480_6550, \9455 );
and \U$16954 ( \26075 , RIfcd2218_7413, \9457 );
and \U$16955 ( \26076 , RIfcb01e0_7026, \9459 );
or \U$16956 ( \26077 , \26013 , \26014 , \26015 , \26016 , \26017 , \26018 , \26019 , \26020 , \26021 , \26022 , \26023 , \26024 , \26025 , \26026 , \26027 , \26028 , \26029 , \26030 , \26031 , \26032 , \26033 , \26034 , \26035 , \26036 , \26037 , \26038 , \26039 , \26040 , \26041 , \26042 , \26043 , \26044 , \26045 , \26046 , \26047 , \26048 , \26049 , \26050 , \26051 , \26052 , \26053 , \26054 , \26055 , \26056 , \26057 , \26058 , \26059 , \26060 , \26061 , \26062 , \26063 , \26064 , \26065 , \26066 , \26067 , \26068 , \26069 , \26070 , \26071 , \26072 , \26073 , \26074 , \26075 , \26076 );
and \U$16957 ( \26078 , RIfc47b40_5838, \9462 );
and \U$16958 ( \26079 , RIfc84158_6525, \9464 );
and \U$16959 ( \26080 , RIfc4b920_5882, \9466 );
and \U$16960 ( \26081 , RIe1fa4d8_4225, \9468 );
and \U$16961 ( \26082 , RIfc4ba88_5883, \9470 );
and \U$16962 ( \26083 , RIfcb7530_7108, \9472 );
and \U$16963 ( \26084 , RIfcd58f0_7452, \9474 );
and \U$16964 ( \26085 , RIe1f5a50_4172, \9476 );
and \U$16965 ( \26086 , RIf153488_5407, \9478 );
and \U$16966 ( \26087 , RIf151ca0_5390, \9480 );
and \U$16967 ( \26088 , RIfc51e60_5954, \9482 );
and \U$16968 ( \26089 , RIe1f3728_4147, \9484 );
and \U$16969 ( \26090 , RIfc9aef8_6785, \9486 );
and \U$16970 ( \26091 , RIfcbaaa0_7146, \9488 );
and \U$16971 ( \26092 , RIfc52130_5956, \9490 );
and \U$16972 ( \26093 , RIe1ee430_4088, \9492 );
and \U$16973 ( \26094 , RIe1ebcd0_4060, \9494 );
and \U$16974 ( \26095 , RIe1e8fd0_4028, \9496 );
and \U$16975 ( \26096 , RIe1e62d0_3996, \9498 );
and \U$16976 ( \26097 , RIe1e35d0_3964, \9500 );
and \U$16977 ( \26098 , RIe1e08d0_3932, \9502 );
and \U$16978 ( \26099 , RIe1ddbd0_3900, \9504 );
and \U$16979 ( \26100 , RIe1daed0_3868, \9506 );
and \U$16980 ( \26101 , RIe1d81d0_3836, \9508 );
and \U$16981 ( \26102 , RIe1d27d0_3772, \9510 );
and \U$16982 ( \26103 , RIe1cfad0_3740, \9512 );
and \U$16983 ( \26104 , RIe1ccdd0_3708, \9514 );
and \U$16984 ( \26105 , RIe1ca0d0_3676, \9516 );
and \U$16985 ( \26106 , RIe1c73d0_3644, \9518 );
and \U$16986 ( \26107 , RIe1c46d0_3612, \9520 );
and \U$16987 ( \26108 , RIe1c19d0_3580, \9522 );
and \U$16988 ( \26109 , RIe1becd0_3548, \9524 );
and \U$16989 ( \26110 , RIfce0b88_7579, \9526 );
and \U$16990 ( \26111 , RIfc82808_6507, \9528 );
and \U$16991 ( \26112 , RIe1b9708_3487, \9530 );
and \U$16992 ( \26113 , RIe1b76b0_3464, \9532 );
and \U$16993 ( \26114 , RIfcd5bc0_7454, \9534 );
and \U$16994 ( \26115 , RIfcb69f0_7100, \9536 );
and \U$16995 ( \26116 , RIe1b54f0_3440, \9538 );
and \U$16996 ( \26117 , RIe1b4140_3426, \9540 );
and \U$16997 ( \26118 , RIfc89f90_6592, \9542 );
and \U$16998 ( \26119 , RIfce9af8_7681, \9544 );
and \U$16999 ( \26120 , RIe1b2958_3409, \9546 );
and \U$17000 ( \26121 , RIe1b0ea0_3390, \9548 );
and \U$17001 ( \26122 , RIfc4a138_5865, \9550 );
and \U$17002 ( \26123 , RIfc8a260_6594, \9552 );
and \U$17003 ( \26124 , RIe1ac850_3340, \9554 );
and \U$17004 ( \26125 , RIe1ab1d0_3324, \9556 );
and \U$17005 ( \26126 , RIe1a9010_3300, \9558 );
and \U$17006 ( \26127 , RIe1a6310_3268, \9560 );
and \U$17007 ( \26128 , RIe1a3610_3236, \9562 );
and \U$17008 ( \26129 , RIe1a0910_3204, \9564 );
and \U$17009 ( \26130 , RIe18ce10_2980, \9566 );
and \U$17010 ( \26131 , RIe179310_2756, \9568 );
and \U$17011 ( \26132 , RIe226c68_4731, \9570 );
and \U$17012 ( \26133 , RIe21b868_4603, \9572 );
and \U$17013 ( \26134 , RIe205068_4347, \9574 );
and \U$17014 ( \26135 , RIe1ff0c8_4279, \9576 );
and \U$17015 ( \26136 , RIe1f8480_4202, \9578 );
and \U$17016 ( \26137 , RIe1f0fc8_4119, \9580 );
and \U$17017 ( \26138 , RIe1d54d0_3804, \9582 );
and \U$17018 ( \26139 , RIe1bbfd0_3516, \9584 );
and \U$17019 ( \26140 , RIe1aee48_3367, \9586 );
and \U$17020 ( \26141 , RIe171480_2666, \9588 );
or \U$17021 ( \26142 , \26078 , \26079 , \26080 , \26081 , \26082 , \26083 , \26084 , \26085 , \26086 , \26087 , \26088 , \26089 , \26090 , \26091 , \26092 , \26093 , \26094 , \26095 , \26096 , \26097 , \26098 , \26099 , \26100 , \26101 , \26102 , \26103 , \26104 , \26105 , \26106 , \26107 , \26108 , \26109 , \26110 , \26111 , \26112 , \26113 , \26114 , \26115 , \26116 , \26117 , \26118 , \26119 , \26120 , \26121 , \26122 , \26123 , \26124 , \26125 , \26126 , \26127 , \26128 , \26129 , \26130 , \26131 , \26132 , \26133 , \26134 , \26135 , \26136 , \26137 , \26138 , \26139 , \26140 , \26141 );
or \U$17022 ( \26143 , \26077 , \26142 );
_DC g3680 ( \26144_nG3680 , \26143 , \9597 );
buf \U$17023 ( \26145 , \26144_nG3680 );
xor \U$17024 ( \26146 , \26012 , \26145 );
and \U$17025 ( \26147 , RIdec5810_711, \9059 );
and \U$17026 ( \26148 , RIdec2b10_679, \9061 );
and \U$17027 ( \26149 , RIfce6f60_7650, \9063 );
and \U$17028 ( \26150 , RIdebfe10_647, \9065 );
and \U$17029 ( \26151 , RIfc95228_6719, \9067 );
and \U$17030 ( \26152 , RIdebd110_615, \9069 );
and \U$17031 ( \26153 , RIdeba410_583, \9071 );
and \U$17032 ( \26154 , RIdeb7710_551, \9073 );
and \U$17033 ( \26155 , RIfe879a8_7887, \9075 );
and \U$17034 ( \26156 , RIdeb1d10_487, \9077 );
and \U$17035 ( \26157 , RIfcc16e8_7223, \9079 );
and \U$17036 ( \26158 , RIdeaf010_455, \9081 );
and \U$17037 ( \26159 , RIfca4f48_6899, \9083 );
and \U$17038 ( \26160 , RIdeaadf8_423, \9085 );
and \U$17039 ( \26161 , RIdea44f8_391, \9087 );
and \U$17040 ( \26162 , RIde9dbf8_359, \9089 );
and \U$17041 ( \26163 , RIee1cf48_4788, \9091 );
and \U$17042 ( \26164 , RIee1bfd0_4777, \9093 );
and \U$17043 ( \26165 , RIfc95660_6722, \9095 );
and \U$17044 ( \26166 , RIfcee148_7731, \9097 );
and \U$17045 ( \26167 , RIfe87840_7886, \9099 );
and \U$17046 ( \26168 , RIfe876d8_7885, \9101 );
and \U$17047 ( \26169 , RIde8a0f8_263, \9103 );
and \U$17048 ( \26170 , RIde85f58_243, \9105 );
and \U$17049 ( \26171 , RIfcb0780_7030, \9107 );
and \U$17050 ( \26172 , RIfcee9b8_7737, \9109 );
and \U$17051 ( \26173 , RIfc5f150_6104, \9111 );
and \U$17052 ( \26174 , RIfcdee00_7558, \9113 );
and \U$17053 ( \26175 , RIfcd8050_7480, \9115 );
and \U$17054 ( \26176 , RIe16ba80_2602, \9117 );
and \U$17055 ( \26177 , RIfca5380_6902, \9119 );
and \U$17056 ( \26178 , RIe1680d8_2561, \9121 );
and \U$17057 ( \26179 , RIe165810_2532, \9123 );
and \U$17058 ( \26180 , RIe162b10_2500, \9125 );
and \U$17059 ( \26181 , RIee377f8_5090, \9127 );
and \U$17060 ( \26182 , RIe15fe10_2468, \9129 );
and \U$17061 ( \26183 , RIee36448_5076, \9131 );
and \U$17062 ( \26184 , RIe15d110_2436, \9133 );
and \U$17063 ( \26185 , RIe157710_2372, \9135 );
and \U$17064 ( \26186 , RIe154a10_2340, \9137 );
and \U$17065 ( \26187 , RIfc3f3c8_5745, \9139 );
and \U$17066 ( \26188 , RIe151d10_2308, \9141 );
and \U$17067 ( \26189 , RIfcde9c8_7555, \9143 );
and \U$17068 ( \26190 , RIe14f010_2276, \9145 );
and \U$17069 ( \26191 , RIfc4a2a0_5866, \9147 );
and \U$17070 ( \26192 , RIe14c310_2244, \9149 );
and \U$17071 ( \26193 , RIe149610_2212, \9151 );
and \U$17072 ( \26194 , RIe146910_2180, \9153 );
and \U$17073 ( \26195 , RIfc62288_6139, \9155 );
and \U$17074 ( \26196 , RIee33478_5042, \9157 );
and \U$17075 ( \26197 , RIfc71b70_6316, \9159 );
and \U$17076 ( \26198 , RIee312b8_5018, \9161 );
and \U$17077 ( \26199 , RIe1411e0_2118, \9163 );
and \U$17078 ( \26200 , RIfe87570_7884, \9165 );
and \U$17079 ( \26201 , RIdf3cf28_2070, \9167 );
and \U$17080 ( \26202 , RIfe87408_7883, \9169 );
and \U$17081 ( \26203 , RIfcc99b0_7316, \9171 );
and \U$17082 ( \26204 , RIfccf0e0_7378, \9173 );
and \U$17083 ( \26205 , RIfcaeb60_7010, \9175 );
and \U$17084 ( \26206 , RIfcca220_7322, \9177 );
and \U$17085 ( \26207 , RIdf35bd8_1988, \9179 );
and \U$17086 ( \26208 , RIdf33748_1962, \9181 );
and \U$17087 ( \26209 , RIdf31588_1938, \9183 );
and \U$17088 ( \26210 , RIdf2f530_1915, \9185 );
or \U$17089 ( \26211 , \26147 , \26148 , \26149 , \26150 , \26151 , \26152 , \26153 , \26154 , \26155 , \26156 , \26157 , \26158 , \26159 , \26160 , \26161 , \26162 , \26163 , \26164 , \26165 , \26166 , \26167 , \26168 , \26169 , \26170 , \26171 , \26172 , \26173 , \26174 , \26175 , \26176 , \26177 , \26178 , \26179 , \26180 , \26181 , \26182 , \26183 , \26184 , \26185 , \26186 , \26187 , \26188 , \26189 , \26190 , \26191 , \26192 , \26193 , \26194 , \26195 , \26196 , \26197 , \26198 , \26199 , \26200 , \26201 , \26202 , \26203 , \26204 , \26205 , \26206 , \26207 , \26208 , \26209 , \26210 );
and \U$17090 ( \26212 , RIee2be58_4958, \9188 );
and \U$17091 ( \26213 , RIee2a508_4940, \9190 );
and \U$17092 ( \26214 , RIee28ff0_4925, \9192 );
and \U$17093 ( \26215 , RIee27da8_4912, \9194 );
and \U$17094 ( \26216 , RIdf2a508_1858, \9196 );
and \U$17095 ( \26217 , RIdf28348_1834, \9198 );
and \U$17096 ( \26218 , RIdf265c0_1813, \9200 );
and \U$17097 ( \26219 , RIdf24b08_1794, \9202 );
and \U$17098 ( \26220 , RIfc74708_6347, \9204 );
and \U$17099 ( \26221 , RIfc42578_5777, \9206 );
and \U$17100 ( \26222 , RIfc43388_5787, \9208 );
and \U$17101 ( \26223 , RIfc745a0_6346, \9210 );
and \U$17102 ( \26224 , RIfcb0078_7025, \9212 );
and \U$17103 ( \26225 , RIdf1fc48_1738, \9214 );
and \U$17104 ( \26226 , RIfcaff10_7024, \9216 );
and \U$17105 ( \26227 , RIdf195a0_1665, \9218 );
and \U$17106 ( \26228 , RIdf173e0_1641, \9220 );
and \U$17107 ( \26229 , RIdf146e0_1609, \9222 );
and \U$17108 ( \26230 , RIdf119e0_1577, \9224 );
and \U$17109 ( \26231 , RIdf0ece0_1545, \9226 );
and \U$17110 ( \26232 , RIdf0bfe0_1513, \9228 );
and \U$17111 ( \26233 , RIdf092e0_1481, \9230 );
and \U$17112 ( \26234 , RIdf065e0_1449, \9232 );
and \U$17113 ( \26235 , RIdf038e0_1417, \9234 );
and \U$17114 ( \26236 , RIdefdee0_1353, \9236 );
and \U$17115 ( \26237 , RIdefb1e0_1321, \9238 );
and \U$17116 ( \26238 , RIdef84e0_1289, \9240 );
and \U$17117 ( \26239 , RIdef57e0_1257, \9242 );
and \U$17118 ( \26240 , RIdef2ae0_1225, \9244 );
and \U$17119 ( \26241 , RIdeefde0_1193, \9246 );
and \U$17120 ( \26242 , RIdeed0e0_1161, \9248 );
and \U$17121 ( \26243 , RIdeea3e0_1129, \9250 );
and \U$17122 ( \26244 , RIee257b0_4885, \9252 );
and \U$17123 ( \26245 , RIfca73d8_6925, \9254 );
and \U$17124 ( \26246 , RIee23e60_4867, \9256 );
and \U$17125 ( \26247 , RIfce66f0_7644, \9258 );
and \U$17126 ( \26248 , RIdee4cb0_1067, \9260 );
and \U$17127 ( \26249 , RIdee2f28_1046, \9262 );
and \U$17128 ( \26250 , RIdee0d68_1022, \9264 );
and \U$17129 ( \26251 , RIdeded10_999, \9266 );
and \U$17130 ( \26252 , RIfcca388_7323, \9268 );
and \U$17131 ( \26253 , RIfce6858_7645, \9270 );
and \U$17132 ( \26254 , RIfcceca8_7375, \9272 );
and \U$17133 ( \26255 , RIfcdc970_7532, \9274 );
and \U$17134 ( \26256 , RIded9b80_941, \9276 );
and \U$17135 ( \26257 , RIfeaaac0_8258, \9278 );
and \U$17136 ( \26258 , RIded5800_893, \9280 );
and \U$17137 ( \26259 , RIded3208_866, \9282 );
and \U$17138 ( \26260 , RIded0c10_839, \9284 );
and \U$17139 ( \26261 , RIdecdf10_807, \9286 );
and \U$17140 ( \26262 , RIdecb210_775, \9288 );
and \U$17141 ( \26263 , RIdec8510_743, \9290 );
and \U$17142 ( \26264 , RIdeb4a10_519, \9292 );
and \U$17143 ( \26265 , RIde972f8_327, \9294 );
and \U$17144 ( \26266 , RIe16e618_2633, \9296 );
and \U$17145 ( \26267 , RIe15a410_2404, \9298 );
and \U$17146 ( \26268 , RIe143c10_2148, \9300 );
and \U$17147 ( \26269 , RIdf38608_2018, \9302 );
and \U$17148 ( \26270 , RIdf2cc68_1886, \9304 );
and \U$17149 ( \26271 , RIdf1d4e8_1710, \9306 );
and \U$17150 ( \26272 , RIdf00be0_1385, \9308 );
and \U$17151 ( \26273 , RIdee76e0_1097, \9310 );
and \U$17152 ( \26274 , RIdedc448_970, \9312 );
and \U$17153 ( \26275 , RIde7d240_200, \9314 );
or \U$17154 ( \26276 , \26212 , \26213 , \26214 , \26215 , \26216 , \26217 , \26218 , \26219 , \26220 , \26221 , \26222 , \26223 , \26224 , \26225 , \26226 , \26227 , \26228 , \26229 , \26230 , \26231 , \26232 , \26233 , \26234 , \26235 , \26236 , \26237 , \26238 , \26239 , \26240 , \26241 , \26242 , \26243 , \26244 , \26245 , \26246 , \26247 , \26248 , \26249 , \26250 , \26251 , \26252 , \26253 , \26254 , \26255 , \26256 , \26257 , \26258 , \26259 , \26260 , \26261 , \26262 , \26263 , \26264 , \26265 , \26266 , \26267 , \26268 , \26269 , \26270 , \26271 , \26272 , \26273 , \26274 , \26275 );
or \U$17155 ( \26277 , \26211 , \26276 );
_DC g25d8 ( \26278_nG25d8 , \26277 , \9323 );
buf \U$17156 ( \26279 , \26278_nG25d8 );
and \U$17157 ( \26280 , RIe19daa8_3171, \9333 );
and \U$17158 ( \26281 , RIe19ada8_3139, \9335 );
and \U$17159 ( \26282 , RIf1457c0_5250, \9337 );
and \U$17160 ( \26283 , RIe1980a8_3107, \9339 );
and \U$17161 ( \26284 , RIf1449b0_5240, \9341 );
and \U$17162 ( \26285 , RIe1953a8_3075, \9343 );
and \U$17163 ( \26286 , RIe1926a8_3043, \9345 );
and \U$17164 ( \26287 , RIe18f9a8_3011, \9347 );
and \U$17165 ( \26288 , RIe189fa8_2947, \9349 );
and \U$17166 ( \26289 , RIe1872a8_2915, \9351 );
and \U$17167 ( \26290 , RIf143ba0_5230, \9353 );
and \U$17168 ( \26291 , RIe1845a8_2883, \9355 );
and \U$17169 ( \26292 , RIfc912e0_6674, \9357 );
and \U$17170 ( \26293 , RIe1818a8_2851, \9359 );
and \U$17171 ( \26294 , RIe17eba8_2819, \9361 );
and \U$17172 ( \26295 , RIe17bea8_2787, \9363 );
and \U$17173 ( \26296 , RIfc915b0_6676, \9365 );
and \U$17174 ( \26297 , RIfcbe5b0_7188, \9367 );
and \U$17175 ( \26298 , RIfce3b58_7613, \9369 );
and \U$17176 ( \26299 , RIe175da0_2718, \9371 );
and \U$17177 ( \26300 , RIfceb448_7699, \9373 );
and \U$17178 ( \26301 , RIfcc7958_7293, \9375 );
and \U$17179 ( \26302 , RIfc42de8_5783, \9377 );
and \U$17180 ( \26303 , RIfc96e48_6739, \9379 );
and \U$17181 ( \26304 , RIfc7a810_6416, \9381 );
and \U$17182 ( \26305 , RIfc96ce0_6738, \9383 );
and \U$17183 ( \26306 , RIfcc7ac0_7294, \9385 );
and \U$17184 ( \26307 , RIe173be0_2694, \9387 );
and \U$17185 ( \26308 , RIfce39f0_7612, \9389 );
and \U$17186 ( \26309 , RIfc7a540_6414, \9391 );
and \U$17187 ( \26310 , RIfc91b50_6680, \9393 );
and \U$17188 ( \26311 , RIfc429b0_5780, \9395 );
and \U$17189 ( \26312 , RIfea9710_8244, \9397 );
and \U$17190 ( \26313 , RIe223e00_4698, \9399 );
and \U$17191 ( \26314 , RIfcd8488_7483, \9401 );
and \U$17192 ( \26315 , RIe221100_4666, \9403 );
and \U$17193 ( \26316 , RIfc920f0_6684, \9405 );
and \U$17194 ( \26317 , RIe21e400_4634, \9407 );
and \U$17195 ( \26318 , RIe218a00_4570, \9409 );
and \U$17196 ( \26319 , RIe215d00_4538, \9411 );
and \U$17197 ( \26320 , RIfc79e38_6409, \9413 );
and \U$17198 ( \26321 , RIe213000_4506, \9415 );
and \U$17199 ( \26322 , RIfcbee20_7194, \9417 );
and \U$17200 ( \26323 , RIe210300_4474, \9419 );
and \U$17201 ( \26324 , RIf168068_5643, \9421 );
and \U$17202 ( \26325 , RIe20d600_4442, \9423 );
and \U$17203 ( \26326 , RIe20a900_4410, \9425 );
and \U$17204 ( \26327 , RIe207c00_4378, \9427 );
and \U$17205 ( \26328 , RIfc5af38_6057, \9429 );
and \U$17206 ( \26329 , RIfcd73a8_7471, \9431 );
and \U$17207 ( \26330 , RIe2027a0_4318, \9433 );
and \U$17208 ( \26331 , RIe200ce8_4299, \9435 );
and \U$17209 ( \26332 , RIfcb2670_7052, \9437 );
and \U$17210 ( \26333 , RIfcdf940_7566, \9439 );
and \U$17211 ( \26334 , RIfc5b208_6059, \9441 );
and \U$17212 ( \26335 , RIfcbf3c0_7198, \9443 );
and \U$17213 ( \26336 , RIf1604a8_5555, \9445 );
and \U$17214 ( \26337 , RIf15e5b8_5533, \9447 );
and \U$17215 ( \26338 , RIfe872a0_7882, \9449 );
and \U$17216 ( \26339 , RIfe87138_7881, \9451 );
and \U$17217 ( \26340 , RIfc78920_6394, \9453 );
and \U$17218 ( \26341 , RIfec1158_8317, \9455 );
and \U$17219 ( \26342 , RIfc93338_6697, \9457 );
and \U$17220 ( \26343 , RIfcea368_7687, \9459 );
or \U$17221 ( \26344 , \26280 , \26281 , \26282 , \26283 , \26284 , \26285 , \26286 , \26287 , \26288 , \26289 , \26290 , \26291 , \26292 , \26293 , \26294 , \26295 , \26296 , \26297 , \26298 , \26299 , \26300 , \26301 , \26302 , \26303 , \26304 , \26305 , \26306 , \26307 , \26308 , \26309 , \26310 , \26311 , \26312 , \26313 , \26314 , \26315 , \26316 , \26317 , \26318 , \26319 , \26320 , \26321 , \26322 , \26323 , \26324 , \26325 , \26326 , \26327 , \26328 , \26329 , \26330 , \26331 , \26332 , \26333 , \26334 , \26335 , \26336 , \26337 , \26338 , \26339 , \26340 , \26341 , \26342 , \26343 );
and \U$17222 ( \26345 , RIfcb23a0_7050, \9462 );
and \U$17223 ( \26346 , RIfc5bbe0_6066, \9464 );
and \U$17224 ( \26347 , RIfcede78_7729, \9466 );
and \U$17225 ( \26348 , RIe1fa370_4224, \9468 );
and \U$17226 ( \26349 , RIfcd4c48_7443, \9470 );
and \U$17227 ( \26350 , RIfce1dd0_7592, \9472 );
and \U$17228 ( \26351 , RIfcbf960_7202, \9474 );
and \U$17229 ( \26352 , RIe1f58e8_4171, \9476 );
and \U$17230 ( \26353 , RIfcbfc30_7204, \9478 );
and \U$17231 ( \26354 , RIfc78380_6390, \9480 );
and \U$17232 ( \26355 , RIfc93770_6700, \9482 );
and \U$17233 ( \26356 , RIe1f35c0_4146, \9484 );
and \U$17234 ( \26357 , RIfcb1f68_7047, \9486 );
and \U$17235 ( \26358 , RIfce1b00_7590, \9488 );
and \U$17236 ( \26359 , RIfc93a40_6702, \9490 );
and \U$17237 ( \26360 , RIe1ee2c8_4087, \9492 );
and \U$17238 ( \26361 , RIe1ebb68_4059, \9494 );
and \U$17239 ( \26362 , RIe1e8e68_4027, \9496 );
and \U$17240 ( \26363 , RIe1e6168_3995, \9498 );
and \U$17241 ( \26364 , RIe1e3468_3963, \9500 );
and \U$17242 ( \26365 , RIe1e0768_3931, \9502 );
and \U$17243 ( \26366 , RIe1dda68_3899, \9504 );
and \U$17244 ( \26367 , RIe1dad68_3867, \9506 );
and \U$17245 ( \26368 , RIe1d8068_3835, \9508 );
and \U$17246 ( \26369 , RIe1d2668_3771, \9510 );
and \U$17247 ( \26370 , RIe1cf968_3739, \9512 );
and \U$17248 ( \26371 , RIe1ccc68_3707, \9514 );
and \U$17249 ( \26372 , RIe1c9f68_3675, \9516 );
and \U$17250 ( \26373 , RIe1c7268_3643, \9518 );
and \U$17251 ( \26374 , RIe1c4568_3611, \9520 );
and \U$17252 ( \26375 , RIe1c1868_3579, \9522 );
and \U$17253 ( \26376 , RIe1beb68_3547, \9524 );
and \U$17254 ( \26377 , RIfcdec98_7557, \9526 );
and \U$17255 ( \26378 , RIfc94148_6707, \9528 );
and \U$17256 ( \26379 , RIe1b95a0_3486, \9530 );
and \U$17257 ( \26380 , RIe1b7548_3463, \9532 );
and \U$17258 ( \26381 , RIfcd12a0_7402, \9534 );
and \U$17259 ( \26382 , RIfceabd8_7693, \9536 );
and \U$17260 ( \26383 , RIe1b5388_3439, \9538 );
and \U$17261 ( \26384 , RIe1b3fd8_3425, \9540 );
and \U$17262 ( \26385 , RIfc94850_6712, \9542 );
and \U$17263 ( \26386 , RIfcd7c18_7477, \9544 );
and \U$17264 ( \26387 , RIe1b27f0_3408, \9546 );
and \U$17265 ( \26388 , RIe1b0d38_3389, \9548 );
and \U$17266 ( \26389 , RIfc76a30_6372, \9550 );
and \U$17267 ( \26390 , RIfce2640_7598, \9552 );
and \U$17268 ( \26391 , RIe1ac6e8_3339, \9554 );
and \U$17269 ( \26392 , RIe1ab068_3323, \9556 );
and \U$17270 ( \26393 , RIe1a8ea8_3299, \9558 );
and \U$17271 ( \26394 , RIe1a61a8_3267, \9560 );
and \U$17272 ( \26395 , RIe1a34a8_3235, \9562 );
and \U$17273 ( \26396 , RIe1a07a8_3203, \9564 );
and \U$17274 ( \26397 , RIe18cca8_2979, \9566 );
and \U$17275 ( \26398 , RIe1791a8_2755, \9568 );
and \U$17276 ( \26399 , RIe226b00_4730, \9570 );
and \U$17277 ( \26400 , RIe21b700_4602, \9572 );
and \U$17278 ( \26401 , RIe204f00_4346, \9574 );
and \U$17279 ( \26402 , RIe1fef60_4278, \9576 );
and \U$17280 ( \26403 , RIe1f8318_4201, \9578 );
and \U$17281 ( \26404 , RIe1f0e60_4118, \9580 );
and \U$17282 ( \26405 , RIe1d5368_3803, \9582 );
and \U$17283 ( \26406 , RIe1bbe68_3515, \9584 );
and \U$17284 ( \26407 , RIe1aece0_3366, \9586 );
and \U$17285 ( \26408 , RIe171318_2665, \9588 );
or \U$17286 ( \26409 , \26345 , \26346 , \26347 , \26348 , \26349 , \26350 , \26351 , \26352 , \26353 , \26354 , \26355 , \26356 , \26357 , \26358 , \26359 , \26360 , \26361 , \26362 , \26363 , \26364 , \26365 , \26366 , \26367 , \26368 , \26369 , \26370 , \26371 , \26372 , \26373 , \26374 , \26375 , \26376 , \26377 , \26378 , \26379 , \26380 , \26381 , \26382 , \26383 , \26384 , \26385 , \26386 , \26387 , \26388 , \26389 , \26390 , \26391 , \26392 , \26393 , \26394 , \26395 , \26396 , \26397 , \26398 , \26399 , \26400 , \26401 , \26402 , \26403 , \26404 , \26405 , \26406 , \26407 , \26408 );
or \U$17287 ( \26410 , \26344 , \26409 );
_DC g3705 ( \26411_nG3705 , \26410 , \9597 );
buf \U$17288 ( \26412 , \26411_nG3705 );
and \U$17289 ( \26413 , \26279 , \26412 );
and \U$17290 ( \26414 , \24373 , \24506 );
and \U$17291 ( \26415 , \24506 , \24781 );
and \U$17292 ( \26416 , \24373 , \24781 );
or \U$17293 ( \26417 , \26414 , \26415 , \26416 );
and \U$17294 ( \26418 , \26412 , \26417 );
and \U$17295 ( \26419 , \26279 , \26417 );
or \U$17296 ( \26420 , \26413 , \26418 , \26419 );
xor \U$17297 ( \26421 , \26146 , \26420 );
buf g440c ( \26422_nG440c , \26421 );
xor \U$17298 ( \26423 , \26279 , \26412 );
xor \U$17299 ( \26424 , \26423 , \26417 );
buf g440f ( \26425_nG440f , \26424 );
nand \U$17300 ( \26426 , \26425_nG440f , \24783_nG4412 );
and \U$17301 ( \26427 , \26422_nG440c , \26426 );
xor \U$17302 ( \26428 , \26425_nG440f , \24783_nG4412 );
not \U$17303 ( \26429 , \26428 );
xor \U$17304 ( \26430 , \26422_nG440c , \26425_nG440f );
and \U$17305 ( \26431 , \26429 , \26430 );
and \U$17307 ( \26432 , \26428 , \10694_nG9c0e );
or \U$17308 ( \26433 , 1'b0 , \26432 );
xor \U$17309 ( \26434 , \26427 , \26433 );
xor \U$17310 ( \26435 , \26427 , \26434 );
buf \U$17311 ( \26436 , \26435 );
buf \U$17312 ( \26437 , \26436 );
xor \U$17313 ( \26438 , \25879 , \26437 );
and \U$17314 ( \26439 , \25449 , \25454 );
and \U$17315 ( \26440 , \25449 , \25867 );
and \U$17316 ( \26441 , \25454 , \25867 );
or \U$17317 ( \26442 , \26439 , \26440 , \26441 );
and \U$17318 ( \26443 , \26438 , \26442 );
and \U$17319 ( \26444 , \25460 , \25465 );
and \U$17320 ( \26445 , \25460 , \25865 );
and \U$17321 ( \26446 , \25465 , \25865 );
or \U$17322 ( \26447 , \26444 , \26445 , \26446 );
buf \U$17323 ( \26448 , \26447 );
and \U$17324 ( \26449 , \25343 , \25349 );
and \U$17325 ( \26450 , \25343 , \25356 );
and \U$17326 ( \26451 , \25349 , \25356 );
or \U$17327 ( \26452 , \26449 , \26450 , \26451 );
buf \U$17328 ( \26453 , \26452 );
and \U$17329 ( \26454 , \24792 , \10995_nG9c0b );
and \U$17330 ( \26455 , \24789 , \11283_nG9c08 );
or \U$17331 ( \26456 , \26454 , \26455 );
xor \U$17332 ( \26457 , \24788 , \26456 );
buf \U$17333 ( \26458 , \26457 );
buf \U$17335 ( \26459 , \26458 );
and \U$17336 ( \26460 , \23201 , \11598_nG9c05 );
and \U$17337 ( \26461 , \23198 , \12470_nG9c02 );
or \U$17338 ( \26462 , \26460 , \26461 );
xor \U$17339 ( \26463 , \23197 , \26462 );
buf \U$17340 ( \26464 , \26463 );
buf \U$17342 ( \26465 , \26464 );
xor \U$17343 ( \26466 , \26459 , \26465 );
buf \U$17344 ( \26467 , \26466 );
xor \U$17345 ( \26468 , \26453 , \26467 );
and \U$17346 ( \26469 , \18702 , \15373_nG9bf3 );
and \U$17347 ( \26470 , \18699 , \16315_nG9bf0 );
or \U$17348 ( \26471 , \26469 , \26470 );
xor \U$17349 ( \26472 , \18698 , \26471 );
buf \U$17350 ( \26473 , \26472 );
buf \U$17352 ( \26474 , \26473 );
xor \U$17353 ( \26475 , \26468 , \26474 );
buf \U$17354 ( \26476 , \26475 );
and \U$17355 ( \26477 , \15940 , \18107_nG9be7 );
and \U$17356 ( \26478 , \15937 , \19091_nG9be4 );
or \U$17357 ( \26479 , \26477 , \26478 );
xor \U$17358 ( \26480 , \15936 , \26479 );
buf \U$17359 ( \26481 , \26480 );
buf \U$17361 ( \26482 , \26481 );
xor \U$17362 ( \26483 , \26476 , \26482 );
and \U$17363 ( \26484 , \14631 , \19586_nG9be1 );
and \U$17364 ( \26485 , \14628 , \20608_nG9bde );
or \U$17365 ( \26486 , \26484 , \26485 );
xor \U$17366 ( \26487 , \14627 , \26486 );
buf \U$17367 ( \26488 , \26487 );
buf \U$17369 ( \26489 , \26488 );
xor \U$17370 ( \26490 , \26483 , \26489 );
buf \U$17371 ( \26491 , \26490 );
and \U$17372 ( \26492 , \25367 , \25373 );
and \U$17373 ( \26493 , \25367 , \25380 );
and \U$17374 ( \26494 , \25373 , \25380 );
or \U$17375 ( \26495 , \26492 , \26493 , \26494 );
buf \U$17376 ( \26496 , \26495 );
xor \U$17377 ( \26497 , \26491 , \26496 );
and \U$17378 ( \26498 , \10707 , \25860_nG9bc9 );
and \U$17379 ( \26499 , \25480 , \25786 );
and \U$17380 ( \26500 , \25786 , \25848 );
and \U$17381 ( \26501 , \25480 , \25848 );
or \U$17382 ( \26502 , \26499 , \26500 , \26501 );
and \U$17383 ( \26503 , \25810 , \25831 );
and \U$17384 ( \26504 , \25831 , \25846 );
and \U$17385 ( \26505 , \25810 , \25846 );
or \U$17386 ( \26506 , \26503 , \26504 , \26505 );
and \U$17387 ( \26507 , \25488 , \25492 );
and \U$17388 ( \26508 , \25492 , \25497 );
and \U$17389 ( \26509 , \25488 , \25497 );
or \U$17390 ( \26510 , \26507 , \26508 , \26509 );
and \U$17391 ( \26511 , \25818 , \25822 );
and \U$17392 ( \26512 , \25822 , \25830 );
and \U$17393 ( \26513 , \25818 , \25830 );
or \U$17394 ( \26514 , \26511 , \26512 , \26513 );
xor \U$17395 ( \26515 , \26510 , \26514 );
and \U$17396 ( \26516 , \22556 , \12790 );
and \U$17397 ( \26517 , \23617 , \12461 );
nor \U$17398 ( \26518 , \26516 , \26517 );
xnor \U$17399 ( \26519 , \26518 , \12780 );
and \U$17400 ( \26520 , \18035 , \16635 );
and \U$17401 ( \26521 , \19032 , \16301 );
nor \U$17402 ( \26522 , \26520 , \26521 );
xnor \U$17403 ( \26523 , \26522 , \16625 );
xor \U$17404 ( \26524 , \26519 , \26523 );
and \U$17405 ( \26525 , \10988 , \25826 );
and \U$17406 ( \26526 , \11270 , \25264 );
nor \U$17407 ( \26527 , \26525 , \26526 );
xnor \U$17408 ( \26528 , \26527 , \25773 );
xor \U$17409 ( \26529 , \26524 , \26528 );
xor \U$17410 ( \26530 , \26515 , \26529 );
xor \U$17411 ( \26531 , \26506 , \26530 );
and \U$17412 ( \26532 , \24199 , \11574 );
and \U$17413 ( \26533 , \25272 , \11278 );
nor \U$17414 ( \26534 , \26532 , \26533 );
xnor \U$17415 ( \26535 , \26534 , \11580 );
and \U$17416 ( \26536 , \21033 , \14054 );
and \U$17417 ( \26537 , \22090 , \13692 );
nor \U$17418 ( \26538 , \26536 , \26537 );
xnor \U$17419 ( \26539 , \26538 , \14035 );
xor \U$17420 ( \26540 , \26535 , \26539 );
and \U$17421 ( \26541 , RIdec5810_711, \9333 );
and \U$17422 ( \26542 , RIdec2b10_679, \9335 );
and \U$17423 ( \26543 , RIfce6f60_7650, \9337 );
and \U$17424 ( \26544 , RIdebfe10_647, \9339 );
and \U$17425 ( \26545 , RIfc95228_6719, \9341 );
and \U$17426 ( \26546 , RIdebd110_615, \9343 );
and \U$17427 ( \26547 , RIdeba410_583, \9345 );
and \U$17428 ( \26548 , RIdeb7710_551, \9347 );
and \U$17429 ( \26549 , RIfe879a8_7887, \9349 );
and \U$17430 ( \26550 , RIdeb1d10_487, \9351 );
and \U$17431 ( \26551 , RIfcc16e8_7223, \9353 );
and \U$17432 ( \26552 , RIdeaf010_455, \9355 );
and \U$17433 ( \26553 , RIfca4f48_6899, \9357 );
and \U$17434 ( \26554 , RIdeaadf8_423, \9359 );
and \U$17435 ( \26555 , RIdea44f8_391, \9361 );
and \U$17436 ( \26556 , RIde9dbf8_359, \9363 );
and \U$17437 ( \26557 , RIee1cf48_4788, \9365 );
and \U$17438 ( \26558 , RIee1bfd0_4777, \9367 );
and \U$17439 ( \26559 , RIfc95660_6722, \9369 );
and \U$17440 ( \26560 , RIfcee148_7731, \9371 );
and \U$17441 ( \26561 , RIfe87840_7886, \9373 );
and \U$17442 ( \26562 , RIfe876d8_7885, \9375 );
and \U$17443 ( \26563 , RIde8a0f8_263, \9377 );
and \U$17444 ( \26564 , RIde85f58_243, \9379 );
and \U$17445 ( \26565 , RIfcb0780_7030, \9381 );
and \U$17446 ( \26566 , RIfcee9b8_7737, \9383 );
and \U$17447 ( \26567 , RIfc5f150_6104, \9385 );
and \U$17448 ( \26568 , RIfcdee00_7558, \9387 );
and \U$17449 ( \26569 , RIfcd8050_7480, \9389 );
and \U$17450 ( \26570 , RIe16ba80_2602, \9391 );
and \U$17451 ( \26571 , RIfca5380_6902, \9393 );
and \U$17452 ( \26572 , RIe1680d8_2561, \9395 );
and \U$17453 ( \26573 , RIe165810_2532, \9397 );
and \U$17454 ( \26574 , RIe162b10_2500, \9399 );
and \U$17455 ( \26575 , RIee377f8_5090, \9401 );
and \U$17456 ( \26576 , RIe15fe10_2468, \9403 );
and \U$17457 ( \26577 , RIee36448_5076, \9405 );
and \U$17458 ( \26578 , RIe15d110_2436, \9407 );
and \U$17459 ( \26579 , RIe157710_2372, \9409 );
and \U$17460 ( \26580 , RIe154a10_2340, \9411 );
and \U$17461 ( \26581 , RIfc3f3c8_5745, \9413 );
and \U$17462 ( \26582 , RIe151d10_2308, \9415 );
and \U$17463 ( \26583 , RIfcde9c8_7555, \9417 );
and \U$17464 ( \26584 , RIe14f010_2276, \9419 );
and \U$17465 ( \26585 , RIfc4a2a0_5866, \9421 );
and \U$17466 ( \26586 , RIe14c310_2244, \9423 );
and \U$17467 ( \26587 , RIe149610_2212, \9425 );
and \U$17468 ( \26588 , RIe146910_2180, \9427 );
and \U$17469 ( \26589 , RIfc62288_6139, \9429 );
and \U$17470 ( \26590 , RIee33478_5042, \9431 );
and \U$17471 ( \26591 , RIfc71b70_6316, \9433 );
and \U$17472 ( \26592 , RIee312b8_5018, \9435 );
and \U$17473 ( \26593 , RIe1411e0_2118, \9437 );
and \U$17474 ( \26594 , RIfe87570_7884, \9439 );
and \U$17475 ( \26595 , RIdf3cf28_2070, \9441 );
and \U$17476 ( \26596 , RIfe87408_7883, \9443 );
and \U$17477 ( \26597 , RIfcc99b0_7316, \9445 );
and \U$17478 ( \26598 , RIfccf0e0_7378, \9447 );
and \U$17479 ( \26599 , RIfcaeb60_7010, \9449 );
and \U$17480 ( \26600 , RIfcca220_7322, \9451 );
and \U$17481 ( \26601 , RIdf35bd8_1988, \9453 );
and \U$17482 ( \26602 , RIdf33748_1962, \9455 );
and \U$17483 ( \26603 , RIdf31588_1938, \9457 );
and \U$17484 ( \26604 , RIdf2f530_1915, \9459 );
or \U$17485 ( \26605 , \26541 , \26542 , \26543 , \26544 , \26545 , \26546 , \26547 , \26548 , \26549 , \26550 , \26551 , \26552 , \26553 , \26554 , \26555 , \26556 , \26557 , \26558 , \26559 , \26560 , \26561 , \26562 , \26563 , \26564 , \26565 , \26566 , \26567 , \26568 , \26569 , \26570 , \26571 , \26572 , \26573 , \26574 , \26575 , \26576 , \26577 , \26578 , \26579 , \26580 , \26581 , \26582 , \26583 , \26584 , \26585 , \26586 , \26587 , \26588 , \26589 , \26590 , \26591 , \26592 , \26593 , \26594 , \26595 , \26596 , \26597 , \26598 , \26599 , \26600 , \26601 , \26602 , \26603 , \26604 );
and \U$17486 ( \26606 , RIee2be58_4958, \9462 );
and \U$17487 ( \26607 , RIee2a508_4940, \9464 );
and \U$17488 ( \26608 , RIee28ff0_4925, \9466 );
and \U$17489 ( \26609 , RIee27da8_4912, \9468 );
and \U$17490 ( \26610 , RIdf2a508_1858, \9470 );
and \U$17491 ( \26611 , RIdf28348_1834, \9472 );
and \U$17492 ( \26612 , RIdf265c0_1813, \9474 );
and \U$17493 ( \26613 , RIdf24b08_1794, \9476 );
and \U$17494 ( \26614 , RIfc74708_6347, \9478 );
and \U$17495 ( \26615 , RIfc42578_5777, \9480 );
and \U$17496 ( \26616 , RIfc43388_5787, \9482 );
and \U$17497 ( \26617 , RIfc745a0_6346, \9484 );
and \U$17498 ( \26618 , RIfcb0078_7025, \9486 );
and \U$17499 ( \26619 , RIdf1fc48_1738, \9488 );
and \U$17500 ( \26620 , RIfcaff10_7024, \9490 );
and \U$17501 ( \26621 , RIdf195a0_1665, \9492 );
and \U$17502 ( \26622 , RIdf173e0_1641, \9494 );
and \U$17503 ( \26623 , RIdf146e0_1609, \9496 );
and \U$17504 ( \26624 , RIdf119e0_1577, \9498 );
and \U$17505 ( \26625 , RIdf0ece0_1545, \9500 );
and \U$17506 ( \26626 , RIdf0bfe0_1513, \9502 );
and \U$17507 ( \26627 , RIdf092e0_1481, \9504 );
and \U$17508 ( \26628 , RIdf065e0_1449, \9506 );
and \U$17509 ( \26629 , RIdf038e0_1417, \9508 );
and \U$17510 ( \26630 , RIdefdee0_1353, \9510 );
and \U$17511 ( \26631 , RIdefb1e0_1321, \9512 );
and \U$17512 ( \26632 , RIdef84e0_1289, \9514 );
and \U$17513 ( \26633 , RIdef57e0_1257, \9516 );
and \U$17514 ( \26634 , RIdef2ae0_1225, \9518 );
and \U$17515 ( \26635 , RIdeefde0_1193, \9520 );
and \U$17516 ( \26636 , RIdeed0e0_1161, \9522 );
and \U$17517 ( \26637 , RIdeea3e0_1129, \9524 );
and \U$17518 ( \26638 , RIee257b0_4885, \9526 );
and \U$17519 ( \26639 , RIfca73d8_6925, \9528 );
and \U$17520 ( \26640 , RIee23e60_4867, \9530 );
and \U$17521 ( \26641 , RIfce66f0_7644, \9532 );
and \U$17522 ( \26642 , RIdee4cb0_1067, \9534 );
and \U$17523 ( \26643 , RIdee2f28_1046, \9536 );
and \U$17524 ( \26644 , RIdee0d68_1022, \9538 );
and \U$17525 ( \26645 , RIdeded10_999, \9540 );
and \U$17526 ( \26646 , RIfcca388_7323, \9542 );
and \U$17527 ( \26647 , RIfce6858_7645, \9544 );
and \U$17528 ( \26648 , RIfcceca8_7375, \9546 );
and \U$17529 ( \26649 , RIfcdc970_7532, \9548 );
and \U$17530 ( \26650 , RIded9b80_941, \9550 );
and \U$17531 ( \26651 , RIfeaaac0_8258, \9552 );
and \U$17532 ( \26652 , RIded5800_893, \9554 );
and \U$17533 ( \26653 , RIded3208_866, \9556 );
and \U$17534 ( \26654 , RIded0c10_839, \9558 );
and \U$17535 ( \26655 , RIdecdf10_807, \9560 );
and \U$17536 ( \26656 , RIdecb210_775, \9562 );
and \U$17537 ( \26657 , RIdec8510_743, \9564 );
and \U$17538 ( \26658 , RIdeb4a10_519, \9566 );
and \U$17539 ( \26659 , RIde972f8_327, \9568 );
and \U$17540 ( \26660 , RIe16e618_2633, \9570 );
and \U$17541 ( \26661 , RIe15a410_2404, \9572 );
and \U$17542 ( \26662 , RIe143c10_2148, \9574 );
and \U$17543 ( \26663 , RIdf38608_2018, \9576 );
and \U$17544 ( \26664 , RIdf2cc68_1886, \9578 );
and \U$17545 ( \26665 , RIdf1d4e8_1710, \9580 );
and \U$17546 ( \26666 , RIdf00be0_1385, \9582 );
and \U$17547 ( \26667 , RIdee76e0_1097, \9584 );
and \U$17548 ( \26668 , RIdedc448_970, \9586 );
and \U$17549 ( \26669 , RIde7d240_200, \9588 );
or \U$17550 ( \26670 , \26606 , \26607 , \26608 , \26609 , \26610 , \26611 , \26612 , \26613 , \26614 , \26615 , \26616 , \26617 , \26618 , \26619 , \26620 , \26621 , \26622 , \26623 , \26624 , \26625 , \26626 , \26627 , \26628 , \26629 , \26630 , \26631 , \26632 , \26633 , \26634 , \26635 , \26636 , \26637 , \26638 , \26639 , \26640 , \26641 , \26642 , \26643 , \26644 , \26645 , \26646 , \26647 , \26648 , \26649 , \26650 , \26651 , \26652 , \26653 , \26654 , \26655 , \26656 , \26657 , \26658 , \26659 , \26660 , \26661 , \26662 , \26663 , \26664 , \26665 , \26666 , \26667 , \26668 , \26669 );
or \U$17551 ( \26671 , \26605 , \26670 );
_DC g5db2 ( \26672_nG5db2 , \26671 , \9597 );
and \U$17552 ( \26673 , RIe19daa8_3171, \9059 );
and \U$17553 ( \26674 , RIe19ada8_3139, \9061 );
and \U$17554 ( \26675 , RIf1457c0_5250, \9063 );
and \U$17555 ( \26676 , RIe1980a8_3107, \9065 );
and \U$17556 ( \26677 , RIf1449b0_5240, \9067 );
and \U$17557 ( \26678 , RIe1953a8_3075, \9069 );
and \U$17558 ( \26679 , RIe1926a8_3043, \9071 );
and \U$17559 ( \26680 , RIe18f9a8_3011, \9073 );
and \U$17560 ( \26681 , RIe189fa8_2947, \9075 );
and \U$17561 ( \26682 , RIe1872a8_2915, \9077 );
and \U$17562 ( \26683 , RIf143ba0_5230, \9079 );
and \U$17563 ( \26684 , RIe1845a8_2883, \9081 );
and \U$17564 ( \26685 , RIfc912e0_6674, \9083 );
and \U$17565 ( \26686 , RIe1818a8_2851, \9085 );
and \U$17566 ( \26687 , RIe17eba8_2819, \9087 );
and \U$17567 ( \26688 , RIe17bea8_2787, \9089 );
and \U$17568 ( \26689 , RIfc915b0_6676, \9091 );
and \U$17569 ( \26690 , RIfcbe5b0_7188, \9093 );
and \U$17570 ( \26691 , RIfce3b58_7613, \9095 );
and \U$17571 ( \26692 , RIe175da0_2718, \9097 );
and \U$17572 ( \26693 , RIfceb448_7699, \9099 );
and \U$17573 ( \26694 , RIfcc7958_7293, \9101 );
and \U$17574 ( \26695 , RIfc42de8_5783, \9103 );
and \U$17575 ( \26696 , RIfc96e48_6739, \9105 );
and \U$17576 ( \26697 , RIfc7a810_6416, \9107 );
and \U$17577 ( \26698 , RIfc96ce0_6738, \9109 );
and \U$17578 ( \26699 , RIfcc7ac0_7294, \9111 );
and \U$17579 ( \26700 , RIe173be0_2694, \9113 );
and \U$17580 ( \26701 , RIfce39f0_7612, \9115 );
and \U$17581 ( \26702 , RIfc7a540_6414, \9117 );
and \U$17582 ( \26703 , RIfc91b50_6680, \9119 );
and \U$17583 ( \26704 , RIfc429b0_5780, \9121 );
and \U$17584 ( \26705 , RIfea9710_8244, \9123 );
and \U$17585 ( \26706 , RIe223e00_4698, \9125 );
and \U$17586 ( \26707 , RIfcd8488_7483, \9127 );
and \U$17587 ( \26708 , RIe221100_4666, \9129 );
and \U$17588 ( \26709 , RIfc920f0_6684, \9131 );
and \U$17589 ( \26710 , RIe21e400_4634, \9133 );
and \U$17590 ( \26711 , RIe218a00_4570, \9135 );
and \U$17591 ( \26712 , RIe215d00_4538, \9137 );
and \U$17592 ( \26713 , RIfc79e38_6409, \9139 );
and \U$17593 ( \26714 , RIe213000_4506, \9141 );
and \U$17594 ( \26715 , RIfcbee20_7194, \9143 );
and \U$17595 ( \26716 , RIe210300_4474, \9145 );
and \U$17596 ( \26717 , RIf168068_5643, \9147 );
and \U$17597 ( \26718 , RIe20d600_4442, \9149 );
and \U$17598 ( \26719 , RIe20a900_4410, \9151 );
and \U$17599 ( \26720 , RIe207c00_4378, \9153 );
and \U$17600 ( \26721 , RIfc5af38_6057, \9155 );
and \U$17601 ( \26722 , RIfcd73a8_7471, \9157 );
and \U$17602 ( \26723 , RIe2027a0_4318, \9159 );
and \U$17603 ( \26724 , RIe200ce8_4299, \9161 );
and \U$17604 ( \26725 , RIfcb2670_7052, \9163 );
and \U$17605 ( \26726 , RIfcdf940_7566, \9165 );
and \U$17606 ( \26727 , RIfc5b208_6059, \9167 );
and \U$17607 ( \26728 , RIfcbf3c0_7198, \9169 );
and \U$17608 ( \26729 , RIf1604a8_5555, \9171 );
and \U$17609 ( \26730 , RIf15e5b8_5533, \9173 );
and \U$17610 ( \26731 , RIfe872a0_7882, \9175 );
and \U$17611 ( \26732 , RIfe87138_7881, \9177 );
and \U$17612 ( \26733 , RIfc78920_6394, \9179 );
and \U$17613 ( \26734 , RIfec1158_8317, \9181 );
and \U$17614 ( \26735 , RIfc93338_6697, \9183 );
and \U$17615 ( \26736 , RIfcea368_7687, \9185 );
or \U$17616 ( \26737 , \26673 , \26674 , \26675 , \26676 , \26677 , \26678 , \26679 , \26680 , \26681 , \26682 , \26683 , \26684 , \26685 , \26686 , \26687 , \26688 , \26689 , \26690 , \26691 , \26692 , \26693 , \26694 , \26695 , \26696 , \26697 , \26698 , \26699 , \26700 , \26701 , \26702 , \26703 , \26704 , \26705 , \26706 , \26707 , \26708 , \26709 , \26710 , \26711 , \26712 , \26713 , \26714 , \26715 , \26716 , \26717 , \26718 , \26719 , \26720 , \26721 , \26722 , \26723 , \26724 , \26725 , \26726 , \26727 , \26728 , \26729 , \26730 , \26731 , \26732 , \26733 , \26734 , \26735 , \26736 );
and \U$17617 ( \26738 , RIfcb23a0_7050, \9188 );
and \U$17618 ( \26739 , RIfc5bbe0_6066, \9190 );
and \U$17619 ( \26740 , RIfcede78_7729, \9192 );
and \U$17620 ( \26741 , RIe1fa370_4224, \9194 );
and \U$17621 ( \26742 , RIfcd4c48_7443, \9196 );
and \U$17622 ( \26743 , RIfce1dd0_7592, \9198 );
and \U$17623 ( \26744 , RIfcbf960_7202, \9200 );
and \U$17624 ( \26745 , RIe1f58e8_4171, \9202 );
and \U$17625 ( \26746 , RIfcbfc30_7204, \9204 );
and \U$17626 ( \26747 , RIfc78380_6390, \9206 );
and \U$17627 ( \26748 , RIfc93770_6700, \9208 );
and \U$17628 ( \26749 , RIe1f35c0_4146, \9210 );
and \U$17629 ( \26750 , RIfcb1f68_7047, \9212 );
and \U$17630 ( \26751 , RIfce1b00_7590, \9214 );
and \U$17631 ( \26752 , RIfc93a40_6702, \9216 );
and \U$17632 ( \26753 , RIe1ee2c8_4087, \9218 );
and \U$17633 ( \26754 , RIe1ebb68_4059, \9220 );
and \U$17634 ( \26755 , RIe1e8e68_4027, \9222 );
and \U$17635 ( \26756 , RIe1e6168_3995, \9224 );
and \U$17636 ( \26757 , RIe1e3468_3963, \9226 );
and \U$17637 ( \26758 , RIe1e0768_3931, \9228 );
and \U$17638 ( \26759 , RIe1dda68_3899, \9230 );
and \U$17639 ( \26760 , RIe1dad68_3867, \9232 );
and \U$17640 ( \26761 , RIe1d8068_3835, \9234 );
and \U$17641 ( \26762 , RIe1d2668_3771, \9236 );
and \U$17642 ( \26763 , RIe1cf968_3739, \9238 );
and \U$17643 ( \26764 , RIe1ccc68_3707, \9240 );
and \U$17644 ( \26765 , RIe1c9f68_3675, \9242 );
and \U$17645 ( \26766 , RIe1c7268_3643, \9244 );
and \U$17646 ( \26767 , RIe1c4568_3611, \9246 );
and \U$17647 ( \26768 , RIe1c1868_3579, \9248 );
and \U$17648 ( \26769 , RIe1beb68_3547, \9250 );
and \U$17649 ( \26770 , RIfcdec98_7557, \9252 );
and \U$17650 ( \26771 , RIfc94148_6707, \9254 );
and \U$17651 ( \26772 , RIe1b95a0_3486, \9256 );
and \U$17652 ( \26773 , RIe1b7548_3463, \9258 );
and \U$17653 ( \26774 , RIfcd12a0_7402, \9260 );
and \U$17654 ( \26775 , RIfceabd8_7693, \9262 );
and \U$17655 ( \26776 , RIe1b5388_3439, \9264 );
and \U$17656 ( \26777 , RIe1b3fd8_3425, \9266 );
and \U$17657 ( \26778 , RIfc94850_6712, \9268 );
and \U$17658 ( \26779 , RIfcd7c18_7477, \9270 );
and \U$17659 ( \26780 , RIe1b27f0_3408, \9272 );
and \U$17660 ( \26781 , RIe1b0d38_3389, \9274 );
and \U$17661 ( \26782 , RIfc76a30_6372, \9276 );
and \U$17662 ( \26783 , RIfce2640_7598, \9278 );
and \U$17663 ( \26784 , RIe1ac6e8_3339, \9280 );
and \U$17664 ( \26785 , RIe1ab068_3323, \9282 );
and \U$17665 ( \26786 , RIe1a8ea8_3299, \9284 );
and \U$17666 ( \26787 , RIe1a61a8_3267, \9286 );
and \U$17667 ( \26788 , RIe1a34a8_3235, \9288 );
and \U$17668 ( \26789 , RIe1a07a8_3203, \9290 );
and \U$17669 ( \26790 , RIe18cca8_2979, \9292 );
and \U$17670 ( \26791 , RIe1791a8_2755, \9294 );
and \U$17671 ( \26792 , RIe226b00_4730, \9296 );
and \U$17672 ( \26793 , RIe21b700_4602, \9298 );
and \U$17673 ( \26794 , RIe204f00_4346, \9300 );
and \U$17674 ( \26795 , RIe1fef60_4278, \9302 );
and \U$17675 ( \26796 , RIe1f8318_4201, \9304 );
and \U$17676 ( \26797 , RIe1f0e60_4118, \9306 );
and \U$17677 ( \26798 , RIe1d5368_3803, \9308 );
and \U$17678 ( \26799 , RIe1bbe68_3515, \9310 );
and \U$17679 ( \26800 , RIe1aece0_3366, \9312 );
and \U$17680 ( \26801 , RIe171318_2665, \9314 );
or \U$17681 ( \26802 , \26738 , \26739 , \26740 , \26741 , \26742 , \26743 , \26744 , \26745 , \26746 , \26747 , \26748 , \26749 , \26750 , \26751 , \26752 , \26753 , \26754 , \26755 , \26756 , \26757 , \26758 , \26759 , \26760 , \26761 , \26762 , \26763 , \26764 , \26765 , \26766 , \26767 , \26768 , \26769 , \26770 , \26771 , \26772 , \26773 , \26774 , \26775 , \26776 , \26777 , \26778 , \26779 , \26780 , \26781 , \26782 , \26783 , \26784 , \26785 , \26786 , \26787 , \26788 , \26789 , \26790 , \26791 , \26792 , \26793 , \26794 , \26795 , \26796 , \26797 , \26798 , \26799 , \26800 , \26801 );
or \U$17682 ( \26803 , \26737 , \26802 );
_DC g5e36 ( \26804_nG5e36 , \26803 , \9323 );
xor g5e37 ( \26805_nG5e37 , \26672_nG5db2 , \26804_nG5e36 );
buf \U$17683 ( \26806 , \26805_nG5e37 );
xor \U$17684 ( \26807 , \26806 , \25770 );
and \U$17685 ( \26808 , \10687 , \26807 );
xor \U$17686 ( \26809 , \26540 , \26808 );
and \U$17687 ( \26810 , \19558 , \15336 );
and \U$17688 ( \26811 , \20544 , \14963 );
nor \U$17689 ( \26812 , \26810 , \26811 );
xnor \U$17690 ( \26813 , \26812 , \15342 );
and \U$17691 ( \26814 , \15321 , \19534 );
and \U$17692 ( \26815 , \16267 , \19045 );
nor \U$17693 ( \26816 , \26814 , \26815 );
xnor \U$17694 ( \26817 , \26816 , \19540 );
xor \U$17695 ( \26818 , \26813 , \26817 );
and \U$17696 ( \26819 , \14024 , \21005 );
and \U$17697 ( \26820 , \14950 , \20557 );
nor \U$17698 ( \26821 , \26819 , \26820 );
xnor \U$17699 ( \26822 , \26821 , \21011 );
xor \U$17700 ( \26823 , \26818 , \26822 );
xor \U$17701 ( \26824 , \26809 , \26823 );
and \U$17702 ( \26825 , \25815 , \10983 );
_DC g65bf ( \26826_nG65bf , \26671 , \9597 );
_DC g65c0 ( \26827_nG65c0 , \26803 , \9323 );
and g65c1 ( \26828_nG65c1 , \26826_nG65bf , \26827_nG65c0 );
buf \U$17703 ( \26829 , \26828_nG65c1 );
and \U$17704 ( \26830 , \26829 , \10691 );
nor \U$17705 ( \26831 , \26825 , \26830 );
xnor \U$17706 ( \26832 , \26831 , \10980 );
and \U$17707 ( \26833 , \12769 , \22542 );
and \U$17708 ( \26834 , \13679 , \22103 );
nor \U$17709 ( \26835 , \26833 , \26834 );
xnor \U$17710 ( \26836 , \26835 , \22548 );
xor \U$17711 ( \26837 , \26832 , \26836 );
and \U$17712 ( \26838 , \11586 , \24138 );
and \U$17713 ( \26839 , \12448 , \23630 );
nor \U$17714 ( \26840 , \26838 , \26839 );
xnor \U$17715 ( \26841 , \26840 , \24144 );
xor \U$17716 ( \26842 , \26837 , \26841 );
xor \U$17717 ( \26843 , \26824 , \26842 );
xor \U$17718 ( \26844 , \26531 , \26843 );
xor \U$17719 ( \26845 , \26502 , \26844 );
and \U$17720 ( \26846 , \25484 , \25498 );
and \U$17721 ( \26847 , \25498 , \25785 );
and \U$17722 ( \26848 , \25484 , \25785 );
or \U$17723 ( \26849 , \26846 , \26847 , \26848 );
and \U$17724 ( \26850 , \25791 , \25805 );
and \U$17725 ( \26851 , \25805 , \25847 );
and \U$17726 ( \26852 , \25791 , \25847 );
or \U$17727 ( \26853 , \26850 , \26851 , \26852 );
xor \U$17728 ( \26854 , \26849 , \26853 );
and \U$17729 ( \26855 , \25795 , \25799 );
and \U$17730 ( \26856 , \25799 , \25804 );
and \U$17731 ( \26857 , \25795 , \25804 );
or \U$17732 ( \26858 , \26855 , \26856 , \26857 );
and \U$17733 ( \26859 , \25775 , \25779 );
and \U$17734 ( \26860 , \25779 , \25784 );
and \U$17735 ( \26861 , \25775 , \25784 );
or \U$17736 ( \26862 , \26859 , \26860 , \26861 );
xor \U$17737 ( \26863 , \26858 , \26862 );
and \U$17738 ( \26864 , \25836 , \25840 );
and \U$17739 ( \26865 , \25840 , \25845 );
and \U$17740 ( \26866 , \25836 , \25845 );
or \U$17741 ( \26867 , \26864 , \26865 , \26866 );
and \U$17742 ( \26868 , \25503 , \25774 );
xor \U$17743 ( \26869 , \26867 , \26868 );
and \U$17744 ( \26870 , \16655 , \18090 );
and \U$17745 ( \26871 , \17627 , \17655 );
nor \U$17746 ( \26872 , \26870 , \26871 );
xnor \U$17747 ( \26873 , \26872 , \18046 );
xor \U$17748 ( \26874 , \26869 , \26873 );
xor \U$17749 ( \26875 , \26863 , \26874 );
xor \U$17750 ( \26876 , \26854 , \26875 );
xor \U$17751 ( \26877 , \26845 , \26876 );
and \U$17752 ( \26878 , \25471 , \25475 );
and \U$17753 ( \26879 , \25475 , \25849 );
and \U$17754 ( \26880 , \25471 , \25849 );
or \U$17755 ( \26881 , \26878 , \26879 , \26880 );
xor \U$17756 ( \26882 , \26877 , \26881 );
and \U$17757 ( \26883 , \25850 , \25854 );
and \U$17758 ( \26884 , \25855 , \25858 );
or \U$17759 ( \26885 , \26883 , \26884 );
xor \U$17760 ( \26886 , \26882 , \26885 );
buf g9bc6 ( \26887_nG9bc6 , \26886 );
and \U$17761 ( \26888 , \10704 , \26887_nG9bc6 );
or \U$17762 ( \26889 , \26498 , \26888 );
xor \U$17763 ( \26890 , \10703 , \26889 );
buf \U$17764 ( \26891 , \26890 );
buf \U$17766 ( \26892 , \26891 );
xor \U$17767 ( \26893 , \26497 , \26892 );
buf \U$17768 ( \26894 , \26893 );
xor \U$17769 ( \26895 , \26448 , \26894 );
and \U$17770 ( \26896 , \25382 , \25413 );
and \U$17771 ( \26897 , \25382 , \25420 );
and \U$17772 ( \26898 , \25413 , \25420 );
or \U$17773 ( \26899 , \26896 , \26897 , \26898 );
buf \U$17774 ( \26900 , \26899 );
xor \U$17775 ( \26901 , \26895 , \26900 );
buf \U$17776 ( \26902 , \26901 );
and \U$17777 ( \26903 , \25433 , \25438 );
and \U$17778 ( \26904 , \25433 , \25445 );
and \U$17779 ( \26905 , \25438 , \25445 );
or \U$17780 ( \26906 , \26903 , \26904 , \26905 );
buf \U$17781 ( \26907 , \26906 );
and \U$17782 ( \26908 , \25387 , \25404 );
and \U$17783 ( \26909 , \25387 , \25411 );
and \U$17784 ( \26910 , \25404 , \25411 );
or \U$17785 ( \26911 , \26908 , \26909 , \26910 );
buf \U$17786 ( \26912 , \26911 );
and \U$17787 ( \26913 , \12157 , \22629_nG9bd5 );
and \U$17788 ( \26914 , \12154 , \23696_nG9bd2 );
or \U$17789 ( \26915 , \26913 , \26914 );
xor \U$17790 ( \26916 , \12153 , \26915 );
buf \U$17791 ( \26917 , \26916 );
buf \U$17793 ( \26918 , \26917 );
xor \U$17794 ( \26919 , \26912 , \26918 );
and \U$17795 ( \26920 , \10421 , \24226_nG9bcf );
and \U$17796 ( \26921 , \10418 , \25298_nG9bcc );
or \U$17797 ( \26922 , \26920 , \26921 );
xor \U$17798 ( \26923 , \10417 , \26922 );
buf \U$17799 ( \26924 , \26923 );
buf \U$17801 ( \26925 , \26924 );
xor \U$17802 ( \26926 , \26919 , \26925 );
buf \U$17803 ( \26927 , \26926 );
xor \U$17804 ( \26928 , \26907 , \26927 );
and \U$17805 ( \26929 , \25389 , \25395 );
and \U$17806 ( \26930 , \25389 , \25402 );
and \U$17807 ( \26931 , \25395 , \25402 );
or \U$17808 ( \26932 , \26929 , \26930 , \26931 );
buf \U$17809 ( \26933 , \26932 );
and \U$17810 ( \26934 , \25335 , \25341 );
buf \U$17811 ( \26935 , \26934 );
and \U$17812 ( \26936 , \21658 , \12801_nG9bff );
and \U$17813 ( \26937 , \21655 , \13705_nG9bfc );
or \U$17814 ( \26938 , \26936 , \26937 );
xor \U$17815 ( \26939 , \21654 , \26938 );
buf \U$17816 ( \26940 , \26939 );
buf \U$17818 ( \26941 , \26940 );
xor \U$17819 ( \26942 , \26935 , \26941 );
and \U$17820 ( \26943 , \20155 , \14070_nG9bf9 );
and \U$17821 ( \26944 , \20152 , \14984_nG9bf6 );
or \U$17822 ( \26945 , \26943 , \26944 );
xor \U$17823 ( \26946 , \20151 , \26945 );
buf \U$17824 ( \26947 , \26946 );
buf \U$17826 ( \26948 , \26947 );
xor \U$17827 ( \26949 , \26942 , \26948 );
buf \U$17828 ( \26950 , \26949 );
xor \U$17829 ( \26951 , \26933 , \26950 );
and \U$17830 ( \26952 , \17297 , \16680_nG9bed );
and \U$17831 ( \26953 , \17294 , \17665_nG9bea );
or \U$17832 ( \26954 , \26952 , \26953 );
xor \U$17833 ( \26955 , \17293 , \26954 );
buf \U$17834 ( \26956 , \26955 );
buf \U$17836 ( \26957 , \26956 );
xor \U$17837 ( \26958 , \26951 , \26957 );
buf \U$17838 ( \26959 , \26958 );
and \U$17839 ( \26960 , \25332 , \25358 );
and \U$17840 ( \26961 , \25332 , \25365 );
and \U$17841 ( \26962 , \25358 , \25365 );
or \U$17842 ( \26963 , \26960 , \26961 , \26962 );
buf \U$17843 ( \26964 , \26963 );
xor \U$17844 ( \26965 , \26959 , \26964 );
and \U$17845 ( \26966 , \13370 , \21086_nG9bdb );
and \U$17846 ( \26967 , \13367 , \22129_nG9bd8 );
or \U$17847 ( \26968 , \26966 , \26967 );
xor \U$17848 ( \26969 , \13366 , \26968 );
buf \U$17849 ( \26970 , \26969 );
buf \U$17851 ( \26971 , \26970 );
xor \U$17852 ( \26972 , \26965 , \26971 );
buf \U$17853 ( \26973 , \26972 );
xor \U$17854 ( \26974 , \26928 , \26973 );
buf \U$17855 ( \26975 , \26974 );
xor \U$17856 ( \26976 , \26902 , \26975 );
and \U$17857 ( \26977 , \25422 , \25427 );
and \U$17858 ( \26978 , \25422 , \25447 );
and \U$17859 ( \26979 , \25427 , \25447 );
or \U$17860 ( \26980 , \26977 , \26978 , \26979 );
buf \U$17861 ( \26981 , \26980 );
xor \U$17862 ( \26982 , \26976 , \26981 );
and \U$17863 ( \26983 , \26438 , \26982 );
and \U$17864 ( \26984 , \26442 , \26982 );
or \U$17865 ( \26985 , \26443 , \26983 , \26984 );
and \U$17866 ( \26986 , \25874 , \25878 );
and \U$17867 ( \26987 , \25874 , \26437 );
and \U$17868 ( \26988 , \25878 , \26437 );
or \U$17869 ( \26989 , \26986 , \26987 , \26988 );
xor \U$17870 ( \26990 , \26985 , \26989 );
and \U$17871 ( \26991 , \26902 , \26975 );
and \U$17872 ( \26992 , \26902 , \26981 );
and \U$17873 ( \26993 , \26975 , \26981 );
or \U$17874 ( \26994 , \26991 , \26992 , \26993 );
xor \U$17875 ( \26995 , \26990 , \26994 );
and \U$17876 ( \26996 , \26907 , \26927 );
and \U$17877 ( \26997 , \26907 , \26973 );
and \U$17878 ( \26998 , \26927 , \26973 );
or \U$17879 ( \26999 , \26996 , \26997 , \26998 );
buf \U$17880 ( \27000 , \26999 );
and \U$17881 ( \27001 , \26959 , \26964 );
and \U$17882 ( \27002 , \26959 , \26971 );
and \U$17883 ( \27003 , \26964 , \26971 );
or \U$17884 ( \27004 , \27001 , \27002 , \27003 );
buf \U$17885 ( \27005 , \27004 );
and \U$17886 ( \27006 , \10421 , \25298_nG9bcc );
and \U$17887 ( \27007 , \10418 , \25860_nG9bc9 );
or \U$17888 ( \27008 , \27006 , \27007 );
xor \U$17889 ( \27009 , \10417 , \27008 );
buf \U$17890 ( \27010 , \27009 );
buf \U$17892 ( \27011 , \27010 );
xor \U$17893 ( \27012 , \27005 , \27011 );
and \U$17894 ( \27013 , \10707 , \26887_nG9bc6 );
and \U$17895 ( \27014 , \26849 , \26853 );
and \U$17896 ( \27015 , \26853 , \26875 );
and \U$17897 ( \27016 , \26849 , \26875 );
or \U$17898 ( \27017 , \27014 , \27015 , \27016 );
and \U$17899 ( \27018 , \26510 , \26514 );
and \U$17900 ( \27019 , \26514 , \26529 );
and \U$17901 ( \27020 , \26510 , \26529 );
or \U$17902 ( \27021 , \27018 , \27019 , \27020 );
and \U$17903 ( \27022 , \25272 , \11574 );
and \U$17904 ( \27023 , \25815 , \11278 );
nor \U$17905 ( \27024 , \27022 , \27023 );
xnor \U$17906 ( \27025 , \27024 , \11580 );
not \U$17907 ( \27026 , \26808 );
and \U$17908 ( \27027 , RIdec5978_712, \9333 );
and \U$17909 ( \27028 , RIdec2c78_680, \9335 );
and \U$17910 ( \27029 , RIfc8aad0_6600, \9337 );
and \U$17911 ( \27030 , RIdebff78_648, \9339 );
and \U$17912 ( \27031 , RIfc8ac38_6601, \9341 );
and \U$17913 ( \27032 , RIdebd278_616, \9343 );
and \U$17914 ( \27033 , RIdeba578_584, \9345 );
and \U$17915 ( \27034 , RIdeb7878_552, \9347 );
and \U$17916 ( \27035 , RIfc40e80_5764, \9349 );
and \U$17917 ( \27036 , RIdeb1e78_488, \9351 );
and \U$17918 ( \27037 , RIfcdaeb8_7513, \9353 );
and \U$17919 ( \27038 , RIdeaf178_456, \9355 );
and \U$17920 ( \27039 , RIee1dbf0_4797, \9357 );
and \U$17921 ( \27040 , RIdeab140_424, \9359 );
and \U$17922 ( \27041 , RIdea4840_392, \9361 );
and \U$17923 ( \27042 , RIde9df40_360, \9363 );
and \U$17924 ( \27043 , RIfc8b070_6604, \9365 );
and \U$17925 ( \27044 , RIfcc38a8_7247, \9367 );
and \U$17926 ( \27045 , RIfc807b0_6484, \9369 );
and \U$17927 ( \27046 , RIfcbb8b0_7156, \9371 );
and \U$17928 ( \27047 , RIde91a60_300, \9373 );
and \U$17929 ( \27048 , RIde8e298_283, \9375 );
and \U$17930 ( \27049 , RIde8a440_264, \9377 );
and \U$17931 ( \27050 , RIde862a0_244, \9379 );
and \U$17932 ( \27051 , RIde82100_224, \9381 );
and \U$17933 ( \27052 , RIfcbbb80_7158, \9383 );
and \U$17934 ( \27053 , RIfc8c150_6616, \9385 );
and \U$17935 ( \27054 , RIfcbbfb8_7161, \9387 );
and \U$17936 ( \27055 , RIfc54458_5981, \9389 );
and \U$17937 ( \27056 , RIe16bbe8_2603, \9391 );
and \U$17938 ( \27057 , RIfc8c2b8_6617, \9393 );
and \U$17939 ( \27058 , RIe168240_2562, \9395 );
and \U$17940 ( \27059 , RIe165978_2533, \9397 );
and \U$17941 ( \27060 , RIe162c78_2501, \9399 );
and \U$17942 ( \27061 , RIee37960_5091, \9401 );
and \U$17943 ( \27062 , RIe15ff78_2469, \9403 );
and \U$17944 ( \27063 , RIfcd6b38_7465, \9405 );
and \U$17945 ( \27064 , RIe15d278_2437, \9407 );
and \U$17946 ( \27065 , RIe157878_2373, \9409 );
and \U$17947 ( \27066 , RIe154b78_2341, \9411 );
and \U$17948 ( \27067 , RIfc8e5e0_6642, \9413 );
and \U$17949 ( \27068 , RIe151e78_2309, \9415 );
and \U$17950 ( \27069 , RIfcb4290_7072, \9417 );
and \U$17951 ( \27070 , RIe14f178_2277, \9419 );
and \U$17952 ( \27071 , RIfc56ff0_6012, \9421 );
and \U$17953 ( \27072 , RIe14c478_2245, \9423 );
and \U$17954 ( \27073 , RIe149778_2213, \9425 );
and \U$17955 ( \27074 , RIe146a78_2181, \9427 );
and \U$17956 ( \27075 , RIee346c0_5055, \9429 );
and \U$17957 ( \27076 , RIee335e0_5043, \9431 );
and \U$17958 ( \27077 , RIee32398_5030, \9433 );
and \U$17959 ( \27078 , RIee31420_5019, \9435 );
and \U$17960 ( \27079 , RIe141348_2119, \9437 );
and \U$17961 ( \27080 , RIe13f020_2094, \9439 );
and \U$17962 ( \27081 , RIfec16f8_8321, \9441 );
and \U$17963 ( \27082 , RIdf3a930_2043, \9443 );
and \U$17964 ( \27083 , RIfce3e28_7615, \9445 );
and \U$17965 ( \27084 , RIfc56780_6006, \9447 );
and \U$17966 ( \27085 , RIfcb4128_7071, \9449 );
and \U$17967 ( \27086 , RIfce2eb0_7604, \9451 );
and \U$17968 ( \27087 , RIdf35d40_1989, \9453 );
and \U$17969 ( \27088 , RIfe88218_7893, \9455 );
and \U$17970 ( \27089 , RIdf316f0_1939, \9457 );
and \U$17971 ( \27090 , RIdf2f698_1916, \9459 );
or \U$17972 ( \27091 , \27027 , \27028 , \27029 , \27030 , \27031 , \27032 , \27033 , \27034 , \27035 , \27036 , \27037 , \27038 , \27039 , \27040 , \27041 , \27042 , \27043 , \27044 , \27045 , \27046 , \27047 , \27048 , \27049 , \27050 , \27051 , \27052 , \27053 , \27054 , \27055 , \27056 , \27057 , \27058 , \27059 , \27060 , \27061 , \27062 , \27063 , \27064 , \27065 , \27066 , \27067 , \27068 , \27069 , \27070 , \27071 , \27072 , \27073 , \27074 , \27075 , \27076 , \27077 , \27078 , \27079 , \27080 , \27081 , \27082 , \27083 , \27084 , \27085 , \27086 , \27087 , \27088 , \27089 , \27090 );
and \U$17973 ( \27092 , RIfc7f9a0_6474, \9462 );
and \U$17974 ( \27093 , RIfce4260_7618, \9464 );
and \U$17975 ( \27094 , RIfcd62c8_7459, \9466 );
and \U$17976 ( \27095 , RIfce9990_7680, \9468 );
and \U$17977 ( \27096 , RIdf2a670_1859, \9470 );
and \U$17978 ( \27097 , RIdf284b0_1835, \9472 );
and \U$17979 ( \27098 , RIdf26728_1814, \9474 );
and \U$17980 ( \27099 , RIdf24c70_1795, \9476 );
and \U$17981 ( \27100 , RIfc7ecf8_6465, \9478 );
and \U$17982 ( \27101 , RIfcc31a0_7242, \9480 );
and \U$17983 ( \27102 , RIfc99008_6763, \9482 );
and \U$17984 ( \27103 , RIfc46e98_5829, \9484 );
and \U$17985 ( \27104 , RIfce2a78_7601, \9486 );
and \U$17986 ( \27105 , RIdf1fdb0_1739, \9488 );
and \U$17987 ( \27106 , RIfcc6e18_7285, \9490 );
and \U$17988 ( \27107 , RIdf19708_1666, \9492 );
and \U$17989 ( \27108 , RIdf17548_1642, \9494 );
and \U$17990 ( \27109 , RIdf14848_1610, \9496 );
and \U$17991 ( \27110 , RIdf11b48_1578, \9498 );
and \U$17992 ( \27111 , RIdf0ee48_1546, \9500 );
and \U$17993 ( \27112 , RIdf0c148_1514, \9502 );
and \U$17994 ( \27113 , RIdf09448_1482, \9504 );
and \U$17995 ( \27114 , RIdf06748_1450, \9506 );
and \U$17996 ( \27115 , RIdf03a48_1418, \9508 );
and \U$17997 ( \27116 , RIdefe048_1354, \9510 );
and \U$17998 ( \27117 , RIdefb348_1322, \9512 );
and \U$17999 ( \27118 , RIdef8648_1290, \9514 );
and \U$18000 ( \27119 , RIdef5948_1258, \9516 );
and \U$18001 ( \27120 , RIdef2c48_1226, \9518 );
and \U$18002 ( \27121 , RIdeeff48_1194, \9520 );
and \U$18003 ( \27122 , RIdeed248_1162, \9522 );
and \U$18004 ( \27123 , RIdeea548_1130, \9524 );
and \U$18005 ( \27124 , RIfcd9130_7492, \9526 );
and \U$18006 ( \27125 , RIfc7cb38_6441, \9528 );
and \U$18007 ( \27126 , RIfc97af0_6748, \9530 );
and \U$18008 ( \27127 , RIfcb3e58_7069, \9532 );
and \U$18009 ( \27128 , RIdee4e18_1068, \9534 );
and \U$18010 ( \27129 , RIdee3090_1047, \9536 );
and \U$18011 ( \27130 , RIdee0ed0_1023, \9538 );
and \U$18012 ( \27131 , RIfe88380_7894, \9540 );
and \U$18013 ( \27132 , RIfc97dc0_6750, \9542 );
and \U$18014 ( \27133 , RIfcc2930_7236, \9544 );
and \U$18015 ( \27134 , RIfcd9298_7493, \9546 );
and \U$18016 ( \27135 , RIfc7c868_6439, \9548 );
and \U$18017 ( \27136 , RIded9ce8_942, \9550 );
and \U$18018 ( \27137 , RIded76f0_915, \9552 );
and \U$18019 ( \27138 , RIded5968_894, \9554 );
and \U$18020 ( \27139 , RIded3370_867, \9556 );
and \U$18021 ( \27140 , RIded0d78_840, \9558 );
and \U$18022 ( \27141 , RIdece078_808, \9560 );
and \U$18023 ( \27142 , RIdecb378_776, \9562 );
and \U$18024 ( \27143 , RIdec8678_744, \9564 );
and \U$18025 ( \27144 , RIdeb4b78_520, \9566 );
and \U$18026 ( \27145 , RIde97640_328, \9568 );
and \U$18027 ( \27146 , RIe16e780_2634, \9570 );
and \U$18028 ( \27147 , RIe15a578_2405, \9572 );
and \U$18029 ( \27148 , RIe143d78_2149, \9574 );
and \U$18030 ( \27149 , RIdf38770_2019, \9576 );
and \U$18031 ( \27150 , RIdf2cdd0_1887, \9578 );
and \U$18032 ( \27151 , RIdf1d650_1711, \9580 );
and \U$18033 ( \27152 , RIdf00d48_1386, \9582 );
and \U$18034 ( \27153 , RIdee7848_1098, \9584 );
and \U$18035 ( \27154 , RIdedc5b0_971, \9586 );
and \U$18036 ( \27155 , RIde7d588_201, \9588 );
or \U$18037 ( \27156 , \27092 , \27093 , \27094 , \27095 , \27096 , \27097 , \27098 , \27099 , \27100 , \27101 , \27102 , \27103 , \27104 , \27105 , \27106 , \27107 , \27108 , \27109 , \27110 , \27111 , \27112 , \27113 , \27114 , \27115 , \27116 , \27117 , \27118 , \27119 , \27120 , \27121 , \27122 , \27123 , \27124 , \27125 , \27126 , \27127 , \27128 , \27129 , \27130 , \27131 , \27132 , \27133 , \27134 , \27135 , \27136 , \27137 , \27138 , \27139 , \27140 , \27141 , \27142 , \27143 , \27144 , \27145 , \27146 , \27147 , \27148 , \27149 , \27150 , \27151 , \27152 , \27153 , \27154 , \27155 );
or \U$18038 ( \27157 , \27091 , \27156 );
_DC g5ebb ( \27158_nG5ebb , \27157 , \9597 );
and \U$18039 ( \27159 , RIe19dc10_3172, \9059 );
and \U$18040 ( \27160 , RIe19af10_3140, \9061 );
and \U$18041 ( \27161 , RIfec1590_8320, \9063 );
and \U$18042 ( \27162 , RIe198210_3108, \9065 );
and \U$18043 ( \27163 , RIfec1428_8319, \9067 );
and \U$18044 ( \27164 , RIe195510_3076, \9069 );
and \U$18045 ( \27165 , RIe192810_3044, \9071 );
and \U$18046 ( \27166 , RIe18fb10_3012, \9073 );
and \U$18047 ( \27167 , RIe18a110_2948, \9075 );
and \U$18048 ( \27168 , RIe187410_2916, \9077 );
and \U$18049 ( \27169 , RIfec12c0_8318, \9079 );
and \U$18050 ( \27170 , RIe184710_2884, \9081 );
and \U$18051 ( \27171 , RIfc88370_6572, \9083 );
and \U$18052 ( \27172 , RIe181a10_2852, \9085 );
and \U$18053 ( \27173 , RIe17ed10_2820, \9087 );
and \U$18054 ( \27174 , RIe17c010_2788, \9089 );
and \U$18055 ( \27175 , RIfc6ccb0_6260, \9091 );
and \U$18056 ( \27176 , RIfc5f858_6109, \9093 );
and \U$18057 ( \27177 , RIfca88f0_6940, \9095 );
and \U$18058 ( \27178 , RIe175f08_2719, \9097 );
and \U$18059 ( \27179 , RIfc81020_6490, \9099 );
and \U$18060 ( \27180 , RIfcc6008_7275, \9101 );
and \U$18061 ( \27181 , RIfc4ea58_5917, \9103 );
and \U$18062 ( \27182 , RIfc42140_5774, \9105 );
and \U$18063 ( \27183 , RIfca3b98_6885, \9107 );
and \U$18064 ( \27184 , RIfc5ac68_6055, \9109 );
and \U$18065 ( \27185 , RIfc984c8_6755, \9111 );
and \U$18066 ( \27186 , RIe173d48_2695, \9113 );
and \U$18067 ( \27187 , RIfc9b330_6788, \9115 );
and \U$18068 ( \27188 , RIf16f688_5727, \9117 );
and \U$18069 ( \27189 , RIfc42410_5776, \9119 );
and \U$18070 ( \27190 , RIfc5f588_6107, \9121 );
and \U$18071 ( \27191 , RIfe880b0_7892, \9123 );
and \U$18072 ( \27192 , RIe223f68_4699, \9125 );
and \U$18073 ( \27193 , RIf16bfb0_5688, \9127 );
and \U$18074 ( \27194 , RIe221268_4667, \9129 );
and \U$18075 ( \27195 , RIfc86cf0_6556, \9131 );
and \U$18076 ( \27196 , RIe21e568_4635, \9133 );
and \U$18077 ( \27197 , RIe218b68_4571, \9135 );
and \U$18078 ( \27198 , RIe215e68_4539, \9137 );
and \U$18079 ( \27199 , RIfe87de0_7890, \9139 );
and \U$18080 ( \27200 , RIe213168_4507, \9141 );
and \U$18081 ( \27201 , RIf1692b0_5656, \9143 );
and \U$18082 ( \27202 , RIe210468_4475, \9145 );
and \U$18083 ( \27203 , RIfcdf670_7564, \9147 );
and \U$18084 ( \27204 , RIe20d768_4443, \9149 );
and \U$18085 ( \27205 , RIe20aa68_4411, \9151 );
and \U$18086 ( \27206 , RIe207d68_4379, \9153 );
and \U$18087 ( \27207 , RIfca6460_6914, \9155 );
and \U$18088 ( \27208 , RIf1662e0_5622, \9157 );
and \U$18089 ( \27209 , RIe202908_4319, \9159 );
and \U$18090 ( \27210 , RIfe87b10_7888, \9161 );
and \U$18091 ( \27211 , RIfc58c10_6032, \9163 );
and \U$18092 ( \27212 , RIfc50ab0_5940, \9165 );
and \U$18093 ( \27213 , RIfccd790_7360, \9167 );
and \U$18094 ( \27214 , RIfccd1f0_7356, \9169 );
and \U$18095 ( \27215 , RIf160610_5556, \9171 );
and \U$18096 ( \27216 , RIf15e720_5534, \9173 );
and \U$18097 ( \27217 , RIfe87c78_7889, \9175 );
and \U$18098 ( \27218 , RIfe87f48_7891, \9177 );
and \U$18099 ( \27219 , RIfce7668_7655, \9179 );
and \U$18100 ( \27220 , RIfc86480_6550, \9181 );
and \U$18101 ( \27221 , RIfcd2218_7413, \9183 );
and \U$18102 ( \27222 , RIfcb01e0_7026, \9185 );
or \U$18103 ( \27223 , \27159 , \27160 , \27161 , \27162 , \27163 , \27164 , \27165 , \27166 , \27167 , \27168 , \27169 , \27170 , \27171 , \27172 , \27173 , \27174 , \27175 , \27176 , \27177 , \27178 , \27179 , \27180 , \27181 , \27182 , \27183 , \27184 , \27185 , \27186 , \27187 , \27188 , \27189 , \27190 , \27191 , \27192 , \27193 , \27194 , \27195 , \27196 , \27197 , \27198 , \27199 , \27200 , \27201 , \27202 , \27203 , \27204 , \27205 , \27206 , \27207 , \27208 , \27209 , \27210 , \27211 , \27212 , \27213 , \27214 , \27215 , \27216 , \27217 , \27218 , \27219 , \27220 , \27221 , \27222 );
and \U$18104 ( \27224 , RIfc47b40_5838, \9188 );
and \U$18105 ( \27225 , RIfc84158_6525, \9190 );
and \U$18106 ( \27226 , RIfc4b920_5882, \9192 );
and \U$18107 ( \27227 , RIe1fa4d8_4225, \9194 );
and \U$18108 ( \27228 , RIfc4ba88_5883, \9196 );
and \U$18109 ( \27229 , RIfcb7530_7108, \9198 );
and \U$18110 ( \27230 , RIfcd58f0_7452, \9200 );
and \U$18111 ( \27231 , RIe1f5a50_4172, \9202 );
and \U$18112 ( \27232 , RIf153488_5407, \9204 );
and \U$18113 ( \27233 , RIf151ca0_5390, \9206 );
and \U$18114 ( \27234 , RIfc51e60_5954, \9208 );
and \U$18115 ( \27235 , RIe1f3728_4147, \9210 );
and \U$18116 ( \27236 , RIfc9aef8_6785, \9212 );
and \U$18117 ( \27237 , RIfcbaaa0_7146, \9214 );
and \U$18118 ( \27238 , RIfc52130_5956, \9216 );
and \U$18119 ( \27239 , RIe1ee430_4088, \9218 );
and \U$18120 ( \27240 , RIe1ebcd0_4060, \9220 );
and \U$18121 ( \27241 , RIe1e8fd0_4028, \9222 );
and \U$18122 ( \27242 , RIe1e62d0_3996, \9224 );
and \U$18123 ( \27243 , RIe1e35d0_3964, \9226 );
and \U$18124 ( \27244 , RIe1e08d0_3932, \9228 );
and \U$18125 ( \27245 , RIe1ddbd0_3900, \9230 );
and \U$18126 ( \27246 , RIe1daed0_3868, \9232 );
and \U$18127 ( \27247 , RIe1d81d0_3836, \9234 );
and \U$18128 ( \27248 , RIe1d27d0_3772, \9236 );
and \U$18129 ( \27249 , RIe1cfad0_3740, \9238 );
and \U$18130 ( \27250 , RIe1ccdd0_3708, \9240 );
and \U$18131 ( \27251 , RIe1ca0d0_3676, \9242 );
and \U$18132 ( \27252 , RIe1c73d0_3644, \9244 );
and \U$18133 ( \27253 , RIe1c46d0_3612, \9246 );
and \U$18134 ( \27254 , RIe1c19d0_3580, \9248 );
and \U$18135 ( \27255 , RIe1becd0_3548, \9250 );
and \U$18136 ( \27256 , RIfce0b88_7579, \9252 );
and \U$18137 ( \27257 , RIfc82808_6507, \9254 );
and \U$18138 ( \27258 , RIe1b9708_3487, \9256 );
and \U$18139 ( \27259 , RIe1b76b0_3464, \9258 );
and \U$18140 ( \27260 , RIfcd5bc0_7454, \9260 );
and \U$18141 ( \27261 , RIfcb69f0_7100, \9262 );
and \U$18142 ( \27262 , RIe1b54f0_3440, \9264 );
and \U$18143 ( \27263 , RIe1b4140_3426, \9266 );
and \U$18144 ( \27264 , RIfc89f90_6592, \9268 );
and \U$18145 ( \27265 , RIfce9af8_7681, \9270 );
and \U$18146 ( \27266 , RIe1b2958_3409, \9272 );
and \U$18147 ( \27267 , RIe1b0ea0_3390, \9274 );
and \U$18148 ( \27268 , RIfc4a138_5865, \9276 );
and \U$18149 ( \27269 , RIfc8a260_6594, \9278 );
and \U$18150 ( \27270 , RIe1ac850_3340, \9280 );
and \U$18151 ( \27271 , RIe1ab1d0_3324, \9282 );
and \U$18152 ( \27272 , RIe1a9010_3300, \9284 );
and \U$18153 ( \27273 , RIe1a6310_3268, \9286 );
and \U$18154 ( \27274 , RIe1a3610_3236, \9288 );
and \U$18155 ( \27275 , RIe1a0910_3204, \9290 );
and \U$18156 ( \27276 , RIe18ce10_2980, \9292 );
and \U$18157 ( \27277 , RIe179310_2756, \9294 );
and \U$18158 ( \27278 , RIe226c68_4731, \9296 );
and \U$18159 ( \27279 , RIe21b868_4603, \9298 );
and \U$18160 ( \27280 , RIe205068_4347, \9300 );
and \U$18161 ( \27281 , RIe1ff0c8_4279, \9302 );
and \U$18162 ( \27282 , RIe1f8480_4202, \9304 );
and \U$18163 ( \27283 , RIe1f0fc8_4119, \9306 );
and \U$18164 ( \27284 , RIe1d54d0_3804, \9308 );
and \U$18165 ( \27285 , RIe1bbfd0_3516, \9310 );
and \U$18166 ( \27286 , RIe1aee48_3367, \9312 );
and \U$18167 ( \27287 , RIe171480_2666, \9314 );
or \U$18168 ( \27288 , \27224 , \27225 , \27226 , \27227 , \27228 , \27229 , \27230 , \27231 , \27232 , \27233 , \27234 , \27235 , \27236 , \27237 , \27238 , \27239 , \27240 , \27241 , \27242 , \27243 , \27244 , \27245 , \27246 , \27247 , \27248 , \27249 , \27250 , \27251 , \27252 , \27253 , \27254 , \27255 , \27256 , \27257 , \27258 , \27259 , \27260 , \27261 , \27262 , \27263 , \27264 , \27265 , \27266 , \27267 , \27268 , \27269 , \27270 , \27271 , \27272 , \27273 , \27274 , \27275 , \27276 , \27277 , \27278 , \27279 , \27280 , \27281 , \27282 , \27283 , \27284 , \27285 , \27286 , \27287 );
or \U$18169 ( \27289 , \27223 , \27288 );
_DC g5f3f ( \27290_nG5f3f , \27289 , \9323 );
xor g5f40 ( \27291_nG5f40 , \27158_nG5ebb , \27290_nG5f3f );
buf \U$18170 ( \27292 , \27291_nG5f40 );
and \U$18171 ( \27293 , \26806 , \25770 );
not \U$18172 ( \27294 , \27293 );
and \U$18173 ( \27295 , \27292 , \27294 );
and \U$18174 ( \27296 , \27026 , \27295 );
xor \U$18175 ( \27297 , \27025 , \27296 );
and \U$18176 ( \27298 , \26813 , \26817 );
and \U$18177 ( \27299 , \26817 , \26822 );
and \U$18178 ( \27300 , \26813 , \26822 );
or \U$18179 ( \27301 , \27298 , \27299 , \27300 );
xor \U$18180 ( \27302 , \27297 , \27301 );
and \U$18181 ( \27303 , \26832 , \26836 );
and \U$18182 ( \27304 , \26836 , \26841 );
and \U$18183 ( \27305 , \26832 , \26841 );
or \U$18184 ( \27306 , \27303 , \27304 , \27305 );
xor \U$18185 ( \27307 , \27302 , \27306 );
xor \U$18186 ( \27308 , \27021 , \27307 );
and \U$18187 ( \27309 , \26829 , \10983 );
_DC g65c2 ( \27310_nG65c2 , \27157 , \9597 );
_DC g65c3 ( \27311_nG65c3 , \27289 , \9323 );
and g65c4 ( \27312_nG65c4 , \27310_nG65c2 , \27311_nG65c3 );
buf \U$18188 ( \27313 , \27312_nG65c4 );
and \U$18189 ( \27314 , \27313 , \10691 );
nor \U$18190 ( \27315 , \27309 , \27314 );
xnor \U$18191 ( \27316 , \27315 , \10980 );
and \U$18192 ( \27317 , \19032 , \16635 );
and \U$18193 ( \27318 , \19558 , \16301 );
nor \U$18194 ( \27319 , \27317 , \27318 );
xnor \U$18195 ( \27320 , \27319 , \16625 );
xor \U$18196 ( \27321 , \27316 , \27320 );
and \U$18197 ( \27322 , \11270 , \25826 );
and \U$18198 ( \27323 , \11586 , \25264 );
nor \U$18199 ( \27324 , \27322 , \27323 );
xnor \U$18200 ( \27325 , \27324 , \25773 );
xor \U$18201 ( \27326 , \27321 , \27325 );
and \U$18202 ( \27327 , \20544 , \15336 );
and \U$18203 ( \27328 , \21033 , \14963 );
nor \U$18204 ( \27329 , \27327 , \27328 );
xnor \U$18205 ( \27330 , \27329 , \15342 );
and \U$18206 ( \27331 , \13679 , \22542 );
and \U$18207 ( \27332 , \14024 , \22103 );
nor \U$18208 ( \27333 , \27331 , \27332 );
xnor \U$18209 ( \27334 , \27333 , \22548 );
xor \U$18210 ( \27335 , \27330 , \27334 );
and \U$18211 ( \27336 , \12448 , \24138 );
and \U$18212 ( \27337 , \12769 , \23630 );
nor \U$18213 ( \27338 , \27336 , \27337 );
xnor \U$18214 ( \27339 , \27338 , \24144 );
xor \U$18215 ( \27340 , \27335 , \27339 );
xor \U$18216 ( \27341 , \27326 , \27340 );
and \U$18217 ( \27342 , \22090 , \14054 );
and \U$18218 ( \27343 , \22556 , \13692 );
nor \U$18219 ( \27344 , \27342 , \27343 );
xnor \U$18220 ( \27345 , \27344 , \14035 );
and \U$18221 ( \27346 , \16267 , \19534 );
and \U$18222 ( \27347 , \16655 , \19045 );
nor \U$18223 ( \27348 , \27346 , \27347 );
xnor \U$18224 ( \27349 , \27348 , \19540 );
xor \U$18225 ( \27350 , \27345 , \27349 );
and \U$18226 ( \27351 , \14950 , \21005 );
and \U$18227 ( \27352 , \15321 , \20557 );
nor \U$18228 ( \27353 , \27351 , \27352 );
xnor \U$18229 ( \27354 , \27353 , \21011 );
xor \U$18230 ( \27355 , \27350 , \27354 );
xor \U$18231 ( \27356 , \27341 , \27355 );
xor \U$18232 ( \27357 , \27308 , \27356 );
xor \U$18233 ( \27358 , \27017 , \27357 );
and \U$18234 ( \27359 , \26858 , \26862 );
and \U$18235 ( \27360 , \26862 , \26874 );
and \U$18236 ( \27361 , \26858 , \26874 );
or \U$18237 ( \27362 , \27359 , \27360 , \27361 );
and \U$18238 ( \27363 , \26506 , \26530 );
and \U$18239 ( \27364 , \26530 , \26843 );
and \U$18240 ( \27365 , \26506 , \26843 );
or \U$18241 ( \27366 , \27363 , \27364 , \27365 );
xor \U$18242 ( \27367 , \27362 , \27366 );
and \U$18243 ( \27368 , \26867 , \26868 );
and \U$18244 ( \27369 , \26868 , \26873 );
and \U$18245 ( \27370 , \26867 , \26873 );
or \U$18246 ( \27371 , \27368 , \27369 , \27370 );
and \U$18247 ( \27372 , \26809 , \26823 );
and \U$18248 ( \27373 , \26823 , \26842 );
and \U$18249 ( \27374 , \26809 , \26842 );
or \U$18250 ( \27375 , \27372 , \27373 , \27374 );
xor \U$18251 ( \27376 , \27371 , \27375 );
and \U$18252 ( \27377 , \26535 , \26539 );
and \U$18253 ( \27378 , \26539 , \26808 );
and \U$18254 ( \27379 , \26535 , \26808 );
or \U$18255 ( \27380 , \27377 , \27378 , \27379 );
and \U$18256 ( \27381 , \26519 , \26523 );
and \U$18257 ( \27382 , \26523 , \26528 );
and \U$18258 ( \27383 , \26519 , \26528 );
or \U$18259 ( \27384 , \27381 , \27382 , \27383 );
xor \U$18260 ( \27385 , \27380 , \27384 );
and \U$18261 ( \27386 , \23617 , \12790 );
and \U$18262 ( \27387 , \24199 , \12461 );
nor \U$18263 ( \27388 , \27386 , \27387 );
xnor \U$18264 ( \27389 , \27388 , \12780 );
and \U$18265 ( \27390 , \17627 , \18090 );
and \U$18266 ( \27391 , \18035 , \17655 );
nor \U$18267 ( \27392 , \27390 , \27391 );
xnor \U$18268 ( \27393 , \27392 , \18046 );
xor \U$18269 ( \27394 , \27389 , \27393 );
xor \U$18270 ( \27395 , \27292 , \26806 );
not \U$18271 ( \27396 , \26807 );
and \U$18272 ( \27397 , \27395 , \27396 );
and \U$18273 ( \27398 , \10687 , \27397 );
and \U$18274 ( \27399 , \10988 , \26807 );
nor \U$18275 ( \27400 , \27398 , \27399 );
xnor \U$18276 ( \27401 , \27400 , \27295 );
xor \U$18277 ( \27402 , \27394 , \27401 );
xor \U$18278 ( \27403 , \27385 , \27402 );
xor \U$18279 ( \27404 , \27376 , \27403 );
xor \U$18280 ( \27405 , \27367 , \27404 );
xor \U$18281 ( \27406 , \27358 , \27405 );
and \U$18282 ( \27407 , \26502 , \26844 );
and \U$18283 ( \27408 , \26844 , \26876 );
and \U$18284 ( \27409 , \26502 , \26876 );
or \U$18285 ( \27410 , \27407 , \27408 , \27409 );
xor \U$18286 ( \27411 , \27406 , \27410 );
and \U$18287 ( \27412 , \26877 , \26881 );
and \U$18288 ( \27413 , \26882 , \26885 );
or \U$18289 ( \27414 , \27412 , \27413 );
xor \U$18290 ( \27415 , \27411 , \27414 );
buf g9bc3 ( \27416_nG9bc3 , \27415 );
and \U$18291 ( \27417 , \10704 , \27416_nG9bc3 );
or \U$18292 ( \27418 , \27013 , \27417 );
xor \U$18293 ( \27419 , \10703 , \27418 );
buf \U$18294 ( \27420 , \27419 );
buf \U$18296 ( \27421 , \27420 );
xor \U$18297 ( \27422 , \27012 , \27421 );
buf \U$18298 ( \27423 , \27422 );
xor \U$18299 ( \27424 , \27000 , \27423 );
and \U$18300 ( \27425 , \26935 , \26941 );
and \U$18301 ( \27426 , \26935 , \26948 );
and \U$18302 ( \27427 , \26941 , \26948 );
or \U$18303 ( \27428 , \27425 , \27426 , \27427 );
buf \U$18304 ( \27429 , \27428 );
and \U$18305 ( \27430 , \26427 , \26434 );
buf \U$18306 ( \27431 , \27430 );
buf \U$18308 ( \27432 , \27431 );
and \U$18309 ( \27433 , \24792 , \11283_nG9c08 );
and \U$18310 ( \27434 , \24789 , \11598_nG9c05 );
or \U$18311 ( \27435 , \27433 , \27434 );
xor \U$18312 ( \27436 , \24788 , \27435 );
buf \U$18313 ( \27437 , \27436 );
buf \U$18315 ( \27438 , \27437 );
xor \U$18316 ( \27439 , \27432 , \27438 );
buf \U$18317 ( \27440 , \27439 );
and \U$18318 ( \27441 , \26431 , \10694_nG9c0e );
and \U$18319 ( \27442 , \26428 , \10995_nG9c0b );
or \U$18320 ( \27443 , \27441 , \27442 );
xor \U$18321 ( \27444 , \26427 , \27443 );
buf \U$18322 ( \27445 , \27444 );
buf \U$18324 ( \27446 , \27445 );
xor \U$18325 ( \27447 , \27440 , \27446 );
and \U$18326 ( \27448 , \23201 , \12470_nG9c02 );
and \U$18327 ( \27449 , \23198 , \12801_nG9bff );
or \U$18328 ( \27450 , \27448 , \27449 );
xor \U$18329 ( \27451 , \23197 , \27450 );
buf \U$18330 ( \27452 , \27451 );
buf \U$18332 ( \27453 , \27452 );
xor \U$18333 ( \27454 , \27447 , \27453 );
buf \U$18334 ( \27455 , \27454 );
xor \U$18335 ( \27456 , \27429 , \27455 );
and \U$18336 ( \27457 , \18702 , \16315_nG9bf0 );
and \U$18337 ( \27458 , \18699 , \16680_nG9bed );
or \U$18338 ( \27459 , \27457 , \27458 );
xor \U$18339 ( \27460 , \18698 , \27459 );
buf \U$18340 ( \27461 , \27460 );
buf \U$18342 ( \27462 , \27461 );
xor \U$18343 ( \27463 , \27456 , \27462 );
buf \U$18344 ( \27464 , \27463 );
and \U$18345 ( \27465 , \15940 , \19091_nG9be4 );
and \U$18346 ( \27466 , \15937 , \19586_nG9be1 );
or \U$18347 ( \27467 , \27465 , \27466 );
xor \U$18348 ( \27468 , \15936 , \27467 );
buf \U$18349 ( \27469 , \27468 );
buf \U$18351 ( \27470 , \27469 );
xor \U$18352 ( \27471 , \27464 , \27470 );
and \U$18353 ( \27472 , \14631 , \20608_nG9bde );
and \U$18354 ( \27473 , \14628 , \21086_nG9bdb );
or \U$18355 ( \27474 , \27472 , \27473 );
xor \U$18356 ( \27475 , \14627 , \27474 );
buf \U$18357 ( \27476 , \27475 );
buf \U$18359 ( \27477 , \27476 );
xor \U$18360 ( \27478 , \27471 , \27477 );
buf \U$18361 ( \27479 , \27478 );
and \U$18362 ( \27480 , \26459 , \26465 );
buf \U$18363 ( \27481 , \27480 );
and \U$18364 ( \27482 , \21658 , \13705_nG9bfc );
and \U$18365 ( \27483 , \21655 , \14070_nG9bf9 );
or \U$18366 ( \27484 , \27482 , \27483 );
xor \U$18367 ( \27485 , \21654 , \27484 );
buf \U$18368 ( \27486 , \27485 );
buf \U$18370 ( \27487 , \27486 );
xor \U$18371 ( \27488 , \27481 , \27487 );
and \U$18372 ( \27489 , \20155 , \14984_nG9bf6 );
and \U$18373 ( \27490 , \20152 , \15373_nG9bf3 );
or \U$18374 ( \27491 , \27489 , \27490 );
xor \U$18375 ( \27492 , \20151 , \27491 );
buf \U$18376 ( \27493 , \27492 );
buf \U$18378 ( \27494 , \27493 );
xor \U$18379 ( \27495 , \27488 , \27494 );
buf \U$18380 ( \27496 , \27495 );
and \U$18381 ( \27497 , \26453 , \26467 );
and \U$18382 ( \27498 , \26453 , \26474 );
and \U$18383 ( \27499 , \26467 , \26474 );
or \U$18384 ( \27500 , \27497 , \27498 , \27499 );
buf \U$18385 ( \27501 , \27500 );
xor \U$18386 ( \27502 , \27496 , \27501 );
and \U$18387 ( \27503 , \17297 , \17665_nG9bea );
and \U$18388 ( \27504 , \17294 , \18107_nG9be7 );
or \U$18389 ( \27505 , \27503 , \27504 );
xor \U$18390 ( \27506 , \17293 , \27505 );
buf \U$18391 ( \27507 , \27506 );
buf \U$18393 ( \27508 , \27507 );
xor \U$18394 ( \27509 , \27502 , \27508 );
buf \U$18395 ( \27510 , \27509 );
xor \U$18396 ( \27511 , \27479 , \27510 );
and \U$18397 ( \27512 , \12157 , \23696_nG9bd2 );
and \U$18398 ( \27513 , \12154 , \24226_nG9bcf );
or \U$18399 ( \27514 , \27512 , \27513 );
xor \U$18400 ( \27515 , \12153 , \27514 );
buf \U$18401 ( \27516 , \27515 );
buf \U$18403 ( \27517 , \27516 );
xor \U$18404 ( \27518 , \27511 , \27517 );
buf \U$18405 ( \27519 , \27518 );
xor \U$18406 ( \27520 , \27424 , \27519 );
buf \U$18407 ( \27521 , \27520 );
and \U$18408 ( \27522 , \26448 , \26894 );
and \U$18409 ( \27523 , \26448 , \26900 );
and \U$18410 ( \27524 , \26894 , \26900 );
or \U$18411 ( \27525 , \27522 , \27523 , \27524 );
buf \U$18412 ( \27526 , \27525 );
xor \U$18413 ( \27527 , \27521 , \27526 );
and \U$18414 ( \27528 , \26912 , \26918 );
and \U$18415 ( \27529 , \26912 , \26925 );
and \U$18416 ( \27530 , \26918 , \26925 );
or \U$18417 ( \27531 , \27528 , \27529 , \27530 );
buf \U$18418 ( \27532 , \27531 );
and \U$18419 ( \27533 , \26476 , \26482 );
and \U$18420 ( \27534 , \26476 , \26489 );
and \U$18421 ( \27535 , \26482 , \26489 );
or \U$18422 ( \27536 , \27533 , \27534 , \27535 );
buf \U$18423 ( \27537 , \27536 );
and \U$18424 ( \27538 , \26933 , \26950 );
and \U$18425 ( \27539 , \26933 , \26957 );
and \U$18426 ( \27540 , \26950 , \26957 );
or \U$18427 ( \27541 , \27538 , \27539 , \27540 );
buf \U$18428 ( \27542 , \27541 );
xor \U$18429 ( \27543 , \27537 , \27542 );
and \U$18430 ( \27544 , \13370 , \22129_nG9bd8 );
and \U$18431 ( \27545 , \13367 , \22629_nG9bd5 );
or \U$18432 ( \27546 , \27544 , \27545 );
xor \U$18433 ( \27547 , \13366 , \27546 );
buf \U$18434 ( \27548 , \27547 );
buf \U$18436 ( \27549 , \27548 );
xor \U$18437 ( \27550 , \27543 , \27549 );
buf \U$18438 ( \27551 , \27550 );
xor \U$18439 ( \27552 , \27532 , \27551 );
and \U$18440 ( \27553 , \26491 , \26496 );
and \U$18441 ( \27554 , \26491 , \26892 );
and \U$18442 ( \27555 , \26496 , \26892 );
or \U$18443 ( \27556 , \27553 , \27554 , \27555 );
buf \U$18444 ( \27557 , \27556 );
xor \U$18445 ( \27558 , \27552 , \27557 );
buf \U$18446 ( \27559 , \27558 );
xor \U$18447 ( \27560 , \27527 , \27559 );
and \U$18448 ( \27561 , \26995 , \27560 );
and \U$18449 ( \27562 , \26985 , \26989 );
and \U$18450 ( \27563 , \26985 , \26994 );
and \U$18451 ( \27564 , \26989 , \26994 );
or \U$18452 ( \27565 , \27562 , \27563 , \27564 );
xor \U$18453 ( \27566 , \27561 , \27565 );
and \U$18454 ( \27567 , RIdec5c48_714, \9059 );
and \U$18455 ( \27568 , RIdec2f48_682, \9061 );
and \U$18456 ( \27569 , RIfc7c160_6434, \9063 );
and \U$18457 ( \27570 , RIdec0248_650, \9065 );
and \U$18458 ( \27571 , RIfcb38b8_7065, \9067 );
and \U$18459 ( \27572 , RIdebd548_618, \9069 );
and \U$18460 ( \27573 , RIdeba848_586, \9071 );
and \U$18461 ( \27574 , RIdeb7b48_554, \9073 );
and \U$18462 ( \27575 , RIfce7c08_7659, \9075 );
and \U$18463 ( \27576 , RIdeb2148_490, \9077 );
and \U$18464 ( \27577 , RIfce7aa0_7658, \9079 );
and \U$18465 ( \27578 , RIdeaf448_458, \9081 );
and \U$18466 ( \27579 , RIfca38c8_6883, \9083 );
and \U$18467 ( \27580 , RIdeab7d0_426, \9085 );
and \U$18468 ( \27581 , RIdea4ed0_394, \9087 );
and \U$18469 ( \27582 , RIde9e5d0_362, \9089 );
and \U$18470 ( \27583 , RIfc41e70_5772, \9091 );
and \U$18471 ( \27584 , RIfc5b0a0_6058, \9093 );
and \U$18472 ( \27585 , RIfcdbb60_7522, \9095 );
and \U$18473 ( \27586 , RIfc78650_6392, \9097 );
and \U$18474 ( \27587 , RIfea92d8_8241, \9099 );
and \U$18475 ( \27588 , RIde8e5e0_284, \9101 );
and \U$18476 ( \27589 , RIfea0d40_8174, \9103 );
and \U$18477 ( \27590 , RIfea0bd8_8173, \9105 );
and \U$18478 ( \27591 , RIfcdf508_7563, \9107 );
and \U$18479 ( \27592 , RIfcb1b30_7044, \9109 );
and \U$18480 ( \27593 , RIfc5ccc0_6078, \9111 );
and \U$18481 ( \27594 , RIfcb16f8_7041, \9113 );
and \U$18482 ( \27595 , RIfc77b10_6384, \9115 );
and \U$18483 ( \27596 , RIe16beb8_2605, \9117 );
and \U$18484 ( \27597 , RIe169e60_2582, \9119 );
and \U$18485 ( \27598 , RIe168510_2564, \9121 );
and \U$18486 ( \27599 , RIe165c48_2535, \9123 );
and \U$18487 ( \27600 , RIe162f48_2503, \9125 );
and \U$18488 ( \27601 , RIfc4f9d0_5928, \9127 );
and \U$18489 ( \27602 , RIe160248_2471, \9129 );
and \U$18490 ( \27603 , RIfc4e8f0_5916, \9131 );
and \U$18491 ( \27604 , RIe15d548_2439, \9133 );
and \U$18492 ( \27605 , RIe157b48_2375, \9135 );
and \U$18493 ( \27606 , RIe154e48_2343, \9137 );
and \U$18494 ( \27607 , RIfc4e1e8_5911, \9139 );
and \U$18495 ( \27608 , RIe152148_2311, \9141 );
and \U$18496 ( \27609 , RIfc868b8_6553, \9143 );
and \U$18497 ( \27610 , RIe14f448_2279, \9145 );
and \U$18498 ( \27611 , RIfc865e8_6551, \9147 );
and \U$18499 ( \27612 , RIe14c748_2247, \9149 );
and \U$18500 ( \27613 , RIe149a48_2215, \9151 );
and \U$18501 ( \27614 , RIe146d48_2183, \9153 );
and \U$18502 ( \27615 , RIfc9eb70_6828, \9155 );
and \U$18503 ( \27616 , RIfc9ecd8_6829, \9157 );
and \U$18504 ( \27617 , RIfcc5630_7268, \9159 );
and \U$18505 ( \27618 , RIfc83bb8_6521, \9161 );
and \U$18506 ( \27619 , RIe141618_2121, \9163 );
and \U$18507 ( \27620 , RIfea0ea8_8175, \9165 );
and \U$18508 ( \27621 , RIdf3d1f8_2072, \9167 );
and \U$18509 ( \27622 , RIdf3ac00_2045, \9169 );
and \U$18510 ( \27623 , RIee308e0_5011, \9171 );
and \U$18511 ( \27624 , RIfcd3cd0_7432, \9173 );
and \U$18512 ( \27625 , RIfc84e00_6534, \9175 );
and \U$18513 ( \27626 , RIfc834b0_6516, \9177 );
and \U$18514 ( \27627 , RIdf36010_1991, \9179 );
and \U$18515 ( \27628 , RIdf33a18_1964, \9181 );
and \U$18516 ( \27629 , RIdf31858_1940, \9183 );
and \U$18517 ( \27630 , RIdf2f968_1918, \9185 );
or \U$18518 ( \27631 , \27567 , \27568 , \27569 , \27570 , \27571 , \27572 , \27573 , \27574 , \27575 , \27576 , \27577 , \27578 , \27579 , \27580 , \27581 , \27582 , \27583 , \27584 , \27585 , \27586 , \27587 , \27588 , \27589 , \27590 , \27591 , \27592 , \27593 , \27594 , \27595 , \27596 , \27597 , \27598 , \27599 , \27600 , \27601 , \27602 , \27603 , \27604 , \27605 , \27606 , \27607 , \27608 , \27609 , \27610 , \27611 , \27612 , \27613 , \27614 , \27615 , \27616 , \27617 , \27618 , \27619 , \27620 , \27621 , \27622 , \27623 , \27624 , \27625 , \27626 , \27627 , \27628 , \27629 , \27630 );
and \U$18519 ( \27632 , RIee2c128_4960, \9188 );
and \U$18520 ( \27633 , RIee2a7d8_4942, \9190 );
and \U$18521 ( \27634 , RIee292c0_4927, \9192 );
and \U$18522 ( \27635 , RIee28078_4914, \9194 );
and \U$18523 ( \27636 , RIdf2a940_1861, \9196 );
and \U$18524 ( \27637 , RIdf28780_1837, \9198 );
and \U$18525 ( \27638 , RIfea0a70_8172, \9200 );
and \U$18526 ( \27639 , RIfea0908_8171, \9202 );
and \U$18527 ( \27640 , RIfcd4f18_7445, \9204 );
and \U$18528 ( \27641 , RIfca0628_6847, \9206 );
and \U$18529 ( \27642 , RIdf23050_1775, \9208 );
and \U$18530 ( \27643 , RIfcd3190_7424, \9210 );
and \U$18531 ( \27644 , RIdf21b38_1760, \9212 );
and \U$18532 ( \27645 , RIdf20080_1741, \9214 );
and \U$18533 ( \27646 , RIdf1b328_1686, \9216 );
and \U$18534 ( \27647 , RIdf199d8_1668, \9218 );
and \U$18535 ( \27648 , RIdf17818_1644, \9220 );
and \U$18536 ( \27649 , RIdf14b18_1612, \9222 );
and \U$18537 ( \27650 , RIdf11e18_1580, \9224 );
and \U$18538 ( \27651 , RIdf0f118_1548, \9226 );
and \U$18539 ( \27652 , RIdf0c418_1516, \9228 );
and \U$18540 ( \27653 , RIdf09718_1484, \9230 );
and \U$18541 ( \27654 , RIdf06a18_1452, \9232 );
and \U$18542 ( \27655 , RIdf03d18_1420, \9234 );
and \U$18543 ( \27656 , RIdefe318_1356, \9236 );
and \U$18544 ( \27657 , RIdefb618_1324, \9238 );
and \U$18545 ( \27658 , RIdef8918_1292, \9240 );
and \U$18546 ( \27659 , RIdef5c18_1260, \9242 );
and \U$18547 ( \27660 , RIdef2f18_1228, \9244 );
and \U$18548 ( \27661 , RIdef0218_1196, \9246 );
and \U$18549 ( \27662 , RIdeed518_1164, \9248 );
and \U$18550 ( \27663 , RIdeea818_1132, \9250 );
and \U$18551 ( \27664 , RIfcdf3a0_7562, \9252 );
and \U$18552 ( \27665 , RIfca5218_6901, \9254 );
and \U$18553 ( \27666 , RIfcdc538_7529, \9256 );
and \U$18554 ( \27667 , RIfcdc6a0_7530, \9258 );
and \U$18555 ( \27668 , RIdee50e8_1070, \9260 );
and \U$18556 ( \27669 , RIdee3360_1049, \9262 );
and \U$18557 ( \27670 , RIfea07a0_8170, \9264 );
and \U$18558 ( \27671 , RIdedefe0_1001, \9266 );
and \U$18559 ( \27672 , RIfcb0d20_7034, \9268 );
and \U$18560 ( \27673 , RIfcd4978_7441, \9270 );
and \U$18561 ( \27674 , RIfca49a8_6895, \9272 );
and \U$18562 ( \27675 , RIfca1708_6859, \9274 );
and \U$18563 ( \27676 , RIded9fb8_944, \9276 );
and \U$18564 ( \27677 , RIded79c0_917, \9278 );
and \U$18565 ( \27678 , RIded5ad0_895, \9280 );
and \U$18566 ( \27679 , RIfeab498_8265, \9282 );
and \U$18567 ( \27680 , RIded1048_842, \9284 );
and \U$18568 ( \27681 , RIdece348_810, \9286 );
and \U$18569 ( \27682 , RIdecb648_778, \9288 );
and \U$18570 ( \27683 , RIdec8948_746, \9290 );
and \U$18571 ( \27684 , RIdeb4e48_522, \9292 );
and \U$18572 ( \27685 , RIde97cd0_330, \9294 );
and \U$18573 ( \27686 , RIe16ea50_2636, \9296 );
and \U$18574 ( \27687 , RIe15a848_2407, \9298 );
and \U$18575 ( \27688 , RIe144048_2151, \9300 );
and \U$18576 ( \27689 , RIdf38a40_2021, \9302 );
and \U$18577 ( \27690 , RIdf2d0a0_1889, \9304 );
and \U$18578 ( \27691 , RIdf1d920_1713, \9306 );
and \U$18579 ( \27692 , RIdf01018_1388, \9308 );
and \U$18580 ( \27693 , RIdee7b18_1100, \9310 );
and \U$18581 ( \27694 , RIdedc880_973, \9312 );
and \U$18582 ( \27695 , RIde7dc18_203, \9314 );
or \U$18583 ( \27696 , \27632 , \27633 , \27634 , \27635 , \27636 , \27637 , \27638 , \27639 , \27640 , \27641 , \27642 , \27643 , \27644 , \27645 , \27646 , \27647 , \27648 , \27649 , \27650 , \27651 , \27652 , \27653 , \27654 , \27655 , \27656 , \27657 , \27658 , \27659 , \27660 , \27661 , \27662 , \27663 , \27664 , \27665 , \27666 , \27667 , \27668 , \27669 , \27670 , \27671 , \27672 , \27673 , \27674 , \27675 , \27676 , \27677 , \27678 , \27679 , \27680 , \27681 , \27682 , \27683 , \27684 , \27685 , \27686 , \27687 , \27688 , \27689 , \27690 , \27691 , \27692 , \27693 , \27694 , \27695 );
or \U$18584 ( \27697 , \27631 , \27696 );
_DC g2449 ( \27698_nG2449 , \27697 , \9323 );
buf \U$18585 ( \27699 , \27698_nG2449 );
and \U$18586 ( \27700 , RIe19dee0_3174, \9333 );
and \U$18587 ( \27701 , RIe19b1e0_3142, \9335 );
and \U$18588 ( \27702 , RIfc67580_6198, \9337 );
and \U$18589 ( \27703 , RIe1984e0_3110, \9339 );
and \U$18590 ( \27704 , RIfccb030_7332, \9341 );
and \U$18591 ( \27705 , RIe1957e0_3078, \9343 );
and \U$18592 ( \27706 , RIe192ae0_3046, \9345 );
and \U$18593 ( \27707 , RIe18fde0_3014, \9347 );
and \U$18594 ( \27708 , RIe18a3e0_2950, \9349 );
and \U$18595 ( \27709 , RIe1876e0_2918, \9351 );
and \U$18596 ( \27710 , RIfc6a550_6232, \9353 );
and \U$18597 ( \27711 , RIe1849e0_2886, \9355 );
and \U$18598 ( \27712 , RIfcaa7e0_6962, \9357 );
and \U$18599 ( \27713 , RIe181ce0_2854, \9359 );
and \U$18600 ( \27714 , RIe17efe0_2822, \9361 );
and \U$18601 ( \27715 , RIe17c2e0_2790, \9363 );
and \U$18602 ( \27716 , RIfc65d98_6181, \9365 );
and \U$18603 ( \27717 , RIfc65690_6176, \9367 );
and \U$18604 ( \27718 , RIe1772b8_2733, \9369 );
and \U$18605 ( \27719 , RIfea0638_8169, \9371 );
and \U$18606 ( \27720 , RIfcca928_7327, \9373 );
and \U$18607 ( \27721 , RIfc607d0_6120, \9375 );
and \U$18608 ( \27722 , RIfc65258_6173, \9377 );
and \U$18609 ( \27723 , RIee3d798_5158, \9379 );
and \U$18610 ( \27724 , RIee3c3e8_5144, \9381 );
and \U$18611 ( \27725 , RIfca9430_6948, \9383 );
and \U$18612 ( \27726 , RIee39f58_5118, \9385 );
and \U$18613 ( \27727 , RIe174018_2697, \9387 );
and \U$18614 ( \27728 , RIfcecf00_7718, \9389 );
and \U$18615 ( \27729 , RIfc650f0_6172, \9391 );
and \U$18616 ( \27730 , RIf16e5a8_5715, \9393 );
and \U$18617 ( \27731 , RIfc43a90_5792, \9395 );
and \U$18618 ( \27732 , RIfc65528_6175, \9397 );
and \U$18619 ( \27733 , RIe224238_4701, \9399 );
and \U$18620 ( \27734 , RIfca9f70_6956, \9401 );
and \U$18621 ( \27735 , RIe221538_4669, \9403 );
and \U$18622 ( \27736 , RIfc6b4c8_6243, \9405 );
and \U$18623 ( \27737 , RIe21e838_4637, \9407 );
and \U$18624 ( \27738 , RIe218e38_4573, \9409 );
and \U$18625 ( \27739 , RIe216138_4541, \9411 );
and \U$18626 ( \27740 , RIfc3fda0_5752, \9413 );
and \U$18627 ( \27741 , RIe213438_4509, \9415 );
and \U$18628 ( \27742 , RIfc61310_6128, \9417 );
and \U$18629 ( \27743 , RIe210738_4477, \9419 );
and \U$18630 ( \27744 , RIfc60c08_6123, \9421 );
and \U$18631 ( \27745 , RIe20da38_4445, \9423 );
and \U$18632 ( \27746 , RIe20ad38_4413, \9425 );
and \U$18633 ( \27747 , RIe208038_4381, \9427 );
and \U$18634 ( \27748 , RIfc66ba8_6191, \9429 );
and \U$18635 ( \27749 , RIfccbcd8_7341, \9431 );
and \U$18636 ( \27750 , RIe202bd8_4321, \9433 );
and \U$18637 ( \27751 , RIe200fb8_4301, \9435 );
and \U$18638 ( \27752 , RIfcadbe8_6999, \9437 );
and \U$18639 ( \27753 , RIfccbe40_7342, \9439 );
and \U$18640 ( \27754 , RIfca7540_6926, \9441 );
and \U$18641 ( \27755 , RIfc6a3e8_6231, \9443 );
and \U$18642 ( \27756 , RIfca6898_6917, \9445 );
and \U$18643 ( \27757 , RIfc73358_6333, \9447 );
and \U$18644 ( \27758 , RIe1fd070_4256, \9449 );
and \U$18645 ( \27759 , RIe1fbe28_4243, \9451 );
and \U$18646 ( \27760 , RIfcc2660_7234, \9453 );
and \U$18647 ( \27761 , RIfc44468_5799, \9455 );
and \U$18648 ( \27762 , RIf15a940_5490, \9457 );
and \U$18649 ( \27763 , RIfca7270_6924, \9459 );
or \U$18650 ( \27764 , \27700 , \27701 , \27702 , \27703 , \27704 , \27705 , \27706 , \27707 , \27708 , \27709 , \27710 , \27711 , \27712 , \27713 , \27714 , \27715 , \27716 , \27717 , \27718 , \27719 , \27720 , \27721 , \27722 , \27723 , \27724 , \27725 , \27726 , \27727 , \27728 , \27729 , \27730 , \27731 , \27732 , \27733 , \27734 , \27735 , \27736 , \27737 , \27738 , \27739 , \27740 , \27741 , \27742 , \27743 , \27744 , \27745 , \27746 , \27747 , \27748 , \27749 , \27750 , \27751 , \27752 , \27753 , \27754 , \27755 , \27756 , \27757 , \27758 , \27759 , \27760 , \27761 , \27762 , \27763 );
and \U$18651 ( \27765 , RIfc5e070_6092, \9462 );
and \U$18652 ( \27766 , RIfc5dda0_6090, \9464 );
and \U$18653 ( \27767 , RIfc7e050_6456, \9466 );
and \U$18654 ( \27768 , RIe1fa7a8_4227, \9468 );
and \U$18655 ( \27769 , RIfc5d968_6087, \9470 );
and \U$18656 ( \27770 , RIfcd9568_7495, \9472 );
and \U$18657 ( \27771 , RIfc8d668_6631, \9474 );
and \U$18658 ( \27772 , RIe1f5d20_4174, \9476 );
and \U$18659 ( \27773 , RIfca4138_6889, \9478 );
and \U$18660 ( \27774 , RIfc8cdf8_6625, \9480 );
and \U$18661 ( \27775 , RIfcc7c28_7295, \9482 );
and \U$18662 ( \27776 , RIe1f39f8_4149, \9484 );
and \U$18663 ( \27777 , RIfc99440_6766, \9486 );
and \U$18664 ( \27778 , RIfcbc3f0_7164, \9488 );
and \U$18665 ( \27779 , RIfc5a128_6047, \9490 );
and \U$18666 ( \27780 , RIe1ee700_4090, \9492 );
and \U$18667 ( \27781 , RIe1ebfa0_4062, \9494 );
and \U$18668 ( \27782 , RIe1e92a0_4030, \9496 );
and \U$18669 ( \27783 , RIe1e65a0_3998, \9498 );
and \U$18670 ( \27784 , RIe1e38a0_3966, \9500 );
and \U$18671 ( \27785 , RIe1e0ba0_3934, \9502 );
and \U$18672 ( \27786 , RIe1ddea0_3902, \9504 );
and \U$18673 ( \27787 , RIe1db1a0_3870, \9506 );
and \U$18674 ( \27788 , RIe1d84a0_3838, \9508 );
and \U$18675 ( \27789 , RIe1d2aa0_3774, \9510 );
and \U$18676 ( \27790 , RIe1cfda0_3742, \9512 );
and \U$18677 ( \27791 , RIe1cd0a0_3710, \9514 );
and \U$18678 ( \27792 , RIe1ca3a0_3678, \9516 );
and \U$18679 ( \27793 , RIe1c76a0_3646, \9518 );
and \U$18680 ( \27794 , RIe1c49a0_3614, \9520 );
and \U$18681 ( \27795 , RIe1c1ca0_3582, \9522 );
and \U$18682 ( \27796 , RIe1befa0_3550, \9524 );
and \U$18683 ( \27797 , RIf14cde0_5334, \9526 );
and \U$18684 ( \27798 , RIf14bb98_5321, \9528 );
and \U$18685 ( \27799 , RIe1b99d8_3489, \9530 );
and \U$18686 ( \27800 , RIe1b7980_3466, \9532 );
and \U$18687 ( \27801 , RIfc4c460_5890, \9534 );
and \U$18688 ( \27802 , RIfc9e738_6825, \9536 );
and \U$18689 ( \27803 , RIe1b5658_3441, \9538 );
and \U$18690 ( \27804 , RIfec54d8_8365, \9540 );
and \U$18691 ( \27805 , RIf149168_5291, \9542 );
and \U$18692 ( \27806 , RIf147f20_5278, \9544 );
and \U$18693 ( \27807 , RIe1b2ac0_3410, \9546 );
and \U$18694 ( \27808 , RIe1b1170_3392, \9548 );
and \U$18695 ( \27809 , RIf1473e0_5270, \9550 );
and \U$18696 ( \27810 , RIf1468a0_5262, \9552 );
and \U$18697 ( \27811 , RIe1acb20_3342, \9554 );
and \U$18698 ( \27812 , RIe1ab338_3325, \9556 );
and \U$18699 ( \27813 , RIe1a92e0_3302, \9558 );
and \U$18700 ( \27814 , RIe1a65e0_3270, \9560 );
and \U$18701 ( \27815 , RIe1a38e0_3238, \9562 );
and \U$18702 ( \27816 , RIe1a0be0_3206, \9564 );
and \U$18703 ( \27817 , RIe18d0e0_2982, \9566 );
and \U$18704 ( \27818 , RIe1795e0_2758, \9568 );
and \U$18705 ( \27819 , RIe226f38_4733, \9570 );
and \U$18706 ( \27820 , RIe21bb38_4605, \9572 );
and \U$18707 ( \27821 , RIe205338_4349, \9574 );
and \U$18708 ( \27822 , RIe1ff398_4281, \9576 );
and \U$18709 ( \27823 , RIe1f8750_4204, \9578 );
and \U$18710 ( \27824 , RIe1f1298_4121, \9580 );
and \U$18711 ( \27825 , RIe1d57a0_3806, \9582 );
and \U$18712 ( \27826 , RIe1bc2a0_3518, \9584 );
and \U$18713 ( \27827 , RIe1af118_3369, \9586 );
and \U$18714 ( \27828 , RIe171750_2668, \9588 );
or \U$18715 ( \27829 , \27765 , \27766 , \27767 , \27768 , \27769 , \27770 , \27771 , \27772 , \27773 , \27774 , \27775 , \27776 , \27777 , \27778 , \27779 , \27780 , \27781 , \27782 , \27783 , \27784 , \27785 , \27786 , \27787 , \27788 , \27789 , \27790 , \27791 , \27792 , \27793 , \27794 , \27795 , \27796 , \27797 , \27798 , \27799 , \27800 , \27801 , \27802 , \27803 , \27804 , \27805 , \27806 , \27807 , \27808 , \27809 , \27810 , \27811 , \27812 , \27813 , \27814 , \27815 , \27816 , \27817 , \27818 , \27819 , \27820 , \27821 , \27822 , \27823 , \27824 , \27825 , \27826 , \27827 , \27828 );
or \U$18716 ( \27830 , \27764 , \27829 );
_DC g3576 ( \27831_nG3576 , \27830 , \9597 );
buf \U$18717 ( \27832 , \27831_nG3576 );
xor \U$18718 ( \27833 , \27699 , \27832 );
and \U$18719 ( \27834 , RIdec5ae0_713, \9059 );
and \U$18720 ( \27835 , RIdec2de0_681, \9061 );
and \U$18721 ( \27836 , RIfc82268_6503, \9063 );
and \U$18722 ( \27837 , RIdec00e0_649, \9065 );
and \U$18723 ( \27838 , RIfcb8d18_7125, \9067 );
and \U$18724 ( \27839 , RIdebd3e0_617, \9069 );
and \U$18725 ( \27840 , RIdeba6e0_585, \9071 );
and \U$18726 ( \27841 , RIdeb79e0_553, \9073 );
and \U$18727 ( \27842 , RIfcb9858_7133, \9075 );
and \U$18728 ( \27843 , RIdeb1fe0_489, \9077 );
and \U$18729 ( \27844 , RIfc9efa8_6831, \9079 );
and \U$18730 ( \27845 , RIdeaf2e0_457, \9081 );
and \U$18731 ( \27846 , RIfce0750_7576, \9083 );
and \U$18732 ( \27847 , RIdeab488_425, \9085 );
and \U$18733 ( \27848 , RIdea4b88_393, \9087 );
and \U$18734 ( \27849 , RIde9e288_361, \9089 );
and \U$18735 ( \27850 , RIee1d0b0_4789, \9091 );
and \U$18736 ( \27851 , RIee1c138_4778, \9093 );
and \U$18737 ( \27852 , RIfcd0e68_7399, \9095 );
and \U$18738 ( \27853 , RIfc76d00_6374, \9097 );
and \U$18739 ( \27854 , RIfe89028_7903, \9099 );
and \U$18740 ( \27855 , RIfe88d58_7901, \9101 );
and \U$18741 ( \27856 , RIfe88ec0_7902, \9103 );
and \U$18742 ( \27857 , RIfe88bf0_7900, \9105 );
and \U$18743 ( \27858 , RIfcda7b0_7508, \9107 );
and \U$18744 ( \27859 , RIfc4d810_5904, \9109 );
and \U$18745 ( \27860 , RIfc52dd8_5965, \9111 );
and \U$18746 ( \27861 , RIfcde590_7552, \9113 );
and \U$18747 ( \27862 , RIfc4f868_5927, \9115 );
and \U$18748 ( \27863 , RIe16bd50_2604, \9117 );
and \U$18749 ( \27864 , RIfc68930_6212, \9119 );
and \U$18750 ( \27865 , RIe1683a8_2563, \9121 );
and \U$18751 ( \27866 , RIe165ae0_2534, \9123 );
and \U$18752 ( \27867 , RIe162de0_2502, \9125 );
and \U$18753 ( \27868 , RIfe88a88_7899, \9127 );
and \U$18754 ( \27869 , RIe1600e0_2470, \9129 );
and \U$18755 ( \27870 , RIfcc9140_7310, \9131 );
and \U$18756 ( \27871 , RIe15d3e0_2438, \9133 );
and \U$18757 ( \27872 , RIe1579e0_2374, \9135 );
and \U$18758 ( \27873 , RIe154ce0_2342, \9137 );
and \U$18759 ( \27874 , RIfc698a8_6223, \9139 );
and \U$18760 ( \27875 , RIe151fe0_2310, \9141 );
and \U$18761 ( \27876 , RIee35098_5062, \9143 );
and \U$18762 ( \27877 , RIe14f2e0_2278, \9145 );
and \U$18763 ( \27878 , RIfcc0338_7209, \9147 );
and \U$18764 ( \27879 , RIe14c5e0_2246, \9149 );
and \U$18765 ( \27880 , RIe1498e0_2214, \9151 );
and \U$18766 ( \27881 , RIe146be0_2182, \9153 );
and \U$18767 ( \27882 , RIfc88208_6571, \9155 );
and \U$18768 ( \27883 , RIfc85670_6540, \9157 );
and \U$18769 ( \27884 , RIfc81f98_6501, \9159 );
and \U$18770 ( \27885 , RIfcc4f28_7263, \9161 );
and \U$18771 ( \27886 , RIe1414b0_2120, \9163 );
and \U$18772 ( \27887 , RIe13f188_2095, \9165 );
and \U$18773 ( \27888 , RIdf3d090_2071, \9167 );
and \U$18774 ( \27889 , RIdf3aa98_2044, \9169 );
and \U$18775 ( \27890 , RIfcd2920_7418, \9171 );
and \U$18776 ( \27891 , RIfc7d7e0_6450, \9173 );
and \U$18777 ( \27892 , RIfc49760_5858, \9175 );
and \U$18778 ( \27893 , RIfce5a48_7635, \9177 );
and \U$18779 ( \27894 , RIdf35ea8_1990, \9179 );
and \U$18780 ( \27895 , RIdf338b0_1963, \9181 );
and \U$18781 ( \27896 , RIfe88920_7898, \9183 );
and \U$18782 ( \27897 , RIdf2f800_1917, \9185 );
or \U$18783 ( \27898 , \27834 , \27835 , \27836 , \27837 , \27838 , \27839 , \27840 , \27841 , \27842 , \27843 , \27844 , \27845 , \27846 , \27847 , \27848 , \27849 , \27850 , \27851 , \27852 , \27853 , \27854 , \27855 , \27856 , \27857 , \27858 , \27859 , \27860 , \27861 , \27862 , \27863 , \27864 , \27865 , \27866 , \27867 , \27868 , \27869 , \27870 , \27871 , \27872 , \27873 , \27874 , \27875 , \27876 , \27877 , \27878 , \27879 , \27880 , \27881 , \27882 , \27883 , \27884 , \27885 , \27886 , \27887 , \27888 , \27889 , \27890 , \27891 , \27892 , \27893 , \27894 , \27895 , \27896 , \27897 );
and \U$18784 ( \27899 , RIee2bfc0_4959, \9188 );
and \U$18785 ( \27900 , RIee2a670_4941, \9190 );
and \U$18786 ( \27901 , RIee29158_4926, \9192 );
and \U$18787 ( \27902 , RIee27f10_4913, \9194 );
and \U$18788 ( \27903 , RIdf2a7d8_1860, \9196 );
and \U$18789 ( \27904 , RIdf28618_1836, \9198 );
and \U$18790 ( \27905 , RIdf26890_1815, \9200 );
and \U$18791 ( \27906 , RIdf24dd8_1796, \9202 );
and \U$18792 ( \27907 , RIfcad918_6997, \9204 );
and \U$18793 ( \27908 , RIfc69fb0_6228, \9206 );
and \U$18794 ( \27909 , RIfc63368_6151, \9208 );
and \U$18795 ( \27910 , RIfc623f0_6140, \9210 );
and \U$18796 ( \27911 , RIfc60938_6121, \9212 );
and \U$18797 ( \27912 , RIdf1ff18_1740, \9214 );
and \U$18798 ( \27913 , RIfcba500_7142, \9216 );
and \U$18799 ( \27914 , RIdf19870_1667, \9218 );
and \U$18800 ( \27915 , RIdf176b0_1643, \9220 );
and \U$18801 ( \27916 , RIdf149b0_1611, \9222 );
and \U$18802 ( \27917 , RIdf11cb0_1579, \9224 );
and \U$18803 ( \27918 , RIdf0efb0_1547, \9226 );
and \U$18804 ( \27919 , RIdf0c2b0_1515, \9228 );
and \U$18805 ( \27920 , RIdf095b0_1483, \9230 );
and \U$18806 ( \27921 , RIdf068b0_1451, \9232 );
and \U$18807 ( \27922 , RIdf03bb0_1419, \9234 );
and \U$18808 ( \27923 , RIdefe1b0_1355, \9236 );
and \U$18809 ( \27924 , RIdefb4b0_1323, \9238 );
and \U$18810 ( \27925 , RIdef87b0_1291, \9240 );
and \U$18811 ( \27926 , RIdef5ab0_1259, \9242 );
and \U$18812 ( \27927 , RIdef2db0_1227, \9244 );
and \U$18813 ( \27928 , RIdef00b0_1195, \9246 );
and \U$18814 ( \27929 , RIdeed3b0_1163, \9248 );
and \U$18815 ( \27930 , RIdeea6b0_1131, \9250 );
and \U$18816 ( \27931 , RIfcc9848_7315, \9252 );
and \U$18817 ( \27932 , RIfc69a10_6224, \9254 );
and \U$18818 ( \27933 , RIfcacc70_6988, \9256 );
and \U$18819 ( \27934 , RIfccbfa8_7343, \9258 );
and \U$18820 ( \27935 , RIdee4f80_1069, \9260 );
and \U$18821 ( \27936 , RIdee31f8_1048, \9262 );
and \U$18822 ( \27937 , RIdee1038_1024, \9264 );
and \U$18823 ( \27938 , RIdedee78_1000, \9266 );
and \U$18824 ( \27939 , RIfc84590_6528, \9268 );
and \U$18825 ( \27940 , RIfc9bba0_6794, \9270 );
and \U$18826 ( \27941 , RIee21b38_4842, \9272 );
and \U$18827 ( \27942 , RIfc47168_5831, \9274 );
and \U$18828 ( \27943 , RIded9e50_943, \9276 );
and \U$18829 ( \27944 , RIded7858_916, \9278 );
and \U$18830 ( \27945 , RIfe887b8_7897, \9280 );
and \U$18831 ( \27946 , RIded34d8_868, \9282 );
and \U$18832 ( \27947 , RIded0ee0_841, \9284 );
and \U$18833 ( \27948 , RIdece1e0_809, \9286 );
and \U$18834 ( \27949 , RIdecb4e0_777, \9288 );
and \U$18835 ( \27950 , RIdec87e0_745, \9290 );
and \U$18836 ( \27951 , RIdeb4ce0_521, \9292 );
and \U$18837 ( \27952 , RIde97988_329, \9294 );
and \U$18838 ( \27953 , RIe16e8e8_2635, \9296 );
and \U$18839 ( \27954 , RIe15a6e0_2406, \9298 );
and \U$18840 ( \27955 , RIe143ee0_2150, \9300 );
and \U$18841 ( \27956 , RIdf388d8_2020, \9302 );
and \U$18842 ( \27957 , RIdf2cf38_1888, \9304 );
and \U$18843 ( \27958 , RIdf1d7b8_1712, \9306 );
and \U$18844 ( \27959 , RIdf00eb0_1387, \9308 );
and \U$18845 ( \27960 , RIdee79b0_1099, \9310 );
and \U$18846 ( \27961 , RIdedc718_972, \9312 );
and \U$18847 ( \27962 , RIde7d8d0_202, \9314 );
or \U$18848 ( \27963 , \27899 , \27900 , \27901 , \27902 , \27903 , \27904 , \27905 , \27906 , \27907 , \27908 , \27909 , \27910 , \27911 , \27912 , \27913 , \27914 , \27915 , \27916 , \27917 , \27918 , \27919 , \27920 , \27921 , \27922 , \27923 , \27924 , \27925 , \27926 , \27927 , \27928 , \27929 , \27930 , \27931 , \27932 , \27933 , \27934 , \27935 , \27936 , \27937 , \27938 , \27939 , \27940 , \27941 , \27942 , \27943 , \27944 , \27945 , \27946 , \27947 , \27948 , \27949 , \27950 , \27951 , \27952 , \27953 , \27954 , \27955 , \27956 , \27957 , \27958 , \27959 , \27960 , \27961 , \27962 );
or \U$18849 ( \27964 , \27898 , \27963 );
_DC g24ce ( \27965_nG24ce , \27964 , \9323 );
buf \U$18850 ( \27966 , \27965_nG24ce );
and \U$18851 ( \27967 , RIe19dd78_3173, \9333 );
and \U$18852 ( \27968 , RIe19b078_3141, \9335 );
and \U$18853 ( \27969 , RIfca1438_6857, \9337 );
and \U$18854 ( \27970 , RIe198378_3109, \9339 );
and \U$18855 ( \27971 , RIfca35f8_6881, \9341 );
and \U$18856 ( \27972 , RIe195678_3077, \9343 );
and \U$18857 ( \27973 , RIe192978_3045, \9345 );
and \U$18858 ( \27974 , RIe18fc78_3013, \9347 );
and \U$18859 ( \27975 , RIe18a278_2949, \9349 );
and \U$18860 ( \27976 , RIe187578_2917, \9351 );
and \U$18861 ( \27977 , RIfcba230_7140, \9353 );
and \U$18862 ( \27978 , RIe184878_2885, \9355 );
and \U$18863 ( \27979 , RIf142d90_5220, \9357 );
and \U$18864 ( \27980 , RIe181b78_2853, \9359 );
and \U$18865 ( \27981 , RIe17ee78_2821, \9361 );
and \U$18866 ( \27982 , RIe17c178_2789, \9363 );
and \U$18867 ( \27983 , RIfc9be70_6796, \9365 );
and \U$18868 ( \27984 , RIfc9bd08_6795, \9367 );
and \U$18869 ( \27985 , RIfc4ccd0_5896, \9369 );
and \U$18870 ( \27986 , RIe176070_2720, \9371 );
and \U$18871 ( \27987 , RIfc87c68_6567, \9373 );
and \U$18872 ( \27988 , RIfc87b00_6566, \9375 );
and \U$18873 ( \27989 , RIfcc4c58_7261, \9377 );
and \U$18874 ( \27990 , RIfc4fca0_5930, \9379 );
and \U$18875 ( \27991 , RIfc4f598_5925, \9381 );
and \U$18876 ( \27992 , RIfc876c8_6563, \9383 );
and \U$18877 ( \27993 , RIfc4dae0_5906, \9385 );
and \U$18878 ( \27994 , RIe173eb0_2696, \9387 );
and \U$18879 ( \27995 , RIfcb9420_7130, \9389 );
and \U$18880 ( \27996 , RIfc4e080_5910, \9391 );
and \U$18881 ( \27997 , RIfc4e350_5912, \9393 );
and \U$18882 ( \27998 , RIfc9d388_6811, \9395 );
and \U$18883 ( \27999 , RIfc40a48_5761, \9397 );
and \U$18884 ( \28000 , RIe2240d0_4700, \9399 );
and \U$18885 ( \28001 , RIfc85508_6539, \9401 );
and \U$18886 ( \28002 , RIe2213d0_4668, \9403 );
and \U$18887 ( \28003 , RIfc9ba38_6793, \9405 );
and \U$18888 ( \28004 , RIe21e6d0_4636, \9407 );
and \U$18889 ( \28005 , RIe218cd0_4572, \9409 );
and \U$18890 ( \28006 , RIe215fd0_4540, \9411 );
and \U$18891 ( \28007 , RIfc52c70_5964, \9413 );
and \U$18892 ( \28008 , RIe2132d0_4508, \9415 );
and \U$18893 ( \28009 , RIfca3760_6882, \9417 );
and \U$18894 ( \28010 , RIe2105d0_4476, \9419 );
and \U$18895 ( \28011 , RIfc97988_6747, \9421 );
and \U$18896 ( \28012 , RIe20d8d0_4444, \9423 );
and \U$18897 ( \28013 , RIe20abd0_4412, \9425 );
and \U$18898 ( \28014 , RIe207ed0_4380, \9427 );
and \U$18899 ( \28015 , RIfceb5b0_7700, \9429 );
and \U$18900 ( \28016 , RIfcddbb8_7545, \9431 );
and \U$18901 ( \28017 , RIe202a70_4320, \9433 );
and \U$18902 ( \28018 , RIe200e50_4300, \9435 );
and \U$18903 ( \28019 , RIfc73d30_6340, \9437 );
and \U$18904 ( \28020 , RIfcaf100_7014, \9439 );
and \U$18905 ( \28021 , RIfc71468_6311, \9441 );
and \U$18906 ( \28022 , RIfcdcad8_7533, \9443 );
and \U$18907 ( \28023 , RIfcdda50_7544, \9445 );
and \U$18908 ( \28024 , RIfca8620_6938, \9447 );
and \U$18909 ( \28025 , RIe1fcf08_4255, \9449 );
and \U$18910 ( \28026 , RIe1fbcc0_4242, \9451 );
and \U$18911 ( \28027 , RIfc6c008_6251, \9453 );
and \U$18912 ( \28028 , RIfcdd1e0_7538, \9455 );
and \U$18913 ( \28029 , RIfca9700_6950, \9457 );
and \U$18914 ( \28030 , RIfca92c8_6947, \9459 );
or \U$18915 ( \28031 , \27967 , \27968 , \27969 , \27970 , \27971 , \27972 , \27973 , \27974 , \27975 , \27976 , \27977 , \27978 , \27979 , \27980 , \27981 , \27982 , \27983 , \27984 , \27985 , \27986 , \27987 , \27988 , \27989 , \27990 , \27991 , \27992 , \27993 , \27994 , \27995 , \27996 , \27997 , \27998 , \27999 , \28000 , \28001 , \28002 , \28003 , \28004 , \28005 , \28006 , \28007 , \28008 , \28009 , \28010 , \28011 , \28012 , \28013 , \28014 , \28015 , \28016 , \28017 , \28018 , \28019 , \28020 , \28021 , \28022 , \28023 , \28024 , \28025 , \28026 , \28027 , \28028 , \28029 , \28030 );
and \U$18916 ( \28032 , RIfcce5a0_7370, \9462 );
and \U$18917 ( \28033 , RIfc6ba68_6247, \9464 );
and \U$18918 ( \28034 , RIfc6f410_6288, \9466 );
and \U$18919 ( \28035 , RIe1fa640_4226, \9468 );
and \U$18920 ( \28036 , RIfcce000_7366, \9470 );
and \U$18921 ( \28037 , RIfc53918_5973, \9472 );
and \U$18922 ( \28038 , RIfcce708_7371, \9474 );
and \U$18923 ( \28039 , RIe1f5bb8_4173, \9476 );
and \U$18924 ( \28040 , RIf1535f0_5408, \9478 );
and \U$18925 ( \28041 , RIf151e08_5391, \9480 );
and \U$18926 ( \28042 , RIfc72db8_6329, \9482 );
and \U$18927 ( \28043 , RIe1f3890_4148, \9484 );
and \U$18928 ( \28044 , RIf14fc48_5367, \9486 );
and \U$18929 ( \28045 , RIfc72c50_6328, \9488 );
and \U$18930 ( \28046 , RIfc73e98_6341, \9490 );
and \U$18931 ( \28047 , RIe1ee598_4089, \9492 );
and \U$18932 ( \28048 , RIe1ebe38_4061, \9494 );
and \U$18933 ( \28049 , RIe1e9138_4029, \9496 );
and \U$18934 ( \28050 , RIe1e6438_3997, \9498 );
and \U$18935 ( \28051 , RIe1e3738_3965, \9500 );
and \U$18936 ( \28052 , RIe1e0a38_3933, \9502 );
and \U$18937 ( \28053 , RIe1ddd38_3901, \9504 );
and \U$18938 ( \28054 , RIe1db038_3869, \9506 );
and \U$18939 ( \28055 , RIe1d8338_3837, \9508 );
and \U$18940 ( \28056 , RIe1d2938_3773, \9510 );
and \U$18941 ( \28057 , RIe1cfc38_3741, \9512 );
and \U$18942 ( \28058 , RIe1ccf38_3709, \9514 );
and \U$18943 ( \28059 , RIe1ca238_3677, \9516 );
and \U$18944 ( \28060 , RIe1c7538_3645, \9518 );
and \U$18945 ( \28061 , RIe1c4838_3613, \9520 );
and \U$18946 ( \28062 , RIe1c1b38_3581, \9522 );
and \U$18947 ( \28063 , RIe1bee38_3549, \9524 );
and \U$18948 ( \28064 , RIfcb8a48_7123, \9526 );
and \U$18949 ( \28065 , RIfcb84a8_7119, \9528 );
and \U$18950 ( \28066 , RIe1b9870_3488, \9530 );
and \U$18951 ( \28067 , RIe1b7818_3465, \9532 );
and \U$18952 ( \28068 , RIfc85940_6542, \9534 );
and \U$18953 ( \28069 , RIfc9e198_6821, \9536 );
and \U$18954 ( \28070 , RIfeac140_8274, \9538 );
and \U$18955 ( \28071 , RIe1b42a8_3427, \9540 );
and \U$18956 ( \28072 , RIfc518c0_5950, \9542 );
and \U$18957 ( \28073 , RIfc838e8_6519, \9544 );
and \U$18958 ( \28074 , RIfe884e8_7895, \9546 );
and \U$18959 ( \28075 , RIe1b1008_3391, \9548 );
and \U$18960 ( \28076 , RIfcc5900_7270, \9550 );
and \U$18961 ( \28077 , RIfc82ad8_6509, \9552 );
and \U$18962 ( \28078 , RIe1ac9b8_3341, \9554 );
and \U$18963 ( \28079 , RIfe88650_7896, \9556 );
and \U$18964 ( \28080 , RIe1a9178_3301, \9558 );
and \U$18965 ( \28081 , RIe1a6478_3269, \9560 );
and \U$18966 ( \28082 , RIe1a3778_3237, \9562 );
and \U$18967 ( \28083 , RIe1a0a78_3205, \9564 );
and \U$18968 ( \28084 , RIe18cf78_2981, \9566 );
and \U$18969 ( \28085 , RIe179478_2757, \9568 );
and \U$18970 ( \28086 , RIe226dd0_4732, \9570 );
and \U$18971 ( \28087 , RIe21b9d0_4604, \9572 );
and \U$18972 ( \28088 , RIe2051d0_4348, \9574 );
and \U$18973 ( \28089 , RIe1ff230_4280, \9576 );
and \U$18974 ( \28090 , RIe1f85e8_4203, \9578 );
and \U$18975 ( \28091 , RIe1f1130_4120, \9580 );
and \U$18976 ( \28092 , RIe1d5638_3805, \9582 );
and \U$18977 ( \28093 , RIe1bc138_3517, \9584 );
and \U$18978 ( \28094 , RIe1aefb0_3368, \9586 );
and \U$18979 ( \28095 , RIe1715e8_2667, \9588 );
or \U$18980 ( \28096 , \28032 , \28033 , \28034 , \28035 , \28036 , \28037 , \28038 , \28039 , \28040 , \28041 , \28042 , \28043 , \28044 , \28045 , \28046 , \28047 , \28048 , \28049 , \28050 , \28051 , \28052 , \28053 , \28054 , \28055 , \28056 , \28057 , \28058 , \28059 , \28060 , \28061 , \28062 , \28063 , \28064 , \28065 , \28066 , \28067 , \28068 , \28069 , \28070 , \28071 , \28072 , \28073 , \28074 , \28075 , \28076 , \28077 , \28078 , \28079 , \28080 , \28081 , \28082 , \28083 , \28084 , \28085 , \28086 , \28087 , \28088 , \28089 , \28090 , \28091 , \28092 , \28093 , \28094 , \28095 );
or \U$18981 ( \28097 , \28031 , \28096 );
_DC g35fb ( \28098_nG35fb , \28097 , \9597 );
buf \U$18982 ( \28099 , \28098_nG35fb );
and \U$18983 ( \28100 , \27966 , \28099 );
and \U$18984 ( \28101 , \26012 , \26145 );
and \U$18985 ( \28102 , \26145 , \26420 );
and \U$18986 ( \28103 , \26012 , \26420 );
or \U$18987 ( \28104 , \28101 , \28102 , \28103 );
and \U$18988 ( \28105 , \28099 , \28104 );
and \U$18989 ( \28106 , \27966 , \28104 );
or \U$18990 ( \28107 , \28100 , \28105 , \28106 );
xor \U$18991 ( \28108 , \27833 , \28107 );
buf g4406 ( \28109_nG4406 , \28108 );
xor \U$18992 ( \28110 , \27966 , \28099 );
xor \U$18993 ( \28111 , \28110 , \28104 );
buf g4409 ( \28112_nG4409 , \28111 );
nand \U$18994 ( \28113 , \28112_nG4409 , \26422_nG440c );
and \U$18995 ( \28114 , \28109_nG4406 , \28113 );
xor \U$18996 ( \28115 , \28112_nG4409 , \26422_nG440c );
not \U$18997 ( \28116 , \28115 );
xor \U$18998 ( \28117 , \28109_nG4406 , \28112_nG4409 );
and \U$18999 ( \28118 , \28116 , \28117 );
and \U$19001 ( \28119 , \28115 , \10694_nG9c0e );
or \U$19002 ( \28120 , 1'b0 , \28119 );
xor \U$19003 ( \28121 , \28114 , \28120 );
xor \U$19004 ( \28122 , \28114 , \28121 );
buf \U$19005 ( \28123 , \28122 );
buf \U$19006 ( \28124 , \28123 );
xor \U$19007 ( \28125 , \27566 , \28124 );
and \U$19008 ( \28126 , \27521 , \27526 );
and \U$19009 ( \28127 , \27521 , \27559 );
and \U$19010 ( \28128 , \27526 , \27559 );
or \U$19011 ( \28129 , \28126 , \28127 , \28128 );
and \U$19012 ( \28130 , \28125 , \28129 );
and \U$19013 ( \28131 , \27532 , \27551 );
and \U$19014 ( \28132 , \27532 , \27557 );
and \U$19015 ( \28133 , \27551 , \27557 );
or \U$19016 ( \28134 , \28131 , \28132 , \28133 );
buf \U$19017 ( \28135 , \28134 );
and \U$19018 ( \28136 , \27496 , \27501 );
and \U$19019 ( \28137 , \27496 , \27508 );
and \U$19020 ( \28138 , \27501 , \27508 );
or \U$19021 ( \28139 , \28136 , \28137 , \28138 );
buf \U$19022 ( \28140 , \28139 );
and \U$19023 ( \28141 , \13370 , \22629_nG9bd5 );
and \U$19024 ( \28142 , \13367 , \23696_nG9bd2 );
or \U$19025 ( \28143 , \28141 , \28142 );
xor \U$19026 ( \28144 , \13366 , \28143 );
buf \U$19027 ( \28145 , \28144 );
buf \U$19029 ( \28146 , \28145 );
xor \U$19030 ( \28147 , \28140 , \28146 );
and \U$19031 ( \28148 , \12157 , \24226_nG9bcf );
and \U$19032 ( \28149 , \12154 , \25298_nG9bcc );
or \U$19033 ( \28150 , \28148 , \28149 );
xor \U$19034 ( \28151 , \12153 , \28150 );
buf \U$19035 ( \28152 , \28151 );
buf \U$19037 ( \28153 , \28152 );
xor \U$19038 ( \28154 , \28147 , \28153 );
buf \U$19039 ( \28155 , \28154 );
and \U$19040 ( \28156 , \27432 , \27438 );
buf \U$19041 ( \28157 , \28156 );
and \U$19042 ( \28158 , \23201 , \12801_nG9bff );
and \U$19043 ( \28159 , \23198 , \13705_nG9bfc );
or \U$19044 ( \28160 , \28158 , \28159 );
xor \U$19045 ( \28161 , \23197 , \28160 );
buf \U$19046 ( \28162 , \28161 );
buf \U$19048 ( \28163 , \28162 );
xor \U$19049 ( \28164 , \28157 , \28163 );
and \U$19050 ( \28165 , \21658 , \14070_nG9bf9 );
and \U$19051 ( \28166 , \21655 , \14984_nG9bf6 );
or \U$19052 ( \28167 , \28165 , \28166 );
xor \U$19053 ( \28168 , \21654 , \28167 );
buf \U$19054 ( \28169 , \28168 );
buf \U$19056 ( \28170 , \28169 );
xor \U$19057 ( \28171 , \28164 , \28170 );
buf \U$19058 ( \28172 , \28171 );
and \U$19059 ( \28173 , \18702 , \16680_nG9bed );
and \U$19060 ( \28174 , \18699 , \17665_nG9bea );
or \U$19061 ( \28175 , \28173 , \28174 );
xor \U$19062 ( \28176 , \18698 , \28175 );
buf \U$19063 ( \28177 , \28176 );
buf \U$19065 ( \28178 , \28177 );
xor \U$19066 ( \28179 , \28172 , \28178 );
and \U$19067 ( \28180 , \17297 , \18107_nG9be7 );
and \U$19068 ( \28181 , \17294 , \19091_nG9be4 );
or \U$19069 ( \28182 , \28180 , \28181 );
xor \U$19070 ( \28183 , \17293 , \28182 );
buf \U$19071 ( \28184 , \28183 );
buf \U$19073 ( \28185 , \28184 );
xor \U$19074 ( \28186 , \28179 , \28185 );
buf \U$19075 ( \28187 , \28186 );
and \U$19076 ( \28188 , \27429 , \27455 );
and \U$19077 ( \28189 , \27429 , \27462 );
and \U$19078 ( \28190 , \27455 , \27462 );
or \U$19079 ( \28191 , \28188 , \28189 , \28190 );
buf \U$19080 ( \28192 , \28191 );
xor \U$19081 ( \28193 , \28187 , \28192 );
and \U$19082 ( \28194 , \15940 , \19586_nG9be1 );
and \U$19083 ( \28195 , \15937 , \20608_nG9bde );
or \U$19084 ( \28196 , \28194 , \28195 );
xor \U$19085 ( \28197 , \15936 , \28196 );
buf \U$19086 ( \28198 , \28197 );
buf \U$19088 ( \28199 , \28198 );
xor \U$19089 ( \28200 , \28193 , \28199 );
buf \U$19090 ( \28201 , \28200 );
xor \U$19091 ( \28202 , \28155 , \28201 );
and \U$19092 ( \28203 , \10707 , \27416_nG9bc3 );
and \U$19093 ( \28204 , \27362 , \27366 );
and \U$19094 ( \28205 , \27366 , \27404 );
and \U$19095 ( \28206 , \27362 , \27404 );
or \U$19096 ( \28207 , \28204 , \28205 , \28206 );
and \U$19097 ( \28208 , \27371 , \27375 );
and \U$19098 ( \28209 , \27375 , \27403 );
and \U$19099 ( \28210 , \27371 , \27403 );
or \U$19100 ( \28211 , \28208 , \28209 , \28210 );
and \U$19101 ( \28212 , \27021 , \27307 );
and \U$19102 ( \28213 , \27307 , \27356 );
and \U$19103 ( \28214 , \27021 , \27356 );
or \U$19104 ( \28215 , \28212 , \28213 , \28214 );
xor \U$19105 ( \28216 , \28211 , \28215 );
and \U$19106 ( \28217 , \27297 , \27301 );
and \U$19107 ( \28218 , \27301 , \27306 );
and \U$19108 ( \28219 , \27297 , \27306 );
or \U$19109 ( \28220 , \28217 , \28218 , \28219 );
and \U$19110 ( \28221 , \27380 , \27384 );
and \U$19111 ( \28222 , \27384 , \27402 );
and \U$19112 ( \28223 , \27380 , \27402 );
or \U$19113 ( \28224 , \28221 , \28222 , \28223 );
xor \U$19114 ( \28225 , \28220 , \28224 );
and \U$19115 ( \28226 , \27326 , \27340 );
and \U$19116 ( \28227 , \27340 , \27355 );
and \U$19117 ( \28228 , \27326 , \27355 );
or \U$19118 ( \28229 , \28226 , \28227 , \28228 );
xor \U$19119 ( \28230 , \28225 , \28229 );
xor \U$19120 ( \28231 , \28216 , \28230 );
xor \U$19121 ( \28232 , \28207 , \28231 );
and \U$19122 ( \28233 , \27316 , \27320 );
and \U$19123 ( \28234 , \27320 , \27325 );
and \U$19124 ( \28235 , \27316 , \27325 );
or \U$19125 ( \28236 , \28233 , \28234 , \28235 );
and \U$19126 ( \28237 , \27330 , \27334 );
and \U$19127 ( \28238 , \27334 , \27339 );
and \U$19128 ( \28239 , \27330 , \27339 );
or \U$19129 ( \28240 , \28237 , \28238 , \28239 );
xor \U$19130 ( \28241 , \28236 , \28240 );
and \U$19131 ( \28242 , \27345 , \27349 );
and \U$19132 ( \28243 , \27349 , \27354 );
and \U$19133 ( \28244 , \27345 , \27354 );
or \U$19134 ( \28245 , \28242 , \28243 , \28244 );
xor \U$19135 ( \28246 , \28241 , \28245 );
and \U$19136 ( \28247 , \27389 , \27393 );
and \U$19137 ( \28248 , \27393 , \27401 );
and \U$19138 ( \28249 , \27389 , \27401 );
or \U$19139 ( \28250 , \28247 , \28248 , \28249 );
and \U$19140 ( \28251 , \25815 , \11574 );
and \U$19141 ( \28252 , \26829 , \11278 );
nor \U$19142 ( \28253 , \28251 , \28252 );
xnor \U$19143 ( \28254 , \28253 , \11580 );
and \U$19144 ( \28255 , \22556 , \14054 );
and \U$19145 ( \28256 , \23617 , \13692 );
nor \U$19146 ( \28257 , \28255 , \28256 );
xnor \U$19147 ( \28258 , \28257 , \14035 );
xor \U$19148 ( \28259 , \28254 , \28258 );
and \U$19149 ( \28260 , RIdec5ae0_713, \9333 );
and \U$19150 ( \28261 , RIdec2de0_681, \9335 );
and \U$19151 ( \28262 , RIfc82268_6503, \9337 );
and \U$19152 ( \28263 , RIdec00e0_649, \9339 );
and \U$19153 ( \28264 , RIfcb8d18_7125, \9341 );
and \U$19154 ( \28265 , RIdebd3e0_617, \9343 );
and \U$19155 ( \28266 , RIdeba6e0_585, \9345 );
and \U$19156 ( \28267 , RIdeb79e0_553, \9347 );
and \U$19157 ( \28268 , RIfcb9858_7133, \9349 );
and \U$19158 ( \28269 , RIdeb1fe0_489, \9351 );
and \U$19159 ( \28270 , RIfc9efa8_6831, \9353 );
and \U$19160 ( \28271 , RIdeaf2e0_457, \9355 );
and \U$19161 ( \28272 , RIfce0750_7576, \9357 );
and \U$19162 ( \28273 , RIdeab488_425, \9359 );
and \U$19163 ( \28274 , RIdea4b88_393, \9361 );
and \U$19164 ( \28275 , RIde9e288_361, \9363 );
and \U$19165 ( \28276 , RIee1d0b0_4789, \9365 );
and \U$19166 ( \28277 , RIee1c138_4778, \9367 );
and \U$19167 ( \28278 , RIfcd0e68_7399, \9369 );
and \U$19168 ( \28279 , RIfc76d00_6374, \9371 );
and \U$19169 ( \28280 , RIfe89028_7903, \9373 );
and \U$19170 ( \28281 , RIfe88d58_7901, \9375 );
and \U$19171 ( \28282 , RIfe88ec0_7902, \9377 );
and \U$19172 ( \28283 , RIfe88bf0_7900, \9379 );
and \U$19173 ( \28284 , RIfcda7b0_7508, \9381 );
and \U$19174 ( \28285 , RIfc4d810_5904, \9383 );
and \U$19175 ( \28286 , RIfc52dd8_5965, \9385 );
and \U$19176 ( \28287 , RIfcde590_7552, \9387 );
and \U$19177 ( \28288 , RIfc4f868_5927, \9389 );
and \U$19178 ( \28289 , RIe16bd50_2604, \9391 );
and \U$19179 ( \28290 , RIfc68930_6212, \9393 );
and \U$19180 ( \28291 , RIe1683a8_2563, \9395 );
and \U$19181 ( \28292 , RIe165ae0_2534, \9397 );
and \U$19182 ( \28293 , RIe162de0_2502, \9399 );
and \U$19183 ( \28294 , RIfe88a88_7899, \9401 );
and \U$19184 ( \28295 , RIe1600e0_2470, \9403 );
and \U$19185 ( \28296 , RIfcc9140_7310, \9405 );
and \U$19186 ( \28297 , RIe15d3e0_2438, \9407 );
and \U$19187 ( \28298 , RIe1579e0_2374, \9409 );
and \U$19188 ( \28299 , RIe154ce0_2342, \9411 );
and \U$19189 ( \28300 , RIfc698a8_6223, \9413 );
and \U$19190 ( \28301 , RIe151fe0_2310, \9415 );
and \U$19191 ( \28302 , RIee35098_5062, \9417 );
and \U$19192 ( \28303 , RIe14f2e0_2278, \9419 );
and \U$19193 ( \28304 , RIfcc0338_7209, \9421 );
and \U$19194 ( \28305 , RIe14c5e0_2246, \9423 );
and \U$19195 ( \28306 , RIe1498e0_2214, \9425 );
and \U$19196 ( \28307 , RIe146be0_2182, \9427 );
and \U$19197 ( \28308 , RIfc88208_6571, \9429 );
and \U$19198 ( \28309 , RIfc85670_6540, \9431 );
and \U$19199 ( \28310 , RIfc81f98_6501, \9433 );
and \U$19200 ( \28311 , RIfcc4f28_7263, \9435 );
and \U$19201 ( \28312 , RIe1414b0_2120, \9437 );
and \U$19202 ( \28313 , RIe13f188_2095, \9439 );
and \U$19203 ( \28314 , RIdf3d090_2071, \9441 );
and \U$19204 ( \28315 , RIdf3aa98_2044, \9443 );
and \U$19205 ( \28316 , RIfcd2920_7418, \9445 );
and \U$19206 ( \28317 , RIfc7d7e0_6450, \9447 );
and \U$19207 ( \28318 , RIfc49760_5858, \9449 );
and \U$19208 ( \28319 , RIfce5a48_7635, \9451 );
and \U$19209 ( \28320 , RIdf35ea8_1990, \9453 );
and \U$19210 ( \28321 , RIdf338b0_1963, \9455 );
and \U$19211 ( \28322 , RIfe88920_7898, \9457 );
and \U$19212 ( \28323 , RIdf2f800_1917, \9459 );
or \U$19213 ( \28324 , \28260 , \28261 , \28262 , \28263 , \28264 , \28265 , \28266 , \28267 , \28268 , \28269 , \28270 , \28271 , \28272 , \28273 , \28274 , \28275 , \28276 , \28277 , \28278 , \28279 , \28280 , \28281 , \28282 , \28283 , \28284 , \28285 , \28286 , \28287 , \28288 , \28289 , \28290 , \28291 , \28292 , \28293 , \28294 , \28295 , \28296 , \28297 , \28298 , \28299 , \28300 , \28301 , \28302 , \28303 , \28304 , \28305 , \28306 , \28307 , \28308 , \28309 , \28310 , \28311 , \28312 , \28313 , \28314 , \28315 , \28316 , \28317 , \28318 , \28319 , \28320 , \28321 , \28322 , \28323 );
and \U$19214 ( \28325 , RIee2bfc0_4959, \9462 );
and \U$19215 ( \28326 , RIee2a670_4941, \9464 );
and \U$19216 ( \28327 , RIee29158_4926, \9466 );
and \U$19217 ( \28328 , RIee27f10_4913, \9468 );
and \U$19218 ( \28329 , RIdf2a7d8_1860, \9470 );
and \U$19219 ( \28330 , RIdf28618_1836, \9472 );
and \U$19220 ( \28331 , RIdf26890_1815, \9474 );
and \U$19221 ( \28332 , RIdf24dd8_1796, \9476 );
and \U$19222 ( \28333 , RIfcad918_6997, \9478 );
and \U$19223 ( \28334 , RIfc69fb0_6228, \9480 );
and \U$19224 ( \28335 , RIfc63368_6151, \9482 );
and \U$19225 ( \28336 , RIfc623f0_6140, \9484 );
and \U$19226 ( \28337 , RIfc60938_6121, \9486 );
and \U$19227 ( \28338 , RIdf1ff18_1740, \9488 );
and \U$19228 ( \28339 , RIfcba500_7142, \9490 );
and \U$19229 ( \28340 , RIdf19870_1667, \9492 );
and \U$19230 ( \28341 , RIdf176b0_1643, \9494 );
and \U$19231 ( \28342 , RIdf149b0_1611, \9496 );
and \U$19232 ( \28343 , RIdf11cb0_1579, \9498 );
and \U$19233 ( \28344 , RIdf0efb0_1547, \9500 );
and \U$19234 ( \28345 , RIdf0c2b0_1515, \9502 );
and \U$19235 ( \28346 , RIdf095b0_1483, \9504 );
and \U$19236 ( \28347 , RIdf068b0_1451, \9506 );
and \U$19237 ( \28348 , RIdf03bb0_1419, \9508 );
and \U$19238 ( \28349 , RIdefe1b0_1355, \9510 );
and \U$19239 ( \28350 , RIdefb4b0_1323, \9512 );
and \U$19240 ( \28351 , RIdef87b0_1291, \9514 );
and \U$19241 ( \28352 , RIdef5ab0_1259, \9516 );
and \U$19242 ( \28353 , RIdef2db0_1227, \9518 );
and \U$19243 ( \28354 , RIdef00b0_1195, \9520 );
and \U$19244 ( \28355 , RIdeed3b0_1163, \9522 );
and \U$19245 ( \28356 , RIdeea6b0_1131, \9524 );
and \U$19246 ( \28357 , RIfcc9848_7315, \9526 );
and \U$19247 ( \28358 , RIfc69a10_6224, \9528 );
and \U$19248 ( \28359 , RIfcacc70_6988, \9530 );
and \U$19249 ( \28360 , RIfccbfa8_7343, \9532 );
and \U$19250 ( \28361 , RIdee4f80_1069, \9534 );
and \U$19251 ( \28362 , RIdee31f8_1048, \9536 );
and \U$19252 ( \28363 , RIdee1038_1024, \9538 );
and \U$19253 ( \28364 , RIdedee78_1000, \9540 );
and \U$19254 ( \28365 , RIfc84590_6528, \9542 );
and \U$19255 ( \28366 , RIfc9bba0_6794, \9544 );
and \U$19256 ( \28367 , RIee21b38_4842, \9546 );
and \U$19257 ( \28368 , RIfc47168_5831, \9548 );
and \U$19258 ( \28369 , RIded9e50_943, \9550 );
and \U$19259 ( \28370 , RIded7858_916, \9552 );
and \U$19260 ( \28371 , RIfe887b8_7897, \9554 );
and \U$19261 ( \28372 , RIded34d8_868, \9556 );
and \U$19262 ( \28373 , RIded0ee0_841, \9558 );
and \U$19263 ( \28374 , RIdece1e0_809, \9560 );
and \U$19264 ( \28375 , RIdecb4e0_777, \9562 );
and \U$19265 ( \28376 , RIdec87e0_745, \9564 );
and \U$19266 ( \28377 , RIdeb4ce0_521, \9566 );
and \U$19267 ( \28378 , RIde97988_329, \9568 );
and \U$19268 ( \28379 , RIe16e8e8_2635, \9570 );
and \U$19269 ( \28380 , RIe15a6e0_2406, \9572 );
and \U$19270 ( \28381 , RIe143ee0_2150, \9574 );
and \U$19271 ( \28382 , RIdf388d8_2020, \9576 );
and \U$19272 ( \28383 , RIdf2cf38_1888, \9578 );
and \U$19273 ( \28384 , RIdf1d7b8_1712, \9580 );
and \U$19274 ( \28385 , RIdf00eb0_1387, \9582 );
and \U$19275 ( \28386 , RIdee79b0_1099, \9584 );
and \U$19276 ( \28387 , RIdedc718_972, \9586 );
and \U$19277 ( \28388 , RIde7d8d0_202, \9588 );
or \U$19278 ( \28389 , \28325 , \28326 , \28327 , \28328 , \28329 , \28330 , \28331 , \28332 , \28333 , \28334 , \28335 , \28336 , \28337 , \28338 , \28339 , \28340 , \28341 , \28342 , \28343 , \28344 , \28345 , \28346 , \28347 , \28348 , \28349 , \28350 , \28351 , \28352 , \28353 , \28354 , \28355 , \28356 , \28357 , \28358 , \28359 , \28360 , \28361 , \28362 , \28363 , \28364 , \28365 , \28366 , \28367 , \28368 , \28369 , \28370 , \28371 , \28372 , \28373 , \28374 , \28375 , \28376 , \28377 , \28378 , \28379 , \28380 , \28381 , \28382 , \28383 , \28384 , \28385 , \28386 , \28387 , \28388 );
or \U$19279 ( \28390 , \28324 , \28389 );
_DC g5fc4 ( \28391_nG5fc4 , \28390 , \9597 );
and \U$19280 ( \28392 , RIe19dd78_3173, \9059 );
and \U$19281 ( \28393 , RIe19b078_3141, \9061 );
and \U$19282 ( \28394 , RIfca1438_6857, \9063 );
and \U$19283 ( \28395 , RIe198378_3109, \9065 );
and \U$19284 ( \28396 , RIfca35f8_6881, \9067 );
and \U$19285 ( \28397 , RIe195678_3077, \9069 );
and \U$19286 ( \28398 , RIe192978_3045, \9071 );
and \U$19287 ( \28399 , RIe18fc78_3013, \9073 );
and \U$19288 ( \28400 , RIe18a278_2949, \9075 );
and \U$19289 ( \28401 , RIe187578_2917, \9077 );
and \U$19290 ( \28402 , RIfcba230_7140, \9079 );
and \U$19291 ( \28403 , RIe184878_2885, \9081 );
and \U$19292 ( \28404 , RIf142d90_5220, \9083 );
and \U$19293 ( \28405 , RIe181b78_2853, \9085 );
and \U$19294 ( \28406 , RIe17ee78_2821, \9087 );
and \U$19295 ( \28407 , RIe17c178_2789, \9089 );
and \U$19296 ( \28408 , RIfc9be70_6796, \9091 );
and \U$19297 ( \28409 , RIfc9bd08_6795, \9093 );
and \U$19298 ( \28410 , RIfc4ccd0_5896, \9095 );
and \U$19299 ( \28411 , RIe176070_2720, \9097 );
and \U$19300 ( \28412 , RIfc87c68_6567, \9099 );
and \U$19301 ( \28413 , RIfc87b00_6566, \9101 );
and \U$19302 ( \28414 , RIfcc4c58_7261, \9103 );
and \U$19303 ( \28415 , RIfc4fca0_5930, \9105 );
and \U$19304 ( \28416 , RIfc4f598_5925, \9107 );
and \U$19305 ( \28417 , RIfc876c8_6563, \9109 );
and \U$19306 ( \28418 , RIfc4dae0_5906, \9111 );
and \U$19307 ( \28419 , RIe173eb0_2696, \9113 );
and \U$19308 ( \28420 , RIfcb9420_7130, \9115 );
and \U$19309 ( \28421 , RIfc4e080_5910, \9117 );
and \U$19310 ( \28422 , RIfc4e350_5912, \9119 );
and \U$19311 ( \28423 , RIfc9d388_6811, \9121 );
and \U$19312 ( \28424 , RIfc40a48_5761, \9123 );
and \U$19313 ( \28425 , RIe2240d0_4700, \9125 );
and \U$19314 ( \28426 , RIfc85508_6539, \9127 );
and \U$19315 ( \28427 , RIe2213d0_4668, \9129 );
and \U$19316 ( \28428 , RIfc9ba38_6793, \9131 );
and \U$19317 ( \28429 , RIe21e6d0_4636, \9133 );
and \U$19318 ( \28430 , RIe218cd0_4572, \9135 );
and \U$19319 ( \28431 , RIe215fd0_4540, \9137 );
and \U$19320 ( \28432 , RIfc52c70_5964, \9139 );
and \U$19321 ( \28433 , RIe2132d0_4508, \9141 );
and \U$19322 ( \28434 , RIfca3760_6882, \9143 );
and \U$19323 ( \28435 , RIe2105d0_4476, \9145 );
and \U$19324 ( \28436 , RIfc97988_6747, \9147 );
and \U$19325 ( \28437 , RIe20d8d0_4444, \9149 );
and \U$19326 ( \28438 , RIe20abd0_4412, \9151 );
and \U$19327 ( \28439 , RIe207ed0_4380, \9153 );
and \U$19328 ( \28440 , RIfceb5b0_7700, \9155 );
and \U$19329 ( \28441 , RIfcddbb8_7545, \9157 );
and \U$19330 ( \28442 , RIe202a70_4320, \9159 );
and \U$19331 ( \28443 , RIe200e50_4300, \9161 );
and \U$19332 ( \28444 , RIfc73d30_6340, \9163 );
and \U$19333 ( \28445 , RIfcaf100_7014, \9165 );
and \U$19334 ( \28446 , RIfc71468_6311, \9167 );
and \U$19335 ( \28447 , RIfcdcad8_7533, \9169 );
and \U$19336 ( \28448 , RIfcdda50_7544, \9171 );
and \U$19337 ( \28449 , RIfca8620_6938, \9173 );
and \U$19338 ( \28450 , RIe1fcf08_4255, \9175 );
and \U$19339 ( \28451 , RIe1fbcc0_4242, \9177 );
and \U$19340 ( \28452 , RIfc6c008_6251, \9179 );
and \U$19341 ( \28453 , RIfcdd1e0_7538, \9181 );
and \U$19342 ( \28454 , RIfca9700_6950, \9183 );
and \U$19343 ( \28455 , RIfca92c8_6947, \9185 );
or \U$19344 ( \28456 , \28392 , \28393 , \28394 , \28395 , \28396 , \28397 , \28398 , \28399 , \28400 , \28401 , \28402 , \28403 , \28404 , \28405 , \28406 , \28407 , \28408 , \28409 , \28410 , \28411 , \28412 , \28413 , \28414 , \28415 , \28416 , \28417 , \28418 , \28419 , \28420 , \28421 , \28422 , \28423 , \28424 , \28425 , \28426 , \28427 , \28428 , \28429 , \28430 , \28431 , \28432 , \28433 , \28434 , \28435 , \28436 , \28437 , \28438 , \28439 , \28440 , \28441 , \28442 , \28443 , \28444 , \28445 , \28446 , \28447 , \28448 , \28449 , \28450 , \28451 , \28452 , \28453 , \28454 , \28455 );
and \U$19345 ( \28457 , RIfcce5a0_7370, \9188 );
and \U$19346 ( \28458 , RIfc6ba68_6247, \9190 );
and \U$19347 ( \28459 , RIfc6f410_6288, \9192 );
and \U$19348 ( \28460 , RIe1fa640_4226, \9194 );
and \U$19349 ( \28461 , RIfcce000_7366, \9196 );
and \U$19350 ( \28462 , RIfc53918_5973, \9198 );
and \U$19351 ( \28463 , RIfcce708_7371, \9200 );
and \U$19352 ( \28464 , RIe1f5bb8_4173, \9202 );
and \U$19353 ( \28465 , RIf1535f0_5408, \9204 );
and \U$19354 ( \28466 , RIf151e08_5391, \9206 );
and \U$19355 ( \28467 , RIfc72db8_6329, \9208 );
and \U$19356 ( \28468 , RIe1f3890_4148, \9210 );
and \U$19357 ( \28469 , RIf14fc48_5367, \9212 );
and \U$19358 ( \28470 , RIfc72c50_6328, \9214 );
and \U$19359 ( \28471 , RIfc73e98_6341, \9216 );
and \U$19360 ( \28472 , RIe1ee598_4089, \9218 );
and \U$19361 ( \28473 , RIe1ebe38_4061, \9220 );
and \U$19362 ( \28474 , RIe1e9138_4029, \9222 );
and \U$19363 ( \28475 , RIe1e6438_3997, \9224 );
and \U$19364 ( \28476 , RIe1e3738_3965, \9226 );
and \U$19365 ( \28477 , RIe1e0a38_3933, \9228 );
and \U$19366 ( \28478 , RIe1ddd38_3901, \9230 );
and \U$19367 ( \28479 , RIe1db038_3869, \9232 );
and \U$19368 ( \28480 , RIe1d8338_3837, \9234 );
and \U$19369 ( \28481 , RIe1d2938_3773, \9236 );
and \U$19370 ( \28482 , RIe1cfc38_3741, \9238 );
and \U$19371 ( \28483 , RIe1ccf38_3709, \9240 );
and \U$19372 ( \28484 , RIe1ca238_3677, \9242 );
and \U$19373 ( \28485 , RIe1c7538_3645, \9244 );
and \U$19374 ( \28486 , RIe1c4838_3613, \9246 );
and \U$19375 ( \28487 , RIe1c1b38_3581, \9248 );
and \U$19376 ( \28488 , RIe1bee38_3549, \9250 );
and \U$19377 ( \28489 , RIfcb8a48_7123, \9252 );
and \U$19378 ( \28490 , RIfcb84a8_7119, \9254 );
and \U$19379 ( \28491 , RIe1b9870_3488, \9256 );
and \U$19380 ( \28492 , RIe1b7818_3465, \9258 );
and \U$19381 ( \28493 , RIfc85940_6542, \9260 );
and \U$19382 ( \28494 , RIfc9e198_6821, \9262 );
and \U$19383 ( \28495 , RIfeac140_8274, \9264 );
and \U$19384 ( \28496 , RIe1b42a8_3427, \9266 );
and \U$19385 ( \28497 , RIfc518c0_5950, \9268 );
and \U$19386 ( \28498 , RIfc838e8_6519, \9270 );
and \U$19387 ( \28499 , RIfe884e8_7895, \9272 );
and \U$19388 ( \28500 , RIe1b1008_3391, \9274 );
and \U$19389 ( \28501 , RIfcc5900_7270, \9276 );
and \U$19390 ( \28502 , RIfc82ad8_6509, \9278 );
and \U$19391 ( \28503 , RIe1ac9b8_3341, \9280 );
and \U$19392 ( \28504 , RIfe88650_7896, \9282 );
and \U$19393 ( \28505 , RIe1a9178_3301, \9284 );
and \U$19394 ( \28506 , RIe1a6478_3269, \9286 );
and \U$19395 ( \28507 , RIe1a3778_3237, \9288 );
and \U$19396 ( \28508 , RIe1a0a78_3205, \9290 );
and \U$19397 ( \28509 , RIe18cf78_2981, \9292 );
and \U$19398 ( \28510 , RIe179478_2757, \9294 );
and \U$19399 ( \28511 , RIe226dd0_4732, \9296 );
and \U$19400 ( \28512 , RIe21b9d0_4604, \9298 );
and \U$19401 ( \28513 , RIe2051d0_4348, \9300 );
and \U$19402 ( \28514 , RIe1ff230_4280, \9302 );
and \U$19403 ( \28515 , RIe1f85e8_4203, \9304 );
and \U$19404 ( \28516 , RIe1f1130_4120, \9306 );
and \U$19405 ( \28517 , RIe1d5638_3805, \9308 );
and \U$19406 ( \28518 , RIe1bc138_3517, \9310 );
and \U$19407 ( \28519 , RIe1aefb0_3368, \9312 );
and \U$19408 ( \28520 , RIe1715e8_2667, \9314 );
or \U$19409 ( \28521 , \28457 , \28458 , \28459 , \28460 , \28461 , \28462 , \28463 , \28464 , \28465 , \28466 , \28467 , \28468 , \28469 , \28470 , \28471 , \28472 , \28473 , \28474 , \28475 , \28476 , \28477 , \28478 , \28479 , \28480 , \28481 , \28482 , \28483 , \28484 , \28485 , \28486 , \28487 , \28488 , \28489 , \28490 , \28491 , \28492 , \28493 , \28494 , \28495 , \28496 , \28497 , \28498 , \28499 , \28500 , \28501 , \28502 , \28503 , \28504 , \28505 , \28506 , \28507 , \28508 , \28509 , \28510 , \28511 , \28512 , \28513 , \28514 , \28515 , \28516 , \28517 , \28518 , \28519 , \28520 );
or \U$19410 ( \28522 , \28456 , \28521 );
_DC g6048 ( \28523_nG6048 , \28522 , \9323 );
xor g6049 ( \28524_nG6049 , \28391_nG5fc4 , \28523_nG6048 );
buf \U$19411 ( \28525 , \28524_nG6049 );
xor \U$19412 ( \28526 , \28525 , \27292 );
and \U$19413 ( \28527 , \10687 , \28526 );
xor \U$19414 ( \28528 , \28259 , \28527 );
xor \U$19415 ( \28529 , \28250 , \28528 );
and \U$19416 ( \28530 , \27313 , \10983 );
_DC g65c5 ( \28531_nG65c5 , \28390 , \9597 );
_DC g65c6 ( \28532_nG65c6 , \28522 , \9323 );
and g65c7 ( \28533_nG65c7 , \28531_nG65c5 , \28532_nG65c6 );
buf \U$19417 ( \28534 , \28533_nG65c7 );
and \U$19418 ( \28535 , \28534 , \10691 );
nor \U$19419 ( \28536 , \28530 , \28535 );
xnor \U$19420 ( \28537 , \28536 , \10980 );
and \U$19421 ( \28538 , \14024 , \22542 );
and \U$19422 ( \28539 , \14950 , \22103 );
nor \U$19423 ( \28540 , \28538 , \28539 );
xnor \U$19424 ( \28541 , \28540 , \22548 );
xor \U$19425 ( \28542 , \28537 , \28541 );
and \U$19426 ( \28543 , \12769 , \24138 );
and \U$19427 ( \28544 , \13679 , \23630 );
nor \U$19428 ( \28545 , \28543 , \28544 );
xnor \U$19429 ( \28546 , \28545 , \24144 );
xor \U$19430 ( \28547 , \28542 , \28546 );
xor \U$19431 ( \28548 , \28529 , \28547 );
xor \U$19432 ( \28549 , \28246 , \28548 );
and \U$19433 ( \28550 , \19558 , \16635 );
and \U$19434 ( \28551 , \20544 , \16301 );
nor \U$19435 ( \28552 , \28550 , \28551 );
xnor \U$19436 ( \28553 , \28552 , \16625 );
and \U$19437 ( \28554 , \11586 , \25826 );
and \U$19438 ( \28555 , \12448 , \25264 );
nor \U$19439 ( \28556 , \28554 , \28555 );
xnor \U$19440 ( \28557 , \28556 , \25773 );
xor \U$19441 ( \28558 , \28553 , \28557 );
and \U$19442 ( \28559 , \10988 , \27397 );
and \U$19443 ( \28560 , \11270 , \26807 );
nor \U$19444 ( \28561 , \28559 , \28560 );
xnor \U$19445 ( \28562 , \28561 , \27295 );
xor \U$19446 ( \28563 , \28558 , \28562 );
and \U$19447 ( \28564 , \21033 , \15336 );
and \U$19448 ( \28565 , \22090 , \14963 );
nor \U$19449 ( \28566 , \28564 , \28565 );
xnor \U$19450 ( \28567 , \28566 , \15342 );
and \U$19451 ( \28568 , \16655 , \19534 );
and \U$19452 ( \28569 , \17627 , \19045 );
nor \U$19453 ( \28570 , \28568 , \28569 );
xnor \U$19454 ( \28571 , \28570 , \19540 );
xor \U$19455 ( \28572 , \28567 , \28571 );
and \U$19456 ( \28573 , \15321 , \21005 );
and \U$19457 ( \28574 , \16267 , \20557 );
nor \U$19458 ( \28575 , \28573 , \28574 );
xnor \U$19459 ( \28576 , \28575 , \21011 );
xor \U$19460 ( \28577 , \28572 , \28576 );
xor \U$19461 ( \28578 , \28563 , \28577 );
and \U$19462 ( \28579 , \27025 , \27296 );
and \U$19463 ( \28580 , \24199 , \12790 );
and \U$19464 ( \28581 , \25272 , \12461 );
nor \U$19465 ( \28582 , \28580 , \28581 );
xnor \U$19466 ( \28583 , \28582 , \12780 );
xor \U$19467 ( \28584 , \28579 , \28583 );
and \U$19468 ( \28585 , \18035 , \18090 );
and \U$19469 ( \28586 , \19032 , \17655 );
nor \U$19470 ( \28587 , \28585 , \28586 );
xnor \U$19471 ( \28588 , \28587 , \18046 );
xor \U$19472 ( \28589 , \28584 , \28588 );
xor \U$19473 ( \28590 , \28578 , \28589 );
xor \U$19474 ( \28591 , \28549 , \28590 );
xor \U$19475 ( \28592 , \28232 , \28591 );
and \U$19476 ( \28593 , \27017 , \27357 );
and \U$19477 ( \28594 , \27357 , \27405 );
and \U$19478 ( \28595 , \27017 , \27405 );
or \U$19479 ( \28596 , \28593 , \28594 , \28595 );
xor \U$19480 ( \28597 , \28592 , \28596 );
and \U$19481 ( \28598 , \27406 , \27410 );
and \U$19482 ( \28599 , \27411 , \27414 );
or \U$19483 ( \28600 , \28598 , \28599 );
xor \U$19484 ( \28601 , \28597 , \28600 );
buf g9bc0 ( \28602_nG9bc0 , \28601 );
and \U$19485 ( \28603 , \10704 , \28602_nG9bc0 );
or \U$19486 ( \28604 , \28203 , \28603 );
xor \U$19487 ( \28605 , \10703 , \28604 );
buf \U$19488 ( \28606 , \28605 );
buf \U$19490 ( \28607 , \28606 );
xor \U$19491 ( \28608 , \28202 , \28607 );
buf \U$19492 ( \28609 , \28608 );
xor \U$19493 ( \28610 , \28135 , \28609 );
and \U$19494 ( \28611 , \27005 , \27011 );
and \U$19495 ( \28612 , \27005 , \27421 );
and \U$19496 ( \28613 , \27011 , \27421 );
or \U$19497 ( \28614 , \28611 , \28612 , \28613 );
buf \U$19498 ( \28615 , \28614 );
xor \U$19499 ( \28616 , \28610 , \28615 );
buf \U$19500 ( \28617 , \28616 );
and \U$19501 ( \28618 , \27464 , \27470 );
and \U$19502 ( \28619 , \27464 , \27477 );
and \U$19503 ( \28620 , \27470 , \27477 );
or \U$19504 ( \28621 , \28618 , \28619 , \28620 );
buf \U$19505 ( \28622 , \28621 );
and \U$19506 ( \28623 , \27440 , \27446 );
and \U$19507 ( \28624 , \27440 , \27453 );
and \U$19508 ( \28625 , \27446 , \27453 );
or \U$19509 ( \28626 , \28623 , \28624 , \28625 );
buf \U$19510 ( \28627 , \28626 );
and \U$19511 ( \28628 , \26431 , \10995_nG9c0b );
and \U$19512 ( \28629 , \26428 , \11283_nG9c08 );
or \U$19513 ( \28630 , \28628 , \28629 );
xor \U$19514 ( \28631 , \26427 , \28630 );
buf \U$19515 ( \28632 , \28631 );
buf \U$19517 ( \28633 , \28632 );
and \U$19518 ( \28634 , \24792 , \11598_nG9c05 );
and \U$19519 ( \28635 , \24789 , \12470_nG9c02 );
or \U$19520 ( \28636 , \28634 , \28635 );
xor \U$19521 ( \28637 , \24788 , \28636 );
buf \U$19522 ( \28638 , \28637 );
buf \U$19524 ( \28639 , \28638 );
xor \U$19525 ( \28640 , \28633 , \28639 );
buf \U$19526 ( \28641 , \28640 );
xor \U$19527 ( \28642 , \28627 , \28641 );
and \U$19528 ( \28643 , \20155 , \15373_nG9bf3 );
and \U$19529 ( \28644 , \20152 , \16315_nG9bf0 );
or \U$19530 ( \28645 , \28643 , \28644 );
xor \U$19531 ( \28646 , \20151 , \28645 );
buf \U$19532 ( \28647 , \28646 );
buf \U$19534 ( \28648 , \28647 );
xor \U$19535 ( \28649 , \28642 , \28648 );
buf \U$19536 ( \28650 , \28649 );
and \U$19537 ( \28651 , \27481 , \27487 );
and \U$19538 ( \28652 , \27481 , \27494 );
and \U$19539 ( \28653 , \27487 , \27494 );
or \U$19540 ( \28654 , \28651 , \28652 , \28653 );
buf \U$19541 ( \28655 , \28654 );
xor \U$19542 ( \28656 , \28650 , \28655 );
and \U$19543 ( \28657 , \14631 , \21086_nG9bdb );
and \U$19544 ( \28658 , \14628 , \22129_nG9bd8 );
or \U$19545 ( \28659 , \28657 , \28658 );
xor \U$19546 ( \28660 , \14627 , \28659 );
buf \U$19547 ( \28661 , \28660 );
buf \U$19549 ( \28662 , \28661 );
xor \U$19550 ( \28663 , \28656 , \28662 );
buf \U$19551 ( \28664 , \28663 );
xor \U$19552 ( \28665 , \28622 , \28664 );
and \U$19553 ( \28666 , \10421 , \25860_nG9bc9 );
and \U$19554 ( \28667 , \10418 , \26887_nG9bc6 );
or \U$19555 ( \28668 , \28666 , \28667 );
xor \U$19556 ( \28669 , \10417 , \28668 );
buf \U$19557 ( \28670 , \28669 );
buf \U$19559 ( \28671 , \28670 );
xor \U$19560 ( \28672 , \28665 , \28671 );
buf \U$19561 ( \28673 , \28672 );
and \U$19562 ( \28674 , \27479 , \27510 );
and \U$19563 ( \28675 , \27479 , \27517 );
and \U$19564 ( \28676 , \27510 , \27517 );
or \U$19565 ( \28677 , \28674 , \28675 , \28676 );
buf \U$19566 ( \28678 , \28677 );
xor \U$19567 ( \28679 , \28673 , \28678 );
and \U$19568 ( \28680 , \27537 , \27542 );
and \U$19569 ( \28681 , \27537 , \27549 );
and \U$19570 ( \28682 , \27542 , \27549 );
or \U$19571 ( \28683 , \28680 , \28681 , \28682 );
buf \U$19572 ( \28684 , \28683 );
xor \U$19573 ( \28685 , \28679 , \28684 );
buf \U$19574 ( \28686 , \28685 );
xor \U$19575 ( \28687 , \28617 , \28686 );
and \U$19576 ( \28688 , \27000 , \27423 );
and \U$19577 ( \28689 , \27000 , \27519 );
and \U$19578 ( \28690 , \27423 , \27519 );
or \U$19579 ( \28691 , \28688 , \28689 , \28690 );
buf \U$19580 ( \28692 , \28691 );
xor \U$19581 ( \28693 , \28687 , \28692 );
and \U$19582 ( \28694 , \28125 , \28693 );
and \U$19583 ( \28695 , \28129 , \28693 );
or \U$19584 ( \28696 , \28130 , \28694 , \28695 );
and \U$19585 ( \28697 , \27561 , \27565 );
and \U$19586 ( \28698 , \27561 , \28124 );
and \U$19587 ( \28699 , \27565 , \28124 );
or \U$19588 ( \28700 , \28697 , \28698 , \28699 );
xor \U$19589 ( \28701 , \28696 , \28700 );
and \U$19590 ( \28702 , \28617 , \28686 );
and \U$19591 ( \28703 , \28617 , \28692 );
and \U$19592 ( \28704 , \28686 , \28692 );
or \U$19593 ( \28705 , \28702 , \28703 , \28704 );
xor \U$19594 ( \28706 , \28701 , \28705 );
and \U$19595 ( \28707 , \28673 , \28678 );
and \U$19596 ( \28708 , \28673 , \28684 );
and \U$19597 ( \28709 , \28678 , \28684 );
or \U$19598 ( \28710 , \28707 , \28708 , \28709 );
buf \U$19599 ( \28711 , \28710 );
and \U$19600 ( \28712 , \28187 , \28192 );
and \U$19601 ( \28713 , \28187 , \28199 );
and \U$19602 ( \28714 , \28192 , \28199 );
or \U$19603 ( \28715 , \28712 , \28713 , \28714 );
buf \U$19604 ( \28716 , \28715 );
and \U$19605 ( \28717 , \28172 , \28178 );
and \U$19606 ( \28718 , \28172 , \28185 );
and \U$19607 ( \28719 , \28178 , \28185 );
or \U$19608 ( \28720 , \28717 , \28718 , \28719 );
buf \U$19609 ( \28721 , \28720 );
and \U$19610 ( \28722 , \14631 , \22129_nG9bd8 );
and \U$19611 ( \28723 , \14628 , \22629_nG9bd5 );
or \U$19612 ( \28724 , \28722 , \28723 );
xor \U$19613 ( \28725 , \14627 , \28724 );
buf \U$19614 ( \28726 , \28725 );
buf \U$19616 ( \28727 , \28726 );
xor \U$19617 ( \28728 , \28721 , \28727 );
and \U$19618 ( \28729 , \13370 , \23696_nG9bd2 );
and \U$19619 ( \28730 , \13367 , \24226_nG9bcf );
or \U$19620 ( \28731 , \28729 , \28730 );
xor \U$19621 ( \28732 , \13366 , \28731 );
buf \U$19622 ( \28733 , \28732 );
buf \U$19624 ( \28734 , \28733 );
xor \U$19625 ( \28735 , \28728 , \28734 );
buf \U$19626 ( \28736 , \28735 );
xor \U$19627 ( \28737 , \28716 , \28736 );
and \U$19628 ( \28738 , \28140 , \28146 );
and \U$19629 ( \28739 , \28140 , \28153 );
and \U$19630 ( \28740 , \28146 , \28153 );
or \U$19631 ( \28741 , \28738 , \28739 , \28740 );
buf \U$19632 ( \28742 , \28741 );
xor \U$19633 ( \28743 , \28737 , \28742 );
buf \U$19634 ( \28744 , \28743 );
xor \U$19635 ( \28745 , \28711 , \28744 );
and \U$19636 ( \28746 , \28155 , \28201 );
and \U$19637 ( \28747 , \28155 , \28607 );
and \U$19638 ( \28748 , \28201 , \28607 );
or \U$19639 ( \28749 , \28746 , \28747 , \28748 );
buf \U$19640 ( \28750 , \28749 );
xor \U$19641 ( \28751 , \28745 , \28750 );
buf \U$19642 ( \28752 , \28751 );
and \U$19643 ( \28753 , \12157 , \25298_nG9bcc );
and \U$19644 ( \28754 , \12154 , \25860_nG9bc9 );
or \U$19645 ( \28755 , \28753 , \28754 );
xor \U$19646 ( \28756 , \12153 , \28755 );
buf \U$19647 ( \28757 , \28756 );
buf \U$19649 ( \28758 , \28757 );
and \U$19650 ( \28759 , \10421 , \26887_nG9bc6 );
and \U$19651 ( \28760 , \10418 , \27416_nG9bc3 );
or \U$19652 ( \28761 , \28759 , \28760 );
xor \U$19653 ( \28762 , \10417 , \28761 );
buf \U$19654 ( \28763 , \28762 );
buf \U$19656 ( \28764 , \28763 );
xor \U$19657 ( \28765 , \28758 , \28764 );
and \U$19658 ( \28766 , \10707 , \28602_nG9bc0 );
and \U$19659 ( \28767 , \28207 , \28231 );
and \U$19660 ( \28768 , \28231 , \28591 );
and \U$19661 ( \28769 , \28207 , \28591 );
or \U$19662 ( \28770 , \28767 , \28768 , \28769 );
and \U$19663 ( \28771 , \28211 , \28215 );
and \U$19664 ( \28772 , \28215 , \28230 );
and \U$19665 ( \28773 , \28211 , \28230 );
or \U$19666 ( \28774 , \28771 , \28772 , \28773 );
and \U$19667 ( \28775 , \28563 , \28577 );
and \U$19668 ( \28776 , \28577 , \28589 );
and \U$19669 ( \28777 , \28563 , \28589 );
or \U$19670 ( \28778 , \28775 , \28776 , \28777 );
and \U$19671 ( \28779 , \23617 , \14054 );
and \U$19672 ( \28780 , \24199 , \13692 );
nor \U$19673 ( \28781 , \28779 , \28780 );
xnor \U$19674 ( \28782 , \28781 , \14035 );
and \U$19675 ( \28783 , \17627 , \19534 );
and \U$19676 ( \28784 , \18035 , \19045 );
nor \U$19677 ( \28785 , \28783 , \28784 );
xnor \U$19678 ( \28786 , \28785 , \19540 );
xor \U$19679 ( \28787 , \28782 , \28786 );
and \U$19680 ( \28788 , \16267 , \21005 );
and \U$19681 ( \28789 , \16655 , \20557 );
nor \U$19682 ( \28790 , \28788 , \28789 );
xnor \U$19683 ( \28791 , \28790 , \21011 );
xor \U$19684 ( \28792 , \28787 , \28791 );
and \U$19685 ( \28793 , \25272 , \12790 );
and \U$19686 ( \28794 , \25815 , \12461 );
nor \U$19687 ( \28795 , \28793 , \28794 );
xnor \U$19688 ( \28796 , \28795 , \12780 );
and \U$19689 ( \28797 , \11270 , \27397 );
and \U$19690 ( \28798 , \11586 , \26807 );
nor \U$19691 ( \28799 , \28797 , \28798 );
xnor \U$19692 ( \28800 , \28799 , \27295 );
xor \U$19693 ( \28801 , \28796 , \28800 );
and \U$19694 ( \28802 , RIdec5c48_714, \9333 );
and \U$19695 ( \28803 , RIdec2f48_682, \9335 );
and \U$19696 ( \28804 , RIfc7c160_6434, \9337 );
and \U$19697 ( \28805 , RIdec0248_650, \9339 );
and \U$19698 ( \28806 , RIfcb38b8_7065, \9341 );
and \U$19699 ( \28807 , RIdebd548_618, \9343 );
and \U$19700 ( \28808 , RIdeba848_586, \9345 );
and \U$19701 ( \28809 , RIdeb7b48_554, \9347 );
and \U$19702 ( \28810 , RIfce7c08_7659, \9349 );
and \U$19703 ( \28811 , RIdeb2148_490, \9351 );
and \U$19704 ( \28812 , RIfce7aa0_7658, \9353 );
and \U$19705 ( \28813 , RIdeaf448_458, \9355 );
and \U$19706 ( \28814 , RIfca38c8_6883, \9357 );
and \U$19707 ( \28815 , RIdeab7d0_426, \9359 );
and \U$19708 ( \28816 , RIdea4ed0_394, \9361 );
and \U$19709 ( \28817 , RIde9e5d0_362, \9363 );
and \U$19710 ( \28818 , RIfc41e70_5772, \9365 );
and \U$19711 ( \28819 , RIfc5b0a0_6058, \9367 );
and \U$19712 ( \28820 , RIfcdbb60_7522, \9369 );
and \U$19713 ( \28821 , RIfc78650_6392, \9371 );
and \U$19714 ( \28822 , RIfea92d8_8241, \9373 );
and \U$19715 ( \28823 , RIde8e5e0_284, \9375 );
and \U$19716 ( \28824 , RIfea0d40_8174, \9377 );
and \U$19717 ( \28825 , RIfea0bd8_8173, \9379 );
and \U$19718 ( \28826 , RIfcdf508_7563, \9381 );
and \U$19719 ( \28827 , RIfcb1b30_7044, \9383 );
and \U$19720 ( \28828 , RIfc5ccc0_6078, \9385 );
and \U$19721 ( \28829 , RIfcb16f8_7041, \9387 );
and \U$19722 ( \28830 , RIfc77b10_6384, \9389 );
and \U$19723 ( \28831 , RIe16beb8_2605, \9391 );
and \U$19724 ( \28832 , RIe169e60_2582, \9393 );
and \U$19725 ( \28833 , RIe168510_2564, \9395 );
and \U$19726 ( \28834 , RIe165c48_2535, \9397 );
and \U$19727 ( \28835 , RIe162f48_2503, \9399 );
and \U$19728 ( \28836 , RIfc4f9d0_5928, \9401 );
and \U$19729 ( \28837 , RIe160248_2471, \9403 );
and \U$19730 ( \28838 , RIfc4e8f0_5916, \9405 );
and \U$19731 ( \28839 , RIe15d548_2439, \9407 );
and \U$19732 ( \28840 , RIe157b48_2375, \9409 );
and \U$19733 ( \28841 , RIe154e48_2343, \9411 );
and \U$19734 ( \28842 , RIfc4e1e8_5911, \9413 );
and \U$19735 ( \28843 , RIe152148_2311, \9415 );
and \U$19736 ( \28844 , RIfc868b8_6553, \9417 );
and \U$19737 ( \28845 , RIe14f448_2279, \9419 );
and \U$19738 ( \28846 , RIfc865e8_6551, \9421 );
and \U$19739 ( \28847 , RIe14c748_2247, \9423 );
and \U$19740 ( \28848 , RIe149a48_2215, \9425 );
and \U$19741 ( \28849 , RIe146d48_2183, \9427 );
and \U$19742 ( \28850 , RIfc9eb70_6828, \9429 );
and \U$19743 ( \28851 , RIfc9ecd8_6829, \9431 );
and \U$19744 ( \28852 , RIfcc5630_7268, \9433 );
and \U$19745 ( \28853 , RIfc83bb8_6521, \9435 );
and \U$19746 ( \28854 , RIe141618_2121, \9437 );
and \U$19747 ( \28855 , RIfea0ea8_8175, \9439 );
and \U$19748 ( \28856 , RIdf3d1f8_2072, \9441 );
and \U$19749 ( \28857 , RIdf3ac00_2045, \9443 );
and \U$19750 ( \28858 , RIee308e0_5011, \9445 );
and \U$19751 ( \28859 , RIfcd3cd0_7432, \9447 );
and \U$19752 ( \28860 , RIfc84e00_6534, \9449 );
and \U$19753 ( \28861 , RIfc834b0_6516, \9451 );
and \U$19754 ( \28862 , RIdf36010_1991, \9453 );
and \U$19755 ( \28863 , RIdf33a18_1964, \9455 );
and \U$19756 ( \28864 , RIdf31858_1940, \9457 );
and \U$19757 ( \28865 , RIdf2f968_1918, \9459 );
or \U$19758 ( \28866 , \28802 , \28803 , \28804 , \28805 , \28806 , \28807 , \28808 , \28809 , \28810 , \28811 , \28812 , \28813 , \28814 , \28815 , \28816 , \28817 , \28818 , \28819 , \28820 , \28821 , \28822 , \28823 , \28824 , \28825 , \28826 , \28827 , \28828 , \28829 , \28830 , \28831 , \28832 , \28833 , \28834 , \28835 , \28836 , \28837 , \28838 , \28839 , \28840 , \28841 , \28842 , \28843 , \28844 , \28845 , \28846 , \28847 , \28848 , \28849 , \28850 , \28851 , \28852 , \28853 , \28854 , \28855 , \28856 , \28857 , \28858 , \28859 , \28860 , \28861 , \28862 , \28863 , \28864 , \28865 );
and \U$19759 ( \28867 , RIee2c128_4960, \9462 );
and \U$19760 ( \28868 , RIee2a7d8_4942, \9464 );
and \U$19761 ( \28869 , RIee292c0_4927, \9466 );
and \U$19762 ( \28870 , RIee28078_4914, \9468 );
and \U$19763 ( \28871 , RIdf2a940_1861, \9470 );
and \U$19764 ( \28872 , RIdf28780_1837, \9472 );
and \U$19765 ( \28873 , RIfea0a70_8172, \9474 );
and \U$19766 ( \28874 , RIfea0908_8171, \9476 );
and \U$19767 ( \28875 , RIfcd4f18_7445, \9478 );
and \U$19768 ( \28876 , RIfca0628_6847, \9480 );
and \U$19769 ( \28877 , RIdf23050_1775, \9482 );
and \U$19770 ( \28878 , RIfcd3190_7424, \9484 );
and \U$19771 ( \28879 , RIdf21b38_1760, \9486 );
and \U$19772 ( \28880 , RIdf20080_1741, \9488 );
and \U$19773 ( \28881 , RIdf1b328_1686, \9490 );
and \U$19774 ( \28882 , RIdf199d8_1668, \9492 );
and \U$19775 ( \28883 , RIdf17818_1644, \9494 );
and \U$19776 ( \28884 , RIdf14b18_1612, \9496 );
and \U$19777 ( \28885 , RIdf11e18_1580, \9498 );
and \U$19778 ( \28886 , RIdf0f118_1548, \9500 );
and \U$19779 ( \28887 , RIdf0c418_1516, \9502 );
and \U$19780 ( \28888 , RIdf09718_1484, \9504 );
and \U$19781 ( \28889 , RIdf06a18_1452, \9506 );
and \U$19782 ( \28890 , RIdf03d18_1420, \9508 );
and \U$19783 ( \28891 , RIdefe318_1356, \9510 );
and \U$19784 ( \28892 , RIdefb618_1324, \9512 );
and \U$19785 ( \28893 , RIdef8918_1292, \9514 );
and \U$19786 ( \28894 , RIdef5c18_1260, \9516 );
and \U$19787 ( \28895 , RIdef2f18_1228, \9518 );
and \U$19788 ( \28896 , RIdef0218_1196, \9520 );
and \U$19789 ( \28897 , RIdeed518_1164, \9522 );
and \U$19790 ( \28898 , RIdeea818_1132, \9524 );
and \U$19791 ( \28899 , RIfcdf3a0_7562, \9526 );
and \U$19792 ( \28900 , RIfca5218_6901, \9528 );
and \U$19793 ( \28901 , RIfcdc538_7529, \9530 );
and \U$19794 ( \28902 , RIfcdc6a0_7530, \9532 );
and \U$19795 ( \28903 , RIdee50e8_1070, \9534 );
and \U$19796 ( \28904 , RIdee3360_1049, \9536 );
and \U$19797 ( \28905 , RIfea07a0_8170, \9538 );
and \U$19798 ( \28906 , RIdedefe0_1001, \9540 );
and \U$19799 ( \28907 , RIfcb0d20_7034, \9542 );
and \U$19800 ( \28908 , RIfcd4978_7441, \9544 );
and \U$19801 ( \28909 , RIfca49a8_6895, \9546 );
and \U$19802 ( \28910 , RIfca1708_6859, \9548 );
and \U$19803 ( \28911 , RIded9fb8_944, \9550 );
and \U$19804 ( \28912 , RIded79c0_917, \9552 );
and \U$19805 ( \28913 , RIded5ad0_895, \9554 );
and \U$19806 ( \28914 , RIfeab498_8265, \9556 );
and \U$19807 ( \28915 , RIded1048_842, \9558 );
and \U$19808 ( \28916 , RIdece348_810, \9560 );
and \U$19809 ( \28917 , RIdecb648_778, \9562 );
and \U$19810 ( \28918 , RIdec8948_746, \9564 );
and \U$19811 ( \28919 , RIdeb4e48_522, \9566 );
and \U$19812 ( \28920 , RIde97cd0_330, \9568 );
and \U$19813 ( \28921 , RIe16ea50_2636, \9570 );
and \U$19814 ( \28922 , RIe15a848_2407, \9572 );
and \U$19815 ( \28923 , RIe144048_2151, \9574 );
and \U$19816 ( \28924 , RIdf38a40_2021, \9576 );
and \U$19817 ( \28925 , RIdf2d0a0_1889, \9578 );
and \U$19818 ( \28926 , RIdf1d920_1713, \9580 );
and \U$19819 ( \28927 , RIdf01018_1388, \9582 );
and \U$19820 ( \28928 , RIdee7b18_1100, \9584 );
and \U$19821 ( \28929 , RIdedc880_973, \9586 );
and \U$19822 ( \28930 , RIde7dc18_203, \9588 );
or \U$19823 ( \28931 , \28867 , \28868 , \28869 , \28870 , \28871 , \28872 , \28873 , \28874 , \28875 , \28876 , \28877 , \28878 , \28879 , \28880 , \28881 , \28882 , \28883 , \28884 , \28885 , \28886 , \28887 , \28888 , \28889 , \28890 , \28891 , \28892 , \28893 , \28894 , \28895 , \28896 , \28897 , \28898 , \28899 , \28900 , \28901 , \28902 , \28903 , \28904 , \28905 , \28906 , \28907 , \28908 , \28909 , \28910 , \28911 , \28912 , \28913 , \28914 , \28915 , \28916 , \28917 , \28918 , \28919 , \28920 , \28921 , \28922 , \28923 , \28924 , \28925 , \28926 , \28927 , \28928 , \28929 , \28930 );
or \U$19824 ( \28932 , \28866 , \28931 );
_DC g60cd ( \28933_nG60cd , \28932 , \9597 );
and \U$19825 ( \28934 , RIe19dee0_3174, \9059 );
and \U$19826 ( \28935 , RIe19b1e0_3142, \9061 );
and \U$19827 ( \28936 , RIfc67580_6198, \9063 );
and \U$19828 ( \28937 , RIe1984e0_3110, \9065 );
and \U$19829 ( \28938 , RIfccb030_7332, \9067 );
and \U$19830 ( \28939 , RIe1957e0_3078, \9069 );
and \U$19831 ( \28940 , RIe192ae0_3046, \9071 );
and \U$19832 ( \28941 , RIe18fde0_3014, \9073 );
and \U$19833 ( \28942 , RIe18a3e0_2950, \9075 );
and \U$19834 ( \28943 , RIe1876e0_2918, \9077 );
and \U$19835 ( \28944 , RIfc6a550_6232, \9079 );
and \U$19836 ( \28945 , RIe1849e0_2886, \9081 );
and \U$19837 ( \28946 , RIfcaa7e0_6962, \9083 );
and \U$19838 ( \28947 , RIe181ce0_2854, \9085 );
and \U$19839 ( \28948 , RIe17efe0_2822, \9087 );
and \U$19840 ( \28949 , RIe17c2e0_2790, \9089 );
and \U$19841 ( \28950 , RIfc65d98_6181, \9091 );
and \U$19842 ( \28951 , RIfc65690_6176, \9093 );
and \U$19843 ( \28952 , RIe1772b8_2733, \9095 );
and \U$19844 ( \28953 , RIfea0638_8169, \9097 );
and \U$19845 ( \28954 , RIfcca928_7327, \9099 );
and \U$19846 ( \28955 , RIfc607d0_6120, \9101 );
and \U$19847 ( \28956 , RIfc65258_6173, \9103 );
and \U$19848 ( \28957 , RIee3d798_5158, \9105 );
and \U$19849 ( \28958 , RIee3c3e8_5144, \9107 );
and \U$19850 ( \28959 , RIfca9430_6948, \9109 );
and \U$19851 ( \28960 , RIee39f58_5118, \9111 );
and \U$19852 ( \28961 , RIe174018_2697, \9113 );
and \U$19853 ( \28962 , RIfcecf00_7718, \9115 );
and \U$19854 ( \28963 , RIfc650f0_6172, \9117 );
and \U$19855 ( \28964 , RIf16e5a8_5715, \9119 );
and \U$19856 ( \28965 , RIfc43a90_5792, \9121 );
and \U$19857 ( \28966 , RIfc65528_6175, \9123 );
and \U$19858 ( \28967 , RIe224238_4701, \9125 );
and \U$19859 ( \28968 , RIfca9f70_6956, \9127 );
and \U$19860 ( \28969 , RIe221538_4669, \9129 );
and \U$19861 ( \28970 , RIfc6b4c8_6243, \9131 );
and \U$19862 ( \28971 , RIe21e838_4637, \9133 );
and \U$19863 ( \28972 , RIe218e38_4573, \9135 );
and \U$19864 ( \28973 , RIe216138_4541, \9137 );
and \U$19865 ( \28974 , RIfc3fda0_5752, \9139 );
and \U$19866 ( \28975 , RIe213438_4509, \9141 );
and \U$19867 ( \28976 , RIfc61310_6128, \9143 );
and \U$19868 ( \28977 , RIe210738_4477, \9145 );
and \U$19869 ( \28978 , RIfc60c08_6123, \9147 );
and \U$19870 ( \28979 , RIe20da38_4445, \9149 );
and \U$19871 ( \28980 , RIe20ad38_4413, \9151 );
and \U$19872 ( \28981 , RIe208038_4381, \9153 );
and \U$19873 ( \28982 , RIfc66ba8_6191, \9155 );
and \U$19874 ( \28983 , RIfccbcd8_7341, \9157 );
and \U$19875 ( \28984 , RIe202bd8_4321, \9159 );
and \U$19876 ( \28985 , RIe200fb8_4301, \9161 );
and \U$19877 ( \28986 , RIfcadbe8_6999, \9163 );
and \U$19878 ( \28987 , RIfccbe40_7342, \9165 );
and \U$19879 ( \28988 , RIfca7540_6926, \9167 );
and \U$19880 ( \28989 , RIfc6a3e8_6231, \9169 );
and \U$19881 ( \28990 , RIfca6898_6917, \9171 );
and \U$19882 ( \28991 , RIfc73358_6333, \9173 );
and \U$19883 ( \28992 , RIe1fd070_4256, \9175 );
and \U$19884 ( \28993 , RIe1fbe28_4243, \9177 );
and \U$19885 ( \28994 , RIfcc2660_7234, \9179 );
and \U$19886 ( \28995 , RIfc44468_5799, \9181 );
and \U$19887 ( \28996 , RIf15a940_5490, \9183 );
and \U$19888 ( \28997 , RIfca7270_6924, \9185 );
or \U$19889 ( \28998 , \28934 , \28935 , \28936 , \28937 , \28938 , \28939 , \28940 , \28941 , \28942 , \28943 , \28944 , \28945 , \28946 , \28947 , \28948 , \28949 , \28950 , \28951 , \28952 , \28953 , \28954 , \28955 , \28956 , \28957 , \28958 , \28959 , \28960 , \28961 , \28962 , \28963 , \28964 , \28965 , \28966 , \28967 , \28968 , \28969 , \28970 , \28971 , \28972 , \28973 , \28974 , \28975 , \28976 , \28977 , \28978 , \28979 , \28980 , \28981 , \28982 , \28983 , \28984 , \28985 , \28986 , \28987 , \28988 , \28989 , \28990 , \28991 , \28992 , \28993 , \28994 , \28995 , \28996 , \28997 );
and \U$19890 ( \28999 , RIfc5e070_6092, \9188 );
and \U$19891 ( \29000 , RIfc5dda0_6090, \9190 );
and \U$19892 ( \29001 , RIfc7e050_6456, \9192 );
and \U$19893 ( \29002 , RIe1fa7a8_4227, \9194 );
and \U$19894 ( \29003 , RIfc5d968_6087, \9196 );
and \U$19895 ( \29004 , RIfcd9568_7495, \9198 );
and \U$19896 ( \29005 , RIfc8d668_6631, \9200 );
and \U$19897 ( \29006 , RIe1f5d20_4174, \9202 );
and \U$19898 ( \29007 , RIfca4138_6889, \9204 );
and \U$19899 ( \29008 , RIfc8cdf8_6625, \9206 );
and \U$19900 ( \29009 , RIfcc7c28_7295, \9208 );
and \U$19901 ( \29010 , RIe1f39f8_4149, \9210 );
and \U$19902 ( \29011 , RIfc99440_6766, \9212 );
and \U$19903 ( \29012 , RIfcbc3f0_7164, \9214 );
and \U$19904 ( \29013 , RIfc5a128_6047, \9216 );
and \U$19905 ( \29014 , RIe1ee700_4090, \9218 );
and \U$19906 ( \29015 , RIe1ebfa0_4062, \9220 );
and \U$19907 ( \29016 , RIe1e92a0_4030, \9222 );
and \U$19908 ( \29017 , RIe1e65a0_3998, \9224 );
and \U$19909 ( \29018 , RIe1e38a0_3966, \9226 );
and \U$19910 ( \29019 , RIe1e0ba0_3934, \9228 );
and \U$19911 ( \29020 , RIe1ddea0_3902, \9230 );
and \U$19912 ( \29021 , RIe1db1a0_3870, \9232 );
and \U$19913 ( \29022 , RIe1d84a0_3838, \9234 );
and \U$19914 ( \29023 , RIe1d2aa0_3774, \9236 );
and \U$19915 ( \29024 , RIe1cfda0_3742, \9238 );
and \U$19916 ( \29025 , RIe1cd0a0_3710, \9240 );
and \U$19917 ( \29026 , RIe1ca3a0_3678, \9242 );
and \U$19918 ( \29027 , RIe1c76a0_3646, \9244 );
and \U$19919 ( \29028 , RIe1c49a0_3614, \9246 );
and \U$19920 ( \29029 , RIe1c1ca0_3582, \9248 );
and \U$19921 ( \29030 , RIe1befa0_3550, \9250 );
and \U$19922 ( \29031 , RIf14cde0_5334, \9252 );
and \U$19923 ( \29032 , RIf14bb98_5321, \9254 );
and \U$19924 ( \29033 , RIe1b99d8_3489, \9256 );
and \U$19925 ( \29034 , RIe1b7980_3466, \9258 );
and \U$19926 ( \29035 , RIfc4c460_5890, \9260 );
and \U$19927 ( \29036 , RIfc9e738_6825, \9262 );
and \U$19928 ( \29037 , RIe1b5658_3441, \9264 );
and \U$19929 ( \29038 , RIfec54d8_8365, \9266 );
and \U$19930 ( \29039 , RIf149168_5291, \9268 );
and \U$19931 ( \29040 , RIf147f20_5278, \9270 );
and \U$19932 ( \29041 , RIe1b2ac0_3410, \9272 );
and \U$19933 ( \29042 , RIe1b1170_3392, \9274 );
and \U$19934 ( \29043 , RIf1473e0_5270, \9276 );
and \U$19935 ( \29044 , RIf1468a0_5262, \9278 );
and \U$19936 ( \29045 , RIe1acb20_3342, \9280 );
and \U$19937 ( \29046 , RIe1ab338_3325, \9282 );
and \U$19938 ( \29047 , RIe1a92e0_3302, \9284 );
and \U$19939 ( \29048 , RIe1a65e0_3270, \9286 );
and \U$19940 ( \29049 , RIe1a38e0_3238, \9288 );
and \U$19941 ( \29050 , RIe1a0be0_3206, \9290 );
and \U$19942 ( \29051 , RIe18d0e0_2982, \9292 );
and \U$19943 ( \29052 , RIe1795e0_2758, \9294 );
and \U$19944 ( \29053 , RIe226f38_4733, \9296 );
and \U$19945 ( \29054 , RIe21bb38_4605, \9298 );
and \U$19946 ( \29055 , RIe205338_4349, \9300 );
and \U$19947 ( \29056 , RIe1ff398_4281, \9302 );
and \U$19948 ( \29057 , RIe1f8750_4204, \9304 );
and \U$19949 ( \29058 , RIe1f1298_4121, \9306 );
and \U$19950 ( \29059 , RIe1d57a0_3806, \9308 );
and \U$19951 ( \29060 , RIe1bc2a0_3518, \9310 );
and \U$19952 ( \29061 , RIe1af118_3369, \9312 );
and \U$19953 ( \29062 , RIe171750_2668, \9314 );
or \U$19954 ( \29063 , \28999 , \29000 , \29001 , \29002 , \29003 , \29004 , \29005 , \29006 , \29007 , \29008 , \29009 , \29010 , \29011 , \29012 , \29013 , \29014 , \29015 , \29016 , \29017 , \29018 , \29019 , \29020 , \29021 , \29022 , \29023 , \29024 , \29025 , \29026 , \29027 , \29028 , \29029 , \29030 , \29031 , \29032 , \29033 , \29034 , \29035 , \29036 , \29037 , \29038 , \29039 , \29040 , \29041 , \29042 , \29043 , \29044 , \29045 , \29046 , \29047 , \29048 , \29049 , \29050 , \29051 , \29052 , \29053 , \29054 , \29055 , \29056 , \29057 , \29058 , \29059 , \29060 , \29061 , \29062 );
or \U$19955 ( \29064 , \28998 , \29063 );
_DC g6151 ( \29065_nG6151 , \29064 , \9323 );
xor g6152 ( \29066_nG6152 , \28933_nG60cd , \29065_nG6151 );
buf \U$19956 ( \29067 , \29066_nG6152 );
xor \U$19957 ( \29068 , \29067 , \28525 );
not \U$19958 ( \29069 , \28526 );
and \U$19959 ( \29070 , \29068 , \29069 );
and \U$19960 ( \29071 , \10687 , \29070 );
and \U$19961 ( \29072 , \10988 , \28526 );
nor \U$19962 ( \29073 , \29071 , \29072 );
and \U$19963 ( \29074 , \28525 , \27292 );
not \U$19964 ( \29075 , \29074 );
and \U$19965 ( \29076 , \29067 , \29075 );
xnor \U$19966 ( \29077 , \29073 , \29076 );
xor \U$19967 ( \29078 , \28801 , \29077 );
xor \U$19968 ( \29079 , \28792 , \29078 );
and \U$19969 ( \29080 , \28534 , \10983 );
_DC g65c8 ( \29081_nG65c8 , \28932 , \9597 );
_DC g65c9 ( \29082_nG65c9 , \29064 , \9323 );
and g65ca ( \29083_nG65ca , \29081_nG65c8 , \29082_nG65c9 );
buf \U$19970 ( \29084 , \29083_nG65ca );
and \U$19971 ( \29085 , \29084 , \10691 );
nor \U$19972 ( \29086 , \29080 , \29085 );
xnor \U$19973 ( \29087 , \29086 , \10980 );
and \U$19974 ( \29088 , \20544 , \16635 );
and \U$19975 ( \29089 , \21033 , \16301 );
nor \U$19976 ( \29090 , \29088 , \29089 );
xnor \U$19977 ( \29091 , \29090 , \16625 );
xor \U$19978 ( \29092 , \29087 , \29091 );
and \U$19979 ( \29093 , \12448 , \25826 );
and \U$19980 ( \29094 , \12769 , \25264 );
nor \U$19981 ( \29095 , \29093 , \29094 );
xnor \U$19982 ( \29096 , \29095 , \25773 );
xor \U$19983 ( \29097 , \29092 , \29096 );
xor \U$19984 ( \29098 , \29079 , \29097 );
xor \U$19985 ( \29099 , \28778 , \29098 );
and \U$19986 ( \29100 , \28579 , \28583 );
and \U$19987 ( \29101 , \28583 , \28588 );
and \U$19988 ( \29102 , \28579 , \28588 );
or \U$19989 ( \29103 , \29100 , \29101 , \29102 );
and \U$19990 ( \29104 , \22090 , \15336 );
and \U$19991 ( \29105 , \22556 , \14963 );
nor \U$19992 ( \29106 , \29104 , \29105 );
xnor \U$19993 ( \29107 , \29106 , \15342 );
and \U$19994 ( \29108 , \14950 , \22542 );
and \U$19995 ( \29109 , \15321 , \22103 );
nor \U$19996 ( \29110 , \29108 , \29109 );
xnor \U$19997 ( \29111 , \29110 , \22548 );
xor \U$19998 ( \29112 , \29107 , \29111 );
and \U$19999 ( \29113 , \13679 , \24138 );
and \U$20000 ( \29114 , \14024 , \23630 );
nor \U$20001 ( \29115 , \29113 , \29114 );
xnor \U$20002 ( \29116 , \29115 , \24144 );
xor \U$20003 ( \29117 , \29112 , \29116 );
xor \U$20004 ( \29118 , \29103 , \29117 );
and \U$20005 ( \29119 , \26829 , \11574 );
and \U$20006 ( \29120 , \27313 , \11278 );
nor \U$20007 ( \29121 , \29119 , \29120 );
xnor \U$20008 ( \29122 , \29121 , \11580 );
not \U$20009 ( \29123 , \28527 );
and \U$20010 ( \29124 , \29123 , \29076 );
xor \U$20011 ( \29125 , \29122 , \29124 );
and \U$20012 ( \29126 , \28254 , \28258 );
and \U$20013 ( \29127 , \28258 , \28527 );
and \U$20014 ( \29128 , \28254 , \28527 );
or \U$20015 ( \29129 , \29126 , \29127 , \29128 );
xor \U$20016 ( \29130 , \29125 , \29129 );
and \U$20017 ( \29131 , \19032 , \18090 );
and \U$20018 ( \29132 , \19558 , \17655 );
nor \U$20019 ( \29133 , \29131 , \29132 );
xnor \U$20020 ( \29134 , \29133 , \18046 );
xor \U$20021 ( \29135 , \29130 , \29134 );
xor \U$20022 ( \29136 , \29118 , \29135 );
xor \U$20023 ( \29137 , \29099 , \29136 );
xor \U$20024 ( \29138 , \28774 , \29137 );
and \U$20025 ( \29139 , \28220 , \28224 );
and \U$20026 ( \29140 , \28224 , \28229 );
and \U$20027 ( \29141 , \28220 , \28229 );
or \U$20028 ( \29142 , \29139 , \29140 , \29141 );
and \U$20029 ( \29143 , \28246 , \28548 );
and \U$20030 ( \29144 , \28548 , \28590 );
and \U$20031 ( \29145 , \28246 , \28590 );
or \U$20032 ( \29146 , \29143 , \29144 , \29145 );
xor \U$20033 ( \29147 , \29142 , \29146 );
and \U$20034 ( \29148 , \28236 , \28240 );
and \U$20035 ( \29149 , \28240 , \28245 );
and \U$20036 ( \29150 , \28236 , \28245 );
or \U$20037 ( \29151 , \29148 , \29149 , \29150 );
and \U$20038 ( \29152 , \28250 , \28528 );
and \U$20039 ( \29153 , \28528 , \28547 );
and \U$20040 ( \29154 , \28250 , \28547 );
or \U$20041 ( \29155 , \29152 , \29153 , \29154 );
xor \U$20042 ( \29156 , \29151 , \29155 );
and \U$20043 ( \29157 , \28537 , \28541 );
and \U$20044 ( \29158 , \28541 , \28546 );
and \U$20045 ( \29159 , \28537 , \28546 );
or \U$20046 ( \29160 , \29157 , \29158 , \29159 );
and \U$20047 ( \29161 , \28553 , \28557 );
and \U$20048 ( \29162 , \28557 , \28562 );
and \U$20049 ( \29163 , \28553 , \28562 );
or \U$20050 ( \29164 , \29161 , \29162 , \29163 );
xor \U$20051 ( \29165 , \29160 , \29164 );
and \U$20052 ( \29166 , \28567 , \28571 );
and \U$20053 ( \29167 , \28571 , \28576 );
and \U$20054 ( \29168 , \28567 , \28576 );
or \U$20055 ( \29169 , \29166 , \29167 , \29168 );
xor \U$20056 ( \29170 , \29165 , \29169 );
xor \U$20057 ( \29171 , \29156 , \29170 );
xor \U$20058 ( \29172 , \29147 , \29171 );
xor \U$20059 ( \29173 , \29138 , \29172 );
xor \U$20060 ( \29174 , \28770 , \29173 );
and \U$20061 ( \29175 , \28592 , \28596 );
and \U$20062 ( \29176 , \28597 , \28600 );
or \U$20063 ( \29177 , \29175 , \29176 );
xor \U$20064 ( \29178 , \29174 , \29177 );
buf g9bbd ( \29179_nG9bbd , \29178 );
and \U$20065 ( \29180 , \10704 , \29179_nG9bbd );
or \U$20066 ( \29181 , \28766 , \29180 );
xor \U$20067 ( \29182 , \10703 , \29181 );
buf \U$20068 ( \29183 , \29182 );
buf \U$20070 ( \29184 , \29183 );
xor \U$20071 ( \29185 , \28765 , \29184 );
buf \U$20072 ( \29186 , \29185 );
and \U$20073 ( \29187 , \28622 , \28664 );
and \U$20074 ( \29188 , \28622 , \28671 );
and \U$20075 ( \29189 , \28664 , \28671 );
or \U$20076 ( \29190 , \29187 , \29188 , \29189 );
buf \U$20077 ( \29191 , \29190 );
xor \U$20078 ( \29192 , \29186 , \29191 );
and \U$20079 ( \29193 , \28650 , \28655 );
and \U$20080 ( \29194 , \28650 , \28662 );
and \U$20081 ( \29195 , \28655 , \28662 );
or \U$20082 ( \29196 , \29193 , \29194 , \29195 );
buf \U$20083 ( \29197 , \29196 );
and \U$20084 ( \29198 , \28627 , \28641 );
and \U$20085 ( \29199 , \28627 , \28648 );
and \U$20086 ( \29200 , \28641 , \28648 );
or \U$20087 ( \29201 , \29198 , \29199 , \29200 );
buf \U$20088 ( \29202 , \29201 );
and \U$20089 ( \29203 , \28633 , \28639 );
buf \U$20090 ( \29204 , \29203 );
and \U$20091 ( \29205 , \23201 , \13705_nG9bfc );
and \U$20092 ( \29206 , \23198 , \14070_nG9bf9 );
or \U$20093 ( \29207 , \29205 , \29206 );
xor \U$20094 ( \29208 , \23197 , \29207 );
buf \U$20095 ( \29209 , \29208 );
buf \U$20097 ( \29210 , \29209 );
xor \U$20098 ( \29211 , \29204 , \29210 );
and \U$20099 ( \29212 , \21658 , \14984_nG9bf6 );
and \U$20100 ( \29213 , \21655 , \15373_nG9bf3 );
or \U$20101 ( \29214 , \29212 , \29213 );
xor \U$20102 ( \29215 , \21654 , \29214 );
buf \U$20103 ( \29216 , \29215 );
buf \U$20105 ( \29217 , \29216 );
xor \U$20106 ( \29218 , \29211 , \29217 );
buf \U$20107 ( \29219 , \29218 );
xor \U$20108 ( \29220 , \29202 , \29219 );
and \U$20109 ( \29221 , \18702 , \17665_nG9bea );
and \U$20110 ( \29222 , \18699 , \18107_nG9be7 );
or \U$20111 ( \29223 , \29221 , \29222 );
xor \U$20112 ( \29224 , \18698 , \29223 );
buf \U$20113 ( \29225 , \29224 );
buf \U$20115 ( \29226 , \29225 );
xor \U$20116 ( \29227 , \29220 , \29226 );
buf \U$20117 ( \29228 , \29227 );
xor \U$20118 ( \29229 , \29197 , \29228 );
and \U$20119 ( \29230 , \28157 , \28163 );
and \U$20120 ( \29231 , \28157 , \28170 );
and \U$20121 ( \29232 , \28163 , \28170 );
or \U$20122 ( \29233 , \29230 , \29231 , \29232 );
buf \U$20123 ( \29234 , \29233 );
and \U$20124 ( \29235 , \28114 , \28121 );
buf \U$20125 ( \29236 , \29235 );
buf \U$20127 ( \29237 , \29236 );
and \U$20128 ( \29238 , \26431 , \11283_nG9c08 );
and \U$20129 ( \29239 , \26428 , \11598_nG9c05 );
or \U$20130 ( \29240 , \29238 , \29239 );
xor \U$20131 ( \29241 , \26427 , \29240 );
buf \U$20132 ( \29242 , \29241 );
buf \U$20134 ( \29243 , \29242 );
xor \U$20135 ( \29244 , \29237 , \29243 );
buf \U$20136 ( \29245 , \29244 );
and \U$20137 ( \29246 , \28118 , \10694_nG9c0e );
and \U$20138 ( \29247 , \28115 , \10995_nG9c0b );
or \U$20139 ( \29248 , \29246 , \29247 );
xor \U$20140 ( \29249 , \28114 , \29248 );
buf \U$20141 ( \29250 , \29249 );
buf \U$20143 ( \29251 , \29250 );
xor \U$20144 ( \29252 , \29245 , \29251 );
and \U$20145 ( \29253 , \24792 , \12470_nG9c02 );
and \U$20146 ( \29254 , \24789 , \12801_nG9bff );
or \U$20147 ( \29255 , \29253 , \29254 );
xor \U$20148 ( \29256 , \24788 , \29255 );
buf \U$20149 ( \29257 , \29256 );
buf \U$20151 ( \29258 , \29257 );
xor \U$20152 ( \29259 , \29252 , \29258 );
buf \U$20153 ( \29260 , \29259 );
xor \U$20154 ( \29261 , \29234 , \29260 );
and \U$20155 ( \29262 , \20155 , \16315_nG9bf0 );
and \U$20156 ( \29263 , \20152 , \16680_nG9bed );
or \U$20157 ( \29264 , \29262 , \29263 );
xor \U$20158 ( \29265 , \20151 , \29264 );
buf \U$20159 ( \29266 , \29265 );
buf \U$20161 ( \29267 , \29266 );
xor \U$20162 ( \29268 , \29261 , \29267 );
buf \U$20163 ( \29269 , \29268 );
and \U$20164 ( \29270 , \17297 , \19091_nG9be4 );
and \U$20165 ( \29271 , \17294 , \19586_nG9be1 );
or \U$20166 ( \29272 , \29270 , \29271 );
xor \U$20167 ( \29273 , \17293 , \29272 );
buf \U$20168 ( \29274 , \29273 );
buf \U$20170 ( \29275 , \29274 );
xor \U$20171 ( \29276 , \29269 , \29275 );
and \U$20172 ( \29277 , \15940 , \20608_nG9bde );
and \U$20173 ( \29278 , \15937 , \21086_nG9bdb );
or \U$20174 ( \29279 , \29277 , \29278 );
xor \U$20175 ( \29280 , \15936 , \29279 );
buf \U$20176 ( \29281 , \29280 );
buf \U$20178 ( \29282 , \29281 );
xor \U$20179 ( \29283 , \29276 , \29282 );
buf \U$20180 ( \29284 , \29283 );
xor \U$20181 ( \29285 , \29229 , \29284 );
buf \U$20182 ( \29286 , \29285 );
xor \U$20183 ( \29287 , \29192 , \29286 );
buf \U$20184 ( \29288 , \29287 );
xor \U$20185 ( \29289 , \28752 , \29288 );
and \U$20186 ( \29290 , \28135 , \28609 );
and \U$20187 ( \29291 , \28135 , \28615 );
and \U$20188 ( \29292 , \28609 , \28615 );
or \U$20189 ( \29293 , \29290 , \29291 , \29292 );
buf \U$20190 ( \29294 , \29293 );
xor \U$20191 ( \29295 , \29289 , \29294 );
and \U$20192 ( \29296 , \28706 , \29295 );
and \U$20193 ( \29297 , \28696 , \28700 );
and \U$20194 ( \29298 , \28696 , \28705 );
and \U$20195 ( \29299 , \28700 , \28705 );
or \U$20196 ( \29300 , \29297 , \29298 , \29299 );
xor \U$20197 ( \29301 , \29296 , \29300 );
and \U$20198 ( \29302 , RIdec5f18_716, \9059 );
and \U$20199 ( \29303 , RIdec3218_684, \9061 );
and \U$20200 ( \29304 , RIee20350_4825, \9063 );
and \U$20201 ( \29305 , RIdec0518_652, \9065 );
and \U$20202 ( \29306 , RIee1f6a8_4816, \9067 );
and \U$20203 ( \29307 , RIdebd818_620, \9069 );
and \U$20204 ( \29308 , RIdebab18_588, \9071 );
and \U$20205 ( \29309 , RIdeb7e18_556, \9073 );
and \U$20206 ( \29310 , RIfce4da0_7626, \9075 );
and \U$20207 ( \29311 , RIdeb2418_492, \9077 );
and \U$20208 ( \29312 , RIfcea908_7691, \9079 );
and \U$20209 ( \29313 , RIdeaf718_460, \9081 );
and \U$20210 ( \29314 , RIfce20a0_7594, \9083 );
and \U$20211 ( \29315 , RIdeabe60_428, \9085 );
and \U$20212 ( \29316 , RIdea5560_396, \9087 );
and \U$20213 ( \29317 , RIde9ec60_364, \9089 );
and \U$20214 ( \29318 , RIfce6420_7642, \9091 );
and \U$20215 ( \29319 , RIee1c2a0_4779, \9093 );
and \U$20216 ( \29320 , RIfc75950_6360, \9095 );
and \U$20217 ( \29321 , RIee1ad88_4764, \9097 );
and \U$20218 ( \29322 , RIde920f0_302, \9099 );
and \U$20219 ( \29323 , RIfea4148_8211, \9101 );
and \U$20220 ( \29324 , RIfeaa688_8255, \9103 );
and \U$20221 ( \29325 , RIfea3fe0_8210, \9105 );
and \U$20222 ( \29326 , RIde82790_226, \9107 );
and \U$20223 ( \29327 , RIfc6f848_6291, \9109 );
and \U$20224 ( \29328 , RIfc5dc38_6089, \9111 );
and \U$20225 ( \29329 , RIfc76b98_6373, \9113 );
and \U$20226 ( \29330 , RIfcae2f0_7004, \9115 );
and \U$20227 ( \29331 , RIe16c020_2606, \9117 );
and \U$20228 ( \29332 , RIe16a130_2584, \9119 );
and \U$20229 ( \29333 , RIe1687e0_2566, \9121 );
and \U$20230 ( \29334 , RIe165f18_2537, \9123 );
and \U$20231 ( \29335 , RIe163218_2505, \9125 );
and \U$20232 ( \29336 , RIfcadd50_7000, \9127 );
and \U$20233 ( \29337 , RIe160518_2473, \9129 );
and \U$20234 ( \29338 , RIfc55268_5991, \9131 );
and \U$20235 ( \29339 , RIe15d818_2441, \9133 );
and \U$20236 ( \29340 , RIe157e18_2377, \9135 );
and \U$20237 ( \29341 , RIe155118_2345, \9137 );
and \U$20238 ( \29342 , RIfc45548_5811, \9139 );
and \U$20239 ( \29343 , RIe152418_2313, \9141 );
and \U$20240 ( \29344 , RIfc498c8_5859, \9143 );
and \U$20241 ( \29345 , RIe14f718_2281, \9145 );
and \U$20242 ( \29346 , RIfcbda70_7180, \9147 );
and \U$20243 ( \29347 , RIe14ca18_2249, \9149 );
and \U$20244 ( \29348 , RIe149d18_2217, \9151 );
and \U$20245 ( \29349 , RIe147018_2185, \9153 );
and \U$20246 ( \29350 , RIee34828_5056, \9155 );
and \U$20247 ( \29351 , RIee33748_5044, \9157 );
and \U$20248 ( \29352 , RIee32668_5032, \9159 );
and \U$20249 ( \29353 , RIee31588_5020, \9161 );
and \U$20250 ( \29354 , RIe1418e8_2123, \9163 );
and \U$20251 ( \29355 , RIe13f458_2097, \9165 );
and \U$20252 ( \29356 , RIdf3d360_2073, \9167 );
and \U$20253 ( \29357 , RIdf3aed0_2047, \9169 );
and \U$20254 ( \29358 , RIfc526d0_5960, \9171 );
and \U$20255 ( \29359 , RIfc42848_5779, \9173 );
and \U$20256 ( \29360 , RIfcae9f8_7009, \9175 );
and \U$20257 ( \29361 , RIfcb7260_7106, \9177 );
and \U$20258 ( \29362 , RIfea42b0_8212, \9179 );
and \U$20259 ( \29363 , RIdf33ce8_1966, \9181 );
and \U$20260 ( \29364 , RIdf31b28_1942, \9183 );
and \U$20261 ( \29365 , RIdf2fc38_1920, \9185 );
or \U$20262 ( \29366 , \29302 , \29303 , \29304 , \29305 , \29306 , \29307 , \29308 , \29309 , \29310 , \29311 , \29312 , \29313 , \29314 , \29315 , \29316 , \29317 , \29318 , \29319 , \29320 , \29321 , \29322 , \29323 , \29324 , \29325 , \29326 , \29327 , \29328 , \29329 , \29330 , \29331 , \29332 , \29333 , \29334 , \29335 , \29336 , \29337 , \29338 , \29339 , \29340 , \29341 , \29342 , \29343 , \29344 , \29345 , \29346 , \29347 , \29348 , \29349 , \29350 , \29351 , \29352 , \29353 , \29354 , \29355 , \29356 , \29357 , \29358 , \29359 , \29360 , \29361 , \29362 , \29363 , \29364 , \29365 );
and \U$20263 ( \29367 , RIee2c3f8_4962, \9188 );
and \U$20264 ( \29368 , RIfc4cfa0_5898, \9190 );
and \U$20265 ( \29369 , RIfc572c0_6014, \9192 );
and \U$20266 ( \29370 , RIfc4f430_5924, \9194 );
and \U$20267 ( \29371 , RIfea3e78_8209, \9196 );
and \U$20268 ( \29372 , RIdf28a50_1839, \9198 );
and \U$20269 ( \29373 , RIdf26b60_1817, \9200 );
and \U$20270 ( \29374 , RIdf250a8_1798, \9202 );
and \U$20271 ( \29375 , RIfc9b600_6790, \9204 );
and \U$20272 ( \29376 , RIfcb9df8_7137, \9206 );
and \U$20273 ( \29377 , RIdf23320_1777, \9208 );
and \U$20274 ( \29378 , RIfc86318_6549, \9210 );
and \U$20275 ( \29379 , RIfeabfd8_8273, \9212 );
and \U$20276 ( \29380 , RIdf201e8_1742, \9214 );
and \U$20277 ( \29381 , RIdf1b5f8_1688, \9216 );
and \U$20278 ( \29382 , RIdf19ca8_1670, \9218 );
and \U$20279 ( \29383 , RIdf17ae8_1646, \9220 );
and \U$20280 ( \29384 , RIdf14de8_1614, \9222 );
and \U$20281 ( \29385 , RIdf120e8_1582, \9224 );
and \U$20282 ( \29386 , RIdf0f3e8_1550, \9226 );
and \U$20283 ( \29387 , RIdf0c6e8_1518, \9228 );
and \U$20284 ( \29388 , RIdf099e8_1486, \9230 );
and \U$20285 ( \29389 , RIdf06ce8_1454, \9232 );
and \U$20286 ( \29390 , RIdf03fe8_1422, \9234 );
and \U$20287 ( \29391 , RIdefe5e8_1358, \9236 );
and \U$20288 ( \29392 , RIdefb8e8_1326, \9238 );
and \U$20289 ( \29393 , RIdef8be8_1294, \9240 );
and \U$20290 ( \29394 , RIdef5ee8_1262, \9242 );
and \U$20291 ( \29395 , RIdef31e8_1230, \9244 );
and \U$20292 ( \29396 , RIdef04e8_1198, \9246 );
and \U$20293 ( \29397 , RIdeed7e8_1166, \9248 );
and \U$20294 ( \29398 , RIdeeaae8_1134, \9250 );
and \U$20295 ( \29399 , RIfc89018_6581, \9252 );
and \U$20296 ( \29400 , RIfcc54c8_7267, \9254 );
and \U$20297 ( \29401 , RIfc89180_6582, \9256 );
and \U$20298 ( \29402 , RIfc4b380_5878, \9258 );
and \U$20299 ( \29403 , RIdee53b8_1072, \9260 );
and \U$20300 ( \29404 , RIdee34c8_1050, \9262 );
and \U$20301 ( \29405 , RIfea3d10_8208, \9264 );
and \U$20302 ( \29406 , RIdedf148_1002, \9266 );
and \U$20303 ( \29407 , RIfcae188_7003, \9268 );
and \U$20304 ( \29408 , RIfc4b0b0_5876, \9270 );
and \U$20305 ( \29409 , RIfc74870_6348, \9272 );
and \U$20306 ( \29410 , RIfce4968_7623, \9274 );
and \U$20307 ( \29411 , RIdeda288_946, \9276 );
and \U$20308 ( \29412 , RIded7c90_919, \9278 );
and \U$20309 ( \29413 , RIded5da0_897, \9280 );
and \U$20310 ( \29414 , RIded3640_869, \9282 );
and \U$20311 ( \29415 , RIded1318_844, \9284 );
and \U$20312 ( \29416 , RIdece618_812, \9286 );
and \U$20313 ( \29417 , RIdecb918_780, \9288 );
and \U$20314 ( \29418 , RIdec8c18_748, \9290 );
and \U$20315 ( \29419 , RIdeb5118_524, \9292 );
and \U$20316 ( \29420 , RIde98360_332, \9294 );
and \U$20317 ( \29421 , RIe16ed20_2638, \9296 );
and \U$20318 ( \29422 , RIe15ab18_2409, \9298 );
and \U$20319 ( \29423 , RIe144318_2153, \9300 );
and \U$20320 ( \29424 , RIdf38d10_2023, \9302 );
and \U$20321 ( \29425 , RIdf2d370_1891, \9304 );
and \U$20322 ( \29426 , RIdf1dbf0_1715, \9306 );
and \U$20323 ( \29427 , RIdf012e8_1390, \9308 );
and \U$20324 ( \29428 , RIdee7de8_1102, \9310 );
and \U$20325 ( \29429 , RIdedcb50_975, \9312 );
and \U$20326 ( \29430 , RIde7e2a8_205, \9314 );
or \U$20327 ( \29431 , \29367 , \29368 , \29369 , \29370 , \29371 , \29372 , \29373 , \29374 , \29375 , \29376 , \29377 , \29378 , \29379 , \29380 , \29381 , \29382 , \29383 , \29384 , \29385 , \29386 , \29387 , \29388 , \29389 , \29390 , \29391 , \29392 , \29393 , \29394 , \29395 , \29396 , \29397 , \29398 , \29399 , \29400 , \29401 , \29402 , \29403 , \29404 , \29405 , \29406 , \29407 , \29408 , \29409 , \29410 , \29411 , \29412 , \29413 , \29414 , \29415 , \29416 , \29417 , \29418 , \29419 , \29420 , \29421 , \29422 , \29423 , \29424 , \29425 , \29426 , \29427 , \29428 , \29429 , \29430 );
or \U$20328 ( \29432 , \29366 , \29431 );
_DC g233f ( \29433_nG233f , \29432 , \9323 );
buf \U$20329 ( \29434 , \29433_nG233f );
and \U$20330 ( \29435 , RIe19e1b0_3176, \9333 );
and \U$20331 ( \29436 , RIe19b4b0_3144, \9335 );
and \U$20332 ( \29437 , RIfc9cf50_6808, \9337 );
and \U$20333 ( \29438 , RIe1987b0_3112, \9339 );
and \U$20334 ( \29439 , RIfc87290_6560, \9341 );
and \U$20335 ( \29440 , RIe195ab0_3080, \9343 );
and \U$20336 ( \29441 , RIe192db0_3048, \9345 );
and \U$20337 ( \29442 , RIe1900b0_3016, \9347 );
and \U$20338 ( \29443 , RIe18a6b0_2952, \9349 );
and \U$20339 ( \29444 , RIe1879b0_2920, \9351 );
and \U$20340 ( \29445 , RIfc842c0_6526, \9353 );
and \U$20341 ( \29446 , RIe184cb0_2888, \9355 );
and \U$20342 ( \29447 , RIfc83a50_6520, \9357 );
and \U$20343 ( \29448 , RIe181fb0_2856, \9359 );
and \U$20344 ( \29449 , RIe17f2b0_2824, \9361 );
and \U$20345 ( \29450 , RIe17c5b0_2792, \9363 );
and \U$20346 ( \29451 , RIfc9d0b8_6809, \9365 );
and \U$20347 ( \29452 , RIfc9e030_6820, \9367 );
and \U$20348 ( \29453 , RIe177420_2734, \9369 );
and \U$20349 ( \29454 , RIe176340_2722, \9371 );
and \U$20350 ( \29455 , RIfc4f700_5926, \9373 );
and \U$20351 ( \29456 , RIfcc4820_7258, \9375 );
and \U$20352 ( \29457 , RIfc4fb38_5929, \9377 );
and \U$20353 ( \29458 , RIfce8040_7662, \9379 );
and \U$20354 ( \29459 , RIee3c6b8_5146, \9381 );
and \U$20355 ( \29460 , RIee3b308_5132, \9383 );
and \U$20356 ( \29461 , RIfc812f0_6492, \9385 );
and \U$20357 ( \29462 , RIe174180_2698, \9387 );
and \U$20358 ( \29463 , RIfcd3028_7423, \9389 );
and \U$20359 ( \29464 , RIfc7f400_6470, \9391 );
and \U$20360 ( \29465 , RIfc46a60_5826, \9393 );
and \U$20361 ( \29466 , RIfc472d0_5832, \9395 );
and \U$20362 ( \29467 , RIf16cc58_5697, \9397 );
and \U$20363 ( \29468 , RIe224508_4703, \9399 );
and \U$20364 ( \29469 , RIfc7d3a8_6447, \9401 );
and \U$20365 ( \29470 , RIe221808_4671, \9403 );
and \U$20366 ( \29471 , RIfc97c58_6749, \9405 );
and \U$20367 ( \29472 , RIe21eb08_4639, \9407 );
and \U$20368 ( \29473 , RIe219108_4575, \9409 );
and \U$20369 ( \29474 , RIe216408_4543, \9411 );
and \U$20370 ( \29475 , RIfcdbe30_7524, \9413 );
and \U$20371 ( \29476 , RIe213708_4511, \9415 );
and \U$20372 ( \29477 , RIf169580_5658, \9417 );
and \U$20373 ( \29478 , RIe210a08_4479, \9419 );
and \U$20374 ( \29479 , RIfca4570_6892, \9421 );
and \U$20375 ( \29480 , RIe20dd08_4447, \9423 );
and \U$20376 ( \29481 , RIe20b008_4415, \9425 );
and \U$20377 ( \29482 , RIe208308_4383, \9427 );
and \U$20378 ( \29483 , RIfc7b080_6422, \9429 );
and \U$20379 ( \29484 , RIfc59cf0_6044, \9431 );
and \U$20380 ( \29485 , RIfea9b48_8247, \9433 );
and \U$20381 ( \29486 , RIfea4418_8213, \9435 );
and \U$20382 ( \29487 , RIfc79cd0_6408, \9437 );
and \U$20383 ( \29488 , RIfcd19a8_7407, \9439 );
and \U$20384 ( \29489 , RIfcc81c8_7299, \9441 );
and \U$20385 ( \29490 , RIf162230_5576, \9443 );
and \U$20386 ( \29491 , RIf160778_5557, \9445 );
and \U$20387 ( \29492 , RIf15e888_5535, \9447 );
and \U$20388 ( \29493 , RIfea4580_8214, \9449 );
and \U$20389 ( \29494 , RIfea46e8_8215, \9451 );
and \U$20390 ( \29495 , RIfc77f48_6387, \9453 );
and \U$20391 ( \29496 , RIfc41fd8_5773, \9455 );
and \U$20392 ( \29497 , RIf15aaa8_5491, \9457 );
and \U$20393 ( \29498 , RIfc7c430_6436, \9459 );
or \U$20394 ( \29499 , \29435 , \29436 , \29437 , \29438 , \29439 , \29440 , \29441 , \29442 , \29443 , \29444 , \29445 , \29446 , \29447 , \29448 , \29449 , \29450 , \29451 , \29452 , \29453 , \29454 , \29455 , \29456 , \29457 , \29458 , \29459 , \29460 , \29461 , \29462 , \29463 , \29464 , \29465 , \29466 , \29467 , \29468 , \29469 , \29470 , \29471 , \29472 , \29473 , \29474 , \29475 , \29476 , \29477 , \29478 , \29479 , \29480 , \29481 , \29482 , \29483 , \29484 , \29485 , \29486 , \29487 , \29488 , \29489 , \29490 , \29491 , \29492 , \29493 , \29494 , \29495 , \29496 , \29497 , \29498 );
and \U$20395 ( \29500 , RIf159158_5473, \9462 );
and \U$20396 ( \29501 , RIf157f10_5460, \9464 );
and \U$20397 ( \29502 , RIfcae890_7008, \9466 );
and \U$20398 ( \29503 , RIe1faa78_4229, \9468 );
and \U$20399 ( \29504 , RIfc4a840_5870, \9470 );
and \U$20400 ( \29505 , RIfc4ed28_5919, \9472 );
and \U$20401 ( \29506 , RIfce0e58_7581, \9474 );
and \U$20402 ( \29507 , RIe1f5ff0_4176, \9476 );
and \U$20403 ( \29508 , RIf153758_5409, \9478 );
and \U$20404 ( \29509 , RIf151f70_5392, \9480 );
and \U$20405 ( \29510 , RIfccb468_7335, \9482 );
and \U$20406 ( \29511 , RIe1f3cc8_4151, \9484 );
and \U$20407 ( \29512 , RIfc68ed0_6216, \9486 );
and \U$20408 ( \29513 , RIfc6d250_6264, \9488 );
and \U$20409 ( \29514 , RIfca9ca0_6954, \9490 );
and \U$20410 ( \29515 , RIe1ee9d0_4092, \9492 );
and \U$20411 ( \29516 , RIe1ec270_4064, \9494 );
and \U$20412 ( \29517 , RIe1e9570_4032, \9496 );
and \U$20413 ( \29518 , RIe1e6870_4000, \9498 );
and \U$20414 ( \29519 , RIe1e3b70_3968, \9500 );
and \U$20415 ( \29520 , RIe1e0e70_3936, \9502 );
and \U$20416 ( \29521 , RIe1de170_3904, \9504 );
and \U$20417 ( \29522 , RIe1db470_3872, \9506 );
and \U$20418 ( \29523 , RIe1d8770_3840, \9508 );
and \U$20419 ( \29524 , RIe1d2d70_3776, \9510 );
and \U$20420 ( \29525 , RIe1d0070_3744, \9512 );
and \U$20421 ( \29526 , RIe1cd370_3712, \9514 );
and \U$20422 ( \29527 , RIe1ca670_3680, \9516 );
and \U$20423 ( \29528 , RIe1c7970_3648, \9518 );
and \U$20424 ( \29529 , RIe1c4c70_3616, \9520 );
and \U$20425 ( \29530 , RIe1c1f70_3584, \9522 );
and \U$20426 ( \29531 , RIe1bf270_3552, \9524 );
and \U$20427 ( \29532 , RIfc784e8_6391, \9526 );
and \U$20428 ( \29533 , RIfcbef88_7195, \9528 );
and \U$20429 ( \29534 , RIe1b9ca8_3491, \9530 );
and \U$20430 ( \29535 , RIe1b7ae8_3467, \9532 );
and \U$20431 ( \29536 , RIfcc20c0_7230, \9534 );
and \U$20432 ( \29537 , RIfca6190_6912, \9536 );
and \U$20433 ( \29538 , RIe1b5928_3443, \9538 );
and \U$20434 ( \29539 , RIe1b4410_3428, \9540 );
and \U$20435 ( \29540 , RIfcb81d8_7117, \9542 );
and \U$20436 ( \29541 , RIfcc5090_7264, \9544 );
and \U$20437 ( \29542 , RIe1b2d90_3412, \9546 );
and \U$20438 ( \29543 , RIe1b1440_3394, \9548 );
and \U$20439 ( \29544 , RIfcd5350_7448, \9550 );
and \U$20440 ( \29545 , RIfcb9588_7131, \9552 );
and \U$20441 ( \29546 , RIe1acc88_3343, \9554 );
and \U$20442 ( \29547 , RIe1ab4a0_3326, \9556 );
and \U$20443 ( \29548 , RIe1a95b0_3304, \9558 );
and \U$20444 ( \29549 , RIe1a68b0_3272, \9560 );
and \U$20445 ( \29550 , RIe1a3bb0_3240, \9562 );
and \U$20446 ( \29551 , RIe1a0eb0_3208, \9564 );
and \U$20447 ( \29552 , RIe18d3b0_2984, \9566 );
and \U$20448 ( \29553 , RIe1798b0_2760, \9568 );
and \U$20449 ( \29554 , RIe227208_4735, \9570 );
and \U$20450 ( \29555 , RIe21be08_4607, \9572 );
and \U$20451 ( \29556 , RIe205608_4351, \9574 );
and \U$20452 ( \29557 , RIe1ff668_4283, \9576 );
and \U$20453 ( \29558 , RIe1f8a20_4206, \9578 );
and \U$20454 ( \29559 , RIe1f1568_4123, \9580 );
and \U$20455 ( \29560 , RIe1d5a70_3808, \9582 );
and \U$20456 ( \29561 , RIe1bc570_3520, \9584 );
and \U$20457 ( \29562 , RIe1af3e8_3371, \9586 );
and \U$20458 ( \29563 , RIe171a20_2670, \9588 );
or \U$20459 ( \29564 , \29500 , \29501 , \29502 , \29503 , \29504 , \29505 , \29506 , \29507 , \29508 , \29509 , \29510 , \29511 , \29512 , \29513 , \29514 , \29515 , \29516 , \29517 , \29518 , \29519 , \29520 , \29521 , \29522 , \29523 , \29524 , \29525 , \29526 , \29527 , \29528 , \29529 , \29530 , \29531 , \29532 , \29533 , \29534 , \29535 , \29536 , \29537 , \29538 , \29539 , \29540 , \29541 , \29542 , \29543 , \29544 , \29545 , \29546 , \29547 , \29548 , \29549 , \29550 , \29551 , \29552 , \29553 , \29554 , \29555 , \29556 , \29557 , \29558 , \29559 , \29560 , \29561 , \29562 , \29563 );
or \U$20460 ( \29565 , \29499 , \29564 );
_DC g346c ( \29566_nG346c , \29565 , \9597 );
buf \U$20461 ( \29567 , \29566_nG346c );
xor \U$20462 ( \29568 , \29434 , \29567 );
and \U$20463 ( \29569 , RIdec5db0_715, \9059 );
and \U$20464 ( \29570 , RIdec30b0_683, \9061 );
and \U$20465 ( \29571 , RIee201e8_4824, \9063 );
and \U$20466 ( \29572 , RIdec03b0_651, \9065 );
and \U$20467 ( \29573 , RIfcaf538_7017, \9067 );
and \U$20468 ( \29574 , RIdebd6b0_619, \9069 );
and \U$20469 ( \29575 , RIdeba9b0_587, \9071 );
and \U$20470 ( \29576 , RIdeb7cb0_555, \9073 );
and \U$20471 ( \29577 , RIfc40fe8_5765, \9075 );
and \U$20472 ( \29578 , RIdeb22b0_491, \9077 );
and \U$20473 ( \29579 , RIfcd08c8_7395, \9079 );
and \U$20474 ( \29580 , RIdeaf5b0_459, \9081 );
and \U$20475 ( \29581 , RIee1dd58_4798, \9083 );
and \U$20476 ( \29582 , RIdeabb18_427, \9085 );
and \U$20477 ( \29583 , RIdea5218_395, \9087 );
and \U$20478 ( \29584 , RIde9e918_363, \9089 );
and \U$20479 ( \29585 , RIee1d218_4790, \9091 );
and \U$20480 ( \29586 , RIfcedd10_7728, \9093 );
and \U$20481 ( \29587 , RIfce62b8_7641, \9095 );
and \U$20482 ( \29588 , RIfcc92a8_7311, \9097 );
and \U$20483 ( \29589 , RIde91da8_301, \9099 );
and \U$20484 ( \29590 , RIde8e928_285, \9101 );
and \U$20485 ( \29591 , RIde8a788_265, \9103 );
and \U$20486 ( \29592 , RIde865e8_245, \9105 );
and \U$20487 ( \29593 , RIde82448_225, \9107 );
and \U$20488 ( \29594 , RIfea1448_8179, \9109 );
and \U$20489 ( \29595 , RIfc750e0_6354, \9111 );
and \U$20490 ( \29596 , RIfcc19b8_7225, \9113 );
and \U$20491 ( \29597 , RIfced8d8_7725, \9115 );
and \U$20492 ( \29598 , RIfec5eb0_8372, \9117 );
and \U$20493 ( \29599 , RIe169fc8_2583, \9119 );
and \U$20494 ( \29600 , RIe168678_2565, \9121 );
and \U$20495 ( \29601 , RIe165db0_2536, \9123 );
and \U$20496 ( \29602 , RIe1630b0_2504, \9125 );
and \U$20497 ( \29603 , RIfccfc20_7386, \9127 );
and \U$20498 ( \29604 , RIe1603b0_2472, \9129 );
and \U$20499 ( \29605 , RIee365b0_5077, \9131 );
and \U$20500 ( \29606 , RIe15d6b0_2440, \9133 );
and \U$20501 ( \29607 , RIe157cb0_2376, \9135 );
and \U$20502 ( \29608 , RIe154fb0_2344, \9137 );
and \U$20503 ( \29609 , RIfea1718_8181, \9139 );
and \U$20504 ( \29610 , RIe1522b0_2312, \9141 );
and \U$20505 ( \29611 , RIee35200_5063, \9143 );
and \U$20506 ( \29612 , RIe14f5b0_2280, \9145 );
and \U$20507 ( \29613 , RIfcb0348_7027, \9147 );
and \U$20508 ( \29614 , RIe14c8b0_2248, \9149 );
and \U$20509 ( \29615 , RIe149bb0_2216, \9151 );
and \U$20510 ( \29616 , RIe146eb0_2184, \9153 );
and \U$20511 ( \29617 , RIfc73790_6336, \9155 );
and \U$20512 ( \29618 , RIfcdf238_7561, \9157 );
and \U$20513 ( \29619 , RIee32500_5031, \9159 );
and \U$20514 ( \29620 , RIfc94f58_6717, \9161 );
and \U$20515 ( \29621 , RIe141780_2122, \9163 );
and \U$20516 ( \29622 , RIe13f2f0_2096, \9165 );
and \U$20517 ( \29623 , RIfec5be0_8370, \9167 );
and \U$20518 ( \29624 , RIdf3ad68_2046, \9169 );
and \U$20519 ( \29625 , RIfea15b0_8180, \9171 );
and \U$20520 ( \29626 , RIfc5fb28_6111, \9173 );
and \U$20521 ( \29627 , RIfcae728_7007, \9175 );
and \U$20522 ( \29628 , RIfc74438_6345, \9177 );
and \U$20523 ( \29629 , RIdf36178_1992, \9179 );
and \U$20524 ( \29630 , RIdf33b80_1965, \9181 );
and \U$20525 ( \29631 , RIdf319c0_1941, \9183 );
and \U$20526 ( \29632 , RIdf2fad0_1919, \9185 );
or \U$20527 ( \29633 , \29569 , \29570 , \29571 , \29572 , \29573 , \29574 , \29575 , \29576 , \29577 , \29578 , \29579 , \29580 , \29581 , \29582 , \29583 , \29584 , \29585 , \29586 , \29587 , \29588 , \29589 , \29590 , \29591 , \29592 , \29593 , \29594 , \29595 , \29596 , \29597 , \29598 , \29599 , \29600 , \29601 , \29602 , \29603 , \29604 , \29605 , \29606 , \29607 , \29608 , \29609 , \29610 , \29611 , \29612 , \29613 , \29614 , \29615 , \29616 , \29617 , \29618 , \29619 , \29620 , \29621 , \29622 , \29623 , \29624 , \29625 , \29626 , \29627 , \29628 , \29629 , \29630 , \29631 , \29632 );
and \U$20528 ( \29634 , RIee2c290_4961, \9188 );
and \U$20529 ( \29635 , RIee2a940_4943, \9190 );
and \U$20530 ( \29636 , RIfc70658_6301, \9192 );
and \U$20531 ( \29637 , RIfc704f0_6300, \9194 );
and \U$20532 ( \29638 , RIdf2aaa8_1862, \9196 );
and \U$20533 ( \29639 , RIdf288e8_1838, \9198 );
and \U$20534 ( \29640 , RIdf269f8_1816, \9200 );
and \U$20535 ( \29641 , RIdf24f40_1797, \9202 );
and \U$20536 ( \29642 , RIfc64b50_6168, \9204 );
and \U$20537 ( \29643 , RIfccaa90_7328, \9206 );
and \U$20538 ( \29644 , RIdf231b8_1776, \9208 );
and \U$20539 ( \29645 , RIfcad4e0_6994, \9210 );
and \U$20540 ( \29646 , RIdf21ca0_1761, \9212 );
and \U$20541 ( \29647 , RIfeaad90_8260, \9214 );
and \U$20542 ( \29648 , RIdf1b490_1687, \9216 );
and \U$20543 ( \29649 , RIdf19b40_1669, \9218 );
and \U$20544 ( \29650 , RIdf17980_1645, \9220 );
and \U$20545 ( \29651 , RIdf14c80_1613, \9222 );
and \U$20546 ( \29652 , RIdf11f80_1581, \9224 );
and \U$20547 ( \29653 , RIdf0f280_1549, \9226 );
and \U$20548 ( \29654 , RIdf0c580_1517, \9228 );
and \U$20549 ( \29655 , RIdf09880_1485, \9230 );
and \U$20550 ( \29656 , RIdf06b80_1453, \9232 );
and \U$20551 ( \29657 , RIdf03e80_1421, \9234 );
and \U$20552 ( \29658 , RIdefe480_1357, \9236 );
and \U$20553 ( \29659 , RIdefb780_1325, \9238 );
and \U$20554 ( \29660 , RIdef8a80_1293, \9240 );
and \U$20555 ( \29661 , RIdef5d80_1261, \9242 );
and \U$20556 ( \29662 , RIdef3080_1229, \9244 );
and \U$20557 ( \29663 , RIdef0380_1197, \9246 );
and \U$20558 ( \29664 , RIdeed680_1165, \9248 );
and \U$20559 ( \29665 , RIdeea980_1133, \9250 );
and \U$20560 ( \29666 , RIfc595e8_6039, \9252 );
and \U$20561 ( \29667 , RIfcac568_6983, \9254 );
and \U$20562 ( \29668 , RIfcccf20_7354, \9256 );
and \U$20563 ( \29669 , RIfccd358_7357, \9258 );
and \U$20564 ( \29670 , RIdee5250_1071, \9260 );
and \U$20565 ( \29671 , RIfea7f28_8227, \9262 );
and \U$20566 ( \29672 , RIdee11a0_1025, \9264 );
and \U$20567 ( \29673 , RIfea12e0_8178, \9266 );
and \U$20568 ( \29674 , RIfc679b8_6201, \9268 );
and \U$20569 ( \29675 , RIee22510_4849, \9270 );
and \U$20570 ( \29676 , RIfc6dd90_6272, \9272 );
and \U$20571 ( \29677 , RIfc6cb48_6259, \9274 );
and \U$20572 ( \29678 , RIdeda120_945, \9276 );
and \U$20573 ( \29679 , RIded7b28_918, \9278 );
and \U$20574 ( \29680 , RIded5c38_896, \9280 );
and \U$20575 ( \29681 , RIfec5d48_8371, \9282 );
and \U$20576 ( \29682 , RIded11b0_843, \9284 );
and \U$20577 ( \29683 , RIdece4b0_811, \9286 );
and \U$20578 ( \29684 , RIdecb7b0_779, \9288 );
and \U$20579 ( \29685 , RIdec8ab0_747, \9290 );
and \U$20580 ( \29686 , RIdeb4fb0_523, \9292 );
and \U$20581 ( \29687 , RIde98018_331, \9294 );
and \U$20582 ( \29688 , RIe16ebb8_2637, \9296 );
and \U$20583 ( \29689 , RIe15a9b0_2408, \9298 );
and \U$20584 ( \29690 , RIe1441b0_2152, \9300 );
and \U$20585 ( \29691 , RIdf38ba8_2022, \9302 );
and \U$20586 ( \29692 , RIdf2d208_1890, \9304 );
and \U$20587 ( \29693 , RIdf1da88_1714, \9306 );
and \U$20588 ( \29694 , RIdf01180_1389, \9308 );
and \U$20589 ( \29695 , RIdee7c80_1101, \9310 );
and \U$20590 ( \29696 , RIdedc9e8_974, \9312 );
and \U$20591 ( \29697 , RIde7df60_204, \9314 );
or \U$20592 ( \29698 , \29634 , \29635 , \29636 , \29637 , \29638 , \29639 , \29640 , \29641 , \29642 , \29643 , \29644 , \29645 , \29646 , \29647 , \29648 , \29649 , \29650 , \29651 , \29652 , \29653 , \29654 , \29655 , \29656 , \29657 , \29658 , \29659 , \29660 , \29661 , \29662 , \29663 , \29664 , \29665 , \29666 , \29667 , \29668 , \29669 , \29670 , \29671 , \29672 , \29673 , \29674 , \29675 , \29676 , \29677 , \29678 , \29679 , \29680 , \29681 , \29682 , \29683 , \29684 , \29685 , \29686 , \29687 , \29688 , \29689 , \29690 , \29691 , \29692 , \29693 , \29694 , \29695 , \29696 , \29697 );
or \U$20593 ( \29699 , \29633 , \29698 );
_DC g23c4 ( \29700_nG23c4 , \29699 , \9323 );
buf \U$20594 ( \29701 , \29700_nG23c4 );
and \U$20595 ( \29702 , RIe19e048_3175, \9333 );
and \U$20596 ( \29703 , RIe19b348_3143, \9335 );
and \U$20597 ( \29704 , RIfcc3ce0_7250, \9337 );
and \U$20598 ( \29705 , RIe198648_3111, \9339 );
and \U$20599 ( \29706 , RIfc7efc8_6467, \9341 );
and \U$20600 ( \29707 , RIe195948_3079, \9343 );
and \U$20601 ( \29708 , RIe192c48_3047, \9345 );
and \U$20602 ( \29709 , RIe18ff48_3015, \9347 );
and \U$20603 ( \29710 , RIe18a548_2951, \9349 );
and \U$20604 ( \29711 , RIe187848_2919, \9351 );
and \U$20605 ( \29712 , RIfc46790_5824, \9353 );
and \U$20606 ( \29713 , RIe184b48_2887, \9355 );
and \U$20607 ( \29714 , RIfc98d38_6761, \9357 );
and \U$20608 ( \29715 , RIe181e48_2855, \9359 );
and \U$20609 ( \29716 , RIe17f148_2823, \9361 );
and \U$20610 ( \29717 , RIe17c448_2791, \9363 );
and \U$20611 ( \29718 , RIfcb5d48_7091, \9365 );
and \U$20612 ( \29719 , RIfc995a8_6767, \9367 );
and \U$20613 ( \29720 , RIfc9a3b8_6777, \9369 );
and \U$20614 ( \29721 , RIe1761d8_2721, \9371 );
and \U$20615 ( \29722 , RIfc54188_5979, \9373 );
and \U$20616 ( \29723 , RIfcd2bf0_7420, \9375 );
and \U$20617 ( \29724 , RIfc8b778_6609, \9377 );
and \U$20618 ( \29725 , RIfc7dee8_6455, \9379 );
and \U$20619 ( \29726 , RIee3c550_5145, \9381 );
and \U$20620 ( \29727 , RIfc8c420_6618, \9383 );
and \U$20621 ( \29728 , RIee3a0c0_5119, \9385 );
and \U$20622 ( \29729 , RIfeaba38_8269, \9387 );
and \U$20623 ( \29730 , RIfc46628_5823, \9389 );
and \U$20624 ( \29731 , RIfcbc288_7163, \9391 );
and \U$20625 ( \29732 , RIf16e710_5716, \9393 );
and \U$20626 ( \29733 , RIfc8fdc8_6659, \9395 );
and \U$20627 ( \29734 , RIfc48c20_5850, \9397 );
and \U$20628 ( \29735 , RIe2243a0_4702, \9399 );
and \U$20629 ( \29736 , RIfca0358_6845, \9401 );
and \U$20630 ( \29737 , RIe2216a0_4670, \9403 );
and \U$20631 ( \29738 , RIfc9a688_6779, \9405 );
and \U$20632 ( \29739 , RIe21e9a0_4638, \9407 );
and \U$20633 ( \29740 , RIe218fa0_4574, \9409 );
and \U$20634 ( \29741 , RIe2162a0_4542, \9411 );
and \U$20635 ( \29742 , RIfc456b0_5812, \9413 );
and \U$20636 ( \29743 , RIe2135a0_4510, \9415 );
and \U$20637 ( \29744 , RIf169418_5657, \9417 );
and \U$20638 ( \29745 , RIe2108a0_4478, \9419 );
and \U$20639 ( \29746 , RIfc8bfe8_6615, \9421 );
and \U$20640 ( \29747 , RIe20dba0_4446, \9423 );
and \U$20641 ( \29748 , RIe20aea0_4414, \9425 );
and \U$20642 ( \29749 , RIe2081a0_4382, \9427 );
and \U$20643 ( \29750 , RIfc8c9c0_6622, \9429 );
and \U$20644 ( \29751 , RIfc7f568_6471, \9431 );
and \U$20645 ( \29752 , RIe202d40_4322, \9433 );
and \U$20646 ( \29753 , RIe201120_4302, \9435 );
and \U$20647 ( \29754 , RIfce2910_7600, \9437 );
and \U$20648 ( \29755 , RIfc487e8_5847, \9439 );
and \U$20649 ( \29756 , RIfc46d30_5828, \9441 );
and \U$20650 ( \29757 , RIfc992d8_6765, \9443 );
and \U$20651 ( \29758 , RIfca2680_6870, \9445 );
and \U$20652 ( \29759 , RIfc44a08_5803, \9447 );
and \U$20653 ( \29760 , RIe1fd1d8_4257, \9449 );
and \U$20654 ( \29761 , RIe1fbf90_4244, \9451 );
and \U$20655 ( \29762 , RIfc580d0_6024, \9453 );
and \U$20656 ( \29763 , RIfcbdbd8_7181, \9455 );
and \U$20657 ( \29764 , RIfc8dd70_6636, \9457 );
and \U$20658 ( \29765 , RIfce01b0_7572, \9459 );
or \U$20659 ( \29766 , \29702 , \29703 , \29704 , \29705 , \29706 , \29707 , \29708 , \29709 , \29710 , \29711 , \29712 , \29713 , \29714 , \29715 , \29716 , \29717 , \29718 , \29719 , \29720 , \29721 , \29722 , \29723 , \29724 , \29725 , \29726 , \29727 , \29728 , \29729 , \29730 , \29731 , \29732 , \29733 , \29734 , \29735 , \29736 , \29737 , \29738 , \29739 , \29740 , \29741 , \29742 , \29743 , \29744 , \29745 , \29746 , \29747 , \29748 , \29749 , \29750 , \29751 , \29752 , \29753 , \29754 , \29755 , \29756 , \29757 , \29758 , \29759 , \29760 , \29761 , \29762 , \29763 , \29764 , \29765 );
and \U$20660 ( \29767 , RIfc7bbc0_6430, \9462 );
and \U$20661 ( \29768 , RIfc90368_6663, \9464 );
and \U$20662 ( \29769 , RIfc7b8f0_6428, \9466 );
and \U$20663 ( \29770 , RIe1fa910_4228, \9468 );
and \U$20664 ( \29771 , RIfcd8b90_7488, \9470 );
and \U$20665 ( \29772 , RIfc43ec8_5795, \9472 );
and \U$20666 ( \29773 , RIfc7b788_6427, \9474 );
and \U$20667 ( \29774 , RIe1f5e88_4175, \9476 );
and \U$20668 ( \29775 , RIfc7b350_6424, \9478 );
and \U$20669 ( \29776 , RIfc90d40_6670, \9480 );
and \U$20670 ( \29777 , RIfca3490_6880, \9482 );
and \U$20671 ( \29778 , RIe1f3b60_4150, \9484 );
and \U$20672 ( \29779 , RIfc91010_6672, \9486 );
and \U$20673 ( \29780 , RIfcdb728_7519, \9488 );
and \U$20674 ( \29781 , RIfcd8758_7485, \9490 );
and \U$20675 ( \29782 , RIe1ee868_4091, \9492 );
and \U$20676 ( \29783 , RIe1ec108_4063, \9494 );
and \U$20677 ( \29784 , RIe1e9408_4031, \9496 );
and \U$20678 ( \29785 , RIe1e6708_3999, \9498 );
and \U$20679 ( \29786 , RIe1e3a08_3967, \9500 );
and \U$20680 ( \29787 , RIe1e0d08_3935, \9502 );
and \U$20681 ( \29788 , RIe1de008_3903, \9504 );
and \U$20682 ( \29789 , RIe1db308_3871, \9506 );
and \U$20683 ( \29790 , RIe1d8608_3839, \9508 );
and \U$20684 ( \29791 , RIe1d2c08_3775, \9510 );
and \U$20685 ( \29792 , RIe1cff08_3743, \9512 );
and \U$20686 ( \29793 , RIe1cd208_3711, \9514 );
and \U$20687 ( \29794 , RIe1ca508_3679, \9516 );
and \U$20688 ( \29795 , RIe1c7808_3647, \9518 );
and \U$20689 ( \29796 , RIe1c4b08_3615, \9520 );
and \U$20690 ( \29797 , RIe1c1e08_3583, \9522 );
and \U$20691 ( \29798 , RIe1bf108_3551, \9524 );
and \U$20692 ( \29799 , RIf14cf48_5335, \9526 );
and \U$20693 ( \29800 , RIfc78d58_6397, \9528 );
and \U$20694 ( \29801 , RIe1b9b40_3490, \9530 );
and \U$20695 ( \29802 , RIfec5910_8368, \9532 );
and \U$20696 ( \29803 , RIfc78a88_6395, \9534 );
and \U$20697 ( \29804 , RIfcd51e8_7447, \9536 );
and \U$20698 ( \29805 , RIe1b57c0_3442, \9538 );
and \U$20699 ( \29806 , RIfea1010_8176, \9540 );
and \U$20700 ( \29807 , RIf1492d0_5292, \9542 );
and \U$20701 ( \29808 , RIfec5a78_8369, \9544 );
and \U$20702 ( \29809 , RIe1b2c28_3411, \9546 );
and \U$20703 ( \29810 , RIe1b12d8_3393, \9548 );
and \U$20704 ( \29811 , RIfec5640_8366, \9550 );
and \U$20705 ( \29812 , RIf146a08_5263, \9552 );
and \U$20706 ( \29813 , RIfec57a8_8367, \9554 );
and \U$20707 ( \29814 , RIfea1178_8177, \9556 );
and \U$20708 ( \29815 , RIe1a9448_3303, \9558 );
and \U$20709 ( \29816 , RIe1a6748_3271, \9560 );
and \U$20710 ( \29817 , RIe1a3a48_3239, \9562 );
and \U$20711 ( \29818 , RIe1a0d48_3207, \9564 );
and \U$20712 ( \29819 , RIe18d248_2983, \9566 );
and \U$20713 ( \29820 , RIe179748_2759, \9568 );
and \U$20714 ( \29821 , RIe2270a0_4734, \9570 );
and \U$20715 ( \29822 , RIe21bca0_4606, \9572 );
and \U$20716 ( \29823 , RIe2054a0_4350, \9574 );
and \U$20717 ( \29824 , RIe1ff500_4282, \9576 );
and \U$20718 ( \29825 , RIe1f88b8_4205, \9578 );
and \U$20719 ( \29826 , RIe1f1400_4122, \9580 );
and \U$20720 ( \29827 , RIe1d5908_3807, \9582 );
and \U$20721 ( \29828 , RIe1bc408_3519, \9584 );
and \U$20722 ( \29829 , RIe1af280_3370, \9586 );
and \U$20723 ( \29830 , RIe1718b8_2669, \9588 );
or \U$20724 ( \29831 , \29767 , \29768 , \29769 , \29770 , \29771 , \29772 , \29773 , \29774 , \29775 , \29776 , \29777 , \29778 , \29779 , \29780 , \29781 , \29782 , \29783 , \29784 , \29785 , \29786 , \29787 , \29788 , \29789 , \29790 , \29791 , \29792 , \29793 , \29794 , \29795 , \29796 , \29797 , \29798 , \29799 , \29800 , \29801 , \29802 , \29803 , \29804 , \29805 , \29806 , \29807 , \29808 , \29809 , \29810 , \29811 , \29812 , \29813 , \29814 , \29815 , \29816 , \29817 , \29818 , \29819 , \29820 , \29821 , \29822 , \29823 , \29824 , \29825 , \29826 , \29827 , \29828 , \29829 , \29830 );
or \U$20725 ( \29832 , \29766 , \29831 );
_DC g34f1 ( \29833_nG34f1 , \29832 , \9597 );
buf \U$20726 ( \29834 , \29833_nG34f1 );
and \U$20727 ( \29835 , \29701 , \29834 );
and \U$20728 ( \29836 , \27699 , \27832 );
and \U$20729 ( \29837 , \27832 , \28107 );
and \U$20730 ( \29838 , \27699 , \28107 );
or \U$20731 ( \29839 , \29836 , \29837 , \29838 );
and \U$20732 ( \29840 , \29834 , \29839 );
and \U$20733 ( \29841 , \29701 , \29839 );
or \U$20734 ( \29842 , \29835 , \29840 , \29841 );
xor \U$20735 ( \29843 , \29568 , \29842 );
buf g4400 ( \29844_nG4400 , \29843 );
xor \U$20736 ( \29845 , \29701 , \29834 );
xor \U$20737 ( \29846 , \29845 , \29839 );
buf g4403 ( \29847_nG4403 , \29846 );
nand \U$20738 ( \29848 , \29847_nG4403 , \28109_nG4406 );
and \U$20739 ( \29849 , \29844_nG4400 , \29848 );
xor \U$20740 ( \29850 , \29847_nG4403 , \28109_nG4406 );
not \U$20741 ( \29851 , \29850 );
xor \U$20742 ( \29852 , \29844_nG4400 , \29847_nG4403 );
and \U$20743 ( \29853 , \29851 , \29852 );
and \U$20745 ( \29854 , \29850 , \10694_nG9c0e );
or \U$20746 ( \29855 , 1'b0 , \29854 );
xor \U$20747 ( \29856 , \29849 , \29855 );
xor \U$20748 ( \29857 , \29849 , \29856 );
buf \U$20749 ( \29858 , \29857 );
buf \U$20750 ( \29859 , \29858 );
xor \U$20751 ( \29860 , \29301 , \29859 );
and \U$20752 ( \29861 , \28752 , \29288 );
and \U$20753 ( \29862 , \28752 , \29294 );
and \U$20754 ( \29863 , \29288 , \29294 );
or \U$20755 ( \29864 , \29861 , \29862 , \29863 );
and \U$20756 ( \29865 , \29860 , \29864 );
and \U$20757 ( \29866 , \29186 , \29191 );
and \U$20758 ( \29867 , \29186 , \29286 );
and \U$20759 ( \29868 , \29191 , \29286 );
or \U$20760 ( \29869 , \29866 , \29867 , \29868 );
buf \U$20761 ( \29870 , \29869 );
and \U$20762 ( \29871 , \29197 , \29228 );
and \U$20763 ( \29872 , \29197 , \29284 );
and \U$20764 ( \29873 , \29228 , \29284 );
or \U$20765 ( \29874 , \29871 , \29872 , \29873 );
buf \U$20766 ( \29875 , \29874 );
and \U$20767 ( \29876 , \29202 , \29219 );
and \U$20768 ( \29877 , \29202 , \29226 );
and \U$20769 ( \29878 , \29219 , \29226 );
or \U$20770 ( \29879 , \29876 , \29877 , \29878 );
buf \U$20771 ( \29880 , \29879 );
and \U$20772 ( \29881 , \14631 , \22629_nG9bd5 );
and \U$20773 ( \29882 , \14628 , \23696_nG9bd2 );
or \U$20774 ( \29883 , \29881 , \29882 );
xor \U$20775 ( \29884 , \14627 , \29883 );
buf \U$20776 ( \29885 , \29884 );
buf \U$20778 ( \29886 , \29885 );
xor \U$20779 ( \29887 , \29880 , \29886 );
and \U$20780 ( \29888 , \13370 , \24226_nG9bcf );
and \U$20781 ( \29889 , \13367 , \25298_nG9bcc );
or \U$20782 ( \29890 , \29888 , \29889 );
xor \U$20783 ( \29891 , \13366 , \29890 );
buf \U$20784 ( \29892 , \29891 );
buf \U$20786 ( \29893 , \29892 );
xor \U$20787 ( \29894 , \29887 , \29893 );
buf \U$20788 ( \29895 , \29894 );
xor \U$20789 ( \29896 , \29875 , \29895 );
and \U$20790 ( \29897 , \28721 , \28727 );
and \U$20791 ( \29898 , \28721 , \28734 );
and \U$20792 ( \29899 , \28727 , \28734 );
or \U$20793 ( \29900 , \29897 , \29898 , \29899 );
buf \U$20794 ( \29901 , \29900 );
xor \U$20795 ( \29902 , \29896 , \29901 );
buf \U$20796 ( \29903 , \29902 );
xor \U$20797 ( \29904 , \29870 , \29903 );
and \U$20798 ( \29905 , \29234 , \29260 );
and \U$20799 ( \29906 , \29234 , \29267 );
and \U$20800 ( \29907 , \29260 , \29267 );
or \U$20801 ( \29908 , \29905 , \29906 , \29907 );
buf \U$20802 ( \29909 , \29908 );
and \U$20803 ( \29910 , \29204 , \29210 );
and \U$20804 ( \29911 , \29204 , \29217 );
and \U$20805 ( \29912 , \29210 , \29217 );
or \U$20806 ( \29913 , \29910 , \29911 , \29912 );
buf \U$20807 ( \29914 , \29913 );
and \U$20808 ( \29915 , \29237 , \29243 );
buf \U$20809 ( \29916 , \29915 );
and \U$20810 ( \29917 , \24792 , \12801_nG9bff );
and \U$20811 ( \29918 , \24789 , \13705_nG9bfc );
or \U$20812 ( \29919 , \29917 , \29918 );
xor \U$20813 ( \29920 , \24788 , \29919 );
buf \U$20814 ( \29921 , \29920 );
buf \U$20816 ( \29922 , \29921 );
xor \U$20817 ( \29923 , \29916 , \29922 );
and \U$20818 ( \29924 , \23201 , \14070_nG9bf9 );
and \U$20819 ( \29925 , \23198 , \14984_nG9bf6 );
or \U$20820 ( \29926 , \29924 , \29925 );
xor \U$20821 ( \29927 , \23197 , \29926 );
buf \U$20822 ( \29928 , \29927 );
buf \U$20824 ( \29929 , \29928 );
xor \U$20825 ( \29930 , \29923 , \29929 );
buf \U$20826 ( \29931 , \29930 );
xor \U$20827 ( \29932 , \29914 , \29931 );
and \U$20828 ( \29933 , \20155 , \16680_nG9bed );
and \U$20829 ( \29934 , \20152 , \17665_nG9bea );
or \U$20830 ( \29935 , \29933 , \29934 );
xor \U$20831 ( \29936 , \20151 , \29935 );
buf \U$20832 ( \29937 , \29936 );
buf \U$20834 ( \29938 , \29937 );
xor \U$20835 ( \29939 , \29932 , \29938 );
buf \U$20836 ( \29940 , \29939 );
xor \U$20837 ( \29941 , \29909 , \29940 );
and \U$20838 ( \29942 , \17297 , \19586_nG9be1 );
and \U$20839 ( \29943 , \17294 , \20608_nG9bde );
or \U$20840 ( \29944 , \29942 , \29943 );
xor \U$20841 ( \29945 , \17293 , \29944 );
buf \U$20842 ( \29946 , \29945 );
buf \U$20844 ( \29947 , \29946 );
xor \U$20845 ( \29948 , \29941 , \29947 );
buf \U$20846 ( \29949 , \29948 );
and \U$20847 ( \29950 , \12157 , \25860_nG9bc9 );
and \U$20848 ( \29951 , \12154 , \26887_nG9bc6 );
or \U$20849 ( \29952 , \29950 , \29951 );
xor \U$20850 ( \29953 , \12153 , \29952 );
buf \U$20851 ( \29954 , \29953 );
buf \U$20853 ( \29955 , \29954 );
xor \U$20854 ( \29956 , \29949 , \29955 );
and \U$20855 ( \29957 , \10707 , \29179_nG9bbd );
and \U$20856 ( \29958 , \29142 , \29146 );
and \U$20857 ( \29959 , \29146 , \29171 );
and \U$20858 ( \29960 , \29142 , \29171 );
or \U$20859 ( \29961 , \29958 , \29959 , \29960 );
and \U$20860 ( \29962 , \29103 , \29117 );
and \U$20861 ( \29963 , \29117 , \29135 );
and \U$20862 ( \29964 , \29103 , \29135 );
or \U$20863 ( \29965 , \29962 , \29963 , \29964 );
and \U$20864 ( \29966 , \29151 , \29155 );
and \U$20865 ( \29967 , \29155 , \29170 );
and \U$20866 ( \29968 , \29151 , \29170 );
or \U$20867 ( \29969 , \29966 , \29967 , \29968 );
xor \U$20868 ( \29970 , \29965 , \29969 );
and \U$20869 ( \29971 , \27313 , \11574 );
and \U$20870 ( \29972 , \28534 , \11278 );
nor \U$20871 ( \29973 , \29971 , \29972 );
xnor \U$20872 ( \29974 , \29973 , \11580 );
and \U$20873 ( \29975 , \24199 , \14054 );
and \U$20874 ( \29976 , \25272 , \13692 );
nor \U$20875 ( \29977 , \29975 , \29976 );
xnor \U$20876 ( \29978 , \29977 , \14035 );
xor \U$20877 ( \29979 , \29974 , \29978 );
and \U$20878 ( \29980 , RIdec5db0_715, \9333 );
and \U$20879 ( \29981 , RIdec30b0_683, \9335 );
and \U$20880 ( \29982 , RIee201e8_4824, \9337 );
and \U$20881 ( \29983 , RIdec03b0_651, \9339 );
and \U$20882 ( \29984 , RIfcaf538_7017, \9341 );
and \U$20883 ( \29985 , RIdebd6b0_619, \9343 );
and \U$20884 ( \29986 , RIdeba9b0_587, \9345 );
and \U$20885 ( \29987 , RIdeb7cb0_555, \9347 );
and \U$20886 ( \29988 , RIfc40fe8_5765, \9349 );
and \U$20887 ( \29989 , RIdeb22b0_491, \9351 );
and \U$20888 ( \29990 , RIfcd08c8_7395, \9353 );
and \U$20889 ( \29991 , RIdeaf5b0_459, \9355 );
and \U$20890 ( \29992 , RIee1dd58_4798, \9357 );
and \U$20891 ( \29993 , RIdeabb18_427, \9359 );
and \U$20892 ( \29994 , RIdea5218_395, \9361 );
and \U$20893 ( \29995 , RIde9e918_363, \9363 );
and \U$20894 ( \29996 , RIee1d218_4790, \9365 );
and \U$20895 ( \29997 , RIfcedd10_7728, \9367 );
and \U$20896 ( \29998 , RIfce62b8_7641, \9369 );
and \U$20897 ( \29999 , RIfcc92a8_7311, \9371 );
and \U$20898 ( \30000 , RIde91da8_301, \9373 );
and \U$20899 ( \30001 , RIde8e928_285, \9375 );
and \U$20900 ( \30002 , RIde8a788_265, \9377 );
and \U$20901 ( \30003 , RIde865e8_245, \9379 );
and \U$20902 ( \30004 , RIde82448_225, \9381 );
and \U$20903 ( \30005 , RIfea1448_8179, \9383 );
and \U$20904 ( \30006 , RIfc750e0_6354, \9385 );
and \U$20905 ( \30007 , RIfcc19b8_7225, \9387 );
and \U$20906 ( \30008 , RIfced8d8_7725, \9389 );
and \U$20907 ( \30009 , RIfec5eb0_8372, \9391 );
and \U$20908 ( \30010 , RIe169fc8_2583, \9393 );
and \U$20909 ( \30011 , RIe168678_2565, \9395 );
and \U$20910 ( \30012 , RIe165db0_2536, \9397 );
and \U$20911 ( \30013 , RIe1630b0_2504, \9399 );
and \U$20912 ( \30014 , RIfccfc20_7386, \9401 );
and \U$20913 ( \30015 , RIe1603b0_2472, \9403 );
and \U$20914 ( \30016 , RIee365b0_5077, \9405 );
and \U$20915 ( \30017 , RIe15d6b0_2440, \9407 );
and \U$20916 ( \30018 , RIe157cb0_2376, \9409 );
and \U$20917 ( \30019 , RIe154fb0_2344, \9411 );
and \U$20918 ( \30020 , RIfea1718_8181, \9413 );
and \U$20919 ( \30021 , RIe1522b0_2312, \9415 );
and \U$20920 ( \30022 , RIee35200_5063, \9417 );
and \U$20921 ( \30023 , RIe14f5b0_2280, \9419 );
and \U$20922 ( \30024 , RIfcb0348_7027, \9421 );
and \U$20923 ( \30025 , RIe14c8b0_2248, \9423 );
and \U$20924 ( \30026 , RIe149bb0_2216, \9425 );
and \U$20925 ( \30027 , RIe146eb0_2184, \9427 );
and \U$20926 ( \30028 , RIfc73790_6336, \9429 );
and \U$20927 ( \30029 , RIfcdf238_7561, \9431 );
and \U$20928 ( \30030 , RIee32500_5031, \9433 );
and \U$20929 ( \30031 , RIfc94f58_6717, \9435 );
and \U$20930 ( \30032 , RIe141780_2122, \9437 );
and \U$20931 ( \30033 , RIe13f2f0_2096, \9439 );
and \U$20932 ( \30034 , RIfec5be0_8370, \9441 );
and \U$20933 ( \30035 , RIdf3ad68_2046, \9443 );
and \U$20934 ( \30036 , RIfea15b0_8180, \9445 );
and \U$20935 ( \30037 , RIfc5fb28_6111, \9447 );
and \U$20936 ( \30038 , RIfcae728_7007, \9449 );
and \U$20937 ( \30039 , RIfc74438_6345, \9451 );
and \U$20938 ( \30040 , RIdf36178_1992, \9453 );
and \U$20939 ( \30041 , RIdf33b80_1965, \9455 );
and \U$20940 ( \30042 , RIdf319c0_1941, \9457 );
and \U$20941 ( \30043 , RIdf2fad0_1919, \9459 );
or \U$20942 ( \30044 , \29980 , \29981 , \29982 , \29983 , \29984 , \29985 , \29986 , \29987 , \29988 , \29989 , \29990 , \29991 , \29992 , \29993 , \29994 , \29995 , \29996 , \29997 , \29998 , \29999 , \30000 , \30001 , \30002 , \30003 , \30004 , \30005 , \30006 , \30007 , \30008 , \30009 , \30010 , \30011 , \30012 , \30013 , \30014 , \30015 , \30016 , \30017 , \30018 , \30019 , \30020 , \30021 , \30022 , \30023 , \30024 , \30025 , \30026 , \30027 , \30028 , \30029 , \30030 , \30031 , \30032 , \30033 , \30034 , \30035 , \30036 , \30037 , \30038 , \30039 , \30040 , \30041 , \30042 , \30043 );
and \U$20943 ( \30045 , RIee2c290_4961, \9462 );
and \U$20944 ( \30046 , RIee2a940_4943, \9464 );
and \U$20945 ( \30047 , RIfc70658_6301, \9466 );
and \U$20946 ( \30048 , RIfc704f0_6300, \9468 );
and \U$20947 ( \30049 , RIdf2aaa8_1862, \9470 );
and \U$20948 ( \30050 , RIdf288e8_1838, \9472 );
and \U$20949 ( \30051 , RIdf269f8_1816, \9474 );
and \U$20950 ( \30052 , RIdf24f40_1797, \9476 );
and \U$20951 ( \30053 , RIfc64b50_6168, \9478 );
and \U$20952 ( \30054 , RIfccaa90_7328, \9480 );
and \U$20953 ( \30055 , RIdf231b8_1776, \9482 );
and \U$20954 ( \30056 , RIfcad4e0_6994, \9484 );
and \U$20955 ( \30057 , RIdf21ca0_1761, \9486 );
and \U$20956 ( \30058 , RIfeaad90_8260, \9488 );
and \U$20957 ( \30059 , RIdf1b490_1687, \9490 );
and \U$20958 ( \30060 , RIdf19b40_1669, \9492 );
and \U$20959 ( \30061 , RIdf17980_1645, \9494 );
and \U$20960 ( \30062 , RIdf14c80_1613, \9496 );
and \U$20961 ( \30063 , RIdf11f80_1581, \9498 );
and \U$20962 ( \30064 , RIdf0f280_1549, \9500 );
and \U$20963 ( \30065 , RIdf0c580_1517, \9502 );
and \U$20964 ( \30066 , RIdf09880_1485, \9504 );
and \U$20965 ( \30067 , RIdf06b80_1453, \9506 );
and \U$20966 ( \30068 , RIdf03e80_1421, \9508 );
and \U$20967 ( \30069 , RIdefe480_1357, \9510 );
and \U$20968 ( \30070 , RIdefb780_1325, \9512 );
and \U$20969 ( \30071 , RIdef8a80_1293, \9514 );
and \U$20970 ( \30072 , RIdef5d80_1261, \9516 );
and \U$20971 ( \30073 , RIdef3080_1229, \9518 );
and \U$20972 ( \30074 , RIdef0380_1197, \9520 );
and \U$20973 ( \30075 , RIdeed680_1165, \9522 );
and \U$20974 ( \30076 , RIdeea980_1133, \9524 );
and \U$20975 ( \30077 , RIfc595e8_6039, \9526 );
and \U$20976 ( \30078 , RIfcac568_6983, \9528 );
and \U$20977 ( \30079 , RIfcccf20_7354, \9530 );
and \U$20978 ( \30080 , RIfccd358_7357, \9532 );
and \U$20979 ( \30081 , RIdee5250_1071, \9534 );
and \U$20980 ( \30082 , RIfea7f28_8227, \9536 );
and \U$20981 ( \30083 , RIdee11a0_1025, \9538 );
and \U$20982 ( \30084 , RIfea12e0_8178, \9540 );
and \U$20983 ( \30085 , RIfc679b8_6201, \9542 );
and \U$20984 ( \30086 , RIee22510_4849, \9544 );
and \U$20985 ( \30087 , RIfc6dd90_6272, \9546 );
and \U$20986 ( \30088 , RIfc6cb48_6259, \9548 );
and \U$20987 ( \30089 , RIdeda120_945, \9550 );
and \U$20988 ( \30090 , RIded7b28_918, \9552 );
and \U$20989 ( \30091 , RIded5c38_896, \9554 );
and \U$20990 ( \30092 , RIfec5d48_8371, \9556 );
and \U$20991 ( \30093 , RIded11b0_843, \9558 );
and \U$20992 ( \30094 , RIdece4b0_811, \9560 );
and \U$20993 ( \30095 , RIdecb7b0_779, \9562 );
and \U$20994 ( \30096 , RIdec8ab0_747, \9564 );
and \U$20995 ( \30097 , RIdeb4fb0_523, \9566 );
and \U$20996 ( \30098 , RIde98018_331, \9568 );
and \U$20997 ( \30099 , RIe16ebb8_2637, \9570 );
and \U$20998 ( \30100 , RIe15a9b0_2408, \9572 );
and \U$20999 ( \30101 , RIe1441b0_2152, \9574 );
and \U$21000 ( \30102 , RIdf38ba8_2022, \9576 );
and \U$21001 ( \30103 , RIdf2d208_1890, \9578 );
and \U$21002 ( \30104 , RIdf1da88_1714, \9580 );
and \U$21003 ( \30105 , RIdf01180_1389, \9582 );
and \U$21004 ( \30106 , RIdee7c80_1101, \9584 );
and \U$21005 ( \30107 , RIdedc9e8_974, \9586 );
and \U$21006 ( \30108 , RIde7df60_204, \9588 );
or \U$21007 ( \30109 , \30045 , \30046 , \30047 , \30048 , \30049 , \30050 , \30051 , \30052 , \30053 , \30054 , \30055 , \30056 , \30057 , \30058 , \30059 , \30060 , \30061 , \30062 , \30063 , \30064 , \30065 , \30066 , \30067 , \30068 , \30069 , \30070 , \30071 , \30072 , \30073 , \30074 , \30075 , \30076 , \30077 , \30078 , \30079 , \30080 , \30081 , \30082 , \30083 , \30084 , \30085 , \30086 , \30087 , \30088 , \30089 , \30090 , \30091 , \30092 , \30093 , \30094 , \30095 , \30096 , \30097 , \30098 , \30099 , \30100 , \30101 , \30102 , \30103 , \30104 , \30105 , \30106 , \30107 , \30108 );
or \U$21008 ( \30110 , \30044 , \30109 );
_DC g61d6 ( \30111_nG61d6 , \30110 , \9597 );
and \U$21009 ( \30112 , RIe19e048_3175, \9059 );
and \U$21010 ( \30113 , RIe19b348_3143, \9061 );
and \U$21011 ( \30114 , RIfcc3ce0_7250, \9063 );
and \U$21012 ( \30115 , RIe198648_3111, \9065 );
and \U$21013 ( \30116 , RIfc7efc8_6467, \9067 );
and \U$21014 ( \30117 , RIe195948_3079, \9069 );
and \U$21015 ( \30118 , RIe192c48_3047, \9071 );
and \U$21016 ( \30119 , RIe18ff48_3015, \9073 );
and \U$21017 ( \30120 , RIe18a548_2951, \9075 );
and \U$21018 ( \30121 , RIe187848_2919, \9077 );
and \U$21019 ( \30122 , RIfc46790_5824, \9079 );
and \U$21020 ( \30123 , RIe184b48_2887, \9081 );
and \U$21021 ( \30124 , RIfc98d38_6761, \9083 );
and \U$21022 ( \30125 , RIe181e48_2855, \9085 );
and \U$21023 ( \30126 , RIe17f148_2823, \9087 );
and \U$21024 ( \30127 , RIe17c448_2791, \9089 );
and \U$21025 ( \30128 , RIfcb5d48_7091, \9091 );
and \U$21026 ( \30129 , RIfc995a8_6767, \9093 );
and \U$21027 ( \30130 , RIfc9a3b8_6777, \9095 );
and \U$21028 ( \30131 , RIe1761d8_2721, \9097 );
and \U$21029 ( \30132 , RIfc54188_5979, \9099 );
and \U$21030 ( \30133 , RIfcd2bf0_7420, \9101 );
and \U$21031 ( \30134 , RIfc8b778_6609, \9103 );
and \U$21032 ( \30135 , RIfc7dee8_6455, \9105 );
and \U$21033 ( \30136 , RIee3c550_5145, \9107 );
and \U$21034 ( \30137 , RIfc8c420_6618, \9109 );
and \U$21035 ( \30138 , RIee3a0c0_5119, \9111 );
and \U$21036 ( \30139 , RIfeaba38_8269, \9113 );
and \U$21037 ( \30140 , RIfc46628_5823, \9115 );
and \U$21038 ( \30141 , RIfcbc288_7163, \9117 );
and \U$21039 ( \30142 , RIf16e710_5716, \9119 );
and \U$21040 ( \30143 , RIfc8fdc8_6659, \9121 );
and \U$21041 ( \30144 , RIfc48c20_5850, \9123 );
and \U$21042 ( \30145 , RIe2243a0_4702, \9125 );
and \U$21043 ( \30146 , RIfca0358_6845, \9127 );
and \U$21044 ( \30147 , RIe2216a0_4670, \9129 );
and \U$21045 ( \30148 , RIfc9a688_6779, \9131 );
and \U$21046 ( \30149 , RIe21e9a0_4638, \9133 );
and \U$21047 ( \30150 , RIe218fa0_4574, \9135 );
and \U$21048 ( \30151 , RIe2162a0_4542, \9137 );
and \U$21049 ( \30152 , RIfc456b0_5812, \9139 );
and \U$21050 ( \30153 , RIe2135a0_4510, \9141 );
and \U$21051 ( \30154 , RIf169418_5657, \9143 );
and \U$21052 ( \30155 , RIe2108a0_4478, \9145 );
and \U$21053 ( \30156 , RIfc8bfe8_6615, \9147 );
and \U$21054 ( \30157 , RIe20dba0_4446, \9149 );
and \U$21055 ( \30158 , RIe20aea0_4414, \9151 );
and \U$21056 ( \30159 , RIe2081a0_4382, \9153 );
and \U$21057 ( \30160 , RIfc8c9c0_6622, \9155 );
and \U$21058 ( \30161 , RIfc7f568_6471, \9157 );
and \U$21059 ( \30162 , RIe202d40_4322, \9159 );
and \U$21060 ( \30163 , RIe201120_4302, \9161 );
and \U$21061 ( \30164 , RIfce2910_7600, \9163 );
and \U$21062 ( \30165 , RIfc487e8_5847, \9165 );
and \U$21063 ( \30166 , RIfc46d30_5828, \9167 );
and \U$21064 ( \30167 , RIfc992d8_6765, \9169 );
and \U$21065 ( \30168 , RIfca2680_6870, \9171 );
and \U$21066 ( \30169 , RIfc44a08_5803, \9173 );
and \U$21067 ( \30170 , RIe1fd1d8_4257, \9175 );
and \U$21068 ( \30171 , RIe1fbf90_4244, \9177 );
and \U$21069 ( \30172 , RIfc580d0_6024, \9179 );
and \U$21070 ( \30173 , RIfcbdbd8_7181, \9181 );
and \U$21071 ( \30174 , RIfc8dd70_6636, \9183 );
and \U$21072 ( \30175 , RIfce01b0_7572, \9185 );
or \U$21073 ( \30176 , \30112 , \30113 , \30114 , \30115 , \30116 , \30117 , \30118 , \30119 , \30120 , \30121 , \30122 , \30123 , \30124 , \30125 , \30126 , \30127 , \30128 , \30129 , \30130 , \30131 , \30132 , \30133 , \30134 , \30135 , \30136 , \30137 , \30138 , \30139 , \30140 , \30141 , \30142 , \30143 , \30144 , \30145 , \30146 , \30147 , \30148 , \30149 , \30150 , \30151 , \30152 , \30153 , \30154 , \30155 , \30156 , \30157 , \30158 , \30159 , \30160 , \30161 , \30162 , \30163 , \30164 , \30165 , \30166 , \30167 , \30168 , \30169 , \30170 , \30171 , \30172 , \30173 , \30174 , \30175 );
and \U$21074 ( \30177 , RIfc7bbc0_6430, \9188 );
and \U$21075 ( \30178 , RIfc90368_6663, \9190 );
and \U$21076 ( \30179 , RIfc7b8f0_6428, \9192 );
and \U$21077 ( \30180 , RIe1fa910_4228, \9194 );
and \U$21078 ( \30181 , RIfcd8b90_7488, \9196 );
and \U$21079 ( \30182 , RIfc43ec8_5795, \9198 );
and \U$21080 ( \30183 , RIfc7b788_6427, \9200 );
and \U$21081 ( \30184 , RIe1f5e88_4175, \9202 );
and \U$21082 ( \30185 , RIfc7b350_6424, \9204 );
and \U$21083 ( \30186 , RIfc90d40_6670, \9206 );
and \U$21084 ( \30187 , RIfca3490_6880, \9208 );
and \U$21085 ( \30188 , RIe1f3b60_4150, \9210 );
and \U$21086 ( \30189 , RIfc91010_6672, \9212 );
and \U$21087 ( \30190 , RIfcdb728_7519, \9214 );
and \U$21088 ( \30191 , RIfcd8758_7485, \9216 );
and \U$21089 ( \30192 , RIe1ee868_4091, \9218 );
and \U$21090 ( \30193 , RIe1ec108_4063, \9220 );
and \U$21091 ( \30194 , RIe1e9408_4031, \9222 );
and \U$21092 ( \30195 , RIe1e6708_3999, \9224 );
and \U$21093 ( \30196 , RIe1e3a08_3967, \9226 );
and \U$21094 ( \30197 , RIe1e0d08_3935, \9228 );
and \U$21095 ( \30198 , RIe1de008_3903, \9230 );
and \U$21096 ( \30199 , RIe1db308_3871, \9232 );
and \U$21097 ( \30200 , RIe1d8608_3839, \9234 );
and \U$21098 ( \30201 , RIe1d2c08_3775, \9236 );
and \U$21099 ( \30202 , RIe1cff08_3743, \9238 );
and \U$21100 ( \30203 , RIe1cd208_3711, \9240 );
and \U$21101 ( \30204 , RIe1ca508_3679, \9242 );
and \U$21102 ( \30205 , RIe1c7808_3647, \9244 );
and \U$21103 ( \30206 , RIe1c4b08_3615, \9246 );
and \U$21104 ( \30207 , RIe1c1e08_3583, \9248 );
and \U$21105 ( \30208 , RIe1bf108_3551, \9250 );
and \U$21106 ( \30209 , RIf14cf48_5335, \9252 );
and \U$21107 ( \30210 , RIfc78d58_6397, \9254 );
and \U$21108 ( \30211 , RIe1b9b40_3490, \9256 );
and \U$21109 ( \30212 , RIfec5910_8368, \9258 );
and \U$21110 ( \30213 , RIfc78a88_6395, \9260 );
and \U$21111 ( \30214 , RIfcd51e8_7447, \9262 );
and \U$21112 ( \30215 , RIe1b57c0_3442, \9264 );
and \U$21113 ( \30216 , RIfea1010_8176, \9266 );
and \U$21114 ( \30217 , RIf1492d0_5292, \9268 );
and \U$21115 ( \30218 , RIfec5a78_8369, \9270 );
and \U$21116 ( \30219 , RIe1b2c28_3411, \9272 );
and \U$21117 ( \30220 , RIe1b12d8_3393, \9274 );
and \U$21118 ( \30221 , RIfec5640_8366, \9276 );
and \U$21119 ( \30222 , RIf146a08_5263, \9278 );
and \U$21120 ( \30223 , RIfec57a8_8367, \9280 );
and \U$21121 ( \30224 , RIfea1178_8177, \9282 );
and \U$21122 ( \30225 , RIe1a9448_3303, \9284 );
and \U$21123 ( \30226 , RIe1a6748_3271, \9286 );
and \U$21124 ( \30227 , RIe1a3a48_3239, \9288 );
and \U$21125 ( \30228 , RIe1a0d48_3207, \9290 );
and \U$21126 ( \30229 , RIe18d248_2983, \9292 );
and \U$21127 ( \30230 , RIe179748_2759, \9294 );
and \U$21128 ( \30231 , RIe2270a0_4734, \9296 );
and \U$21129 ( \30232 , RIe21bca0_4606, \9298 );
and \U$21130 ( \30233 , RIe2054a0_4350, \9300 );
and \U$21131 ( \30234 , RIe1ff500_4282, \9302 );
and \U$21132 ( \30235 , RIe1f88b8_4205, \9304 );
and \U$21133 ( \30236 , RIe1f1400_4122, \9306 );
and \U$21134 ( \30237 , RIe1d5908_3807, \9308 );
and \U$21135 ( \30238 , RIe1bc408_3519, \9310 );
and \U$21136 ( \30239 , RIe1af280_3370, \9312 );
and \U$21137 ( \30240 , RIe1718b8_2669, \9314 );
or \U$21138 ( \30241 , \30177 , \30178 , \30179 , \30180 , \30181 , \30182 , \30183 , \30184 , \30185 , \30186 , \30187 , \30188 , \30189 , \30190 , \30191 , \30192 , \30193 , \30194 , \30195 , \30196 , \30197 , \30198 , \30199 , \30200 , \30201 , \30202 , \30203 , \30204 , \30205 , \30206 , \30207 , \30208 , \30209 , \30210 , \30211 , \30212 , \30213 , \30214 , \30215 , \30216 , \30217 , \30218 , \30219 , \30220 , \30221 , \30222 , \30223 , \30224 , \30225 , \30226 , \30227 , \30228 , \30229 , \30230 , \30231 , \30232 , \30233 , \30234 , \30235 , \30236 , \30237 , \30238 , \30239 , \30240 );
or \U$21139 ( \30242 , \30176 , \30241 );
_DC g625a ( \30243_nG625a , \30242 , \9323 );
xor g625b ( \30244_nG625b , \30111_nG61d6 , \30243_nG625a );
buf \U$21140 ( \30245 , \30244_nG625b );
xor \U$21141 ( \30246 , \30245 , \29067 );
and \U$21142 ( \30247 , \10687 , \30246 );
xor \U$21143 ( \30248 , \29979 , \30247 );
and \U$21144 ( \30249 , \25815 , \12790 );
and \U$21145 ( \30250 , \26829 , \12461 );
nor \U$21146 ( \30251 , \30249 , \30250 );
xnor \U$21147 ( \30252 , \30251 , \12780 );
and \U$21148 ( \30253 , \19558 , \18090 );
and \U$21149 ( \30254 , \20544 , \17655 );
nor \U$21150 ( \30255 , \30253 , \30254 );
xnor \U$21151 ( \30256 , \30255 , \18046 );
xor \U$21152 ( \30257 , \30252 , \30256 );
and \U$21153 ( \30258 , \10988 , \29070 );
and \U$21154 ( \30259 , \11270 , \28526 );
nor \U$21155 ( \30260 , \30258 , \30259 );
xnor \U$21156 ( \30261 , \30260 , \29076 );
xor \U$21157 ( \30262 , \30257 , \30261 );
xor \U$21158 ( \30263 , \30248 , \30262 );
and \U$21159 ( \30264 , \29084 , \10983 );
_DC g65cb ( \30265_nG65cb , \30110 , \9597 );
_DC g65cc ( \30266_nG65cc , \30242 , \9323 );
and g65cd ( \30267_nG65cd , \30265_nG65cb , \30266_nG65cc );
buf \U$21160 ( \30268 , \30267_nG65cd );
and \U$21161 ( \30269 , \30268 , \10691 );
nor \U$21162 ( \30270 , \30264 , \30269 );
xnor \U$21163 ( \30271 , \30270 , \10980 );
and \U$21164 ( \30272 , \15321 , \22542 );
and \U$21165 ( \30273 , \16267 , \22103 );
nor \U$21166 ( \30274 , \30272 , \30273 );
xnor \U$21167 ( \30275 , \30274 , \22548 );
xor \U$21168 ( \30276 , \30271 , \30275 );
and \U$21169 ( \30277 , \14024 , \24138 );
and \U$21170 ( \30278 , \14950 , \23630 );
nor \U$21171 ( \30279 , \30277 , \30278 );
xnor \U$21172 ( \30280 , \30279 , \24144 );
xor \U$21173 ( \30281 , \30276 , \30280 );
xor \U$21174 ( \30282 , \30263 , \30281 );
xor \U$21175 ( \30283 , \29970 , \30282 );
xor \U$21176 ( \30284 , \29961 , \30283 );
and \U$21177 ( \30285 , \28778 , \29098 );
and \U$21178 ( \30286 , \29098 , \29136 );
and \U$21179 ( \30287 , \28778 , \29136 );
or \U$21180 ( \30288 , \30285 , \30286 , \30287 );
and \U$21181 ( \30289 , \29160 , \29164 );
and \U$21182 ( \30290 , \29164 , \29169 );
and \U$21183 ( \30291 , \29160 , \29169 );
or \U$21184 ( \30292 , \30289 , \30290 , \30291 );
and \U$21185 ( \30293 , \29125 , \29129 );
and \U$21186 ( \30294 , \29129 , \29134 );
and \U$21187 ( \30295 , \29125 , \29134 );
or \U$21188 ( \30296 , \30293 , \30294 , \30295 );
xor \U$21189 ( \30297 , \30292 , \30296 );
and \U$21190 ( \30298 , \21033 , \16635 );
and \U$21191 ( \30299 , \22090 , \16301 );
nor \U$21192 ( \30300 , \30298 , \30299 );
xnor \U$21193 ( \30301 , \30300 , \16625 );
and \U$21194 ( \30302 , \12769 , \25826 );
and \U$21195 ( \30303 , \13679 , \25264 );
nor \U$21196 ( \30304 , \30302 , \30303 );
xnor \U$21197 ( \30305 , \30304 , \25773 );
xor \U$21198 ( \30306 , \30301 , \30305 );
and \U$21199 ( \30307 , \11586 , \27397 );
and \U$21200 ( \30308 , \12448 , \26807 );
nor \U$21201 ( \30309 , \30307 , \30308 );
xnor \U$21202 ( \30310 , \30309 , \27295 );
xor \U$21203 ( \30311 , \30306 , \30310 );
xor \U$21204 ( \30312 , \30297 , \30311 );
xor \U$21205 ( \30313 , \30288 , \30312 );
and \U$21206 ( \30314 , \28792 , \29078 );
and \U$21207 ( \30315 , \29078 , \29097 );
and \U$21208 ( \30316 , \28792 , \29097 );
or \U$21209 ( \30317 , \30314 , \30315 , \30316 );
and \U$21210 ( \30318 , \28782 , \28786 );
and \U$21211 ( \30319 , \28786 , \28791 );
and \U$21212 ( \30320 , \28782 , \28791 );
or \U$21213 ( \30321 , \30318 , \30319 , \30320 );
and \U$21214 ( \30322 , \29107 , \29111 );
and \U$21215 ( \30323 , \29111 , \29116 );
and \U$21216 ( \30324 , \29107 , \29116 );
or \U$21217 ( \30325 , \30322 , \30323 , \30324 );
xor \U$21218 ( \30326 , \30321 , \30325 );
and \U$21219 ( \30327 , \29122 , \29124 );
xor \U$21220 ( \30328 , \30326 , \30327 );
xor \U$21221 ( \30329 , \30317 , \30328 );
and \U$21222 ( \30330 , \28796 , \28800 );
and \U$21223 ( \30331 , \28800 , \29077 );
and \U$21224 ( \30332 , \28796 , \29077 );
or \U$21225 ( \30333 , \30330 , \30331 , \30332 );
and \U$21226 ( \30334 , \29087 , \29091 );
and \U$21227 ( \30335 , \29091 , \29096 );
and \U$21228 ( \30336 , \29087 , \29096 );
or \U$21229 ( \30337 , \30334 , \30335 , \30336 );
xor \U$21230 ( \30338 , \30333 , \30337 );
and \U$21231 ( \30339 , \22556 , \15336 );
and \U$21232 ( \30340 , \23617 , \14963 );
nor \U$21233 ( \30341 , \30339 , \30340 );
xnor \U$21234 ( \30342 , \30341 , \15342 );
and \U$21235 ( \30343 , \18035 , \19534 );
and \U$21236 ( \30344 , \19032 , \19045 );
nor \U$21237 ( \30345 , \30343 , \30344 );
xnor \U$21238 ( \30346 , \30345 , \19540 );
xor \U$21239 ( \30347 , \30342 , \30346 );
and \U$21240 ( \30348 , \16655 , \21005 );
and \U$21241 ( \30349 , \17627 , \20557 );
nor \U$21242 ( \30350 , \30348 , \30349 );
xnor \U$21243 ( \30351 , \30350 , \21011 );
xor \U$21244 ( \30352 , \30347 , \30351 );
xor \U$21245 ( \30353 , \30338 , \30352 );
xor \U$21246 ( \30354 , \30329 , \30353 );
xor \U$21247 ( \30355 , \30313 , \30354 );
xor \U$21248 ( \30356 , \30284 , \30355 );
and \U$21249 ( \30357 , \28774 , \29137 );
and \U$21250 ( \30358 , \29137 , \29172 );
and \U$21251 ( \30359 , \28774 , \29172 );
or \U$21252 ( \30360 , \30357 , \30358 , \30359 );
xor \U$21253 ( \30361 , \30356 , \30360 );
and \U$21254 ( \30362 , \28770 , \29173 );
and \U$21255 ( \30363 , \29174 , \29177 );
or \U$21256 ( \30364 , \30362 , \30363 );
xor \U$21257 ( \30365 , \30361 , \30364 );
buf g9bba ( \30366_nG9bba , \30365 );
and \U$21258 ( \30367 , \10704 , \30366_nG9bba );
or \U$21259 ( \30368 , \29957 , \30367 );
xor \U$21260 ( \30369 , \10703 , \30368 );
buf \U$21261 ( \30370 , \30369 );
buf \U$21263 ( \30371 , \30370 );
xor \U$21264 ( \30372 , \29956 , \30371 );
buf \U$21265 ( \30373 , \30372 );
xor \U$21266 ( \30374 , \29904 , \30373 );
buf \U$21267 ( \30375 , \30374 );
and \U$21268 ( \30376 , \28711 , \28744 );
and \U$21269 ( \30377 , \28711 , \28750 );
and \U$21270 ( \30378 , \28744 , \28750 );
or \U$21271 ( \30379 , \30376 , \30377 , \30378 );
buf \U$21272 ( \30380 , \30379 );
xor \U$21273 ( \30381 , \30375 , \30380 );
and \U$21274 ( \30382 , \28716 , \28736 );
and \U$21275 ( \30383 , \28716 , \28742 );
and \U$21276 ( \30384 , \28736 , \28742 );
or \U$21277 ( \30385 , \30382 , \30383 , \30384 );
buf \U$21278 ( \30386 , \30385 );
and \U$21279 ( \30387 , \29269 , \29275 );
and \U$21280 ( \30388 , \29269 , \29282 );
and \U$21281 ( \30389 , \29275 , \29282 );
or \U$21282 ( \30390 , \30387 , \30388 , \30389 );
buf \U$21283 ( \30391 , \30390 );
and \U$21284 ( \30392 , \29245 , \29251 );
and \U$21285 ( \30393 , \29245 , \29258 );
and \U$21286 ( \30394 , \29251 , \29258 );
or \U$21287 ( \30395 , \30392 , \30393 , \30394 );
buf \U$21288 ( \30396 , \30395 );
and \U$21289 ( \30397 , \28118 , \10995_nG9c0b );
and \U$21290 ( \30398 , \28115 , \11283_nG9c08 );
or \U$21291 ( \30399 , \30397 , \30398 );
xor \U$21292 ( \30400 , \28114 , \30399 );
buf \U$21293 ( \30401 , \30400 );
buf \U$21295 ( \30402 , \30401 );
and \U$21296 ( \30403 , \26431 , \11598_nG9c05 );
and \U$21297 ( \30404 , \26428 , \12470_nG9c02 );
or \U$21298 ( \30405 , \30403 , \30404 );
xor \U$21299 ( \30406 , \26427 , \30405 );
buf \U$21300 ( \30407 , \30406 );
buf \U$21302 ( \30408 , \30407 );
xor \U$21303 ( \30409 , \30402 , \30408 );
buf \U$21304 ( \30410 , \30409 );
xor \U$21305 ( \30411 , \30396 , \30410 );
and \U$21306 ( \30412 , \21658 , \15373_nG9bf3 );
and \U$21307 ( \30413 , \21655 , \16315_nG9bf0 );
or \U$21308 ( \30414 , \30412 , \30413 );
xor \U$21309 ( \30415 , \21654 , \30414 );
buf \U$21310 ( \30416 , \30415 );
buf \U$21312 ( \30417 , \30416 );
xor \U$21313 ( \30418 , \30411 , \30417 );
buf \U$21314 ( \30419 , \30418 );
and \U$21315 ( \30420 , \18702 , \18107_nG9be7 );
and \U$21316 ( \30421 , \18699 , \19091_nG9be4 );
or \U$21317 ( \30422 , \30420 , \30421 );
xor \U$21318 ( \30423 , \18698 , \30422 );
buf \U$21319 ( \30424 , \30423 );
buf \U$21321 ( \30425 , \30424 );
xor \U$21322 ( \30426 , \30419 , \30425 );
and \U$21323 ( \30427 , \15940 , \21086_nG9bdb );
and \U$21324 ( \30428 , \15937 , \22129_nG9bd8 );
or \U$21325 ( \30429 , \30427 , \30428 );
xor \U$21326 ( \30430 , \15936 , \30429 );
buf \U$21327 ( \30431 , \30430 );
buf \U$21329 ( \30432 , \30431 );
xor \U$21330 ( \30433 , \30426 , \30432 );
buf \U$21331 ( \30434 , \30433 );
xor \U$21332 ( \30435 , \30391 , \30434 );
and \U$21333 ( \30436 , \10421 , \27416_nG9bc3 );
and \U$21334 ( \30437 , \10418 , \28602_nG9bc0 );
or \U$21335 ( \30438 , \30436 , \30437 );
xor \U$21336 ( \30439 , \10417 , \30438 );
buf \U$21337 ( \30440 , \30439 );
buf \U$21339 ( \30441 , \30440 );
xor \U$21340 ( \30442 , \30435 , \30441 );
buf \U$21341 ( \30443 , \30442 );
xor \U$21342 ( \30444 , \30386 , \30443 );
and \U$21343 ( \30445 , \28758 , \28764 );
and \U$21344 ( \30446 , \28758 , \29184 );
and \U$21345 ( \30447 , \28764 , \29184 );
or \U$21346 ( \30448 , \30445 , \30446 , \30447 );
buf \U$21347 ( \30449 , \30448 );
xor \U$21348 ( \30450 , \30444 , \30449 );
buf \U$21349 ( \30451 , \30450 );
xor \U$21350 ( \30452 , \30381 , \30451 );
and \U$21351 ( \30453 , \29860 , \30452 );
and \U$21352 ( \30454 , \29864 , \30452 );
or \U$21353 ( \30455 , \29865 , \30453 , \30454 );
and \U$21354 ( \30456 , \29296 , \29300 );
and \U$21355 ( \30457 , \29296 , \29859 );
and \U$21356 ( \30458 , \29300 , \29859 );
or \U$21357 ( \30459 , \30456 , \30457 , \30458 );
xor \U$21358 ( \30460 , \30455 , \30459 );
and \U$21359 ( \30461 , \30375 , \30380 );
and \U$21360 ( \30462 , \30375 , \30451 );
and \U$21361 ( \30463 , \30380 , \30451 );
or \U$21362 ( \30464 , \30461 , \30462 , \30463 );
xor \U$21363 ( \30465 , \30460 , \30464 );
and \U$21364 ( \30466 , \30396 , \30410 );
and \U$21365 ( \30467 , \30396 , \30417 );
and \U$21366 ( \30468 , \30410 , \30417 );
or \U$21367 ( \30469 , \30466 , \30467 , \30468 );
buf \U$21368 ( \30470 , \30469 );
and \U$21369 ( \30471 , \30402 , \30408 );
buf \U$21370 ( \30472 , \30471 );
and \U$21371 ( \30473 , \24792 , \13705_nG9bfc );
and \U$21372 ( \30474 , \24789 , \14070_nG9bf9 );
or \U$21373 ( \30475 , \30473 , \30474 );
xor \U$21374 ( \30476 , \24788 , \30475 );
buf \U$21375 ( \30477 , \30476 );
buf \U$21377 ( \30478 , \30477 );
xor \U$21378 ( \30479 , \30472 , \30478 );
and \U$21379 ( \30480 , \23201 , \14984_nG9bf6 );
and \U$21380 ( \30481 , \23198 , \15373_nG9bf3 );
or \U$21381 ( \30482 , \30480 , \30481 );
xor \U$21382 ( \30483 , \23197 , \30482 );
buf \U$21383 ( \30484 , \30483 );
buf \U$21385 ( \30485 , \30484 );
xor \U$21386 ( \30486 , \30479 , \30485 );
buf \U$21387 ( \30487 , \30486 );
xor \U$21388 ( \30488 , \30470 , \30487 );
and \U$21389 ( \30489 , \20155 , \17665_nG9bea );
and \U$21390 ( \30490 , \20152 , \18107_nG9be7 );
or \U$21391 ( \30491 , \30489 , \30490 );
xor \U$21392 ( \30492 , \20151 , \30491 );
buf \U$21393 ( \30493 , \30492 );
buf \U$21395 ( \30494 , \30493 );
xor \U$21396 ( \30495 , \30488 , \30494 );
buf \U$21397 ( \30496 , \30495 );
and \U$21398 ( \30497 , \29914 , \29931 );
and \U$21399 ( \30498 , \29914 , \29938 );
and \U$21400 ( \30499 , \29931 , \29938 );
or \U$21401 ( \30500 , \30497 , \30498 , \30499 );
buf \U$21402 ( \30501 , \30500 );
xor \U$21403 ( \30502 , \30496 , \30501 );
and \U$21404 ( \30503 , \15940 , \22129_nG9bd8 );
and \U$21405 ( \30504 , \15937 , \22629_nG9bd5 );
or \U$21406 ( \30505 , \30503 , \30504 );
xor \U$21407 ( \30506 , \15936 , \30505 );
buf \U$21408 ( \30507 , \30506 );
buf \U$21410 ( \30508 , \30507 );
xor \U$21411 ( \30509 , \30502 , \30508 );
buf \U$21412 ( \30510 , \30509 );
and \U$21413 ( \30511 , \29909 , \29940 );
and \U$21414 ( \30512 , \29909 , \29947 );
and \U$21415 ( \30513 , \29940 , \29947 );
or \U$21416 ( \30514 , \30511 , \30512 , \30513 );
buf \U$21417 ( \30515 , \30514 );
xor \U$21418 ( \30516 , \30510 , \30515 );
and \U$21419 ( \30517 , \10707 , \30366_nG9bba );
and \U$21420 ( \30518 , \29965 , \29969 );
and \U$21421 ( \30519 , \29969 , \30282 );
and \U$21422 ( \30520 , \29965 , \30282 );
or \U$21423 ( \30521 , \30518 , \30519 , \30520 );
and \U$21424 ( \30522 , \30288 , \30312 );
and \U$21425 ( \30523 , \30312 , \30354 );
and \U$21426 ( \30524 , \30288 , \30354 );
or \U$21427 ( \30525 , \30522 , \30523 , \30524 );
xor \U$21428 ( \30526 , \30521 , \30525 );
and \U$21429 ( \30527 , \30321 , \30325 );
and \U$21430 ( \30528 , \30325 , \30327 );
and \U$21431 ( \30529 , \30321 , \30327 );
or \U$21432 ( \30530 , \30527 , \30528 , \30529 );
and \U$21433 ( \30531 , \30248 , \30262 );
and \U$21434 ( \30532 , \30262 , \30281 );
and \U$21435 ( \30533 , \30248 , \30281 );
or \U$21436 ( \30534 , \30531 , \30532 , \30533 );
xor \U$21437 ( \30535 , \30530 , \30534 );
and \U$21438 ( \30536 , \30268 , \10983 );
and \U$21439 ( \30537 , RIdec5f18_716, \9333 );
and \U$21440 ( \30538 , RIdec3218_684, \9335 );
and \U$21441 ( \30539 , RIee20350_4825, \9337 );
and \U$21442 ( \30540 , RIdec0518_652, \9339 );
and \U$21443 ( \30541 , RIee1f6a8_4816, \9341 );
and \U$21444 ( \30542 , RIdebd818_620, \9343 );
and \U$21445 ( \30543 , RIdebab18_588, \9345 );
and \U$21446 ( \30544 , RIdeb7e18_556, \9347 );
and \U$21447 ( \30545 , RIfce4da0_7626, \9349 );
and \U$21448 ( \30546 , RIdeb2418_492, \9351 );
and \U$21449 ( \30547 , RIfcea908_7691, \9353 );
and \U$21450 ( \30548 , RIdeaf718_460, \9355 );
and \U$21451 ( \30549 , RIfce20a0_7594, \9357 );
and \U$21452 ( \30550 , RIdeabe60_428, \9359 );
and \U$21453 ( \30551 , RIdea5560_396, \9361 );
and \U$21454 ( \30552 , RIde9ec60_364, \9363 );
and \U$21455 ( \30553 , RIfce6420_7642, \9365 );
and \U$21456 ( \30554 , RIee1c2a0_4779, \9367 );
and \U$21457 ( \30555 , RIfc75950_6360, \9369 );
and \U$21458 ( \30556 , RIee1ad88_4764, \9371 );
and \U$21459 ( \30557 , RIde920f0_302, \9373 );
and \U$21460 ( \30558 , RIfea4148_8211, \9375 );
and \U$21461 ( \30559 , RIfeaa688_8255, \9377 );
and \U$21462 ( \30560 , RIfea3fe0_8210, \9379 );
and \U$21463 ( \30561 , RIde82790_226, \9381 );
and \U$21464 ( \30562 , RIfc6f848_6291, \9383 );
and \U$21465 ( \30563 , RIfc5dc38_6089, \9385 );
and \U$21466 ( \30564 , RIfc76b98_6373, \9387 );
and \U$21467 ( \30565 , RIfcae2f0_7004, \9389 );
and \U$21468 ( \30566 , RIe16c020_2606, \9391 );
and \U$21469 ( \30567 , RIe16a130_2584, \9393 );
and \U$21470 ( \30568 , RIe1687e0_2566, \9395 );
and \U$21471 ( \30569 , RIe165f18_2537, \9397 );
and \U$21472 ( \30570 , RIe163218_2505, \9399 );
and \U$21473 ( \30571 , RIfcadd50_7000, \9401 );
and \U$21474 ( \30572 , RIe160518_2473, \9403 );
and \U$21475 ( \30573 , RIfc55268_5991, \9405 );
and \U$21476 ( \30574 , RIe15d818_2441, \9407 );
and \U$21477 ( \30575 , RIe157e18_2377, \9409 );
and \U$21478 ( \30576 , RIe155118_2345, \9411 );
and \U$21479 ( \30577 , RIfc45548_5811, \9413 );
and \U$21480 ( \30578 , RIe152418_2313, \9415 );
and \U$21481 ( \30579 , RIfc498c8_5859, \9417 );
and \U$21482 ( \30580 , RIe14f718_2281, \9419 );
and \U$21483 ( \30581 , RIfcbda70_7180, \9421 );
and \U$21484 ( \30582 , RIe14ca18_2249, \9423 );
and \U$21485 ( \30583 , RIe149d18_2217, \9425 );
and \U$21486 ( \30584 , RIe147018_2185, \9427 );
and \U$21487 ( \30585 , RIee34828_5056, \9429 );
and \U$21488 ( \30586 , RIee33748_5044, \9431 );
and \U$21489 ( \30587 , RIee32668_5032, \9433 );
and \U$21490 ( \30588 , RIee31588_5020, \9435 );
and \U$21491 ( \30589 , RIe1418e8_2123, \9437 );
and \U$21492 ( \30590 , RIe13f458_2097, \9439 );
and \U$21493 ( \30591 , RIdf3d360_2073, \9441 );
and \U$21494 ( \30592 , RIdf3aed0_2047, \9443 );
and \U$21495 ( \30593 , RIfc526d0_5960, \9445 );
and \U$21496 ( \30594 , RIfc42848_5779, \9447 );
and \U$21497 ( \30595 , RIfcae9f8_7009, \9449 );
and \U$21498 ( \30596 , RIfcb7260_7106, \9451 );
and \U$21499 ( \30597 , RIfea42b0_8212, \9453 );
and \U$21500 ( \30598 , RIdf33ce8_1966, \9455 );
and \U$21501 ( \30599 , RIdf31b28_1942, \9457 );
and \U$21502 ( \30600 , RIdf2fc38_1920, \9459 );
or \U$21503 ( \30601 , \30537 , \30538 , \30539 , \30540 , \30541 , \30542 , \30543 , \30544 , \30545 , \30546 , \30547 , \30548 , \30549 , \30550 , \30551 , \30552 , \30553 , \30554 , \30555 , \30556 , \30557 , \30558 , \30559 , \30560 , \30561 , \30562 , \30563 , \30564 , \30565 , \30566 , \30567 , \30568 , \30569 , \30570 , \30571 , \30572 , \30573 , \30574 , \30575 , \30576 , \30577 , \30578 , \30579 , \30580 , \30581 , \30582 , \30583 , \30584 , \30585 , \30586 , \30587 , \30588 , \30589 , \30590 , \30591 , \30592 , \30593 , \30594 , \30595 , \30596 , \30597 , \30598 , \30599 , \30600 );
and \U$21504 ( \30602 , RIee2c3f8_4962, \9462 );
and \U$21505 ( \30603 , RIfc4cfa0_5898, \9464 );
and \U$21506 ( \30604 , RIfc572c0_6014, \9466 );
and \U$21507 ( \30605 , RIfc4f430_5924, \9468 );
and \U$21508 ( \30606 , RIfea3e78_8209, \9470 );
and \U$21509 ( \30607 , RIdf28a50_1839, \9472 );
and \U$21510 ( \30608 , RIdf26b60_1817, \9474 );
and \U$21511 ( \30609 , RIdf250a8_1798, \9476 );
and \U$21512 ( \30610 , RIfc9b600_6790, \9478 );
and \U$21513 ( \30611 , RIfcb9df8_7137, \9480 );
and \U$21514 ( \30612 , RIdf23320_1777, \9482 );
and \U$21515 ( \30613 , RIfc86318_6549, \9484 );
and \U$21516 ( \30614 , RIfeabfd8_8273, \9486 );
and \U$21517 ( \30615 , RIdf201e8_1742, \9488 );
and \U$21518 ( \30616 , RIdf1b5f8_1688, \9490 );
and \U$21519 ( \30617 , RIdf19ca8_1670, \9492 );
and \U$21520 ( \30618 , RIdf17ae8_1646, \9494 );
and \U$21521 ( \30619 , RIdf14de8_1614, \9496 );
and \U$21522 ( \30620 , RIdf120e8_1582, \9498 );
and \U$21523 ( \30621 , RIdf0f3e8_1550, \9500 );
and \U$21524 ( \30622 , RIdf0c6e8_1518, \9502 );
and \U$21525 ( \30623 , RIdf099e8_1486, \9504 );
and \U$21526 ( \30624 , RIdf06ce8_1454, \9506 );
and \U$21527 ( \30625 , RIdf03fe8_1422, \9508 );
and \U$21528 ( \30626 , RIdefe5e8_1358, \9510 );
and \U$21529 ( \30627 , RIdefb8e8_1326, \9512 );
and \U$21530 ( \30628 , RIdef8be8_1294, \9514 );
and \U$21531 ( \30629 , RIdef5ee8_1262, \9516 );
and \U$21532 ( \30630 , RIdef31e8_1230, \9518 );
and \U$21533 ( \30631 , RIdef04e8_1198, \9520 );
and \U$21534 ( \30632 , RIdeed7e8_1166, \9522 );
and \U$21535 ( \30633 , RIdeeaae8_1134, \9524 );
and \U$21536 ( \30634 , RIfc89018_6581, \9526 );
and \U$21537 ( \30635 , RIfcc54c8_7267, \9528 );
and \U$21538 ( \30636 , RIfc89180_6582, \9530 );
and \U$21539 ( \30637 , RIfc4b380_5878, \9532 );
and \U$21540 ( \30638 , RIdee53b8_1072, \9534 );
and \U$21541 ( \30639 , RIdee34c8_1050, \9536 );
and \U$21542 ( \30640 , RIfea3d10_8208, \9538 );
and \U$21543 ( \30641 , RIdedf148_1002, \9540 );
and \U$21544 ( \30642 , RIfcae188_7003, \9542 );
and \U$21545 ( \30643 , RIfc4b0b0_5876, \9544 );
and \U$21546 ( \30644 , RIfc74870_6348, \9546 );
and \U$21547 ( \30645 , RIfce4968_7623, \9548 );
and \U$21548 ( \30646 , RIdeda288_946, \9550 );
and \U$21549 ( \30647 , RIded7c90_919, \9552 );
and \U$21550 ( \30648 , RIded5da0_897, \9554 );
and \U$21551 ( \30649 , RIded3640_869, \9556 );
and \U$21552 ( \30650 , RIded1318_844, \9558 );
and \U$21553 ( \30651 , RIdece618_812, \9560 );
and \U$21554 ( \30652 , RIdecb918_780, \9562 );
and \U$21555 ( \30653 , RIdec8c18_748, \9564 );
and \U$21556 ( \30654 , RIdeb5118_524, \9566 );
and \U$21557 ( \30655 , RIde98360_332, \9568 );
and \U$21558 ( \30656 , RIe16ed20_2638, \9570 );
and \U$21559 ( \30657 , RIe15ab18_2409, \9572 );
and \U$21560 ( \30658 , RIe144318_2153, \9574 );
and \U$21561 ( \30659 , RIdf38d10_2023, \9576 );
and \U$21562 ( \30660 , RIdf2d370_1891, \9578 );
and \U$21563 ( \30661 , RIdf1dbf0_1715, \9580 );
and \U$21564 ( \30662 , RIdf012e8_1390, \9582 );
and \U$21565 ( \30663 , RIdee7de8_1102, \9584 );
and \U$21566 ( \30664 , RIdedcb50_975, \9586 );
and \U$21567 ( \30665 , RIde7e2a8_205, \9588 );
or \U$21568 ( \30666 , \30602 , \30603 , \30604 , \30605 , \30606 , \30607 , \30608 , \30609 , \30610 , \30611 , \30612 , \30613 , \30614 , \30615 , \30616 , \30617 , \30618 , \30619 , \30620 , \30621 , \30622 , \30623 , \30624 , \30625 , \30626 , \30627 , \30628 , \30629 , \30630 , \30631 , \30632 , \30633 , \30634 , \30635 , \30636 , \30637 , \30638 , \30639 , \30640 , \30641 , \30642 , \30643 , \30644 , \30645 , \30646 , \30647 , \30648 , \30649 , \30650 , \30651 , \30652 , \30653 , \30654 , \30655 , \30656 , \30657 , \30658 , \30659 , \30660 , \30661 , \30662 , \30663 , \30664 , \30665 );
or \U$21569 ( \30667 , \30601 , \30666 );
_DC g65ce ( \30668_nG65ce , \30667 , \9597 );
and \U$21570 ( \30669 , RIe19e1b0_3176, \9059 );
and \U$21571 ( \30670 , RIe19b4b0_3144, \9061 );
and \U$21572 ( \30671 , RIfc9cf50_6808, \9063 );
and \U$21573 ( \30672 , RIe1987b0_3112, \9065 );
and \U$21574 ( \30673 , RIfc87290_6560, \9067 );
and \U$21575 ( \30674 , RIe195ab0_3080, \9069 );
and \U$21576 ( \30675 , RIe192db0_3048, \9071 );
and \U$21577 ( \30676 , RIe1900b0_3016, \9073 );
and \U$21578 ( \30677 , RIe18a6b0_2952, \9075 );
and \U$21579 ( \30678 , RIe1879b0_2920, \9077 );
and \U$21580 ( \30679 , RIfc842c0_6526, \9079 );
and \U$21581 ( \30680 , RIe184cb0_2888, \9081 );
and \U$21582 ( \30681 , RIfc83a50_6520, \9083 );
and \U$21583 ( \30682 , RIe181fb0_2856, \9085 );
and \U$21584 ( \30683 , RIe17f2b0_2824, \9087 );
and \U$21585 ( \30684 , RIe17c5b0_2792, \9089 );
and \U$21586 ( \30685 , RIfc9d0b8_6809, \9091 );
and \U$21587 ( \30686 , RIfc9e030_6820, \9093 );
and \U$21588 ( \30687 , RIe177420_2734, \9095 );
and \U$21589 ( \30688 , RIe176340_2722, \9097 );
and \U$21590 ( \30689 , RIfc4f700_5926, \9099 );
and \U$21591 ( \30690 , RIfcc4820_7258, \9101 );
and \U$21592 ( \30691 , RIfc4fb38_5929, \9103 );
and \U$21593 ( \30692 , RIfce8040_7662, \9105 );
and \U$21594 ( \30693 , RIee3c6b8_5146, \9107 );
and \U$21595 ( \30694 , RIee3b308_5132, \9109 );
and \U$21596 ( \30695 , RIfc812f0_6492, \9111 );
and \U$21597 ( \30696 , RIe174180_2698, \9113 );
and \U$21598 ( \30697 , RIfcd3028_7423, \9115 );
and \U$21599 ( \30698 , RIfc7f400_6470, \9117 );
and \U$21600 ( \30699 , RIfc46a60_5826, \9119 );
and \U$21601 ( \30700 , RIfc472d0_5832, \9121 );
and \U$21602 ( \30701 , RIf16cc58_5697, \9123 );
and \U$21603 ( \30702 , RIe224508_4703, \9125 );
and \U$21604 ( \30703 , RIfc7d3a8_6447, \9127 );
and \U$21605 ( \30704 , RIe221808_4671, \9129 );
and \U$21606 ( \30705 , RIfc97c58_6749, \9131 );
and \U$21607 ( \30706 , RIe21eb08_4639, \9133 );
and \U$21608 ( \30707 , RIe219108_4575, \9135 );
and \U$21609 ( \30708 , RIe216408_4543, \9137 );
and \U$21610 ( \30709 , RIfcdbe30_7524, \9139 );
and \U$21611 ( \30710 , RIe213708_4511, \9141 );
and \U$21612 ( \30711 , RIf169580_5658, \9143 );
and \U$21613 ( \30712 , RIe210a08_4479, \9145 );
and \U$21614 ( \30713 , RIfca4570_6892, \9147 );
and \U$21615 ( \30714 , RIe20dd08_4447, \9149 );
and \U$21616 ( \30715 , RIe20b008_4415, \9151 );
and \U$21617 ( \30716 , RIe208308_4383, \9153 );
and \U$21618 ( \30717 , RIfc7b080_6422, \9155 );
and \U$21619 ( \30718 , RIfc59cf0_6044, \9157 );
and \U$21620 ( \30719 , RIfea9b48_8247, \9159 );
and \U$21621 ( \30720 , RIfea4418_8213, \9161 );
and \U$21622 ( \30721 , RIfc79cd0_6408, \9163 );
and \U$21623 ( \30722 , RIfcd19a8_7407, \9165 );
and \U$21624 ( \30723 , RIfcc81c8_7299, \9167 );
and \U$21625 ( \30724 , RIf162230_5576, \9169 );
and \U$21626 ( \30725 , RIf160778_5557, \9171 );
and \U$21627 ( \30726 , RIf15e888_5535, \9173 );
and \U$21628 ( \30727 , RIfea4580_8214, \9175 );
and \U$21629 ( \30728 , RIfea46e8_8215, \9177 );
and \U$21630 ( \30729 , RIfc77f48_6387, \9179 );
and \U$21631 ( \30730 , RIfc41fd8_5773, \9181 );
and \U$21632 ( \30731 , RIf15aaa8_5491, \9183 );
and \U$21633 ( \30732 , RIfc7c430_6436, \9185 );
or \U$21634 ( \30733 , \30669 , \30670 , \30671 , \30672 , \30673 , \30674 , \30675 , \30676 , \30677 , \30678 , \30679 , \30680 , \30681 , \30682 , \30683 , \30684 , \30685 , \30686 , \30687 , \30688 , \30689 , \30690 , \30691 , \30692 , \30693 , \30694 , \30695 , \30696 , \30697 , \30698 , \30699 , \30700 , \30701 , \30702 , \30703 , \30704 , \30705 , \30706 , \30707 , \30708 , \30709 , \30710 , \30711 , \30712 , \30713 , \30714 , \30715 , \30716 , \30717 , \30718 , \30719 , \30720 , \30721 , \30722 , \30723 , \30724 , \30725 , \30726 , \30727 , \30728 , \30729 , \30730 , \30731 , \30732 );
and \U$21635 ( \30734 , RIf159158_5473, \9188 );
and \U$21636 ( \30735 , RIf157f10_5460, \9190 );
and \U$21637 ( \30736 , RIfcae890_7008, \9192 );
and \U$21638 ( \30737 , RIe1faa78_4229, \9194 );
and \U$21639 ( \30738 , RIfc4a840_5870, \9196 );
and \U$21640 ( \30739 , RIfc4ed28_5919, \9198 );
and \U$21641 ( \30740 , RIfce0e58_7581, \9200 );
and \U$21642 ( \30741 , RIe1f5ff0_4176, \9202 );
and \U$21643 ( \30742 , RIf153758_5409, \9204 );
and \U$21644 ( \30743 , RIf151f70_5392, \9206 );
and \U$21645 ( \30744 , RIfccb468_7335, \9208 );
and \U$21646 ( \30745 , RIe1f3cc8_4151, \9210 );
and \U$21647 ( \30746 , RIfc68ed0_6216, \9212 );
and \U$21648 ( \30747 , RIfc6d250_6264, \9214 );
and \U$21649 ( \30748 , RIfca9ca0_6954, \9216 );
and \U$21650 ( \30749 , RIe1ee9d0_4092, \9218 );
and \U$21651 ( \30750 , RIe1ec270_4064, \9220 );
and \U$21652 ( \30751 , RIe1e9570_4032, \9222 );
and \U$21653 ( \30752 , RIe1e6870_4000, \9224 );
and \U$21654 ( \30753 , RIe1e3b70_3968, \9226 );
and \U$21655 ( \30754 , RIe1e0e70_3936, \9228 );
and \U$21656 ( \30755 , RIe1de170_3904, \9230 );
and \U$21657 ( \30756 , RIe1db470_3872, \9232 );
and \U$21658 ( \30757 , RIe1d8770_3840, \9234 );
and \U$21659 ( \30758 , RIe1d2d70_3776, \9236 );
and \U$21660 ( \30759 , RIe1d0070_3744, \9238 );
and \U$21661 ( \30760 , RIe1cd370_3712, \9240 );
and \U$21662 ( \30761 , RIe1ca670_3680, \9242 );
and \U$21663 ( \30762 , RIe1c7970_3648, \9244 );
and \U$21664 ( \30763 , RIe1c4c70_3616, \9246 );
and \U$21665 ( \30764 , RIe1c1f70_3584, \9248 );
and \U$21666 ( \30765 , RIe1bf270_3552, \9250 );
and \U$21667 ( \30766 , RIfc784e8_6391, \9252 );
and \U$21668 ( \30767 , RIfcbef88_7195, \9254 );
and \U$21669 ( \30768 , RIe1b9ca8_3491, \9256 );
and \U$21670 ( \30769 , RIe1b7ae8_3467, \9258 );
and \U$21671 ( \30770 , RIfcc20c0_7230, \9260 );
and \U$21672 ( \30771 , RIfca6190_6912, \9262 );
and \U$21673 ( \30772 , RIe1b5928_3443, \9264 );
and \U$21674 ( \30773 , RIe1b4410_3428, \9266 );
and \U$21675 ( \30774 , RIfcb81d8_7117, \9268 );
and \U$21676 ( \30775 , RIfcc5090_7264, \9270 );
and \U$21677 ( \30776 , RIe1b2d90_3412, \9272 );
and \U$21678 ( \30777 , RIe1b1440_3394, \9274 );
and \U$21679 ( \30778 , RIfcd5350_7448, \9276 );
and \U$21680 ( \30779 , RIfcb9588_7131, \9278 );
and \U$21681 ( \30780 , RIe1acc88_3343, \9280 );
and \U$21682 ( \30781 , RIe1ab4a0_3326, \9282 );
and \U$21683 ( \30782 , RIe1a95b0_3304, \9284 );
and \U$21684 ( \30783 , RIe1a68b0_3272, \9286 );
and \U$21685 ( \30784 , RIe1a3bb0_3240, \9288 );
and \U$21686 ( \30785 , RIe1a0eb0_3208, \9290 );
and \U$21687 ( \30786 , RIe18d3b0_2984, \9292 );
and \U$21688 ( \30787 , RIe1798b0_2760, \9294 );
and \U$21689 ( \30788 , RIe227208_4735, \9296 );
and \U$21690 ( \30789 , RIe21be08_4607, \9298 );
and \U$21691 ( \30790 , RIe205608_4351, \9300 );
and \U$21692 ( \30791 , RIe1ff668_4283, \9302 );
and \U$21693 ( \30792 , RIe1f8a20_4206, \9304 );
and \U$21694 ( \30793 , RIe1f1568_4123, \9306 );
and \U$21695 ( \30794 , RIe1d5a70_3808, \9308 );
and \U$21696 ( \30795 , RIe1bc570_3520, \9310 );
and \U$21697 ( \30796 , RIe1af3e8_3371, \9312 );
and \U$21698 ( \30797 , RIe171a20_2670, \9314 );
or \U$21699 ( \30798 , \30734 , \30735 , \30736 , \30737 , \30738 , \30739 , \30740 , \30741 , \30742 , \30743 , \30744 , \30745 , \30746 , \30747 , \30748 , \30749 , \30750 , \30751 , \30752 , \30753 , \30754 , \30755 , \30756 , \30757 , \30758 , \30759 , \30760 , \30761 , \30762 , \30763 , \30764 , \30765 , \30766 , \30767 , \30768 , \30769 , \30770 , \30771 , \30772 , \30773 , \30774 , \30775 , \30776 , \30777 , \30778 , \30779 , \30780 , \30781 , \30782 , \30783 , \30784 , \30785 , \30786 , \30787 , \30788 , \30789 , \30790 , \30791 , \30792 , \30793 , \30794 , \30795 , \30796 , \30797 );
or \U$21700 ( \30799 , \30733 , \30798 );
_DC g65cf ( \30800_nG65cf , \30799 , \9323 );
and g65d0 ( \30801_nG65d0 , \30668_nG65ce , \30800_nG65cf );
buf \U$21701 ( \30802 , \30801_nG65d0 );
and \U$21702 ( \30803 , \30802 , \10691 );
nor \U$21703 ( \30804 , \30536 , \30803 );
xnor \U$21704 ( \30805 , \30804 , \10980 );
not \U$21705 ( \30806 , \30247 );
_DC g62df ( \30807_nG62df , \30667 , \9597 );
_DC g6363 ( \30808_nG6363 , \30799 , \9323 );
xor g6364 ( \30809_nG6364 , \30807_nG62df , \30808_nG6363 );
buf \U$21706 ( \30810 , \30809_nG6364 );
and \U$21707 ( \30811 , \30245 , \29067 );
not \U$21708 ( \30812 , \30811 );
and \U$21709 ( \30813 , \30810 , \30812 );
and \U$21710 ( \30814 , \30806 , \30813 );
xor \U$21711 ( \30815 , \30805 , \30814 );
and \U$21712 ( \30816 , \11270 , \29070 );
and \U$21713 ( \30817 , \11586 , \28526 );
nor \U$21714 ( \30818 , \30816 , \30817 );
xnor \U$21715 ( \30819 , \30818 , \29076 );
xor \U$21716 ( \30820 , \30815 , \30819 );
xor \U$21717 ( \30821 , \30810 , \30245 );
not \U$21718 ( \30822 , \30246 );
and \U$21719 ( \30823 , \30821 , \30822 );
and \U$21720 ( \30824 , \10687 , \30823 );
and \U$21721 ( \30825 , \10988 , \30246 );
nor \U$21722 ( \30826 , \30824 , \30825 );
xnor \U$21723 ( \30827 , \30826 , \30813 );
xor \U$21724 ( \30828 , \30820 , \30827 );
xor \U$21725 ( \30829 , \30535 , \30828 );
and \U$21726 ( \30830 , \30333 , \30337 );
and \U$21727 ( \30831 , \30337 , \30352 );
and \U$21728 ( \30832 , \30333 , \30352 );
or \U$21729 ( \30833 , \30830 , \30831 , \30832 );
and \U$21730 ( \30834 , \29974 , \29978 );
and \U$21731 ( \30835 , \29978 , \30247 );
and \U$21732 ( \30836 , \29974 , \30247 );
or \U$21733 ( \30837 , \30834 , \30835 , \30836 );
and \U$21734 ( \30838 , \30271 , \30275 );
and \U$21735 ( \30839 , \30275 , \30280 );
and \U$21736 ( \30840 , \30271 , \30280 );
or \U$21737 ( \30841 , \30838 , \30839 , \30840 );
xor \U$21738 ( \30842 , \30837 , \30841 );
and \U$21739 ( \30843 , \30342 , \30346 );
and \U$21740 ( \30844 , \30346 , \30351 );
and \U$21741 ( \30845 , \30342 , \30351 );
or \U$21742 ( \30846 , \30843 , \30844 , \30845 );
xor \U$21743 ( \30847 , \30842 , \30846 );
xor \U$21744 ( \30848 , \30833 , \30847 );
and \U$21745 ( \30849 , \30252 , \30256 );
and \U$21746 ( \30850 , \30256 , \30261 );
and \U$21747 ( \30851 , \30252 , \30261 );
or \U$21748 ( \30852 , \30849 , \30850 , \30851 );
and \U$21749 ( \30853 , \30301 , \30305 );
and \U$21750 ( \30854 , \30305 , \30310 );
and \U$21751 ( \30855 , \30301 , \30310 );
or \U$21752 ( \30856 , \30853 , \30854 , \30855 );
xor \U$21753 ( \30857 , \30852 , \30856 );
and \U$21754 ( \30858 , \28534 , \11574 );
and \U$21755 ( \30859 , \29084 , \11278 );
nor \U$21756 ( \30860 , \30858 , \30859 );
xnor \U$21757 ( \30861 , \30860 , \11580 );
and \U$21758 ( \30862 , \25272 , \14054 );
and \U$21759 ( \30863 , \25815 , \13692 );
nor \U$21760 ( \30864 , \30862 , \30863 );
xnor \U$21761 ( \30865 , \30864 , \14035 );
xor \U$21762 ( \30866 , \30861 , \30865 );
and \U$21763 ( \30867 , \19032 , \19534 );
and \U$21764 ( \30868 , \19558 , \19045 );
nor \U$21765 ( \30869 , \30867 , \30868 );
xnor \U$21766 ( \30870 , \30869 , \19540 );
xor \U$21767 ( \30871 , \30866 , \30870 );
xor \U$21768 ( \30872 , \30857 , \30871 );
xor \U$21769 ( \30873 , \30848 , \30872 );
xor \U$21770 ( \30874 , \30829 , \30873 );
and \U$21771 ( \30875 , \30292 , \30296 );
and \U$21772 ( \30876 , \30296 , \30311 );
and \U$21773 ( \30877 , \30292 , \30311 );
or \U$21774 ( \30878 , \30875 , \30876 , \30877 );
and \U$21775 ( \30879 , \30317 , \30328 );
and \U$21776 ( \30880 , \30328 , \30353 );
and \U$21777 ( \30881 , \30317 , \30353 );
or \U$21778 ( \30882 , \30879 , \30880 , \30881 );
xor \U$21779 ( \30883 , \30878 , \30882 );
and \U$21780 ( \30884 , \23617 , \15336 );
and \U$21781 ( \30885 , \24199 , \14963 );
nor \U$21782 ( \30886 , \30884 , \30885 );
xnor \U$21783 ( \30887 , \30886 , \15342 );
and \U$21784 ( \30888 , \17627 , \21005 );
and \U$21785 ( \30889 , \18035 , \20557 );
nor \U$21786 ( \30890 , \30888 , \30889 );
xnor \U$21787 ( \30891 , \30890 , \21011 );
xor \U$21788 ( \30892 , \30887 , \30891 );
and \U$21789 ( \30893 , \16267 , \22542 );
and \U$21790 ( \30894 , \16655 , \22103 );
nor \U$21791 ( \30895 , \30893 , \30894 );
xnor \U$21792 ( \30896 , \30895 , \22548 );
xor \U$21793 ( \30897 , \30892 , \30896 );
and \U$21794 ( \30898 , \26829 , \12790 );
and \U$21795 ( \30899 , \27313 , \12461 );
nor \U$21796 ( \30900 , \30898 , \30899 );
xnor \U$21797 ( \30901 , \30900 , \12780 );
and \U$21798 ( \30902 , \22090 , \16635 );
and \U$21799 ( \30903 , \22556 , \16301 );
nor \U$21800 ( \30904 , \30902 , \30903 );
xnor \U$21801 ( \30905 , \30904 , \16625 );
xor \U$21802 ( \30906 , \30901 , \30905 );
and \U$21803 ( \30907 , \14950 , \24138 );
and \U$21804 ( \30908 , \15321 , \23630 );
nor \U$21805 ( \30909 , \30907 , \30908 );
xnor \U$21806 ( \30910 , \30909 , \24144 );
xor \U$21807 ( \30911 , \30906 , \30910 );
xor \U$21808 ( \30912 , \30897 , \30911 );
and \U$21809 ( \30913 , \20544 , \18090 );
and \U$21810 ( \30914 , \21033 , \17655 );
nor \U$21811 ( \30915 , \30913 , \30914 );
xnor \U$21812 ( \30916 , \30915 , \18046 );
and \U$21813 ( \30917 , \13679 , \25826 );
and \U$21814 ( \30918 , \14024 , \25264 );
nor \U$21815 ( \30919 , \30917 , \30918 );
xnor \U$21816 ( \30920 , \30919 , \25773 );
xor \U$21817 ( \30921 , \30916 , \30920 );
and \U$21818 ( \30922 , \12448 , \27397 );
and \U$21819 ( \30923 , \12769 , \26807 );
nor \U$21820 ( \30924 , \30922 , \30923 );
xnor \U$21821 ( \30925 , \30924 , \27295 );
xor \U$21822 ( \30926 , \30921 , \30925 );
xor \U$21823 ( \30927 , \30912 , \30926 );
xor \U$21824 ( \30928 , \30883 , \30927 );
xor \U$21825 ( \30929 , \30874 , \30928 );
xor \U$21826 ( \30930 , \30526 , \30929 );
and \U$21827 ( \30931 , \29961 , \30283 );
and \U$21828 ( \30932 , \30283 , \30355 );
and \U$21829 ( \30933 , \29961 , \30355 );
or \U$21830 ( \30934 , \30931 , \30932 , \30933 );
xor \U$21831 ( \30935 , \30930 , \30934 );
and \U$21832 ( \30936 , \30356 , \30360 );
and \U$21833 ( \30937 , \30361 , \30364 );
or \U$21834 ( \30938 , \30936 , \30937 );
xor \U$21835 ( \30939 , \30935 , \30938 );
buf g9bb7 ( \30940_nG9bb7 , \30939 );
and \U$21836 ( \30941 , \10704 , \30940_nG9bb7 );
or \U$21837 ( \30942 , \30517 , \30941 );
xor \U$21838 ( \30943 , \10703 , \30942 );
buf \U$21839 ( \30944 , \30943 );
buf \U$21841 ( \30945 , \30944 );
xor \U$21842 ( \30946 , \30516 , \30945 );
buf \U$21843 ( \30947 , \30946 );
and \U$21844 ( \30948 , \29949 , \29955 );
and \U$21845 ( \30949 , \29949 , \30371 );
and \U$21846 ( \30950 , \29955 , \30371 );
or \U$21847 ( \30951 , \30948 , \30949 , \30950 );
buf \U$21848 ( \30952 , \30951 );
xor \U$21849 ( \30953 , \30947 , \30952 );
and \U$21850 ( \30954 , \29916 , \29922 );
and \U$21851 ( \30955 , \29916 , \29929 );
and \U$21852 ( \30956 , \29922 , \29929 );
or \U$21853 ( \30957 , \30954 , \30955 , \30956 );
buf \U$21854 ( \30958 , \30957 );
and \U$21855 ( \30959 , \29849 , \29856 );
buf \U$21856 ( \30960 , \30959 );
buf \U$21858 ( \30961 , \30960 );
and \U$21859 ( \30962 , \28118 , \11283_nG9c08 );
and \U$21860 ( \30963 , \28115 , \11598_nG9c05 );
or \U$21861 ( \30964 , \30962 , \30963 );
xor \U$21862 ( \30965 , \28114 , \30964 );
buf \U$21863 ( \30966 , \30965 );
buf \U$21865 ( \30967 , \30966 );
xor \U$21866 ( \30968 , \30961 , \30967 );
buf \U$21867 ( \30969 , \30968 );
and \U$21868 ( \30970 , \29853 , \10694_nG9c0e );
and \U$21869 ( \30971 , \29850 , \10995_nG9c0b );
or \U$21870 ( \30972 , \30970 , \30971 );
xor \U$21871 ( \30973 , \29849 , \30972 );
buf \U$21872 ( \30974 , \30973 );
buf \U$21874 ( \30975 , \30974 );
xor \U$21875 ( \30976 , \30969 , \30975 );
and \U$21876 ( \30977 , \26431 , \12470_nG9c02 );
and \U$21877 ( \30978 , \26428 , \12801_nG9bff );
or \U$21878 ( \30979 , \30977 , \30978 );
xor \U$21879 ( \30980 , \26427 , \30979 );
buf \U$21880 ( \30981 , \30980 );
buf \U$21882 ( \30982 , \30981 );
xor \U$21883 ( \30983 , \30976 , \30982 );
buf \U$21884 ( \30984 , \30983 );
xor \U$21885 ( \30985 , \30958 , \30984 );
and \U$21886 ( \30986 , \21658 , \16315_nG9bf0 );
and \U$21887 ( \30987 , \21655 , \16680_nG9bed );
or \U$21888 ( \30988 , \30986 , \30987 );
xor \U$21889 ( \30989 , \21654 , \30988 );
buf \U$21890 ( \30990 , \30989 );
buf \U$21892 ( \30991 , \30990 );
xor \U$21893 ( \30992 , \30985 , \30991 );
buf \U$21894 ( \30993 , \30992 );
and \U$21895 ( \30994 , \18702 , \19091_nG9be4 );
and \U$21896 ( \30995 , \18699 , \19586_nG9be1 );
or \U$21897 ( \30996 , \30994 , \30995 );
xor \U$21898 ( \30997 , \18698 , \30996 );
buf \U$21899 ( \30998 , \30997 );
buf \U$21901 ( \30999 , \30998 );
xor \U$21902 ( \31000 , \30993 , \30999 );
and \U$21903 ( \31001 , \17297 , \20608_nG9bde );
and \U$21904 ( \31002 , \17294 , \21086_nG9bdb );
or \U$21905 ( \31003 , \31001 , \31002 );
xor \U$21906 ( \31004 , \17293 , \31003 );
buf \U$21907 ( \31005 , \31004 );
buf \U$21909 ( \31006 , \31005 );
xor \U$21910 ( \31007 , \31000 , \31006 );
buf \U$21911 ( \31008 , \31007 );
and \U$21912 ( \31009 , \13370 , \25298_nG9bcc );
and \U$21913 ( \31010 , \13367 , \25860_nG9bc9 );
or \U$21914 ( \31011 , \31009 , \31010 );
xor \U$21915 ( \31012 , \13366 , \31011 );
buf \U$21916 ( \31013 , \31012 );
buf \U$21918 ( \31014 , \31013 );
xor \U$21919 ( \31015 , \31008 , \31014 );
and \U$21920 ( \31016 , \10421 , \28602_nG9bc0 );
and \U$21921 ( \31017 , \10418 , \29179_nG9bbd );
or \U$21922 ( \31018 , \31016 , \31017 );
xor \U$21923 ( \31019 , \10417 , \31018 );
buf \U$21924 ( \31020 , \31019 );
buf \U$21926 ( \31021 , \31020 );
xor \U$21927 ( \31022 , \31015 , \31021 );
buf \U$21928 ( \31023 , \31022 );
xor \U$21929 ( \31024 , \30953 , \31023 );
buf \U$21930 ( \31025 , \31024 );
and \U$21931 ( \31026 , \29870 , \29903 );
and \U$21932 ( \31027 , \29870 , \30373 );
and \U$21933 ( \31028 , \29903 , \30373 );
or \U$21934 ( \31029 , \31026 , \31027 , \31028 );
buf \U$21935 ( \31030 , \31029 );
xor \U$21936 ( \31031 , \31025 , \31030 );
and \U$21937 ( \31032 , \30419 , \30425 );
and \U$21938 ( \31033 , \30419 , \30432 );
and \U$21939 ( \31034 , \30425 , \30432 );
or \U$21940 ( \31035 , \31032 , \31033 , \31034 );
buf \U$21941 ( \31036 , \31035 );
and \U$21942 ( \31037 , \14631 , \23696_nG9bd2 );
and \U$21943 ( \31038 , \14628 , \24226_nG9bcf );
or \U$21944 ( \31039 , \31037 , \31038 );
xor \U$21945 ( \31040 , \14627 , \31039 );
buf \U$21946 ( \31041 , \31040 );
buf \U$21948 ( \31042 , \31041 );
xor \U$21949 ( \31043 , \31036 , \31042 );
and \U$21950 ( \31044 , \12157 , \26887_nG9bc6 );
and \U$21951 ( \31045 , \12154 , \27416_nG9bc3 );
or \U$21952 ( \31046 , \31044 , \31045 );
xor \U$21953 ( \31047 , \12153 , \31046 );
buf \U$21954 ( \31048 , \31047 );
buf \U$21956 ( \31049 , \31048 );
xor \U$21957 ( \31050 , \31043 , \31049 );
buf \U$21958 ( \31051 , \31050 );
and \U$21959 ( \31052 , \30391 , \30434 );
and \U$21960 ( \31053 , \30391 , \30441 );
and \U$21961 ( \31054 , \30434 , \30441 );
or \U$21962 ( \31055 , \31052 , \31053 , \31054 );
buf \U$21963 ( \31056 , \31055 );
xor \U$21964 ( \31057 , \31051 , \31056 );
and \U$21965 ( \31058 , \29880 , \29886 );
and \U$21966 ( \31059 , \29880 , \29893 );
and \U$21967 ( \31060 , \29886 , \29893 );
or \U$21968 ( \31061 , \31058 , \31059 , \31060 );
buf \U$21969 ( \31062 , \31061 );
xor \U$21970 ( \31063 , \31057 , \31062 );
buf \U$21971 ( \31064 , \31063 );
and \U$21972 ( \31065 , \30386 , \30443 );
and \U$21973 ( \31066 , \30386 , \30449 );
and \U$21974 ( \31067 , \30443 , \30449 );
or \U$21975 ( \31068 , \31065 , \31066 , \31067 );
buf \U$21976 ( \31069 , \31068 );
xor \U$21977 ( \31070 , \31064 , \31069 );
and \U$21978 ( \31071 , \29875 , \29895 );
and \U$21979 ( \31072 , \29875 , \29901 );
and \U$21980 ( \31073 , \29895 , \29901 );
or \U$21981 ( \31074 , \31071 , \31072 , \31073 );
buf \U$21982 ( \31075 , \31074 );
xor \U$21983 ( \31076 , \31070 , \31075 );
buf \U$21984 ( \31077 , \31076 );
xor \U$21985 ( \31078 , \31031 , \31077 );
and \U$21986 ( \31079 , \30465 , \31078 );
and \U$21987 ( \31080 , \30455 , \30459 );
and \U$21988 ( \31081 , \30455 , \30464 );
and \U$21989 ( \31082 , \30459 , \30464 );
or \U$21990 ( \31083 , \31080 , \31081 , \31082 );
xor \U$21991 ( \31084 , \31079 , \31083 );
and \U$21992 ( \31085 , RIdec6350_719, \9059 );
and \U$21993 ( \31086 , RIdec3650_687, \9061 );
and \U$21994 ( \31087 , RIfcaf3d0_7016, \9063 );
and \U$21995 ( \31088 , RIdec0950_655, \9065 );
and \U$21996 ( \31089 , RIfc6a280_6230, \9067 );
and \U$21997 ( \31090 , RIdebdc50_623, \9069 );
and \U$21998 ( \31091 , RIdebaf50_591, \9071 );
and \U$21999 ( \31092 , RIdeb8250_559, \9073 );
and \U$22000 ( \31093 , RIfc42f50_5784, \9075 );
and \U$22001 ( \31094 , RIdeb2850_495, \9077 );
and \U$22002 ( \31095 , RIfc981f8_6753, \9079 );
and \U$22003 ( \31096 , RIdeafb50_463, \9081 );
and \U$22004 ( \31097 , RIfc8c6f0_6620, \9083 );
and \U$22005 ( \31098 , RIdeac838_431, \9085 );
and \U$22006 ( \31099 , RIdea5f38_399, \9087 );
and \U$22007 ( \31100 , RIde9f638_367, \9089 );
and \U$22008 ( \31101 , RIee1d4e8_4792, \9091 );
and \U$22009 ( \31102 , RIfcda648_7507, \9093 );
and \U$22010 ( \31103 , RIfcc6440_7278, \9095 );
and \U$22011 ( \31104 , RIfcd5620_7450, \9097 );
and \U$22012 ( \31105 , RIde92ac8_305, \9099 );
and \U$22013 ( \31106 , RIfea34a0_8202, \9101 );
and \U$22014 ( \31107 , RIfea31d0_8200, \9103 );
and \U$22015 ( \31108 , RIfea3338_8201, \9105 );
and \U$22016 ( \31109 , RIfcb6b58_7101, \9107 );
and \U$22017 ( \31110 , RIfcb6888_7099, \9109 );
and \U$22018 ( \31111 , RIfc9dd60_6818, \9111 );
and \U$22019 ( \31112 , RIee19708_4748, \9113 );
and \U$22020 ( \31113 , RIfc50c18_5941, \9115 );
and \U$22021 ( \31114 , RIe16c458_2609, \9117 );
and \U$22022 ( \31115 , RIfc80a80_6486, \9119 );
and \U$22023 ( \31116 , RIfec62e8_8375, \9121 );
and \U$22024 ( \31117 , RIe166350_2540, \9123 );
and \U$22025 ( \31118 , RIe163650_2508, \9125 );
and \U$22026 ( \31119 , RIee37d98_5094, \9127 );
and \U$22027 ( \31120 , RIe160950_2476, \9129 );
and \U$22028 ( \31121 , RIfcaa678_6961, \9131 );
and \U$22029 ( \31122 , RIe15dc50_2444, \9133 );
and \U$22030 ( \31123 , RIe158250_2380, \9135 );
and \U$22031 ( \31124 , RIe155550_2348, \9137 );
and \U$22032 ( \31125 , RIfea3ba8_8207, \9139 );
and \U$22033 ( \31126 , RIe152850_2316, \9141 );
and \U$22034 ( \31127 , RIee35638_5066, \9143 );
and \U$22035 ( \31128 , RIe14fb50_2284, \9145 );
and \U$22036 ( \31129 , RIfc62f30_6148, \9147 );
and \U$22037 ( \31130 , RIe14ce50_2252, \9149 );
and \U$22038 ( \31131 , RIe14a150_2220, \9151 );
and \U$22039 ( \31132 , RIe147450_2188, \9153 );
and \U$22040 ( \31133 , RIfc97f28_6751, \9155 );
and \U$22041 ( \31134 , RIfc89888_6587, \9157 );
and \U$22042 ( \31135 , RIfc8f558_6653, \9159 );
and \U$22043 ( \31136 , RIfc52838_5961, \9161 );
and \U$22044 ( \31137 , RIe141bb8_2125, \9163 );
and \U$22045 ( \31138 , RIe13f890_2100, \9165 );
and \U$22046 ( \31139 , RIdf3d798_2076, \9167 );
and \U$22047 ( \31140 , RIdf3b308_2050, \9169 );
and \U$22048 ( \31141 , RIee30a48_5012, \9171 );
and \U$22049 ( \31142 , RIfc568e8_6007, \9173 );
and \U$22050 ( \31143 , RIee2e9f0_4989, \9175 );
and \U$22051 ( \31144 , RIee2dbe0_4979, \9177 );
and \U$22052 ( \31145 , RIdf365b0_1995, \9179 );
and \U$22053 ( \31146 , RIfea38d8_8205, \9181 );
and \U$22054 ( \31147 , RIfea3a40_8206, \9183 );
and \U$22055 ( \31148 , RIdf2ff08_1922, \9185 );
or \U$22056 ( \31149 , \31085 , \31086 , \31087 , \31088 , \31089 , \31090 , \31091 , \31092 , \31093 , \31094 , \31095 , \31096 , \31097 , \31098 , \31099 , \31100 , \31101 , \31102 , \31103 , \31104 , \31105 , \31106 , \31107 , \31108 , \31109 , \31110 , \31111 , \31112 , \31113 , \31114 , \31115 , \31116 , \31117 , \31118 , \31119 , \31120 , \31121 , \31122 , \31123 , \31124 , \31125 , \31126 , \31127 , \31128 , \31129 , \31130 , \31131 , \31132 , \31133 , \31134 , \31135 , \31136 , \31137 , \31138 , \31139 , \31140 , \31141 , \31142 , \31143 , \31144 , \31145 , \31146 , \31147 , \31148 );
and \U$22057 ( \31150 , RIee2c6c8_4964, \9188 );
and \U$22058 ( \31151 , RIee2ac10_4945, \9190 );
and \U$22059 ( \31152 , RIee29590_4929, \9192 );
and \U$22060 ( \31153 , RIee28348_4916, \9194 );
and \U$22061 ( \31154 , RIdf2ad78_1864, \9196 );
and \U$22062 ( \31155 , RIdf28e88_1842, \9198 );
and \U$22063 ( \31156 , RIfea3608_8203, \9200 );
and \U$22064 ( \31157 , RIfea3770_8204, \9202 );
and \U$22065 ( \31158 , RIfcc0d10_7216, \9204 );
and \U$22066 ( \31159 , RIfc75c20_6362, \9206 );
and \U$22067 ( \31160 , RIfca50b0_6900, \9208 );
and \U$22068 ( \31161 , RIfc74e10_6352, \9210 );
and \U$22069 ( \31162 , RIfcc9410_7312, \9212 );
and \U$22070 ( \31163 , RIdf20620_1745, \9214 );
and \U$22071 ( \31164 , RIfc73628_6335, \9216 );
and \U$22072 ( \31165 , RIdf1a0e0_1673, \9218 );
and \U$22073 ( \31166 , RIdf17f20_1649, \9220 );
and \U$22074 ( \31167 , RIdf15220_1617, \9222 );
and \U$22075 ( \31168 , RIdf12520_1585, \9224 );
and \U$22076 ( \31169 , RIdf0f820_1553, \9226 );
and \U$22077 ( \31170 , RIdf0cb20_1521, \9228 );
and \U$22078 ( \31171 , RIdf09e20_1489, \9230 );
and \U$22079 ( \31172 , RIdf07120_1457, \9232 );
and \U$22080 ( \31173 , RIdf04420_1425, \9234 );
and \U$22081 ( \31174 , RIdefea20_1361, \9236 );
and \U$22082 ( \31175 , RIdefbd20_1329, \9238 );
and \U$22083 ( \31176 , RIdef9020_1297, \9240 );
and \U$22084 ( \31177 , RIdef6320_1265, \9242 );
and \U$22085 ( \31178 , RIdef3620_1233, \9244 );
and \U$22086 ( \31179 , RIdef0920_1201, \9246 );
and \U$22087 ( \31180 , RIdeedc20_1169, \9248 );
and \U$22088 ( \31181 , RIdeeaf20_1137, \9250 );
and \U$22089 ( \31182 , RIfcab8c0_6974, \9252 );
and \U$22090 ( \31183 , RIfc7c598_6437, \9254 );
and \U$22091 ( \31184 , RIfc5beb0_6068, \9256 );
and \U$22092 ( \31185 , RIfc58ee0_6034, \9258 );
and \U$22093 ( \31186 , RIdee5688_1074, \9260 );
and \U$22094 ( \31187 , RIdee3798_1052, \9262 );
and \U$22095 ( \31188 , RIdee15d8_1028, \9264 );
and \U$22096 ( \31189 , RIdedf580_1005, \9266 );
and \U$22097 ( \31190 , RIfcb3048_7059, \9268 );
and \U$22098 ( \31191 , RIfc72ae8_6327, \9270 );
and \U$22099 ( \31192 , RIfca3d00_6886, \9272 );
and \U$22100 ( \31193 , RIfcb6450_7096, \9274 );
and \U$22101 ( \31194 , RIdeda558_948, \9276 );
and \U$22102 ( \31195 , RIded7f60_921, \9278 );
and \U$22103 ( \31196 , RIfea3068_8199, \9280 );
and \U$22104 ( \31197 , RIded3a78_872, \9282 );
and \U$22105 ( \31198 , RIded1750_847, \9284 );
and \U$22106 ( \31199 , RIdecea50_815, \9286 );
and \U$22107 ( \31200 , RIdecbd50_783, \9288 );
and \U$22108 ( \31201 , RIdec9050_751, \9290 );
and \U$22109 ( \31202 , RIdeb5550_527, \9292 );
and \U$22110 ( \31203 , RIde98d38_335, \9294 );
and \U$22111 ( \31204 , RIe16f158_2641, \9296 );
and \U$22112 ( \31205 , RIe15af50_2412, \9298 );
and \U$22113 ( \31206 , RIe144750_2156, \9300 );
and \U$22114 ( \31207 , RIdf39148_2026, \9302 );
and \U$22115 ( \31208 , RIdf2d7a8_1894, \9304 );
and \U$22116 ( \31209 , RIdf1e028_1718, \9306 );
and \U$22117 ( \31210 , RIdf01720_1393, \9308 );
and \U$22118 ( \31211 , RIdee8220_1105, \9310 );
and \U$22119 ( \31212 , RIdedcf88_978, \9312 );
and \U$22120 ( \31213 , RIde7ec80_208, \9314 );
or \U$22121 ( \31214 , \31150 , \31151 , \31152 , \31153 , \31154 , \31155 , \31156 , \31157 , \31158 , \31159 , \31160 , \31161 , \31162 , \31163 , \31164 , \31165 , \31166 , \31167 , \31168 , \31169 , \31170 , \31171 , \31172 , \31173 , \31174 , \31175 , \31176 , \31177 , \31178 , \31179 , \31180 , \31181 , \31182 , \31183 , \31184 , \31185 , \31186 , \31187 , \31188 , \31189 , \31190 , \31191 , \31192 , \31193 , \31194 , \31195 , \31196 , \31197 , \31198 , \31199 , \31200 , \31201 , \31202 , \31203 , \31204 , \31205 , \31206 , \31207 , \31208 , \31209 , \31210 , \31211 , \31212 , \31213 );
or \U$22122 ( \31215 , \31149 , \31214 );
_DC g2235 ( \31216_nG2235 , \31215 , \9323 );
buf \U$22123 ( \31217 , \31216_nG2235 );
and \U$22124 ( \31218 , RIe19e5e8_3179, \9333 );
and \U$22125 ( \31219 , RIe19b8e8_3147, \9335 );
and \U$22126 ( \31220 , RIfca84b8_6937, \9337 );
and \U$22127 ( \31221 , RIe198be8_3115, \9339 );
and \U$22128 ( \31222 , RIfc846f8_6529, \9341 );
and \U$22129 ( \31223 , RIe195ee8_3083, \9343 );
and \U$22130 ( \31224 , RIe1931e8_3051, \9345 );
and \U$22131 ( \31225 , RIe1904e8_3019, \9347 );
and \U$22132 ( \31226 , RIe18aae8_2955, \9349 );
and \U$22133 ( \31227 , RIe187de8_2923, \9351 );
and \U$22134 ( \31228 , RIfce2be0_7602, \9353 );
and \U$22135 ( \31229 , RIe1850e8_2891, \9355 );
and \U$22136 ( \31230 , RIfc8e310_6640, \9357 );
and \U$22137 ( \31231 , RIe1823e8_2859, \9359 );
and \U$22138 ( \31232 , RIe17f6e8_2827, \9361 );
and \U$22139 ( \31233 , RIe17c9e8_2795, \9363 );
and \U$22140 ( \31234 , RIfcd1570_7404, \9365 );
and \U$22141 ( \31235 , RIfccc278_7345, \9367 );
and \U$22142 ( \31236 , RIf1404c8_5191, \9369 );
and \U$22143 ( \31237 , RIfea2d98_8197, \9371 );
and \U$22144 ( \31238 , RIfcc1b20_7226, \9373 );
and \U$22145 ( \31239 , RIfc60398_6117, \9375 );
and \U$22146 ( \31240 , RIee3e5a8_5168, \9377 );
and \U$22147 ( \31241 , RIee3da68_5160, \9379 );
and \U$22148 ( \31242 , RIfc642e0_6162, \9381 );
and \U$22149 ( \31243 , RIfca7f18_6933, \9383 );
and \U$22150 ( \31244 , RIee3a228_5120, \9385 );
and \U$22151 ( \31245 , RIfec6180_8374, \9387 );
and \U$22152 ( \31246 , RIfca9598_6949, \9389 );
and \U$22153 ( \31247 , RIfc5c720_6074, \9391 );
and \U$22154 ( \31248 , RIfc6bea0_6250, \9393 );
and \U$22155 ( \31249 , RIfccaec8_7331, \9395 );
and \U$22156 ( \31250 , RIfc44cd8_5805, \9397 );
and \U$22157 ( \31251 , RIe224940_4706, \9399 );
and \U$22158 ( \31252 , RIfcb6180_7094, \9401 );
and \U$22159 ( \31253 , RIe221c40_4674, \9403 );
and \U$22160 ( \31254 , RIfc55ad8_5997, \9405 );
and \U$22161 ( \31255 , RIe21ef40_4642, \9407 );
and \U$22162 ( \31256 , RIe219540_4578, \9409 );
and \U$22163 ( \31257 , RIe216840_4546, \9411 );
and \U$22164 ( \31258 , RIfc4dc48_5907, \9413 );
and \U$22165 ( \31259 , RIe213b40_4514, \9415 );
and \U$22166 ( \31260 , RIfcdcf10_7536, \9417 );
and \U$22167 ( \31261 , RIe210e40_4482, \9419 );
and \U$22168 ( \31262 , RIfcab1b8_6969, \9421 );
and \U$22169 ( \31263 , RIe20e140_4450, \9423 );
and \U$22170 ( \31264 , RIe20b440_4418, \9425 );
and \U$22171 ( \31265 , RIe208740_4386, \9427 );
and \U$22172 ( \31266 , RIfce3720_7610, \9429 );
and \U$22173 ( \31267 , RIfc64178_6161, \9431 );
and \U$22174 ( \31268 , RIe203178_4325, \9433 );
and \U$22175 ( \31269 , RIe201558_4305, \9435 );
and \U$22176 ( \31270 , RIfcd2ec0_7422, \9437 );
and \U$22177 ( \31271 , RIf164828_5603, \9439 );
and \U$22178 ( \31272 , RIfc7f838_6473, \9441 );
and \U$22179 ( \31273 , RIf162398_5577, \9443 );
and \U$22180 ( \31274 , RIfcc9c80_7318, \9445 );
and \U$22181 ( \31275 , RIfca8bc0_6942, \9447 );
and \U$22182 ( \31276 , RIfea2ac8_8195, \9449 );
and \U$22183 ( \31277 , RIfea2c30_8196, \9451 );
and \U$22184 ( \31278 , RIfc59318_6037, \9453 );
and \U$22185 ( \31279 , RIfc4f160_5922, \9455 );
and \U$22186 ( \31280 , RIf15ac10_5492, \9457 );
and \U$22187 ( \31281 , RIfcebf88_7707, \9459 );
or \U$22188 ( \31282 , \31218 , \31219 , \31220 , \31221 , \31222 , \31223 , \31224 , \31225 , \31226 , \31227 , \31228 , \31229 , \31230 , \31231 , \31232 , \31233 , \31234 , \31235 , \31236 , \31237 , \31238 , \31239 , \31240 , \31241 , \31242 , \31243 , \31244 , \31245 , \31246 , \31247 , \31248 , \31249 , \31250 , \31251 , \31252 , \31253 , \31254 , \31255 , \31256 , \31257 , \31258 , \31259 , \31260 , \31261 , \31262 , \31263 , \31264 , \31265 , \31266 , \31267 , \31268 , \31269 , \31270 , \31271 , \31272 , \31273 , \31274 , \31275 , \31276 , \31277 , \31278 , \31279 , \31280 , \31281 );
and \U$22189 ( \31283 , RIfcbb040_7150, \9462 );
and \U$22190 ( \31284 , RIfca1870_6860, \9464 );
and \U$22191 ( \31285 , RIfc93d10_6704, \9466 );
and \U$22192 ( \31286 , RIe1faeb0_4232, \9468 );
and \U$22193 ( \31287 , RIf1565c0_5442, \9470 );
and \U$22194 ( \31288 , RIf155a80_5434, \9472 );
and \U$22195 ( \31289 , RIfc45c50_5816, \9474 );
and \U$22196 ( \31290 , RIe1f6428_4179, \9476 );
and \U$22197 ( \31291 , RIfccdbc8_7363, \9478 );
and \U$22198 ( \31292 , RIfcccae8_7351, \9480 );
and \U$22199 ( \31293 , RIfca6cd0_6920, \9482 );
and \U$22200 ( \31294 , RIfec6018_8373, \9484 );
and \U$22201 ( \31295 , RIfc64010_6160, \9486 );
and \U$22202 ( \31296 , RIfc434f0_5788, \9488 );
and \U$22203 ( \31297 , RIfc4c028_5887, \9490 );
and \U$22204 ( \31298 , RIe1eee08_4095, \9492 );
and \U$22205 ( \31299 , RIe1ec6a8_4067, \9494 );
and \U$22206 ( \31300 , RIe1e99a8_4035, \9496 );
and \U$22207 ( \31301 , RIe1e6ca8_4003, \9498 );
and \U$22208 ( \31302 , RIe1e3fa8_3971, \9500 );
and \U$22209 ( \31303 , RIe1e12a8_3939, \9502 );
and \U$22210 ( \31304 , RIe1de5a8_3907, \9504 );
and \U$22211 ( \31305 , RIe1db8a8_3875, \9506 );
and \U$22212 ( \31306 , RIe1d8ba8_3843, \9508 );
and \U$22213 ( \31307 , RIe1d31a8_3779, \9510 );
and \U$22214 ( \31308 , RIe1d04a8_3747, \9512 );
and \U$22215 ( \31309 , RIe1cd7a8_3715, \9514 );
and \U$22216 ( \31310 , RIe1caaa8_3683, \9516 );
and \U$22217 ( \31311 , RIe1c7da8_3651, \9518 );
and \U$22218 ( \31312 , RIe1c50a8_3619, \9520 );
and \U$22219 ( \31313 , RIe1c23a8_3587, \9522 );
and \U$22220 ( \31314 , RIe1bf6a8_3555, \9524 );
and \U$22221 ( \31315 , RIfc63908_6155, \9526 );
and \U$22222 ( \31316 , RIfc6bd38_6249, \9528 );
and \U$22223 ( \31317 , RIe1ba0e0_3494, \9530 );
and \U$22224 ( \31318 , RIe1b7f20_3470, \9532 );
and \U$22225 ( \31319 , RIfc66fe0_6194, \9534 );
and \U$22226 ( \31320 , RIfc92ac8_6691, \9536 );
and \U$22227 ( \31321 , RIe1b5d60_3446, \9538 );
and \U$22228 ( \31322 , RIfea2f00_8198, \9540 );
and \U$22229 ( \31323 , RIfc9bfd8_6797, \9542 );
and \U$22230 ( \31324 , RIfc50d80_5942, \9544 );
and \U$22231 ( \31325 , RIe1b31c8_3415, \9546 );
and \U$22232 ( \31326 , RIe1b1878_3397, \9548 );
and \U$22233 ( \31327 , RIfc4df18_5909, \9550 );
and \U$22234 ( \31328 , RIfc9d658_6813, \9552 );
and \U$22235 ( \31329 , RIe1ad0c0_3346, \9554 );
and \U$22236 ( \31330 , RIe1ab8d8_3329, \9556 );
and \U$22237 ( \31331 , RIe1a99e8_3307, \9558 );
and \U$22238 ( \31332 , RIe1a6ce8_3275, \9560 );
and \U$22239 ( \31333 , RIe1a3fe8_3243, \9562 );
and \U$22240 ( \31334 , RIe1a12e8_3211, \9564 );
and \U$22241 ( \31335 , RIe18d7e8_2987, \9566 );
and \U$22242 ( \31336 , RIe179ce8_2763, \9568 );
and \U$22243 ( \31337 , RIe227640_4738, \9570 );
and \U$22244 ( \31338 , RIe21c240_4610, \9572 );
and \U$22245 ( \31339 , RIe205a40_4354, \9574 );
and \U$22246 ( \31340 , RIe1ffaa0_4286, \9576 );
and \U$22247 ( \31341 , RIe1f8e58_4209, \9578 );
and \U$22248 ( \31342 , RIe1f19a0_4126, \9580 );
and \U$22249 ( \31343 , RIe1d5ea8_3811, \9582 );
and \U$22250 ( \31344 , RIe1bc9a8_3523, \9584 );
and \U$22251 ( \31345 , RIe1af820_3374, \9586 );
and \U$22252 ( \31346 , RIe171e58_2673, \9588 );
or \U$22253 ( \31347 , \31283 , \31284 , \31285 , \31286 , \31287 , \31288 , \31289 , \31290 , \31291 , \31292 , \31293 , \31294 , \31295 , \31296 , \31297 , \31298 , \31299 , \31300 , \31301 , \31302 , \31303 , \31304 , \31305 , \31306 , \31307 , \31308 , \31309 , \31310 , \31311 , \31312 , \31313 , \31314 , \31315 , \31316 , \31317 , \31318 , \31319 , \31320 , \31321 , \31322 , \31323 , \31324 , \31325 , \31326 , \31327 , \31328 , \31329 , \31330 , \31331 , \31332 , \31333 , \31334 , \31335 , \31336 , \31337 , \31338 , \31339 , \31340 , \31341 , \31342 , \31343 , \31344 , \31345 , \31346 );
or \U$22254 ( \31348 , \31282 , \31347 );
_DC g3362 ( \31349_nG3362 , \31348 , \9597 );
buf \U$22255 ( \31350 , \31349_nG3362 );
xor \U$22256 ( \31351 , \31217 , \31350 );
and \U$22257 ( \31352 , RIdec61e8_718, \9059 );
and \U$22258 ( \31353 , RIdec34e8_686, \9061 );
and \U$22259 ( \31354 , RIee20620_4827, \9063 );
and \U$22260 ( \31355 , RIdec07e8_654, \9065 );
and \U$22261 ( \31356 , RIfc4b7b8_5881, \9067 );
and \U$22262 ( \31357 , RIdebdae8_622, \9069 );
and \U$22263 ( \31358 , RIdebade8_590, \9071 );
and \U$22264 ( \31359 , RIdeb80e8_558, \9073 );
and \U$22265 ( \31360 , RIfc41150_5766, \9075 );
and \U$22266 ( \31361 , RIdeb26e8_494, \9077 );
and \U$22267 ( \31362 , RIfc87830_6564, \9079 );
and \U$22268 ( \31363 , RIdeaf9e8_462, \9081 );
and \U$22269 ( \31364 , RIee1dec0_4799, \9083 );
and \U$22270 ( \31365 , RIdeac4f0_430, \9085 );
and \U$22271 ( \31366 , RIdea5bf0_398, \9087 );
and \U$22272 ( \31367 , RIde9f2f0_366, \9089 );
and \U$22273 ( \31368 , RIee1d380_4791, \9091 );
and \U$22274 ( \31369 , RIfc77c78_6385, \9093 );
and \U$22275 ( \31370 , RIfc84f68_6535, \9095 );
and \U$22276 ( \31371 , RIfc6ff50_6296, \9097 );
and \U$22277 ( \31372 , RIde92780_304, \9099 );
and \U$22278 ( \31373 , RIde8efb8_287, \9101 );
and \U$22279 ( \31374 , RIde8ae18_267, \9103 );
and \U$22280 ( \31375 , RIde86c78_247, \9105 );
and \U$22281 ( \31376 , RIee1a680_4759, \9107 );
and \U$22282 ( \31377 , RIee19f78_4754, \9109 );
and \U$22283 ( \31378 , RIfcd7240_7470, \9111 );
and \U$22284 ( \31379 , RIfcbeb50_7192, \9113 );
and \U$22285 ( \31380 , RIfc76328_6367, \9115 );
and \U$22286 ( \31381 , RIe16c2f0_2608, \9117 );
and \U$22287 ( \31382 , RIee388d8_5102, \9119 );
and \U$22288 ( \31383 , RIfea20f0_8188, \9121 );
and \U$22289 ( \31384 , RIe1661e8_2539, \9123 );
and \U$22290 ( \31385 , RIe1634e8_2507, \9125 );
and \U$22291 ( \31386 , RIee37c30_5093, \9127 );
and \U$22292 ( \31387 , RIe1607e8_2475, \9129 );
and \U$22293 ( \31388 , RIfce7500_7654, \9131 );
and \U$22294 ( \31389 , RIe15dae8_2443, \9133 );
and \U$22295 ( \31390 , RIe1580e8_2379, \9135 );
and \U$22296 ( \31391 , RIe1553e8_2347, \9137 );
and \U$22297 ( \31392 , RIfc3f698_5747, \9139 );
and \U$22298 ( \31393 , RIe1526e8_2315, \9141 );
and \U$22299 ( \31394 , RIee354d0_5065, \9143 );
and \U$22300 ( \31395 , RIe14f9e8_2283, \9145 );
and \U$22301 ( \31396 , RIfc83e88_6523, \9147 );
and \U$22302 ( \31397 , RIe14cce8_2251, \9149 );
and \U$22303 ( \31398 , RIe149fe8_2219, \9151 );
and \U$22304 ( \31399 , RIe1472e8_2187, \9153 );
and \U$22305 ( \31400 , RIfcea4d0_7688, \9155 );
and \U$22306 ( \31401 , RIfcb7ad0_7112, \9157 );
and \U$22307 ( \31402 , RIfc695d8_6221, \9159 );
and \U$22308 ( \31403 , RIfc51a28_5951, \9161 );
and \U$22309 ( \31404 , RIe141a50_2124, \9163 );
and \U$22310 ( \31405 , RIe13f728_2099, \9165 );
and \U$22311 ( \31406 , RIdf3d630_2075, \9167 );
and \U$22312 ( \31407 , RIdf3b1a0_2049, \9169 );
and \U$22313 ( \31408 , RIfca9e08_6955, \9171 );
and \U$22314 ( \31409 , RIee2fda0_5003, \9173 );
and \U$22315 ( \31410 , RIfc88a78_6577, \9175 );
and \U$22316 ( \31411 , RIee2da78_4978, \9177 );
and \U$22317 ( \31412 , RIdf36448_1994, \9179 );
and \U$22318 ( \31413 , RIdf33fb8_1968, \9181 );
and \U$22319 ( \31414 , RIdf31df8_1944, \9183 );
and \U$22320 ( \31415 , RIfea2258_8189, \9185 );
or \U$22321 ( \31416 , \31352 , \31353 , \31354 , \31355 , \31356 , \31357 , \31358 , \31359 , \31360 , \31361 , \31362 , \31363 , \31364 , \31365 , \31366 , \31367 , \31368 , \31369 , \31370 , \31371 , \31372 , \31373 , \31374 , \31375 , \31376 , \31377 , \31378 , \31379 , \31380 , \31381 , \31382 , \31383 , \31384 , \31385 , \31386 , \31387 , \31388 , \31389 , \31390 , \31391 , \31392 , \31393 , \31394 , \31395 , \31396 , \31397 , \31398 , \31399 , \31400 , \31401 , \31402 , \31403 , \31404 , \31405 , \31406 , \31407 , \31408 , \31409 , \31410 , \31411 , \31412 , \31413 , \31414 , \31415 );
and \U$22322 ( \31417 , RIee2c560_4963, \9188 );
and \U$22323 ( \31418 , RIee2aaa8_4944, \9190 );
and \U$22324 ( \31419 , RIee29428_4928, \9192 );
and \U$22325 ( \31420 , RIee281e0_4915, \9194 );
and \U$22326 ( \31421 , RIdf2ac10_1863, \9196 );
and \U$22327 ( \31422 , RIdf28d20_1841, \9198 );
and \U$22328 ( \31423 , RIfea27f8_8193, \9200 );
and \U$22329 ( \31424 , RIfea2960_8194, \9202 );
and \U$22330 ( \31425 , RIfcdabe8_7511, \9204 );
and \U$22331 ( \31426 , RIfca08f8_6849, \9206 );
and \U$22332 ( \31427 , RIfc8b1d8_6605, \9208 );
and \U$22333 ( \31428 , RIfc49058_5853, \9210 );
and \U$22334 ( \31429 , RIfca0a60_6850, \9212 );
and \U$22335 ( \31430 , RIdf204b8_1744, \9214 );
and \U$22336 ( \31431 , RIfc99cb0_6772, \9216 );
and \U$22337 ( \31432 , RIdf19f78_1672, \9218 );
and \U$22338 ( \31433 , RIdf17db8_1648, \9220 );
and \U$22339 ( \31434 , RIdf150b8_1616, \9222 );
and \U$22340 ( \31435 , RIdf123b8_1584, \9224 );
and \U$22341 ( \31436 , RIdf0f6b8_1552, \9226 );
and \U$22342 ( \31437 , RIdf0c9b8_1520, \9228 );
and \U$22343 ( \31438 , RIdf09cb8_1488, \9230 );
and \U$22344 ( \31439 , RIdf06fb8_1456, \9232 );
and \U$22345 ( \31440 , RIdf042b8_1424, \9234 );
and \U$22346 ( \31441 , RIdefe8b8_1360, \9236 );
and \U$22347 ( \31442 , RIdefbbb8_1328, \9238 );
and \U$22348 ( \31443 , RIdef8eb8_1296, \9240 );
and \U$22349 ( \31444 , RIdef61b8_1264, \9242 );
and \U$22350 ( \31445 , RIdef34b8_1232, \9244 );
and \U$22351 ( \31446 , RIdef07b8_1200, \9246 );
and \U$22352 ( \31447 , RIdeedab8_1168, \9248 );
and \U$22353 ( \31448 , RIdeeadb8_1136, \9250 );
and \U$22354 ( \31449 , RIfcd1f48_7411, \9252 );
and \U$22355 ( \31450 , RIfc57f68_6023, \9254 );
and \U$22356 ( \31451 , RIfcbe2e0_7186, \9256 );
and \U$22357 ( \31452 , RIfcd8fc8_7491, \9258 );
and \U$22358 ( \31453 , RIdee5520_1073, \9260 );
and \U$22359 ( \31454 , RIfea2690_8192, \9262 );
and \U$22360 ( \31455 , RIdee1470_1027, \9264 );
and \U$22361 ( \31456 , RIdedf418_1004, \9266 );
and \U$22362 ( \31457 , RIfc57b30_6020, \9268 );
and \U$22363 ( \31458 , RIfcb35e8_7063, \9270 );
and \U$22364 ( \31459 , RIfcbd7a0_7178, \9272 );
and \U$22365 ( \31460 , RIfc91178_6673, \9274 );
and \U$22366 ( \31461 , RIfea2528_8191, \9276 );
and \U$22367 ( \31462 , RIded7df8_920, \9278 );
and \U$22368 ( \31463 , RIfea23c0_8190, \9280 );
and \U$22369 ( \31464 , RIded3910_871, \9282 );
and \U$22370 ( \31465 , RIded15e8_846, \9284 );
and \U$22371 ( \31466 , RIdece8e8_814, \9286 );
and \U$22372 ( \31467 , RIdecbbe8_782, \9288 );
and \U$22373 ( \31468 , RIdec8ee8_750, \9290 );
and \U$22374 ( \31469 , RIdeb53e8_526, \9292 );
and \U$22375 ( \31470 , RIde989f0_334, \9294 );
and \U$22376 ( \31471 , RIe16eff0_2640, \9296 );
and \U$22377 ( \31472 , RIe15ade8_2411, \9298 );
and \U$22378 ( \31473 , RIe1445e8_2155, \9300 );
and \U$22379 ( \31474 , RIdf38fe0_2025, \9302 );
and \U$22380 ( \31475 , RIdf2d640_1893, \9304 );
and \U$22381 ( \31476 , RIdf1dec0_1717, \9306 );
and \U$22382 ( \31477 , RIdf015b8_1392, \9308 );
and \U$22383 ( \31478 , RIdee80b8_1104, \9310 );
and \U$22384 ( \31479 , RIdedce20_977, \9312 );
and \U$22385 ( \31480 , RIde7e938_207, \9314 );
or \U$22386 ( \31481 , \31417 , \31418 , \31419 , \31420 , \31421 , \31422 , \31423 , \31424 , \31425 , \31426 , \31427 , \31428 , \31429 , \31430 , \31431 , \31432 , \31433 , \31434 , \31435 , \31436 , \31437 , \31438 , \31439 , \31440 , \31441 , \31442 , \31443 , \31444 , \31445 , \31446 , \31447 , \31448 , \31449 , \31450 , \31451 , \31452 , \31453 , \31454 , \31455 , \31456 , \31457 , \31458 , \31459 , \31460 , \31461 , \31462 , \31463 , \31464 , \31465 , \31466 , \31467 , \31468 , \31469 , \31470 , \31471 , \31472 , \31473 , \31474 , \31475 , \31476 , \31477 , \31478 , \31479 , \31480 );
or \U$22387 ( \31482 , \31416 , \31481 );
_DC g22ba ( \31483_nG22ba , \31482 , \9323 );
buf \U$22388 ( \31484 , \31483_nG22ba );
and \U$22389 ( \31485 , RIe19e480_3178, \9333 );
and \U$22390 ( \31486 , RIe19b780_3146, \9335 );
and \U$22391 ( \31487 , RIfccc980_7350, \9337 );
and \U$22392 ( \31488 , RIe198a80_3114, \9339 );
and \U$22393 ( \31489 , RIfcc1148_7219, \9341 );
and \U$22394 ( \31490 , RIe195d80_3082, \9343 );
and \U$22395 ( \31491 , RIe193080_3050, \9345 );
and \U$22396 ( \31492 , RIe190380_3018, \9347 );
and \U$22397 ( \31493 , RIe18a980_2954, \9349 );
and \U$22398 ( \31494 , RIe187c80_2922, \9351 );
and \U$22399 ( \31495 , RIfcb2ee0_7058, \9353 );
and \U$22400 ( \31496 , RIe184f80_2890, \9355 );
and \U$22401 ( \31497 , RIfc615e0_6130, \9357 );
and \U$22402 ( \31498 , RIe182280_2858, \9359 );
and \U$22403 ( \31499 , RIe17f580_2826, \9361 );
and \U$22404 ( \31500 , RIe17c880_2794, \9363 );
and \U$22405 ( \31501 , RIfc69038_6217, \9365 );
and \U$22406 ( \31502 , RIfc4c898_5893, \9367 );
and \U$22407 ( \31503 , RIfc6f2a8_6287, \9369 );
and \U$22408 ( \31504 , RIe1764a8_2723, \9371 );
and \U$22409 ( \31505 , RIfcad0a8_6991, \9373 );
and \U$22410 ( \31506 , RIfc6adc0_6238, \9375 );
and \U$22411 ( \31507 , RIfc70388_6299, \9377 );
and \U$22412 ( \31508 , RIfea1b50_8184, \9379 );
and \U$22413 ( \31509 , RIfea1f88_8187, \9381 );
and \U$22414 ( \31510 , RIfc56e88_6011, \9383 );
and \U$22415 ( \31511 , RIfea1cb8_8185, \9385 );
and \U$22416 ( \31512 , RIe174450_2700, \9387 );
and \U$22417 ( \31513 , RIfc60d70_6124, \9389 );
and \U$22418 ( \31514 , RIfc6a820_6234, \9391 );
and \U$22419 ( \31515 , RIfea1e20_8186, \9393 );
and \U$22420 ( \31516 , RIf16d798_5705, \9395 );
and \U$22421 ( \31517 , RIfc40bb0_5762, \9397 );
and \U$22422 ( \31518 , RIe2247d8_4705, \9399 );
and \U$22423 ( \31519 , RIfc77138_6377, \9401 );
and \U$22424 ( \31520 , RIe221ad8_4673, \9403 );
and \U$22425 ( \31521 , RIfcd7d80_7478, \9405 );
and \U$22426 ( \31522 , RIe21edd8_4641, \9407 );
and \U$22427 ( \31523 , RIe2193d8_4577, \9409 );
and \U$22428 ( \31524 , RIe2166d8_4545, \9411 );
and \U$22429 ( \31525 , RIfc40070_5754, \9413 );
and \U$22430 ( \31526 , RIe2139d8_4513, \9415 );
and \U$22431 ( \31527 , RIf169850_5660, \9417 );
and \U$22432 ( \31528 , RIe210cd8_4481, \9419 );
and \U$22433 ( \31529 , RIfcc1580_7222, \9421 );
and \U$22434 ( \31530 , RIe20dfd8_4449, \9423 );
and \U$22435 ( \31531 , RIe20b2d8_4417, \9425 );
and \U$22436 ( \31532 , RIe2085d8_4385, \9427 );
and \U$22437 ( \31533 , RIfcd0058_7389, \9429 );
and \U$22438 ( \31534 , RIfc749d8_6349, \9431 );
and \U$22439 ( \31535 , RIe203010_4324, \9433 );
and \U$22440 ( \31536 , RIe2013f0_4304, \9435 );
and \U$22441 ( \31537 , RIfc60230_6116, \9437 );
and \U$22442 ( \31538 , RIfc60668_6119, \9439 );
and \U$22443 ( \31539 , RIfcaf970_7020, \9441 );
and \U$22444 ( \31540 , RIfc45818_5813, \9443 );
and \U$22445 ( \31541 , RIf160a48_5559, \9445 );
and \U$22446 ( \31542 , RIf15eb58_5537, \9447 );
and \U$22447 ( \31543 , RIfea1880_8182, \9449 );
and \U$22448 ( \31544 , RIfea19e8_8183, \9451 );
and \U$22449 ( \31545 , RIfc72110_6320, \9453 );
and \U$22450 ( \31546 , RIfc49b98_5861, \9455 );
and \U$22451 ( \31547 , RIfcca0b8_7321, \9457 );
and \U$22452 ( \31548 , RIfc71738_6313, \9459 );
or \U$22453 ( \31549 , \31485 , \31486 , \31487 , \31488 , \31489 , \31490 , \31491 , \31492 , \31493 , \31494 , \31495 , \31496 , \31497 , \31498 , \31499 , \31500 , \31501 , \31502 , \31503 , \31504 , \31505 , \31506 , \31507 , \31508 , \31509 , \31510 , \31511 , \31512 , \31513 , \31514 , \31515 , \31516 , \31517 , \31518 , \31519 , \31520 , \31521 , \31522 , \31523 , \31524 , \31525 , \31526 , \31527 , \31528 , \31529 , \31530 , \31531 , \31532 , \31533 , \31534 , \31535 , \31536 , \31537 , \31538 , \31539 , \31540 , \31541 , \31542 , \31543 , \31544 , \31545 , \31546 , \31547 , \31548 );
and \U$22454 ( \31550 , RIfc4ca00_5894, \9462 );
and \U$22455 ( \31551 , RIfc71030_6308, \9464 );
and \U$22456 ( \31552 , RIfcde428_7551, \9466 );
and \U$22457 ( \31553 , RIe1fad48_4231, \9468 );
and \U$22458 ( \31554 , RIfc70bf8_6305, \9470 );
and \U$22459 ( \31555 , RIfc63a70_6156, \9472 );
and \U$22460 ( \31556 , RIfca7db0_6932, \9474 );
and \U$22461 ( \31557 , RIe1f62c0_4178, \9476 );
and \U$22462 ( \31558 , RIfcada80_6998, \9478 );
and \U$22463 ( \31559 , RIfc6fde8_6295, \9480 );
and \U$22464 ( \31560 , RIfc6f578_6289, \9482 );
and \U$22465 ( \31561 , RIe1f3f98_4153, \9484 );
and \U$22466 ( \31562 , RIfcde158_7549, \9486 );
and \U$22467 ( \31563 , RIfcad378_6993, \9488 );
and \U$22468 ( \31564 , RIfc65f00_6182, \9490 );
and \U$22469 ( \31565 , RIe1eeca0_4094, \9492 );
and \U$22470 ( \31566 , RIe1ec540_4066, \9494 );
and \U$22471 ( \31567 , RIe1e9840_4034, \9496 );
and \U$22472 ( \31568 , RIe1e6b40_4002, \9498 );
and \U$22473 ( \31569 , RIe1e3e40_3970, \9500 );
and \U$22474 ( \31570 , RIe1e1140_3938, \9502 );
and \U$22475 ( \31571 , RIe1de440_3906, \9504 );
and \U$22476 ( \31572 , RIe1db740_3874, \9506 );
and \U$22477 ( \31573 , RIe1d8a40_3842, \9508 );
and \U$22478 ( \31574 , RIe1d3040_3778, \9510 );
and \U$22479 ( \31575 , RIe1d0340_3746, \9512 );
and \U$22480 ( \31576 , RIe1cd640_3714, \9514 );
and \U$22481 ( \31577 , RIe1ca940_3682, \9516 );
and \U$22482 ( \31578 , RIe1c7c40_3650, \9518 );
and \U$22483 ( \31579 , RIe1c4f40_3618, \9520 );
and \U$22484 ( \31580 , RIe1c2240_3586, \9522 );
and \U$22485 ( \31581 , RIe1bf540_3554, \9524 );
and \U$22486 ( \31582 , RIfc69308_6219, \9526 );
and \U$22487 ( \31583 , RIfccba08_7339, \9528 );
and \U$22488 ( \31584 , RIe1b9f78_3493, \9530 );
and \U$22489 ( \31585 , RIe1b7db8_3469, \9532 );
and \U$22490 ( \31586 , RIfccd628_7359, \9534 );
and \U$22491 ( \31587 , RIfc69740_6222, \9536 );
and \U$22492 ( \31588 , RIe1b5bf8_3445, \9538 );
and \U$22493 ( \31589 , RIe1b4578_3429, \9540 );
and \U$22494 ( \31590 , RIfccf950_7384, \9542 );
and \U$22495 ( \31591 , RIf148088_5279, \9544 );
and \U$22496 ( \31592 , RIe1b3060_3414, \9546 );
and \U$22497 ( \31593 , RIe1b1710_3396, \9548 );
and \U$22498 ( \31594 , RIfc9f818_6837, \9550 );
and \U$22499 ( \31595 , RIfcb9c90_7136, \9552 );
and \U$22500 ( \31596 , RIe1acf58_3345, \9554 );
and \U$22501 ( \31597 , RIe1ab770_3328, \9556 );
and \U$22502 ( \31598 , RIe1a9880_3306, \9558 );
and \U$22503 ( \31599 , RIe1a6b80_3274, \9560 );
and \U$22504 ( \31600 , RIe1a3e80_3242, \9562 );
and \U$22505 ( \31601 , RIe1a1180_3210, \9564 );
and \U$22506 ( \31602 , RIe18d680_2986, \9566 );
and \U$22507 ( \31603 , RIe179b80_2762, \9568 );
and \U$22508 ( \31604 , RIe2274d8_4737, \9570 );
and \U$22509 ( \31605 , RIe21c0d8_4609, \9572 );
and \U$22510 ( \31606 , RIe2058d8_4353, \9574 );
and \U$22511 ( \31607 , RIe1ff938_4285, \9576 );
and \U$22512 ( \31608 , RIe1f8cf0_4208, \9578 );
and \U$22513 ( \31609 , RIe1f1838_4125, \9580 );
and \U$22514 ( \31610 , RIe1d5d40_3810, \9582 );
and \U$22515 ( \31611 , RIe1bc840_3522, \9584 );
and \U$22516 ( \31612 , RIe1af6b8_3373, \9586 );
and \U$22517 ( \31613 , RIe171cf0_2672, \9588 );
or \U$22518 ( \31614 , \31550 , \31551 , \31552 , \31553 , \31554 , \31555 , \31556 , \31557 , \31558 , \31559 , \31560 , \31561 , \31562 , \31563 , \31564 , \31565 , \31566 , \31567 , \31568 , \31569 , \31570 , \31571 , \31572 , \31573 , \31574 , \31575 , \31576 , \31577 , \31578 , \31579 , \31580 , \31581 , \31582 , \31583 , \31584 , \31585 , \31586 , \31587 , \31588 , \31589 , \31590 , \31591 , \31592 , \31593 , \31594 , \31595 , \31596 , \31597 , \31598 , \31599 , \31600 , \31601 , \31602 , \31603 , \31604 , \31605 , \31606 , \31607 , \31608 , \31609 , \31610 , \31611 , \31612 , \31613 );
or \U$22519 ( \31615 , \31549 , \31614 );
_DC g33e7 ( \31616_nG33e7 , \31615 , \9597 );
buf \U$22520 ( \31617 , \31616_nG33e7 );
and \U$22521 ( \31618 , \31484 , \31617 );
and \U$22522 ( \31619 , \29434 , \29567 );
and \U$22523 ( \31620 , \29567 , \29842 );
and \U$22524 ( \31621 , \29434 , \29842 );
or \U$22525 ( \31622 , \31619 , \31620 , \31621 );
and \U$22526 ( \31623 , \31617 , \31622 );
and \U$22527 ( \31624 , \31484 , \31622 );
or \U$22528 ( \31625 , \31618 , \31623 , \31624 );
xor \U$22529 ( \31626 , \31351 , \31625 );
buf g43fa ( \31627_nG43fa , \31626 );
xor \U$22530 ( \31628 , \31484 , \31617 );
xor \U$22531 ( \31629 , \31628 , \31622 );
buf g43fd ( \31630_nG43fd , \31629 );
nand \U$22532 ( \31631 , \31630_nG43fd , \29844_nG4400 );
and \U$22533 ( \31632 , \31627_nG43fa , \31631 );
xor \U$22534 ( \31633 , \31630_nG43fd , \29844_nG4400 );
not \U$22535 ( \31634 , \31633 );
xor \U$22536 ( \31635 , \31627_nG43fa , \31630_nG43fd );
and \U$22537 ( \31636 , \31634 , \31635 );
and \U$22539 ( \31637 , \31633 , \10694_nG9c0e );
or \U$22540 ( \31638 , 1'b0 , \31637 );
xor \U$22541 ( \31639 , \31632 , \31638 );
xor \U$22542 ( \31640 , \31632 , \31639 );
buf \U$22543 ( \31641 , \31640 );
buf \U$22544 ( \31642 , \31641 );
xor \U$22545 ( \31643 , \31084 , \31642 );
and \U$22546 ( \31644 , \31025 , \31030 );
and \U$22547 ( \31645 , \31025 , \31077 );
and \U$22548 ( \31646 , \31030 , \31077 );
or \U$22549 ( \31647 , \31644 , \31645 , \31646 );
and \U$22550 ( \31648 , \31643 , \31647 );
and \U$22551 ( \31649 , \31064 , \31069 );
and \U$22552 ( \31650 , \31064 , \31075 );
and \U$22553 ( \31651 , \31069 , \31075 );
or \U$22554 ( \31652 , \31649 , \31650 , \31651 );
buf \U$22555 ( \31653 , \31652 );
and \U$22556 ( \31654 , \30947 , \30952 );
and \U$22557 ( \31655 , \30947 , \31023 );
and \U$22558 ( \31656 , \30952 , \31023 );
or \U$22559 ( \31657 , \31654 , \31655 , \31656 );
buf \U$22560 ( \31658 , \31657 );
and \U$22561 ( \31659 , \31008 , \31014 );
and \U$22562 ( \31660 , \31008 , \31021 );
and \U$22563 ( \31661 , \31014 , \31021 );
or \U$22564 ( \31662 , \31659 , \31660 , \31661 );
buf \U$22565 ( \31663 , \31662 );
and \U$22566 ( \31664 , \30993 , \30999 );
and \U$22567 ( \31665 , \30993 , \31006 );
and \U$22568 ( \31666 , \30999 , \31006 );
or \U$22569 ( \31667 , \31664 , \31665 , \31666 );
buf \U$22570 ( \31668 , \31667 );
and \U$22571 ( \31669 , \20155 , \18107_nG9be7 );
and \U$22572 ( \31670 , \20152 , \19091_nG9be4 );
or \U$22573 ( \31671 , \31669 , \31670 );
xor \U$22574 ( \31672 , \20151 , \31671 );
buf \U$22575 ( \31673 , \31672 );
buf \U$22577 ( \31674 , \31673 );
and \U$22578 ( \31675 , \18702 , \19586_nG9be1 );
and \U$22579 ( \31676 , \18699 , \20608_nG9bde );
or \U$22580 ( \31677 , \31675 , \31676 );
xor \U$22581 ( \31678 , \18698 , \31677 );
buf \U$22582 ( \31679 , \31678 );
buf \U$22584 ( \31680 , \31679 );
xor \U$22585 ( \31681 , \31674 , \31680 );
and \U$22586 ( \31682 , \17297 , \21086_nG9bdb );
and \U$22587 ( \31683 , \17294 , \22129_nG9bd8 );
or \U$22588 ( \31684 , \31682 , \31683 );
xor \U$22589 ( \31685 , \17293 , \31684 );
buf \U$22590 ( \31686 , \31685 );
buf \U$22592 ( \31687 , \31686 );
xor \U$22593 ( \31688 , \31681 , \31687 );
buf \U$22594 ( \31689 , \31688 );
xor \U$22595 ( \31690 , \31668 , \31689 );
and \U$22596 ( \31691 , \12157 , \27416_nG9bc3 );
and \U$22597 ( \31692 , \12154 , \28602_nG9bc0 );
or \U$22598 ( \31693 , \31691 , \31692 );
xor \U$22599 ( \31694 , \12153 , \31693 );
buf \U$22600 ( \31695 , \31694 );
buf \U$22602 ( \31696 , \31695 );
xor \U$22603 ( \31697 , \31690 , \31696 );
buf \U$22604 ( \31698 , \31697 );
xor \U$22605 ( \31699 , \31663 , \31698 );
and \U$22606 ( \31700 , \31036 , \31042 );
and \U$22607 ( \31701 , \31036 , \31049 );
and \U$22608 ( \31702 , \31042 , \31049 );
or \U$22609 ( \31703 , \31700 , \31701 , \31702 );
buf \U$22610 ( \31704 , \31703 );
xor \U$22611 ( \31705 , \31699 , \31704 );
buf \U$22612 ( \31706 , \31705 );
xor \U$22613 ( \31707 , \31658 , \31706 );
and \U$22614 ( \31708 , \30496 , \30501 );
and \U$22615 ( \31709 , \30496 , \30508 );
and \U$22616 ( \31710 , \30501 , \30508 );
or \U$22617 ( \31711 , \31708 , \31709 , \31710 );
buf \U$22618 ( \31712 , \31711 );
and \U$22619 ( \31713 , \30472 , \30478 );
and \U$22620 ( \31714 , \30472 , \30485 );
and \U$22621 ( \31715 , \30478 , \30485 );
or \U$22622 ( \31716 , \31713 , \31714 , \31715 );
buf \U$22623 ( \31717 , \31716 );
and \U$22624 ( \31718 , \30961 , \30967 );
buf \U$22625 ( \31719 , \31718 );
and \U$22626 ( \31720 , \26431 , \12801_nG9bff );
and \U$22627 ( \31721 , \26428 , \13705_nG9bfc );
or \U$22628 ( \31722 , \31720 , \31721 );
xor \U$22629 ( \31723 , \26427 , \31722 );
buf \U$22630 ( \31724 , \31723 );
buf \U$22632 ( \31725 , \31724 );
xor \U$22633 ( \31726 , \31719 , \31725 );
and \U$22634 ( \31727 , \24792 , \14070_nG9bf9 );
and \U$22635 ( \31728 , \24789 , \14984_nG9bf6 );
or \U$22636 ( \31729 , \31727 , \31728 );
xor \U$22637 ( \31730 , \24788 , \31729 );
buf \U$22638 ( \31731 , \31730 );
buf \U$22640 ( \31732 , \31731 );
xor \U$22641 ( \31733 , \31726 , \31732 );
buf \U$22642 ( \31734 , \31733 );
xor \U$22643 ( \31735 , \31717 , \31734 );
and \U$22644 ( \31736 , \21658 , \16680_nG9bed );
and \U$22645 ( \31737 , \21655 , \17665_nG9bea );
or \U$22646 ( \31738 , \31736 , \31737 );
xor \U$22647 ( \31739 , \21654 , \31738 );
buf \U$22648 ( \31740 , \31739 );
buf \U$22650 ( \31741 , \31740 );
xor \U$22651 ( \31742 , \31735 , \31741 );
buf \U$22652 ( \31743 , \31742 );
and \U$22653 ( \31744 , \15940 , \22629_nG9bd5 );
and \U$22654 ( \31745 , \15937 , \23696_nG9bd2 );
or \U$22655 ( \31746 , \31744 , \31745 );
xor \U$22656 ( \31747 , \15936 , \31746 );
buf \U$22657 ( \31748 , \31747 );
buf \U$22659 ( \31749 , \31748 );
xor \U$22660 ( \31750 , \31743 , \31749 );
and \U$22661 ( \31751 , \14631 , \24226_nG9bcf );
and \U$22662 ( \31752 , \14628 , \25298_nG9bcc );
or \U$22663 ( \31753 , \31751 , \31752 );
xor \U$22664 ( \31754 , \14627 , \31753 );
buf \U$22665 ( \31755 , \31754 );
buf \U$22667 ( \31756 , \31755 );
xor \U$22668 ( \31757 , \31750 , \31756 );
buf \U$22669 ( \31758 , \31757 );
xor \U$22670 ( \31759 , \31712 , \31758 );
and \U$22671 ( \31760 , \10707 , \30940_nG9bb7 );
and \U$22672 ( \31761 , \30829 , \30873 );
and \U$22673 ( \31762 , \30873 , \30928 );
and \U$22674 ( \31763 , \30829 , \30928 );
or \U$22675 ( \31764 , \31761 , \31762 , \31763 );
and \U$22676 ( \31765 , \30530 , \30534 );
and \U$22677 ( \31766 , \30534 , \30828 );
and \U$22678 ( \31767 , \30530 , \30828 );
or \U$22679 ( \31768 , \31765 , \31766 , \31767 );
and \U$22680 ( \31769 , \30833 , \30847 );
and \U$22681 ( \31770 , \30847 , \30872 );
and \U$22682 ( \31771 , \30833 , \30872 );
or \U$22683 ( \31772 , \31769 , \31770 , \31771 );
xor \U$22684 ( \31773 , \31768 , \31772 );
and \U$22685 ( \31774 , \21033 , \18090 );
and \U$22686 ( \31775 , \22090 , \17655 );
nor \U$22687 ( \31776 , \31774 , \31775 );
xnor \U$22688 ( \31777 , \31776 , \18046 );
and \U$22689 ( \31778 , \12769 , \27397 );
and \U$22690 ( \31779 , \13679 , \26807 );
nor \U$22691 ( \31780 , \31778 , \31779 );
xnor \U$22692 ( \31781 , \31780 , \27295 );
xor \U$22693 ( \31782 , \31777 , \31781 );
and \U$22694 ( \31783 , \11586 , \29070 );
and \U$22695 ( \31784 , \12448 , \28526 );
nor \U$22696 ( \31785 , \31783 , \31784 );
xnor \U$22697 ( \31786 , \31785 , \29076 );
xor \U$22698 ( \31787 , \31782 , \31786 );
and \U$22699 ( \31788 , \30802 , \10983 );
and \U$22700 ( \31789 , RIdec61e8_718, \9333 );
and \U$22701 ( \31790 , RIdec34e8_686, \9335 );
and \U$22702 ( \31791 , RIee20620_4827, \9337 );
and \U$22703 ( \31792 , RIdec07e8_654, \9339 );
and \U$22704 ( \31793 , RIfc4b7b8_5881, \9341 );
and \U$22705 ( \31794 , RIdebdae8_622, \9343 );
and \U$22706 ( \31795 , RIdebade8_590, \9345 );
and \U$22707 ( \31796 , RIdeb80e8_558, \9347 );
and \U$22708 ( \31797 , RIfc41150_5766, \9349 );
and \U$22709 ( \31798 , RIdeb26e8_494, \9351 );
and \U$22710 ( \31799 , RIfc87830_6564, \9353 );
and \U$22711 ( \31800 , RIdeaf9e8_462, \9355 );
and \U$22712 ( \31801 , RIee1dec0_4799, \9357 );
and \U$22713 ( \31802 , RIdeac4f0_430, \9359 );
and \U$22714 ( \31803 , RIdea5bf0_398, \9361 );
and \U$22715 ( \31804 , RIde9f2f0_366, \9363 );
and \U$22716 ( \31805 , RIee1d380_4791, \9365 );
and \U$22717 ( \31806 , RIfc77c78_6385, \9367 );
and \U$22718 ( \31807 , RIfc84f68_6535, \9369 );
and \U$22719 ( \31808 , RIfc6ff50_6296, \9371 );
and \U$22720 ( \31809 , RIde92780_304, \9373 );
and \U$22721 ( \31810 , RIde8efb8_287, \9375 );
and \U$22722 ( \31811 , RIde8ae18_267, \9377 );
and \U$22723 ( \31812 , RIde86c78_247, \9379 );
and \U$22724 ( \31813 , RIee1a680_4759, \9381 );
and \U$22725 ( \31814 , RIee19f78_4754, \9383 );
and \U$22726 ( \31815 , RIfcd7240_7470, \9385 );
and \U$22727 ( \31816 , RIfcbeb50_7192, \9387 );
and \U$22728 ( \31817 , RIfc76328_6367, \9389 );
and \U$22729 ( \31818 , RIe16c2f0_2608, \9391 );
and \U$22730 ( \31819 , RIee388d8_5102, \9393 );
and \U$22731 ( \31820 , RIfea20f0_8188, \9395 );
and \U$22732 ( \31821 , RIe1661e8_2539, \9397 );
and \U$22733 ( \31822 , RIe1634e8_2507, \9399 );
and \U$22734 ( \31823 , RIee37c30_5093, \9401 );
and \U$22735 ( \31824 , RIe1607e8_2475, \9403 );
and \U$22736 ( \31825 , RIfce7500_7654, \9405 );
and \U$22737 ( \31826 , RIe15dae8_2443, \9407 );
and \U$22738 ( \31827 , RIe1580e8_2379, \9409 );
and \U$22739 ( \31828 , RIe1553e8_2347, \9411 );
and \U$22740 ( \31829 , RIfc3f698_5747, \9413 );
and \U$22741 ( \31830 , RIe1526e8_2315, \9415 );
and \U$22742 ( \31831 , RIee354d0_5065, \9417 );
and \U$22743 ( \31832 , RIe14f9e8_2283, \9419 );
and \U$22744 ( \31833 , RIfc83e88_6523, \9421 );
and \U$22745 ( \31834 , RIe14cce8_2251, \9423 );
and \U$22746 ( \31835 , RIe149fe8_2219, \9425 );
and \U$22747 ( \31836 , RIe1472e8_2187, \9427 );
and \U$22748 ( \31837 , RIfcea4d0_7688, \9429 );
and \U$22749 ( \31838 , RIfcb7ad0_7112, \9431 );
and \U$22750 ( \31839 , RIfc695d8_6221, \9433 );
and \U$22751 ( \31840 , RIfc51a28_5951, \9435 );
and \U$22752 ( \31841 , RIe141a50_2124, \9437 );
and \U$22753 ( \31842 , RIe13f728_2099, \9439 );
and \U$22754 ( \31843 , RIdf3d630_2075, \9441 );
and \U$22755 ( \31844 , RIdf3b1a0_2049, \9443 );
and \U$22756 ( \31845 , RIfca9e08_6955, \9445 );
and \U$22757 ( \31846 , RIee2fda0_5003, \9447 );
and \U$22758 ( \31847 , RIfc88a78_6577, \9449 );
and \U$22759 ( \31848 , RIee2da78_4978, \9451 );
and \U$22760 ( \31849 , RIdf36448_1994, \9453 );
and \U$22761 ( \31850 , RIdf33fb8_1968, \9455 );
and \U$22762 ( \31851 , RIdf31df8_1944, \9457 );
and \U$22763 ( \31852 , RIfea2258_8189, \9459 );
or \U$22764 ( \31853 , \31789 , \31790 , \31791 , \31792 , \31793 , \31794 , \31795 , \31796 , \31797 , \31798 , \31799 , \31800 , \31801 , \31802 , \31803 , \31804 , \31805 , \31806 , \31807 , \31808 , \31809 , \31810 , \31811 , \31812 , \31813 , \31814 , \31815 , \31816 , \31817 , \31818 , \31819 , \31820 , \31821 , \31822 , \31823 , \31824 , \31825 , \31826 , \31827 , \31828 , \31829 , \31830 , \31831 , \31832 , \31833 , \31834 , \31835 , \31836 , \31837 , \31838 , \31839 , \31840 , \31841 , \31842 , \31843 , \31844 , \31845 , \31846 , \31847 , \31848 , \31849 , \31850 , \31851 , \31852 );
and \U$22765 ( \31854 , RIee2c560_4963, \9462 );
and \U$22766 ( \31855 , RIee2aaa8_4944, \9464 );
and \U$22767 ( \31856 , RIee29428_4928, \9466 );
and \U$22768 ( \31857 , RIee281e0_4915, \9468 );
and \U$22769 ( \31858 , RIdf2ac10_1863, \9470 );
and \U$22770 ( \31859 , RIdf28d20_1841, \9472 );
and \U$22771 ( \31860 , RIfea27f8_8193, \9474 );
and \U$22772 ( \31861 , RIfea2960_8194, \9476 );
and \U$22773 ( \31862 , RIfcdabe8_7511, \9478 );
and \U$22774 ( \31863 , RIfca08f8_6849, \9480 );
and \U$22775 ( \31864 , RIfc8b1d8_6605, \9482 );
and \U$22776 ( \31865 , RIfc49058_5853, \9484 );
and \U$22777 ( \31866 , RIfca0a60_6850, \9486 );
and \U$22778 ( \31867 , RIdf204b8_1744, \9488 );
and \U$22779 ( \31868 , RIfc99cb0_6772, \9490 );
and \U$22780 ( \31869 , RIdf19f78_1672, \9492 );
and \U$22781 ( \31870 , RIdf17db8_1648, \9494 );
and \U$22782 ( \31871 , RIdf150b8_1616, \9496 );
and \U$22783 ( \31872 , RIdf123b8_1584, \9498 );
and \U$22784 ( \31873 , RIdf0f6b8_1552, \9500 );
and \U$22785 ( \31874 , RIdf0c9b8_1520, \9502 );
and \U$22786 ( \31875 , RIdf09cb8_1488, \9504 );
and \U$22787 ( \31876 , RIdf06fb8_1456, \9506 );
and \U$22788 ( \31877 , RIdf042b8_1424, \9508 );
and \U$22789 ( \31878 , RIdefe8b8_1360, \9510 );
and \U$22790 ( \31879 , RIdefbbb8_1328, \9512 );
and \U$22791 ( \31880 , RIdef8eb8_1296, \9514 );
and \U$22792 ( \31881 , RIdef61b8_1264, \9516 );
and \U$22793 ( \31882 , RIdef34b8_1232, \9518 );
and \U$22794 ( \31883 , RIdef07b8_1200, \9520 );
and \U$22795 ( \31884 , RIdeedab8_1168, \9522 );
and \U$22796 ( \31885 , RIdeeadb8_1136, \9524 );
and \U$22797 ( \31886 , RIfcd1f48_7411, \9526 );
and \U$22798 ( \31887 , RIfc57f68_6023, \9528 );
and \U$22799 ( \31888 , RIfcbe2e0_7186, \9530 );
and \U$22800 ( \31889 , RIfcd8fc8_7491, \9532 );
and \U$22801 ( \31890 , RIdee5520_1073, \9534 );
and \U$22802 ( \31891 , RIfea2690_8192, \9536 );
and \U$22803 ( \31892 , RIdee1470_1027, \9538 );
and \U$22804 ( \31893 , RIdedf418_1004, \9540 );
and \U$22805 ( \31894 , RIfc57b30_6020, \9542 );
and \U$22806 ( \31895 , RIfcb35e8_7063, \9544 );
and \U$22807 ( \31896 , RIfcbd7a0_7178, \9546 );
and \U$22808 ( \31897 , RIfc91178_6673, \9548 );
and \U$22809 ( \31898 , RIfea2528_8191, \9550 );
and \U$22810 ( \31899 , RIded7df8_920, \9552 );
and \U$22811 ( \31900 , RIfea23c0_8190, \9554 );
and \U$22812 ( \31901 , RIded3910_871, \9556 );
and \U$22813 ( \31902 , RIded15e8_846, \9558 );
and \U$22814 ( \31903 , RIdece8e8_814, \9560 );
and \U$22815 ( \31904 , RIdecbbe8_782, \9562 );
and \U$22816 ( \31905 , RIdec8ee8_750, \9564 );
and \U$22817 ( \31906 , RIdeb53e8_526, \9566 );
and \U$22818 ( \31907 , RIde989f0_334, \9568 );
and \U$22819 ( \31908 , RIe16eff0_2640, \9570 );
and \U$22820 ( \31909 , RIe15ade8_2411, \9572 );
and \U$22821 ( \31910 , RIe1445e8_2155, \9574 );
and \U$22822 ( \31911 , RIdf38fe0_2025, \9576 );
and \U$22823 ( \31912 , RIdf2d640_1893, \9578 );
and \U$22824 ( \31913 , RIdf1dec0_1717, \9580 );
and \U$22825 ( \31914 , RIdf015b8_1392, \9582 );
and \U$22826 ( \31915 , RIdee80b8_1104, \9584 );
and \U$22827 ( \31916 , RIdedce20_977, \9586 );
and \U$22828 ( \31917 , RIde7e938_207, \9588 );
or \U$22829 ( \31918 , \31854 , \31855 , \31856 , \31857 , \31858 , \31859 , \31860 , \31861 , \31862 , \31863 , \31864 , \31865 , \31866 , \31867 , \31868 , \31869 , \31870 , \31871 , \31872 , \31873 , \31874 , \31875 , \31876 , \31877 , \31878 , \31879 , \31880 , \31881 , \31882 , \31883 , \31884 , \31885 , \31886 , \31887 , \31888 , \31889 , \31890 , \31891 , \31892 , \31893 , \31894 , \31895 , \31896 , \31897 , \31898 , \31899 , \31900 , \31901 , \31902 , \31903 , \31904 , \31905 , \31906 , \31907 , \31908 , \31909 , \31910 , \31911 , \31912 , \31913 , \31914 , \31915 , \31916 , \31917 );
or \U$22830 ( \31919 , \31853 , \31918 );
_DC g65d1 ( \31920_nG65d1 , \31919 , \9597 );
and \U$22831 ( \31921 , RIe19e480_3178, \9059 );
and \U$22832 ( \31922 , RIe19b780_3146, \9061 );
and \U$22833 ( \31923 , RIfccc980_7350, \9063 );
and \U$22834 ( \31924 , RIe198a80_3114, \9065 );
and \U$22835 ( \31925 , RIfcc1148_7219, \9067 );
and \U$22836 ( \31926 , RIe195d80_3082, \9069 );
and \U$22837 ( \31927 , RIe193080_3050, \9071 );
and \U$22838 ( \31928 , RIe190380_3018, \9073 );
and \U$22839 ( \31929 , RIe18a980_2954, \9075 );
and \U$22840 ( \31930 , RIe187c80_2922, \9077 );
and \U$22841 ( \31931 , RIfcb2ee0_7058, \9079 );
and \U$22842 ( \31932 , RIe184f80_2890, \9081 );
and \U$22843 ( \31933 , RIfc615e0_6130, \9083 );
and \U$22844 ( \31934 , RIe182280_2858, \9085 );
and \U$22845 ( \31935 , RIe17f580_2826, \9087 );
and \U$22846 ( \31936 , RIe17c880_2794, \9089 );
and \U$22847 ( \31937 , RIfc69038_6217, \9091 );
and \U$22848 ( \31938 , RIfc4c898_5893, \9093 );
and \U$22849 ( \31939 , RIfc6f2a8_6287, \9095 );
and \U$22850 ( \31940 , RIe1764a8_2723, \9097 );
and \U$22851 ( \31941 , RIfcad0a8_6991, \9099 );
and \U$22852 ( \31942 , RIfc6adc0_6238, \9101 );
and \U$22853 ( \31943 , RIfc70388_6299, \9103 );
and \U$22854 ( \31944 , RIfea1b50_8184, \9105 );
and \U$22855 ( \31945 , RIfea1f88_8187, \9107 );
and \U$22856 ( \31946 , RIfc56e88_6011, \9109 );
and \U$22857 ( \31947 , RIfea1cb8_8185, \9111 );
and \U$22858 ( \31948 , RIe174450_2700, \9113 );
and \U$22859 ( \31949 , RIfc60d70_6124, \9115 );
and \U$22860 ( \31950 , RIfc6a820_6234, \9117 );
and \U$22861 ( \31951 , RIfea1e20_8186, \9119 );
and \U$22862 ( \31952 , RIf16d798_5705, \9121 );
and \U$22863 ( \31953 , RIfc40bb0_5762, \9123 );
and \U$22864 ( \31954 , RIe2247d8_4705, \9125 );
and \U$22865 ( \31955 , RIfc77138_6377, \9127 );
and \U$22866 ( \31956 , RIe221ad8_4673, \9129 );
and \U$22867 ( \31957 , RIfcd7d80_7478, \9131 );
and \U$22868 ( \31958 , RIe21edd8_4641, \9133 );
and \U$22869 ( \31959 , RIe2193d8_4577, \9135 );
and \U$22870 ( \31960 , RIe2166d8_4545, \9137 );
and \U$22871 ( \31961 , RIfc40070_5754, \9139 );
and \U$22872 ( \31962 , RIe2139d8_4513, \9141 );
and \U$22873 ( \31963 , RIf169850_5660, \9143 );
and \U$22874 ( \31964 , RIe210cd8_4481, \9145 );
and \U$22875 ( \31965 , RIfcc1580_7222, \9147 );
and \U$22876 ( \31966 , RIe20dfd8_4449, \9149 );
and \U$22877 ( \31967 , RIe20b2d8_4417, \9151 );
and \U$22878 ( \31968 , RIe2085d8_4385, \9153 );
and \U$22879 ( \31969 , RIfcd0058_7389, \9155 );
and \U$22880 ( \31970 , RIfc749d8_6349, \9157 );
and \U$22881 ( \31971 , RIe203010_4324, \9159 );
and \U$22882 ( \31972 , RIe2013f0_4304, \9161 );
and \U$22883 ( \31973 , RIfc60230_6116, \9163 );
and \U$22884 ( \31974 , RIfc60668_6119, \9165 );
and \U$22885 ( \31975 , RIfcaf970_7020, \9167 );
and \U$22886 ( \31976 , RIfc45818_5813, \9169 );
and \U$22887 ( \31977 , RIf160a48_5559, \9171 );
and \U$22888 ( \31978 , RIf15eb58_5537, \9173 );
and \U$22889 ( \31979 , RIfea1880_8182, \9175 );
and \U$22890 ( \31980 , RIfea19e8_8183, \9177 );
and \U$22891 ( \31981 , RIfc72110_6320, \9179 );
and \U$22892 ( \31982 , RIfc49b98_5861, \9181 );
and \U$22893 ( \31983 , RIfcca0b8_7321, \9183 );
and \U$22894 ( \31984 , RIfc71738_6313, \9185 );
or \U$22895 ( \31985 , \31921 , \31922 , \31923 , \31924 , \31925 , \31926 , \31927 , \31928 , \31929 , \31930 , \31931 , \31932 , \31933 , \31934 , \31935 , \31936 , \31937 , \31938 , \31939 , \31940 , \31941 , \31942 , \31943 , \31944 , \31945 , \31946 , \31947 , \31948 , \31949 , \31950 , \31951 , \31952 , \31953 , \31954 , \31955 , \31956 , \31957 , \31958 , \31959 , \31960 , \31961 , \31962 , \31963 , \31964 , \31965 , \31966 , \31967 , \31968 , \31969 , \31970 , \31971 , \31972 , \31973 , \31974 , \31975 , \31976 , \31977 , \31978 , \31979 , \31980 , \31981 , \31982 , \31983 , \31984 );
and \U$22896 ( \31986 , RIfc4ca00_5894, \9188 );
and \U$22897 ( \31987 , RIfc71030_6308, \9190 );
and \U$22898 ( \31988 , RIfcde428_7551, \9192 );
and \U$22899 ( \31989 , RIe1fad48_4231, \9194 );
and \U$22900 ( \31990 , RIfc70bf8_6305, \9196 );
and \U$22901 ( \31991 , RIfc63a70_6156, \9198 );
and \U$22902 ( \31992 , RIfca7db0_6932, \9200 );
and \U$22903 ( \31993 , RIe1f62c0_4178, \9202 );
and \U$22904 ( \31994 , RIfcada80_6998, \9204 );
and \U$22905 ( \31995 , RIfc6fde8_6295, \9206 );
and \U$22906 ( \31996 , RIfc6f578_6289, \9208 );
and \U$22907 ( \31997 , RIe1f3f98_4153, \9210 );
and \U$22908 ( \31998 , RIfcde158_7549, \9212 );
and \U$22909 ( \31999 , RIfcad378_6993, \9214 );
and \U$22910 ( \32000 , RIfc65f00_6182, \9216 );
and \U$22911 ( \32001 , RIe1eeca0_4094, \9218 );
and \U$22912 ( \32002 , RIe1ec540_4066, \9220 );
and \U$22913 ( \32003 , RIe1e9840_4034, \9222 );
and \U$22914 ( \32004 , RIe1e6b40_4002, \9224 );
and \U$22915 ( \32005 , RIe1e3e40_3970, \9226 );
and \U$22916 ( \32006 , RIe1e1140_3938, \9228 );
and \U$22917 ( \32007 , RIe1de440_3906, \9230 );
and \U$22918 ( \32008 , RIe1db740_3874, \9232 );
and \U$22919 ( \32009 , RIe1d8a40_3842, \9234 );
and \U$22920 ( \32010 , RIe1d3040_3778, \9236 );
and \U$22921 ( \32011 , RIe1d0340_3746, \9238 );
and \U$22922 ( \32012 , RIe1cd640_3714, \9240 );
and \U$22923 ( \32013 , RIe1ca940_3682, \9242 );
and \U$22924 ( \32014 , RIe1c7c40_3650, \9244 );
and \U$22925 ( \32015 , RIe1c4f40_3618, \9246 );
and \U$22926 ( \32016 , RIe1c2240_3586, \9248 );
and \U$22927 ( \32017 , RIe1bf540_3554, \9250 );
and \U$22928 ( \32018 , RIfc69308_6219, \9252 );
and \U$22929 ( \32019 , RIfccba08_7339, \9254 );
and \U$22930 ( \32020 , RIe1b9f78_3493, \9256 );
and \U$22931 ( \32021 , RIe1b7db8_3469, \9258 );
and \U$22932 ( \32022 , RIfccd628_7359, \9260 );
and \U$22933 ( \32023 , RIfc69740_6222, \9262 );
and \U$22934 ( \32024 , RIe1b5bf8_3445, \9264 );
and \U$22935 ( \32025 , RIe1b4578_3429, \9266 );
and \U$22936 ( \32026 , RIfccf950_7384, \9268 );
and \U$22937 ( \32027 , RIf148088_5279, \9270 );
and \U$22938 ( \32028 , RIe1b3060_3414, \9272 );
and \U$22939 ( \32029 , RIe1b1710_3396, \9274 );
and \U$22940 ( \32030 , RIfc9f818_6837, \9276 );
and \U$22941 ( \32031 , RIfcb9c90_7136, \9278 );
and \U$22942 ( \32032 , RIe1acf58_3345, \9280 );
and \U$22943 ( \32033 , RIe1ab770_3328, \9282 );
and \U$22944 ( \32034 , RIe1a9880_3306, \9284 );
and \U$22945 ( \32035 , RIe1a6b80_3274, \9286 );
and \U$22946 ( \32036 , RIe1a3e80_3242, \9288 );
and \U$22947 ( \32037 , RIe1a1180_3210, \9290 );
and \U$22948 ( \32038 , RIe18d680_2986, \9292 );
and \U$22949 ( \32039 , RIe179b80_2762, \9294 );
and \U$22950 ( \32040 , RIe2274d8_4737, \9296 );
and \U$22951 ( \32041 , RIe21c0d8_4609, \9298 );
and \U$22952 ( \32042 , RIe2058d8_4353, \9300 );
and \U$22953 ( \32043 , RIe1ff938_4285, \9302 );
and \U$22954 ( \32044 , RIe1f8cf0_4208, \9304 );
and \U$22955 ( \32045 , RIe1f1838_4125, \9306 );
and \U$22956 ( \32046 , RIe1d5d40_3810, \9308 );
and \U$22957 ( \32047 , RIe1bc840_3522, \9310 );
and \U$22958 ( \32048 , RIe1af6b8_3373, \9312 );
and \U$22959 ( \32049 , RIe171cf0_2672, \9314 );
or \U$22960 ( \32050 , \31986 , \31987 , \31988 , \31989 , \31990 , \31991 , \31992 , \31993 , \31994 , \31995 , \31996 , \31997 , \31998 , \31999 , \32000 , \32001 , \32002 , \32003 , \32004 , \32005 , \32006 , \32007 , \32008 , \32009 , \32010 , \32011 , \32012 , \32013 , \32014 , \32015 , \32016 , \32017 , \32018 , \32019 , \32020 , \32021 , \32022 , \32023 , \32024 , \32025 , \32026 , \32027 , \32028 , \32029 , \32030 , \32031 , \32032 , \32033 , \32034 , \32035 , \32036 , \32037 , \32038 , \32039 , \32040 , \32041 , \32042 , \32043 , \32044 , \32045 , \32046 , \32047 , \32048 , \32049 );
or \U$22961 ( \32051 , \31985 , \32050 );
_DC g65d2 ( \32052_nG65d2 , \32051 , \9323 );
and g65d3 ( \32053_nG65d3 , \31920_nG65d1 , \32052_nG65d2 );
buf \U$22962 ( \32054 , \32053_nG65d3 );
and \U$22963 ( \32055 , \32054 , \10691 );
nor \U$22964 ( \32056 , \31788 , \32055 );
xnor \U$22965 ( \32057 , \32056 , \10980 );
and \U$22966 ( \32058 , \29084 , \11574 );
and \U$22967 ( \32059 , \30268 , \11278 );
nor \U$22968 ( \32060 , \32058 , \32059 );
xnor \U$22969 ( \32061 , \32060 , \11580 );
xor \U$22970 ( \32062 , \32057 , \32061 );
_DC g63e8 ( \32063_nG63e8 , \31919 , \9597 );
_DC g646c ( \32064_nG646c , \32051 , \9323 );
xor g646d ( \32065_nG646d , \32063_nG63e8 , \32064_nG646c );
buf \U$22971 ( \32066 , \32065_nG646d );
xor \U$22972 ( \32067 , \32066 , \30810 );
and \U$22973 ( \32068 , \10687 , \32067 );
xor \U$22974 ( \32069 , \32062 , \32068 );
xor \U$22975 ( \32070 , \31787 , \32069 );
and \U$22976 ( \32071 , \27313 , \12790 );
and \U$22977 ( \32072 , \28534 , \12461 );
nor \U$22978 ( \32073 , \32071 , \32072 );
xnor \U$22979 ( \32074 , \32073 , \12780 );
and \U$22980 ( \32075 , \22556 , \16635 );
and \U$22981 ( \32076 , \23617 , \16301 );
nor \U$22982 ( \32077 , \32075 , \32076 );
xnor \U$22983 ( \32078 , \32077 , \16625 );
xor \U$22984 ( \32079 , \32074 , \32078 );
and \U$22985 ( \32080 , \14024 , \25826 );
and \U$22986 ( \32081 , \14950 , \25264 );
nor \U$22987 ( \32082 , \32080 , \32081 );
xnor \U$22988 ( \32083 , \32082 , \25773 );
xor \U$22989 ( \32084 , \32079 , \32083 );
xor \U$22990 ( \32085 , \32070 , \32084 );
xor \U$22991 ( \32086 , \31773 , \32085 );
xor \U$22992 ( \32087 , \31764 , \32086 );
and \U$22993 ( \32088 , \30878 , \30882 );
and \U$22994 ( \32089 , \30882 , \30927 );
and \U$22995 ( \32090 , \30878 , \30927 );
or \U$22996 ( \32091 , \32088 , \32089 , \32090 );
and \U$22997 ( \32092 , \30837 , \30841 );
and \U$22998 ( \32093 , \30841 , \30846 );
and \U$22999 ( \32094 , \30837 , \30846 );
or \U$23000 ( \32095 , \32092 , \32093 , \32094 );
and \U$23001 ( \32096 , \30897 , \30911 );
and \U$23002 ( \32097 , \30911 , \30926 );
and \U$23003 ( \32098 , \30897 , \30926 );
or \U$23004 ( \32099 , \32096 , \32097 , \32098 );
xor \U$23005 ( \32100 , \32095 , \32099 );
and \U$23006 ( \32101 , \30861 , \30865 );
and \U$23007 ( \32102 , \30865 , \30870 );
and \U$23008 ( \32103 , \30861 , \30870 );
or \U$23009 ( \32104 , \32101 , \32102 , \32103 );
and \U$23010 ( \32105 , \30805 , \30814 );
xor \U$23011 ( \32106 , \32104 , \32105 );
and \U$23012 ( \32107 , \10988 , \30823 );
and \U$23013 ( \32108 , \11270 , \30246 );
nor \U$23014 ( \32109 , \32107 , \32108 );
xnor \U$23015 ( \32110 , \32109 , \30813 );
xor \U$23016 ( \32111 , \32106 , \32110 );
xor \U$23017 ( \32112 , \32100 , \32111 );
xor \U$23018 ( \32113 , \32091 , \32112 );
and \U$23019 ( \32114 , \30852 , \30856 );
and \U$23020 ( \32115 , \30856 , \30871 );
and \U$23021 ( \32116 , \30852 , \30871 );
or \U$23022 ( \32117 , \32114 , \32115 , \32116 );
and \U$23023 ( \32118 , \30887 , \30891 );
and \U$23024 ( \32119 , \30891 , \30896 );
and \U$23025 ( \32120 , \30887 , \30896 );
or \U$23026 ( \32121 , \32118 , \32119 , \32120 );
and \U$23027 ( \32122 , \30901 , \30905 );
and \U$23028 ( \32123 , \30905 , \30910 );
and \U$23029 ( \32124 , \30901 , \30910 );
or \U$23030 ( \32125 , \32122 , \32123 , \32124 );
xor \U$23031 ( \32126 , \32121 , \32125 );
and \U$23032 ( \32127 , \30916 , \30920 );
and \U$23033 ( \32128 , \30920 , \30925 );
and \U$23034 ( \32129 , \30916 , \30925 );
or \U$23035 ( \32130 , \32127 , \32128 , \32129 );
xor \U$23036 ( \32131 , \32126 , \32130 );
xor \U$23037 ( \32132 , \32117 , \32131 );
and \U$23038 ( \32133 , \30815 , \30819 );
and \U$23039 ( \32134 , \30819 , \30827 );
and \U$23040 ( \32135 , \30815 , \30827 );
or \U$23041 ( \32136 , \32133 , \32134 , \32135 );
and \U$23042 ( \32137 , \24199 , \15336 );
and \U$23043 ( \32138 , \25272 , \14963 );
nor \U$23044 ( \32139 , \32137 , \32138 );
xnor \U$23045 ( \32140 , \32139 , \15342 );
and \U$23046 ( \32141 , \16655 , \22542 );
and \U$23047 ( \32142 , \17627 , \22103 );
nor \U$23048 ( \32143 , \32141 , \32142 );
xnor \U$23049 ( \32144 , \32143 , \22548 );
xor \U$23050 ( \32145 , \32140 , \32144 );
and \U$23051 ( \32146 , \15321 , \24138 );
and \U$23052 ( \32147 , \16267 , \23630 );
nor \U$23053 ( \32148 , \32146 , \32147 );
xnor \U$23054 ( \32149 , \32148 , \24144 );
xor \U$23055 ( \32150 , \32145 , \32149 );
xor \U$23056 ( \32151 , \32136 , \32150 );
and \U$23057 ( \32152 , \25815 , \14054 );
and \U$23058 ( \32153 , \26829 , \13692 );
nor \U$23059 ( \32154 , \32152 , \32153 );
xnor \U$23060 ( \32155 , \32154 , \14035 );
and \U$23061 ( \32156 , \19558 , \19534 );
and \U$23062 ( \32157 , \20544 , \19045 );
nor \U$23063 ( \32158 , \32156 , \32157 );
xnor \U$23064 ( \32159 , \32158 , \19540 );
xor \U$23065 ( \32160 , \32155 , \32159 );
and \U$23066 ( \32161 , \18035 , \21005 );
and \U$23067 ( \32162 , \19032 , \20557 );
nor \U$23068 ( \32163 , \32161 , \32162 );
xnor \U$23069 ( \32164 , \32163 , \21011 );
xor \U$23070 ( \32165 , \32160 , \32164 );
xor \U$23071 ( \32166 , \32151 , \32165 );
xor \U$23072 ( \32167 , \32132 , \32166 );
xor \U$23073 ( \32168 , \32113 , \32167 );
xor \U$23074 ( \32169 , \32087 , \32168 );
and \U$23075 ( \32170 , \30521 , \30525 );
and \U$23076 ( \32171 , \30525 , \30929 );
and \U$23077 ( \32172 , \30521 , \30929 );
or \U$23078 ( \32173 , \32170 , \32171 , \32172 );
xor \U$23079 ( \32174 , \32169 , \32173 );
and \U$23080 ( \32175 , \30930 , \30934 );
and \U$23081 ( \32176 , \30935 , \30938 );
or \U$23082 ( \32177 , \32175 , \32176 );
xor \U$23083 ( \32178 , \32174 , \32177 );
buf g9bb4 ( \32179_nG9bb4 , \32178 );
and \U$23084 ( \32180 , \10704 , \32179_nG9bb4 );
or \U$23085 ( \32181 , \31760 , \32180 );
xor \U$23086 ( \32182 , \10703 , \32181 );
buf \U$23087 ( \32183 , \32182 );
buf \U$23089 ( \32184 , \32183 );
xor \U$23090 ( \32185 , \31759 , \32184 );
buf \U$23091 ( \32186 , \32185 );
xor \U$23092 ( \32187 , \31707 , \32186 );
buf \U$23093 ( \32188 , \32187 );
xor \U$23094 ( \32189 , \31653 , \32188 );
and \U$23095 ( \32190 , \31051 , \31056 );
and \U$23096 ( \32191 , \31051 , \31062 );
and \U$23097 ( \32192 , \31056 , \31062 );
or \U$23098 ( \32193 , \32190 , \32191 , \32192 );
buf \U$23099 ( \32194 , \32193 );
and \U$23100 ( \32195 , \30510 , \30515 );
and \U$23101 ( \32196 , \30510 , \30945 );
and \U$23102 ( \32197 , \30515 , \30945 );
or \U$23103 ( \32198 , \32195 , \32196 , \32197 );
buf \U$23104 ( \32199 , \32198 );
xor \U$23105 ( \32200 , \32194 , \32199 );
and \U$23106 ( \32201 , \30470 , \30487 );
and \U$23107 ( \32202 , \30470 , \30494 );
and \U$23108 ( \32203 , \30487 , \30494 );
or \U$23109 ( \32204 , \32201 , \32202 , \32203 );
buf \U$23110 ( \32205 , \32204 );
and \U$23111 ( \32206 , \30958 , \30984 );
and \U$23112 ( \32207 , \30958 , \30991 );
and \U$23113 ( \32208 , \30984 , \30991 );
or \U$23114 ( \32209 , \32206 , \32207 , \32208 );
buf \U$23115 ( \32210 , \32209 );
xor \U$23116 ( \32211 , \32205 , \32210 );
and \U$23117 ( \32212 , \30969 , \30975 );
and \U$23118 ( \32213 , \30969 , \30982 );
and \U$23119 ( \32214 , \30975 , \30982 );
or \U$23120 ( \32215 , \32212 , \32213 , \32214 );
buf \U$23121 ( \32216 , \32215 );
and \U$23122 ( \32217 , \29853 , \10995_nG9c0b );
and \U$23123 ( \32218 , \29850 , \11283_nG9c08 );
or \U$23124 ( \32219 , \32217 , \32218 );
xor \U$23125 ( \32220 , \29849 , \32219 );
buf \U$23126 ( \32221 , \32220 );
buf \U$23128 ( \32222 , \32221 );
and \U$23129 ( \32223 , \28118 , \11598_nG9c05 );
and \U$23130 ( \32224 , \28115 , \12470_nG9c02 );
or \U$23131 ( \32225 , \32223 , \32224 );
xor \U$23132 ( \32226 , \28114 , \32225 );
buf \U$23133 ( \32227 , \32226 );
buf \U$23135 ( \32228 , \32227 );
xor \U$23136 ( \32229 , \32222 , \32228 );
buf \U$23137 ( \32230 , \32229 );
xor \U$23138 ( \32231 , \32216 , \32230 );
and \U$23139 ( \32232 , \23201 , \15373_nG9bf3 );
and \U$23140 ( \32233 , \23198 , \16315_nG9bf0 );
or \U$23141 ( \32234 , \32232 , \32233 );
xor \U$23142 ( \32235 , \23197 , \32234 );
buf \U$23143 ( \32236 , \32235 );
buf \U$23145 ( \32237 , \32236 );
xor \U$23146 ( \32238 , \32231 , \32237 );
buf \U$23147 ( \32239 , \32238 );
xor \U$23148 ( \32240 , \32211 , \32239 );
buf \U$23149 ( \32241 , \32240 );
and \U$23150 ( \32242 , \13370 , \25860_nG9bc9 );
and \U$23151 ( \32243 , \13367 , \26887_nG9bc6 );
or \U$23152 ( \32244 , \32242 , \32243 );
xor \U$23153 ( \32245 , \13366 , \32244 );
buf \U$23154 ( \32246 , \32245 );
buf \U$23156 ( \32247 , \32246 );
xor \U$23157 ( \32248 , \32241 , \32247 );
and \U$23158 ( \32249 , \10421 , \29179_nG9bbd );
and \U$23159 ( \32250 , \10418 , \30366_nG9bba );
or \U$23160 ( \32251 , \32249 , \32250 );
xor \U$23161 ( \32252 , \10417 , \32251 );
buf \U$23162 ( \32253 , \32252 );
buf \U$23164 ( \32254 , \32253 );
xor \U$23165 ( \32255 , \32248 , \32254 );
buf \U$23166 ( \32256 , \32255 );
xor \U$23167 ( \32257 , \32200 , \32256 );
buf \U$23168 ( \32258 , \32257 );
xor \U$23169 ( \32259 , \32189 , \32258 );
and \U$23170 ( \32260 , \31643 , \32259 );
and \U$23171 ( \32261 , \31647 , \32259 );
or \U$23172 ( \32262 , \31648 , \32260 , \32261 );
and \U$23173 ( \32263 , \31079 , \31083 );
and \U$23174 ( \32264 , \31079 , \31642 );
and \U$23175 ( \32265 , \31083 , \31642 );
or \U$23176 ( \32266 , \32263 , \32264 , \32265 );
xor \U$23177 ( \32267 , \32262 , \32266 );
and \U$23178 ( \32268 , \32194 , \32199 );
and \U$23179 ( \32269 , \32194 , \32256 );
and \U$23180 ( \32270 , \32199 , \32256 );
or \U$23181 ( \32271 , \32268 , \32269 , \32270 );
buf \U$23182 ( \32272 , \32271 );
and \U$23183 ( \32273 , \31719 , \31725 );
and \U$23184 ( \32274 , \31719 , \31732 );
and \U$23185 ( \32275 , \31725 , \31732 );
or \U$23186 ( \32276 , \32273 , \32274 , \32275 );
buf \U$23187 ( \32277 , \32276 );
and \U$23188 ( \32278 , \31632 , \31639 );
buf \U$23189 ( \32279 , \32278 );
buf \U$23191 ( \32280 , \32279 );
and \U$23192 ( \32281 , \29853 , \11283_nG9c08 );
and \U$23193 ( \32282 , \29850 , \11598_nG9c05 );
or \U$23194 ( \32283 , \32281 , \32282 );
xor \U$23195 ( \32284 , \29849 , \32283 );
buf \U$23196 ( \32285 , \32284 );
buf \U$23198 ( \32286 , \32285 );
xor \U$23199 ( \32287 , \32280 , \32286 );
buf \U$23200 ( \32288 , \32287 );
and \U$23201 ( \32289 , \31636 , \10694_nG9c0e );
and \U$23202 ( \32290 , \31633 , \10995_nG9c0b );
or \U$23203 ( \32291 , \32289 , \32290 );
xor \U$23204 ( \32292 , \31632 , \32291 );
buf \U$23205 ( \32293 , \32292 );
buf \U$23207 ( \32294 , \32293 );
xor \U$23208 ( \32295 , \32288 , \32294 );
and \U$23209 ( \32296 , \28118 , \12470_nG9c02 );
and \U$23210 ( \32297 , \28115 , \12801_nG9bff );
or \U$23211 ( \32298 , \32296 , \32297 );
xor \U$23212 ( \32299 , \28114 , \32298 );
buf \U$23213 ( \32300 , \32299 );
buf \U$23215 ( \32301 , \32300 );
xor \U$23216 ( \32302 , \32295 , \32301 );
buf \U$23217 ( \32303 , \32302 );
xor \U$23218 ( \32304 , \32277 , \32303 );
and \U$23219 ( \32305 , \23201 , \16315_nG9bf0 );
and \U$23220 ( \32306 , \23198 , \16680_nG9bed );
or \U$23221 ( \32307 , \32305 , \32306 );
xor \U$23222 ( \32308 , \23197 , \32307 );
buf \U$23223 ( \32309 , \32308 );
buf \U$23225 ( \32310 , \32309 );
xor \U$23226 ( \32311 , \32304 , \32310 );
buf \U$23227 ( \32312 , \32311 );
and \U$23228 ( \32313 , \20155 , \19091_nG9be4 );
and \U$23229 ( \32314 , \20152 , \19586_nG9be1 );
or \U$23230 ( \32315 , \32313 , \32314 );
xor \U$23231 ( \32316 , \20151 , \32315 );
buf \U$23232 ( \32317 , \32316 );
buf \U$23234 ( \32318 , \32317 );
xor \U$23235 ( \32319 , \32312 , \32318 );
and \U$23236 ( \32320 , \18702 , \20608_nG9bde );
and \U$23237 ( \32321 , \18699 , \21086_nG9bdb );
or \U$23238 ( \32322 , \32320 , \32321 );
xor \U$23239 ( \32323 , \18698 , \32322 );
buf \U$23240 ( \32324 , \32323 );
buf \U$23242 ( \32325 , \32324 );
xor \U$23243 ( \32326 , \32319 , \32325 );
buf \U$23244 ( \32327 , \32326 );
and \U$23245 ( \32328 , \13370 , \26887_nG9bc6 );
and \U$23246 ( \32329 , \13367 , \27416_nG9bc3 );
or \U$23247 ( \32330 , \32328 , \32329 );
xor \U$23248 ( \32331 , \13366 , \32330 );
buf \U$23249 ( \32332 , \32331 );
buf \U$23251 ( \32333 , \32332 );
xor \U$23252 ( \32334 , \32327 , \32333 );
and \U$23253 ( \32335 , \12157 , \28602_nG9bc0 );
and \U$23254 ( \32336 , \12154 , \29179_nG9bbd );
or \U$23255 ( \32337 , \32335 , \32336 );
xor \U$23256 ( \32338 , \12153 , \32337 );
buf \U$23257 ( \32339 , \32338 );
buf \U$23259 ( \32340 , \32339 );
xor \U$23260 ( \32341 , \32334 , \32340 );
buf \U$23261 ( \32342 , \32341 );
and \U$23262 ( \32343 , \31674 , \31680 );
and \U$23263 ( \32344 , \31674 , \31687 );
and \U$23264 ( \32345 , \31680 , \31687 );
or \U$23265 ( \32346 , \32343 , \32344 , \32345 );
buf \U$23266 ( \32347 , \32346 );
and \U$23267 ( \32348 , \15940 , \23696_nG9bd2 );
and \U$23268 ( \32349 , \15937 , \24226_nG9bcf );
or \U$23269 ( \32350 , \32348 , \32349 );
xor \U$23270 ( \32351 , \15936 , \32350 );
buf \U$23271 ( \32352 , \32351 );
buf \U$23273 ( \32353 , \32352 );
xor \U$23274 ( \32354 , \32347 , \32353 );
and \U$23275 ( \32355 , \14631 , \25298_nG9bcc );
and \U$23276 ( \32356 , \14628 , \25860_nG9bc9 );
or \U$23277 ( \32357 , \32355 , \32356 );
xor \U$23278 ( \32358 , \14627 , \32357 );
buf \U$23279 ( \32359 , \32358 );
buf \U$23281 ( \32360 , \32359 );
xor \U$23282 ( \32361 , \32354 , \32360 );
buf \U$23283 ( \32362 , \32361 );
xor \U$23284 ( \32363 , \32342 , \32362 );
and \U$23285 ( \32364 , \32241 , \32247 );
and \U$23286 ( \32365 , \32241 , \32254 );
and \U$23287 ( \32366 , \32247 , \32254 );
or \U$23288 ( \32367 , \32364 , \32365 , \32366 );
buf \U$23289 ( \32368 , \32367 );
xor \U$23290 ( \32369 , \32363 , \32368 );
buf \U$23291 ( \32370 , \32369 );
xor \U$23292 ( \32371 , \32272 , \32370 );
and \U$23293 ( \32372 , \31663 , \31698 );
and \U$23294 ( \32373 , \31663 , \31704 );
and \U$23295 ( \32374 , \31698 , \31704 );
or \U$23296 ( \32375 , \32372 , \32373 , \32374 );
buf \U$23297 ( \32376 , \32375 );
xor \U$23298 ( \32377 , \32371 , \32376 );
buf \U$23299 ( \32378 , \32377 );
and \U$23300 ( \32379 , \31658 , \31706 );
and \U$23301 ( \32380 , \31658 , \32186 );
and \U$23302 ( \32381 , \31706 , \32186 );
or \U$23303 ( \32382 , \32379 , \32380 , \32381 );
buf \U$23304 ( \32383 , \32382 );
xor \U$23305 ( \32384 , \32378 , \32383 );
and \U$23306 ( \32385 , \32216 , \32230 );
and \U$23307 ( \32386 , \32216 , \32237 );
and \U$23308 ( \32387 , \32230 , \32237 );
or \U$23309 ( \32388 , \32385 , \32386 , \32387 );
buf \U$23310 ( \32389 , \32388 );
and \U$23311 ( \32390 , \32222 , \32228 );
buf \U$23312 ( \32391 , \32390 );
and \U$23313 ( \32392 , \26431 , \13705_nG9bfc );
and \U$23314 ( \32393 , \26428 , \14070_nG9bf9 );
or \U$23315 ( \32394 , \32392 , \32393 );
xor \U$23316 ( \32395 , \26427 , \32394 );
buf \U$23317 ( \32396 , \32395 );
buf \U$23319 ( \32397 , \32396 );
xor \U$23320 ( \32398 , \32391 , \32397 );
and \U$23321 ( \32399 , \24792 , \14984_nG9bf6 );
and \U$23322 ( \32400 , \24789 , \15373_nG9bf3 );
or \U$23323 ( \32401 , \32399 , \32400 );
xor \U$23324 ( \32402 , \24788 , \32401 );
buf \U$23325 ( \32403 , \32402 );
buf \U$23327 ( \32404 , \32403 );
xor \U$23328 ( \32405 , \32398 , \32404 );
buf \U$23329 ( \32406 , \32405 );
xor \U$23330 ( \32407 , \32389 , \32406 );
and \U$23331 ( \32408 , \21658 , \17665_nG9bea );
and \U$23332 ( \32409 , \21655 , \18107_nG9be7 );
or \U$23333 ( \32410 , \32408 , \32409 );
xor \U$23334 ( \32411 , \21654 , \32410 );
buf \U$23335 ( \32412 , \32411 );
buf \U$23337 ( \32413 , \32412 );
xor \U$23338 ( \32414 , \32407 , \32413 );
buf \U$23339 ( \32415 , \32414 );
and \U$23340 ( \32416 , \31717 , \31734 );
and \U$23341 ( \32417 , \31717 , \31741 );
and \U$23342 ( \32418 , \31734 , \31741 );
or \U$23343 ( \32419 , \32416 , \32417 , \32418 );
buf \U$23344 ( \32420 , \32419 );
xor \U$23345 ( \32421 , \32415 , \32420 );
and \U$23346 ( \32422 , \17297 , \22129_nG9bd8 );
and \U$23347 ( \32423 , \17294 , \22629_nG9bd5 );
or \U$23348 ( \32424 , \32422 , \32423 );
xor \U$23349 ( \32425 , \17293 , \32424 );
buf \U$23350 ( \32426 , \32425 );
buf \U$23352 ( \32427 , \32426 );
xor \U$23353 ( \32428 , \32421 , \32427 );
buf \U$23354 ( \32429 , \32428 );
and \U$23355 ( \32430 , \31743 , \31749 );
and \U$23356 ( \32431 , \31743 , \31756 );
and \U$23357 ( \32432 , \31749 , \31756 );
or \U$23358 ( \32433 , \32430 , \32431 , \32432 );
buf \U$23359 ( \32434 , \32433 );
xor \U$23360 ( \32435 , \32429 , \32434 );
and \U$23361 ( \32436 , \31668 , \31689 );
and \U$23362 ( \32437 , \31668 , \31696 );
and \U$23363 ( \32438 , \31689 , \31696 );
or \U$23364 ( \32439 , \32436 , \32437 , \32438 );
buf \U$23365 ( \32440 , \32439 );
xor \U$23366 ( \32441 , \32435 , \32440 );
buf \U$23367 ( \32442 , \32441 );
and \U$23368 ( \32443 , \32205 , \32210 );
and \U$23369 ( \32444 , \32205 , \32239 );
and \U$23370 ( \32445 , \32210 , \32239 );
or \U$23371 ( \32446 , \32443 , \32444 , \32445 );
buf \U$23372 ( \32447 , \32446 );
and \U$23373 ( \32448 , \10421 , \30366_nG9bba );
and \U$23374 ( \32449 , \10418 , \30940_nG9bb7 );
or \U$23375 ( \32450 , \32448 , \32449 );
xor \U$23376 ( \32451 , \10417 , \32450 );
buf \U$23377 ( \32452 , \32451 );
buf \U$23379 ( \32453 , \32452 );
xor \U$23380 ( \32454 , \32447 , \32453 );
and \U$23381 ( \32455 , \10707 , \32179_nG9bb4 );
and \U$23382 ( \32456 , \32091 , \32112 );
and \U$23383 ( \32457 , \32112 , \32167 );
and \U$23384 ( \32458 , \32091 , \32167 );
or \U$23385 ( \32459 , \32456 , \32457 , \32458 );
and \U$23386 ( \32460 , \32095 , \32099 );
and \U$23387 ( \32461 , \32099 , \32111 );
and \U$23388 ( \32462 , \32095 , \32111 );
or \U$23389 ( \32463 , \32460 , \32461 , \32462 );
and \U$23390 ( \32464 , \32117 , \32131 );
and \U$23391 ( \32465 , \32131 , \32166 );
and \U$23392 ( \32466 , \32117 , \32166 );
or \U$23393 ( \32467 , \32464 , \32465 , \32466 );
xor \U$23394 ( \32468 , \32463 , \32467 );
and \U$23395 ( \32469 , \32121 , \32125 );
and \U$23396 ( \32470 , \32125 , \32130 );
and \U$23397 ( \32471 , \32121 , \32130 );
or \U$23398 ( \32472 , \32469 , \32470 , \32471 );
and \U$23399 ( \32473 , \23617 , \16635 );
and \U$23400 ( \32474 , \24199 , \16301 );
nor \U$23401 ( \32475 , \32473 , \32474 );
xnor \U$23402 ( \32476 , \32475 , \16625 );
and \U$23403 ( \32477 , \14950 , \25826 );
and \U$23404 ( \32478 , \15321 , \25264 );
nor \U$23405 ( \32479 , \32477 , \32478 );
xnor \U$23406 ( \32480 , \32479 , \25773 );
xor \U$23407 ( \32481 , \32476 , \32480 );
and \U$23408 ( \32482 , \13679 , \27397 );
and \U$23409 ( \32483 , \14024 , \26807 );
nor \U$23410 ( \32484 , \32482 , \32483 );
xnor \U$23411 ( \32485 , \32484 , \27295 );
xor \U$23412 ( \32486 , \32481 , \32485 );
xor \U$23413 ( \32487 , \32472 , \32486 );
and \U$23414 ( \32488 , \28534 , \12790 );
and \U$23415 ( \32489 , \29084 , \12461 );
nor \U$23416 ( \32490 , \32488 , \32489 );
xnor \U$23417 ( \32491 , \32490 , \12780 );
and \U$23418 ( \32492 , \17627 , \22542 );
and \U$23419 ( \32493 , \18035 , \22103 );
nor \U$23420 ( \32494 , \32492 , \32493 );
xnor \U$23421 ( \32495 , \32494 , \22548 );
xor \U$23422 ( \32496 , \32491 , \32495 );
and \U$23423 ( \32497 , \16267 , \24138 );
and \U$23424 ( \32498 , \16655 , \23630 );
nor \U$23425 ( \32499 , \32497 , \32498 );
xnor \U$23426 ( \32500 , \32499 , \24144 );
xor \U$23427 ( \32501 , \32496 , \32500 );
xor \U$23428 ( \32502 , \32487 , \32501 );
xor \U$23429 ( \32503 , \32468 , \32502 );
xor \U$23430 ( \32504 , \32459 , \32503 );
and \U$23431 ( \32505 , \31768 , \31772 );
and \U$23432 ( \32506 , \31772 , \32085 );
and \U$23433 ( \32507 , \31768 , \32085 );
or \U$23434 ( \32508 , \32505 , \32506 , \32507 );
and \U$23435 ( \32509 , \32104 , \32105 );
and \U$23436 ( \32510 , \32105 , \32110 );
and \U$23437 ( \32511 , \32104 , \32110 );
or \U$23438 ( \32512 , \32509 , \32510 , \32511 );
and \U$23439 ( \32513 , \31777 , \31781 );
and \U$23440 ( \32514 , \31781 , \31786 );
and \U$23441 ( \32515 , \31777 , \31786 );
or \U$23442 ( \32516 , \32513 , \32514 , \32515 );
and \U$23443 ( \32517 , \32074 , \32078 );
and \U$23444 ( \32518 , \32078 , \32083 );
and \U$23445 ( \32519 , \32074 , \32083 );
or \U$23446 ( \32520 , \32517 , \32518 , \32519 );
xor \U$23447 ( \32521 , \32516 , \32520 );
and \U$23448 ( \32522 , \32140 , \32144 );
and \U$23449 ( \32523 , \32144 , \32149 );
and \U$23450 ( \32524 , \32140 , \32149 );
or \U$23451 ( \32525 , \32522 , \32523 , \32524 );
xor \U$23452 ( \32526 , \32521 , \32525 );
xor \U$23453 ( \32527 , \32512 , \32526 );
and \U$23454 ( \32528 , \32054 , \10983 );
and \U$23455 ( \32529 , RIdec6350_719, \9333 );
and \U$23456 ( \32530 , RIdec3650_687, \9335 );
and \U$23457 ( \32531 , RIfcaf3d0_7016, \9337 );
and \U$23458 ( \32532 , RIdec0950_655, \9339 );
and \U$23459 ( \32533 , RIfc6a280_6230, \9341 );
and \U$23460 ( \32534 , RIdebdc50_623, \9343 );
and \U$23461 ( \32535 , RIdebaf50_591, \9345 );
and \U$23462 ( \32536 , RIdeb8250_559, \9347 );
and \U$23463 ( \32537 , RIfc42f50_5784, \9349 );
and \U$23464 ( \32538 , RIdeb2850_495, \9351 );
and \U$23465 ( \32539 , RIfc981f8_6753, \9353 );
and \U$23466 ( \32540 , RIdeafb50_463, \9355 );
and \U$23467 ( \32541 , RIfc8c6f0_6620, \9357 );
and \U$23468 ( \32542 , RIdeac838_431, \9359 );
and \U$23469 ( \32543 , RIdea5f38_399, \9361 );
and \U$23470 ( \32544 , RIde9f638_367, \9363 );
and \U$23471 ( \32545 , RIee1d4e8_4792, \9365 );
and \U$23472 ( \32546 , RIfcda648_7507, \9367 );
and \U$23473 ( \32547 , RIfcc6440_7278, \9369 );
and \U$23474 ( \32548 , RIfcd5620_7450, \9371 );
and \U$23475 ( \32549 , RIde92ac8_305, \9373 );
and \U$23476 ( \32550 , RIfea34a0_8202, \9375 );
and \U$23477 ( \32551 , RIfea31d0_8200, \9377 );
and \U$23478 ( \32552 , RIfea3338_8201, \9379 );
and \U$23479 ( \32553 , RIfcb6b58_7101, \9381 );
and \U$23480 ( \32554 , RIfcb6888_7099, \9383 );
and \U$23481 ( \32555 , RIfc9dd60_6818, \9385 );
and \U$23482 ( \32556 , RIee19708_4748, \9387 );
and \U$23483 ( \32557 , RIfc50c18_5941, \9389 );
and \U$23484 ( \32558 , RIe16c458_2609, \9391 );
and \U$23485 ( \32559 , RIfc80a80_6486, \9393 );
and \U$23486 ( \32560 , RIfec62e8_8375, \9395 );
and \U$23487 ( \32561 , RIe166350_2540, \9397 );
and \U$23488 ( \32562 , RIe163650_2508, \9399 );
and \U$23489 ( \32563 , RIee37d98_5094, \9401 );
and \U$23490 ( \32564 , RIe160950_2476, \9403 );
and \U$23491 ( \32565 , RIfcaa678_6961, \9405 );
and \U$23492 ( \32566 , RIe15dc50_2444, \9407 );
and \U$23493 ( \32567 , RIe158250_2380, \9409 );
and \U$23494 ( \32568 , RIe155550_2348, \9411 );
and \U$23495 ( \32569 , RIfea3ba8_8207, \9413 );
and \U$23496 ( \32570 , RIe152850_2316, \9415 );
and \U$23497 ( \32571 , RIee35638_5066, \9417 );
and \U$23498 ( \32572 , RIe14fb50_2284, \9419 );
and \U$23499 ( \32573 , RIfc62f30_6148, \9421 );
and \U$23500 ( \32574 , RIe14ce50_2252, \9423 );
and \U$23501 ( \32575 , RIe14a150_2220, \9425 );
and \U$23502 ( \32576 , RIe147450_2188, \9427 );
and \U$23503 ( \32577 , RIfc97f28_6751, \9429 );
and \U$23504 ( \32578 , RIfc89888_6587, \9431 );
and \U$23505 ( \32579 , RIfc8f558_6653, \9433 );
and \U$23506 ( \32580 , RIfc52838_5961, \9435 );
and \U$23507 ( \32581 , RIe141bb8_2125, \9437 );
and \U$23508 ( \32582 , RIe13f890_2100, \9439 );
and \U$23509 ( \32583 , RIdf3d798_2076, \9441 );
and \U$23510 ( \32584 , RIdf3b308_2050, \9443 );
and \U$23511 ( \32585 , RIee30a48_5012, \9445 );
and \U$23512 ( \32586 , RIfc568e8_6007, \9447 );
and \U$23513 ( \32587 , RIee2e9f0_4989, \9449 );
and \U$23514 ( \32588 , RIee2dbe0_4979, \9451 );
and \U$23515 ( \32589 , RIdf365b0_1995, \9453 );
and \U$23516 ( \32590 , RIfea38d8_8205, \9455 );
and \U$23517 ( \32591 , RIfea3a40_8206, \9457 );
and \U$23518 ( \32592 , RIdf2ff08_1922, \9459 );
or \U$23519 ( \32593 , \32529 , \32530 , \32531 , \32532 , \32533 , \32534 , \32535 , \32536 , \32537 , \32538 , \32539 , \32540 , \32541 , \32542 , \32543 , \32544 , \32545 , \32546 , \32547 , \32548 , \32549 , \32550 , \32551 , \32552 , \32553 , \32554 , \32555 , \32556 , \32557 , \32558 , \32559 , \32560 , \32561 , \32562 , \32563 , \32564 , \32565 , \32566 , \32567 , \32568 , \32569 , \32570 , \32571 , \32572 , \32573 , \32574 , \32575 , \32576 , \32577 , \32578 , \32579 , \32580 , \32581 , \32582 , \32583 , \32584 , \32585 , \32586 , \32587 , \32588 , \32589 , \32590 , \32591 , \32592 );
and \U$23520 ( \32594 , RIee2c6c8_4964, \9462 );
and \U$23521 ( \32595 , RIee2ac10_4945, \9464 );
and \U$23522 ( \32596 , RIee29590_4929, \9466 );
and \U$23523 ( \32597 , RIee28348_4916, \9468 );
and \U$23524 ( \32598 , RIdf2ad78_1864, \9470 );
and \U$23525 ( \32599 , RIdf28e88_1842, \9472 );
and \U$23526 ( \32600 , RIfea3608_8203, \9474 );
and \U$23527 ( \32601 , RIfea3770_8204, \9476 );
and \U$23528 ( \32602 , RIfcc0d10_7216, \9478 );
and \U$23529 ( \32603 , RIfc75c20_6362, \9480 );
and \U$23530 ( \32604 , RIfca50b0_6900, \9482 );
and \U$23531 ( \32605 , RIfc74e10_6352, \9484 );
and \U$23532 ( \32606 , RIfcc9410_7312, \9486 );
and \U$23533 ( \32607 , RIdf20620_1745, \9488 );
and \U$23534 ( \32608 , RIfc73628_6335, \9490 );
and \U$23535 ( \32609 , RIdf1a0e0_1673, \9492 );
and \U$23536 ( \32610 , RIdf17f20_1649, \9494 );
and \U$23537 ( \32611 , RIdf15220_1617, \9496 );
and \U$23538 ( \32612 , RIdf12520_1585, \9498 );
and \U$23539 ( \32613 , RIdf0f820_1553, \9500 );
and \U$23540 ( \32614 , RIdf0cb20_1521, \9502 );
and \U$23541 ( \32615 , RIdf09e20_1489, \9504 );
and \U$23542 ( \32616 , RIdf07120_1457, \9506 );
and \U$23543 ( \32617 , RIdf04420_1425, \9508 );
and \U$23544 ( \32618 , RIdefea20_1361, \9510 );
and \U$23545 ( \32619 , RIdefbd20_1329, \9512 );
and \U$23546 ( \32620 , RIdef9020_1297, \9514 );
and \U$23547 ( \32621 , RIdef6320_1265, \9516 );
and \U$23548 ( \32622 , RIdef3620_1233, \9518 );
and \U$23549 ( \32623 , RIdef0920_1201, \9520 );
and \U$23550 ( \32624 , RIdeedc20_1169, \9522 );
and \U$23551 ( \32625 , RIdeeaf20_1137, \9524 );
and \U$23552 ( \32626 , RIfcab8c0_6974, \9526 );
and \U$23553 ( \32627 , RIfc7c598_6437, \9528 );
and \U$23554 ( \32628 , RIfc5beb0_6068, \9530 );
and \U$23555 ( \32629 , RIfc58ee0_6034, \9532 );
and \U$23556 ( \32630 , RIdee5688_1074, \9534 );
and \U$23557 ( \32631 , RIdee3798_1052, \9536 );
and \U$23558 ( \32632 , RIdee15d8_1028, \9538 );
and \U$23559 ( \32633 , RIdedf580_1005, \9540 );
and \U$23560 ( \32634 , RIfcb3048_7059, \9542 );
and \U$23561 ( \32635 , RIfc72ae8_6327, \9544 );
and \U$23562 ( \32636 , RIfca3d00_6886, \9546 );
and \U$23563 ( \32637 , RIfcb6450_7096, \9548 );
and \U$23564 ( \32638 , RIdeda558_948, \9550 );
and \U$23565 ( \32639 , RIded7f60_921, \9552 );
and \U$23566 ( \32640 , RIfea3068_8199, \9554 );
and \U$23567 ( \32641 , RIded3a78_872, \9556 );
and \U$23568 ( \32642 , RIded1750_847, \9558 );
and \U$23569 ( \32643 , RIdecea50_815, \9560 );
and \U$23570 ( \32644 , RIdecbd50_783, \9562 );
and \U$23571 ( \32645 , RIdec9050_751, \9564 );
and \U$23572 ( \32646 , RIdeb5550_527, \9566 );
and \U$23573 ( \32647 , RIde98d38_335, \9568 );
and \U$23574 ( \32648 , RIe16f158_2641, \9570 );
and \U$23575 ( \32649 , RIe15af50_2412, \9572 );
and \U$23576 ( \32650 , RIe144750_2156, \9574 );
and \U$23577 ( \32651 , RIdf39148_2026, \9576 );
and \U$23578 ( \32652 , RIdf2d7a8_1894, \9578 );
and \U$23579 ( \32653 , RIdf1e028_1718, \9580 );
and \U$23580 ( \32654 , RIdf01720_1393, \9582 );
and \U$23581 ( \32655 , RIdee8220_1105, \9584 );
and \U$23582 ( \32656 , RIdedcf88_978, \9586 );
and \U$23583 ( \32657 , RIde7ec80_208, \9588 );
or \U$23584 ( \32658 , \32594 , \32595 , \32596 , \32597 , \32598 , \32599 , \32600 , \32601 , \32602 , \32603 , \32604 , \32605 , \32606 , \32607 , \32608 , \32609 , \32610 , \32611 , \32612 , \32613 , \32614 , \32615 , \32616 , \32617 , \32618 , \32619 , \32620 , \32621 , \32622 , \32623 , \32624 , \32625 , \32626 , \32627 , \32628 , \32629 , \32630 , \32631 , \32632 , \32633 , \32634 , \32635 , \32636 , \32637 , \32638 , \32639 , \32640 , \32641 , \32642 , \32643 , \32644 , \32645 , \32646 , \32647 , \32648 , \32649 , \32650 , \32651 , \32652 , \32653 , \32654 , \32655 , \32656 , \32657 );
or \U$23585 ( \32659 , \32593 , \32658 );
_DC g65d4 ( \32660_nG65d4 , \32659 , \9597 );
and \U$23586 ( \32661 , RIe19e5e8_3179, \9059 );
and \U$23587 ( \32662 , RIe19b8e8_3147, \9061 );
and \U$23588 ( \32663 , RIfca84b8_6937, \9063 );
and \U$23589 ( \32664 , RIe198be8_3115, \9065 );
and \U$23590 ( \32665 , RIfc846f8_6529, \9067 );
and \U$23591 ( \32666 , RIe195ee8_3083, \9069 );
and \U$23592 ( \32667 , RIe1931e8_3051, \9071 );
and \U$23593 ( \32668 , RIe1904e8_3019, \9073 );
and \U$23594 ( \32669 , RIe18aae8_2955, \9075 );
and \U$23595 ( \32670 , RIe187de8_2923, \9077 );
and \U$23596 ( \32671 , RIfce2be0_7602, \9079 );
and \U$23597 ( \32672 , RIe1850e8_2891, \9081 );
and \U$23598 ( \32673 , RIfc8e310_6640, \9083 );
and \U$23599 ( \32674 , RIe1823e8_2859, \9085 );
and \U$23600 ( \32675 , RIe17f6e8_2827, \9087 );
and \U$23601 ( \32676 , RIe17c9e8_2795, \9089 );
and \U$23602 ( \32677 , RIfcd1570_7404, \9091 );
and \U$23603 ( \32678 , RIfccc278_7345, \9093 );
and \U$23604 ( \32679 , RIf1404c8_5191, \9095 );
and \U$23605 ( \32680 , RIfea2d98_8197, \9097 );
and \U$23606 ( \32681 , RIfcc1b20_7226, \9099 );
and \U$23607 ( \32682 , RIfc60398_6117, \9101 );
and \U$23608 ( \32683 , RIee3e5a8_5168, \9103 );
and \U$23609 ( \32684 , RIee3da68_5160, \9105 );
and \U$23610 ( \32685 , RIfc642e0_6162, \9107 );
and \U$23611 ( \32686 , RIfca7f18_6933, \9109 );
and \U$23612 ( \32687 , RIee3a228_5120, \9111 );
and \U$23613 ( \32688 , RIfec6180_8374, \9113 );
and \U$23614 ( \32689 , RIfca9598_6949, \9115 );
and \U$23615 ( \32690 , RIfc5c720_6074, \9117 );
and \U$23616 ( \32691 , RIfc6bea0_6250, \9119 );
and \U$23617 ( \32692 , RIfccaec8_7331, \9121 );
and \U$23618 ( \32693 , RIfc44cd8_5805, \9123 );
and \U$23619 ( \32694 , RIe224940_4706, \9125 );
and \U$23620 ( \32695 , RIfcb6180_7094, \9127 );
and \U$23621 ( \32696 , RIe221c40_4674, \9129 );
and \U$23622 ( \32697 , RIfc55ad8_5997, \9131 );
and \U$23623 ( \32698 , RIe21ef40_4642, \9133 );
and \U$23624 ( \32699 , RIe219540_4578, \9135 );
and \U$23625 ( \32700 , RIe216840_4546, \9137 );
and \U$23626 ( \32701 , RIfc4dc48_5907, \9139 );
and \U$23627 ( \32702 , RIe213b40_4514, \9141 );
and \U$23628 ( \32703 , RIfcdcf10_7536, \9143 );
and \U$23629 ( \32704 , RIe210e40_4482, \9145 );
and \U$23630 ( \32705 , RIfcab1b8_6969, \9147 );
and \U$23631 ( \32706 , RIe20e140_4450, \9149 );
and \U$23632 ( \32707 , RIe20b440_4418, \9151 );
and \U$23633 ( \32708 , RIe208740_4386, \9153 );
and \U$23634 ( \32709 , RIfce3720_7610, \9155 );
and \U$23635 ( \32710 , RIfc64178_6161, \9157 );
and \U$23636 ( \32711 , RIe203178_4325, \9159 );
and \U$23637 ( \32712 , RIe201558_4305, \9161 );
and \U$23638 ( \32713 , RIfcd2ec0_7422, \9163 );
and \U$23639 ( \32714 , RIf164828_5603, \9165 );
and \U$23640 ( \32715 , RIfc7f838_6473, \9167 );
and \U$23641 ( \32716 , RIf162398_5577, \9169 );
and \U$23642 ( \32717 , RIfcc9c80_7318, \9171 );
and \U$23643 ( \32718 , RIfca8bc0_6942, \9173 );
and \U$23644 ( \32719 , RIfea2ac8_8195, \9175 );
and \U$23645 ( \32720 , RIfea2c30_8196, \9177 );
and \U$23646 ( \32721 , RIfc59318_6037, \9179 );
and \U$23647 ( \32722 , RIfc4f160_5922, \9181 );
and \U$23648 ( \32723 , RIf15ac10_5492, \9183 );
and \U$23649 ( \32724 , RIfcebf88_7707, \9185 );
or \U$23650 ( \32725 , \32661 , \32662 , \32663 , \32664 , \32665 , \32666 , \32667 , \32668 , \32669 , \32670 , \32671 , \32672 , \32673 , \32674 , \32675 , \32676 , \32677 , \32678 , \32679 , \32680 , \32681 , \32682 , \32683 , \32684 , \32685 , \32686 , \32687 , \32688 , \32689 , \32690 , \32691 , \32692 , \32693 , \32694 , \32695 , \32696 , \32697 , \32698 , \32699 , \32700 , \32701 , \32702 , \32703 , \32704 , \32705 , \32706 , \32707 , \32708 , \32709 , \32710 , \32711 , \32712 , \32713 , \32714 , \32715 , \32716 , \32717 , \32718 , \32719 , \32720 , \32721 , \32722 , \32723 , \32724 );
and \U$23651 ( \32726 , RIfcbb040_7150, \9188 );
and \U$23652 ( \32727 , RIfca1870_6860, \9190 );
and \U$23653 ( \32728 , RIfc93d10_6704, \9192 );
and \U$23654 ( \32729 , RIe1faeb0_4232, \9194 );
and \U$23655 ( \32730 , RIf1565c0_5442, \9196 );
and \U$23656 ( \32731 , RIf155a80_5434, \9198 );
and \U$23657 ( \32732 , RIfc45c50_5816, \9200 );
and \U$23658 ( \32733 , RIe1f6428_4179, \9202 );
and \U$23659 ( \32734 , RIfccdbc8_7363, \9204 );
and \U$23660 ( \32735 , RIfcccae8_7351, \9206 );
and \U$23661 ( \32736 , RIfca6cd0_6920, \9208 );
and \U$23662 ( \32737 , RIfec6018_8373, \9210 );
and \U$23663 ( \32738 , RIfc64010_6160, \9212 );
and \U$23664 ( \32739 , RIfc434f0_5788, \9214 );
and \U$23665 ( \32740 , RIfc4c028_5887, \9216 );
and \U$23666 ( \32741 , RIe1eee08_4095, \9218 );
and \U$23667 ( \32742 , RIe1ec6a8_4067, \9220 );
and \U$23668 ( \32743 , RIe1e99a8_4035, \9222 );
and \U$23669 ( \32744 , RIe1e6ca8_4003, \9224 );
and \U$23670 ( \32745 , RIe1e3fa8_3971, \9226 );
and \U$23671 ( \32746 , RIe1e12a8_3939, \9228 );
and \U$23672 ( \32747 , RIe1de5a8_3907, \9230 );
and \U$23673 ( \32748 , RIe1db8a8_3875, \9232 );
and \U$23674 ( \32749 , RIe1d8ba8_3843, \9234 );
and \U$23675 ( \32750 , RIe1d31a8_3779, \9236 );
and \U$23676 ( \32751 , RIe1d04a8_3747, \9238 );
and \U$23677 ( \32752 , RIe1cd7a8_3715, \9240 );
and \U$23678 ( \32753 , RIe1caaa8_3683, \9242 );
and \U$23679 ( \32754 , RIe1c7da8_3651, \9244 );
and \U$23680 ( \32755 , RIe1c50a8_3619, \9246 );
and \U$23681 ( \32756 , RIe1c23a8_3587, \9248 );
and \U$23682 ( \32757 , RIe1bf6a8_3555, \9250 );
and \U$23683 ( \32758 , RIfc63908_6155, \9252 );
and \U$23684 ( \32759 , RIfc6bd38_6249, \9254 );
and \U$23685 ( \32760 , RIe1ba0e0_3494, \9256 );
and \U$23686 ( \32761 , RIe1b7f20_3470, \9258 );
and \U$23687 ( \32762 , RIfc66fe0_6194, \9260 );
and \U$23688 ( \32763 , RIfc92ac8_6691, \9262 );
and \U$23689 ( \32764 , RIe1b5d60_3446, \9264 );
and \U$23690 ( \32765 , RIfea2f00_8198, \9266 );
and \U$23691 ( \32766 , RIfc9bfd8_6797, \9268 );
and \U$23692 ( \32767 , RIfc50d80_5942, \9270 );
and \U$23693 ( \32768 , RIe1b31c8_3415, \9272 );
and \U$23694 ( \32769 , RIe1b1878_3397, \9274 );
and \U$23695 ( \32770 , RIfc4df18_5909, \9276 );
and \U$23696 ( \32771 , RIfc9d658_6813, \9278 );
and \U$23697 ( \32772 , RIe1ad0c0_3346, \9280 );
and \U$23698 ( \32773 , RIe1ab8d8_3329, \9282 );
and \U$23699 ( \32774 , RIe1a99e8_3307, \9284 );
and \U$23700 ( \32775 , RIe1a6ce8_3275, \9286 );
and \U$23701 ( \32776 , RIe1a3fe8_3243, \9288 );
and \U$23702 ( \32777 , RIe1a12e8_3211, \9290 );
and \U$23703 ( \32778 , RIe18d7e8_2987, \9292 );
and \U$23704 ( \32779 , RIe179ce8_2763, \9294 );
and \U$23705 ( \32780 , RIe227640_4738, \9296 );
and \U$23706 ( \32781 , RIe21c240_4610, \9298 );
and \U$23707 ( \32782 , RIe205a40_4354, \9300 );
and \U$23708 ( \32783 , RIe1ffaa0_4286, \9302 );
and \U$23709 ( \32784 , RIe1f8e58_4209, \9304 );
and \U$23710 ( \32785 , RIe1f19a0_4126, \9306 );
and \U$23711 ( \32786 , RIe1d5ea8_3811, \9308 );
and \U$23712 ( \32787 , RIe1bc9a8_3523, \9310 );
and \U$23713 ( \32788 , RIe1af820_3374, \9312 );
and \U$23714 ( \32789 , RIe171e58_2673, \9314 );
or \U$23715 ( \32790 , \32726 , \32727 , \32728 , \32729 , \32730 , \32731 , \32732 , \32733 , \32734 , \32735 , \32736 , \32737 , \32738 , \32739 , \32740 , \32741 , \32742 , \32743 , \32744 , \32745 , \32746 , \32747 , \32748 , \32749 , \32750 , \32751 , \32752 , \32753 , \32754 , \32755 , \32756 , \32757 , \32758 , \32759 , \32760 , \32761 , \32762 , \32763 , \32764 , \32765 , \32766 , \32767 , \32768 , \32769 , \32770 , \32771 , \32772 , \32773 , \32774 , \32775 , \32776 , \32777 , \32778 , \32779 , \32780 , \32781 , \32782 , \32783 , \32784 , \32785 , \32786 , \32787 , \32788 , \32789 );
or \U$23716 ( \32791 , \32725 , \32790 );
_DC g65d5 ( \32792_nG65d5 , \32791 , \9323 );
and g65d6 ( \32793_nG65d6 , \32660_nG65d4 , \32792_nG65d5 );
buf \U$23717 ( \32794 , \32793_nG65d6 );
and \U$23718 ( \32795 , \32794 , \10691 );
nor \U$23719 ( \32796 , \32528 , \32795 );
xnor \U$23720 ( \32797 , \32796 , \10980 );
not \U$23721 ( \32798 , \32068 );
_DC g64f1 ( \32799_nG64f1 , \32659 , \9597 );
_DC g6575 ( \32800_nG6575 , \32791 , \9323 );
xor g6576 ( \32801_nG6576 , \32799_nG64f1 , \32800_nG6575 );
buf \U$23722 ( \32802 , \32801_nG6576 );
and \U$23723 ( \32803 , \32066 , \30810 );
not \U$23724 ( \32804 , \32803 );
and \U$23725 ( \32805 , \32802 , \32804 );
and \U$23726 ( \32806 , \32798 , \32805 );
xor \U$23727 ( \32807 , \32797 , \32806 );
and \U$23728 ( \32808 , \32057 , \32061 );
and \U$23729 ( \32809 , \32061 , \32068 );
and \U$23730 ( \32810 , \32057 , \32068 );
or \U$23731 ( \32811 , \32808 , \32809 , \32810 );
xor \U$23732 ( \32812 , \32807 , \32811 );
and \U$23733 ( \32813 , \32155 , \32159 );
and \U$23734 ( \32814 , \32159 , \32164 );
and \U$23735 ( \32815 , \32155 , \32164 );
or \U$23736 ( \32816 , \32813 , \32814 , \32815 );
xor \U$23737 ( \32817 , \32812 , \32816 );
xor \U$23738 ( \32818 , \32527 , \32817 );
xor \U$23739 ( \32819 , \32508 , \32818 );
and \U$23740 ( \32820 , \31787 , \32069 );
and \U$23741 ( \32821 , \32069 , \32084 );
and \U$23742 ( \32822 , \31787 , \32084 );
or \U$23743 ( \32823 , \32820 , \32821 , \32822 );
and \U$23744 ( \32824 , \32136 , \32150 );
and \U$23745 ( \32825 , \32150 , \32165 );
and \U$23746 ( \32826 , \32136 , \32165 );
or \U$23747 ( \32827 , \32824 , \32825 , \32826 );
xor \U$23748 ( \32828 , \32823 , \32827 );
and \U$23749 ( \32829 , \22090 , \18090 );
and \U$23750 ( \32830 , \22556 , \17655 );
nor \U$23751 ( \32831 , \32829 , \32830 );
xnor \U$23752 ( \32832 , \32831 , \18046 );
and \U$23753 ( \32833 , \12448 , \29070 );
and \U$23754 ( \32834 , \12769 , \28526 );
nor \U$23755 ( \32835 , \32833 , \32834 );
xnor \U$23756 ( \32836 , \32835 , \29076 );
xor \U$23757 ( \32837 , \32832 , \32836 );
and \U$23758 ( \32838 , \11270 , \30823 );
and \U$23759 ( \32839 , \11586 , \30246 );
nor \U$23760 ( \32840 , \32838 , \32839 );
xnor \U$23761 ( \32841 , \32840 , \30813 );
xor \U$23762 ( \32842 , \32837 , \32841 );
and \U$23763 ( \32843 , \30268 , \11574 );
and \U$23764 ( \32844 , \30802 , \11278 );
nor \U$23765 ( \32845 , \32843 , \32844 );
xnor \U$23766 ( \32846 , \32845 , \11580 );
and \U$23767 ( \32847 , \26829 , \14054 );
and \U$23768 ( \32848 , \27313 , \13692 );
nor \U$23769 ( \32849 , \32847 , \32848 );
xnor \U$23770 ( \32850 , \32849 , \14035 );
xor \U$23771 ( \32851 , \32846 , \32850 );
xor \U$23772 ( \32852 , \32802 , \32066 );
not \U$23773 ( \32853 , \32067 );
and \U$23774 ( \32854 , \32852 , \32853 );
and \U$23775 ( \32855 , \10687 , \32854 );
and \U$23776 ( \32856 , \10988 , \32067 );
nor \U$23777 ( \32857 , \32855 , \32856 );
xnor \U$23778 ( \32858 , \32857 , \32805 );
xor \U$23779 ( \32859 , \32851 , \32858 );
xor \U$23780 ( \32860 , \32842 , \32859 );
and \U$23781 ( \32861 , \25272 , \15336 );
and \U$23782 ( \32862 , \25815 , \14963 );
nor \U$23783 ( \32863 , \32861 , \32862 );
xnor \U$23784 ( \32864 , \32863 , \15342 );
and \U$23785 ( \32865 , \20544 , \19534 );
and \U$23786 ( \32866 , \21033 , \19045 );
nor \U$23787 ( \32867 , \32865 , \32866 );
xnor \U$23788 ( \32868 , \32867 , \19540 );
xor \U$23789 ( \32869 , \32864 , \32868 );
and \U$23790 ( \32870 , \19032 , \21005 );
and \U$23791 ( \32871 , \19558 , \20557 );
nor \U$23792 ( \32872 , \32870 , \32871 );
xnor \U$23793 ( \32873 , \32872 , \21011 );
xor \U$23794 ( \32874 , \32869 , \32873 );
xor \U$23795 ( \32875 , \32860 , \32874 );
xor \U$23796 ( \32876 , \32828 , \32875 );
xor \U$23797 ( \32877 , \32819 , \32876 );
xor \U$23798 ( \32878 , \32504 , \32877 );
and \U$23799 ( \32879 , \31764 , \32086 );
and \U$23800 ( \32880 , \32086 , \32168 );
and \U$23801 ( \32881 , \31764 , \32168 );
or \U$23802 ( \32882 , \32879 , \32880 , \32881 );
xor \U$23803 ( \32883 , \32878 , \32882 );
and \U$23804 ( \32884 , \32169 , \32173 );
and \U$23805 ( \32885 , \32174 , \32177 );
or \U$23806 ( \32886 , \32884 , \32885 );
xor \U$23807 ( \32887 , \32883 , \32886 );
buf g9bb1 ( \32888_nG9bb1 , \32887 );
and \U$23808 ( \32889 , \10704 , \32888_nG9bb1 );
or \U$23809 ( \32890 , \32455 , \32889 );
xor \U$23810 ( \32891 , \10703 , \32890 );
buf \U$23811 ( \32892 , \32891 );
buf \U$23813 ( \32893 , \32892 );
xor \U$23814 ( \32894 , \32454 , \32893 );
buf \U$23815 ( \32895 , \32894 );
xor \U$23816 ( \32896 , \32442 , \32895 );
and \U$23817 ( \32897 , \31712 , \31758 );
and \U$23818 ( \32898 , \31712 , \32184 );
and \U$23819 ( \32899 , \31758 , \32184 );
or \U$23820 ( \32900 , \32897 , \32898 , \32899 );
buf \U$23821 ( \32901 , \32900 );
xor \U$23822 ( \32902 , \32896 , \32901 );
buf \U$23823 ( \32903 , \32902 );
xor \U$23824 ( \32904 , \32384 , \32903 );
xor \U$23825 ( \32905 , \32267 , \32904 );
and \U$23826 ( \32906 , \31653 , \32188 );
and \U$23827 ( \32907 , \31653 , \32258 );
and \U$23828 ( \32908 , \32188 , \32258 );
or \U$23829 ( \32909 , \32906 , \32907 , \32908 );
and \U$23830 ( \32910 , \32905 , \32909 );
and \U$23831 ( \32911 , \32262 , \32266 );
and \U$23832 ( \32912 , \32262 , \32904 );
and \U$23833 ( \32913 , \32266 , \32904 );
or \U$23834 ( \32914 , \32911 , \32912 , \32913 );
xor \U$23835 ( \32915 , \32910 , \32914 );
xor \U$23840 ( \32916 , 1'b0 , \31627_nG43fa );
not \U$23841 ( \32917 , \32916 );
and \U$23845 ( \32918 , \32916 , \10694_nG9c0e );
or \U$23846 ( \32919 , 1'b0 , \32918 );
xor \U$23847 ( \32920 , 1'b0 , \32919 );
xor \U$23848 ( \32921 , 1'b0 , \32920 );
buf \U$23849 ( \32922 , \32921 );
buf \U$23850 ( \32923 , \32922 );
xor \U$23851 ( \32924 , \32915 , \32923 );
and \U$23852 ( \32925 , \32378 , \32383 );
and \U$23853 ( \32926 , \32378 , \32903 );
and \U$23854 ( \32927 , \32383 , \32903 );
or \U$23855 ( \32928 , \32925 , \32926 , \32927 );
and \U$23856 ( \32929 , \32924 , \32928 );
and \U$23857 ( \32930 , \32342 , \32362 );
and \U$23858 ( \32931 , \32342 , \32368 );
and \U$23859 ( \32932 , \32362 , \32368 );
or \U$23860 ( \32933 , \32930 , \32931 , \32932 );
buf \U$23861 ( \32934 , \32933 );
and \U$23862 ( \32935 , \32389 , \32406 );
and \U$23863 ( \32936 , \32389 , \32413 );
and \U$23864 ( \32937 , \32406 , \32413 );
or \U$23865 ( \32938 , \32935 , \32936 , \32937 );
buf \U$23866 ( \32939 , \32938 );
and \U$23867 ( \32940 , \32280 , \32286 );
buf \U$23868 ( \32941 , \32940 );
and \U$23869 ( \32942 , \28118 , \12801_nG9bff );
and \U$23870 ( \32943 , \28115 , \13705_nG9bfc );
or \U$23871 ( \32944 , \32942 , \32943 );
xor \U$23872 ( \32945 , \28114 , \32944 );
buf \U$23873 ( \32946 , \32945 );
buf \U$23875 ( \32947 , \32946 );
xor \U$23876 ( \32948 , \32941 , \32947 );
and \U$23877 ( \32949 , \26431 , \14070_nG9bf9 );
and \U$23878 ( \32950 , \26428 , \14984_nG9bf6 );
or \U$23879 ( \32951 , \32949 , \32950 );
xor \U$23880 ( \32952 , \26427 , \32951 );
buf \U$23881 ( \32953 , \32952 );
buf \U$23883 ( \32954 , \32953 );
xor \U$23884 ( \32955 , \32948 , \32954 );
buf \U$23885 ( \32956 , \32955 );
and \U$23886 ( \32957 , \23201 , \16680_nG9bed );
and \U$23887 ( \32958 , \23198 , \17665_nG9bea );
or \U$23888 ( \32959 , \32957 , \32958 );
xor \U$23889 ( \32960 , \23197 , \32959 );
buf \U$23890 ( \32961 , \32960 );
buf \U$23892 ( \32962 , \32961 );
xor \U$23893 ( \32963 , \32956 , \32962 );
and \U$23894 ( \32964 , \21658 , \18107_nG9be7 );
and \U$23895 ( \32965 , \21655 , \19091_nG9be4 );
or \U$23896 ( \32966 , \32964 , \32965 );
xor \U$23897 ( \32967 , \21654 , \32966 );
buf \U$23898 ( \32968 , \32967 );
buf \U$23900 ( \32969 , \32968 );
xor \U$23901 ( \32970 , \32963 , \32969 );
buf \U$23902 ( \32971 , \32970 );
xor \U$23903 ( \32972 , \32939 , \32971 );
and \U$23904 ( \32973 , \15940 , \24226_nG9bcf );
and \U$23905 ( \32974 , \15937 , \25298_nG9bcc );
or \U$23906 ( \32975 , \32973 , \32974 );
xor \U$23907 ( \32976 , \15936 , \32975 );
buf \U$23908 ( \32977 , \32976 );
buf \U$23910 ( \32978 , \32977 );
xor \U$23911 ( \32979 , \32972 , \32978 );
buf \U$23912 ( \32980 , \32979 );
and \U$23913 ( \32981 , \32277 , \32303 );
and \U$23914 ( \32982 , \32277 , \32310 );
and \U$23915 ( \32983 , \32303 , \32310 );
or \U$23916 ( \32984 , \32981 , \32982 , \32983 );
buf \U$23917 ( \32985 , \32984 );
and \U$23918 ( \32986 , \32288 , \32294 );
and \U$23919 ( \32987 , \32288 , \32301 );
and \U$23920 ( \32988 , \32294 , \32301 );
or \U$23921 ( \32989 , \32986 , \32987 , \32988 );
buf \U$23922 ( \32990 , \32989 );
and \U$23923 ( \32991 , \31636 , \10995_nG9c0b );
and \U$23924 ( \32992 , \31633 , \11283_nG9c08 );
or \U$23925 ( \32993 , \32991 , \32992 );
xor \U$23926 ( \32994 , \31632 , \32993 );
buf \U$23927 ( \32995 , \32994 );
buf \U$23929 ( \32996 , \32995 );
and \U$23930 ( \32997 , \29853 , \11598_nG9c05 );
and \U$23931 ( \32998 , \29850 , \12470_nG9c02 );
or \U$23932 ( \32999 , \32997 , \32998 );
xor \U$23933 ( \33000 , \29849 , \32999 );
buf \U$23934 ( \33001 , \33000 );
buf \U$23936 ( \33002 , \33001 );
xor \U$23937 ( \33003 , \32996 , \33002 );
buf \U$23938 ( \33004 , \33003 );
xor \U$23939 ( \33005 , \32990 , \33004 );
and \U$23940 ( \33006 , \24792 , \15373_nG9bf3 );
and \U$23941 ( \33007 , \24789 , \16315_nG9bf0 );
or \U$23942 ( \33008 , \33006 , \33007 );
xor \U$23943 ( \33009 , \24788 , \33008 );
buf \U$23944 ( \33010 , \33009 );
buf \U$23946 ( \33011 , \33010 );
xor \U$23947 ( \33012 , \33005 , \33011 );
buf \U$23948 ( \33013 , \33012 );
xor \U$23949 ( \33014 , \32985 , \33013 );
and \U$23950 ( \33015 , \17297 , \22629_nG9bd5 );
and \U$23951 ( \33016 , \17294 , \23696_nG9bd2 );
or \U$23952 ( \33017 , \33015 , \33016 );
xor \U$23953 ( \33018 , \17293 , \33017 );
buf \U$23954 ( \33019 , \33018 );
buf \U$23956 ( \33020 , \33019 );
xor \U$23957 ( \33021 , \33014 , \33020 );
buf \U$23958 ( \33022 , \33021 );
xor \U$23959 ( \33023 , \32980 , \33022 );
and \U$23960 ( \33024 , \10707 , \32888_nG9bb1 );
and \U$23961 ( \33025 , \32459 , \32503 );
and \U$23962 ( \33026 , \32503 , \32877 );
and \U$23963 ( \33027 , \32459 , \32877 );
or \U$23964 ( \33028 , \33025 , \33026 , \33027 );
and \U$23965 ( \33029 , \32463 , \32467 );
and \U$23966 ( \33030 , \32467 , \32502 );
and \U$23967 ( \33031 , \32463 , \32502 );
or \U$23968 ( \33032 , \33029 , \33030 , \33031 );
and \U$23969 ( \33033 , \32508 , \32818 );
and \U$23970 ( \33034 , \32818 , \32876 );
and \U$23971 ( \33035 , \32508 , \32876 );
or \U$23972 ( \33036 , \33033 , \33034 , \33035 );
xor \U$23973 ( \33037 , \33032 , \33036 );
and \U$23974 ( \33038 , \32807 , \32811 );
and \U$23975 ( \33039 , \32811 , \32816 );
and \U$23976 ( \33040 , \32807 , \32816 );
or \U$23977 ( \33041 , \33038 , \33039 , \33040 );
and \U$23978 ( \33042 , \32842 , \32859 );
and \U$23979 ( \33043 , \32859 , \32874 );
and \U$23980 ( \33044 , \32842 , \32874 );
or \U$23981 ( \33045 , \33042 , \33043 , \33044 );
xor \U$23982 ( \33046 , \33041 , \33045 );
and \U$23983 ( \33047 , \32832 , \32836 );
and \U$23984 ( \33048 , \32836 , \32841 );
and \U$23985 ( \33049 , \32832 , \32841 );
or \U$23986 ( \33050 , \33047 , \33048 , \33049 );
and \U$23987 ( \33051 , \32476 , \32480 );
and \U$23988 ( \33052 , \32480 , \32485 );
and \U$23989 ( \33053 , \32476 , \32485 );
or \U$23990 ( \33054 , \33051 , \33052 , \33053 );
xor \U$23991 ( \33055 , \33050 , \33054 );
and \U$23992 ( \33056 , \32794 , \10983 );
not \U$23993 ( \33057 , \33056 );
xnor \U$23994 ( \33058 , \33057 , \10980 );
and \U$23995 ( \33059 , \30802 , \11574 );
and \U$23996 ( \33060 , \32054 , \11278 );
nor \U$23997 ( \33061 , \33059 , \33060 );
xnor \U$23998 ( \33062 , \33061 , \11580 );
xor \U$23999 ( \33063 , \33058 , \33062 );
and \U$24000 ( \33064 , \10687 , \32802 );
xor \U$24001 ( \33065 , \33063 , \33064 );
xor \U$24002 ( \33066 , \33055 , \33065 );
xor \U$24003 ( \33067 , \33046 , \33066 );
and \U$24004 ( \33068 , \32472 , \32486 );
and \U$24005 ( \33069 , \32486 , \32501 );
and \U$24006 ( \33070 , \32472 , \32501 );
or \U$24007 ( \33071 , \33068 , \33069 , \33070 );
and \U$24008 ( \33072 , \32846 , \32850 );
and \U$24009 ( \33073 , \32850 , \32858 );
and \U$24010 ( \33074 , \32846 , \32858 );
or \U$24011 ( \33075 , \33072 , \33073 , \33074 );
and \U$24012 ( \33076 , \32864 , \32868 );
and \U$24013 ( \33077 , \32868 , \32873 );
and \U$24014 ( \33078 , \32864 , \32873 );
or \U$24015 ( \33079 , \33076 , \33077 , \33078 );
xor \U$24016 ( \33080 , \33075 , \33079 );
and \U$24017 ( \33081 , \32491 , \32495 );
and \U$24018 ( \33082 , \32495 , \32500 );
and \U$24019 ( \33083 , \32491 , \32500 );
or \U$24020 ( \33084 , \33081 , \33082 , \33083 );
xor \U$24021 ( \33085 , \33080 , \33084 );
xor \U$24022 ( \33086 , \33071 , \33085 );
and \U$24023 ( \33087 , \25815 , \15336 );
and \U$24024 ( \33088 , \26829 , \14963 );
nor \U$24025 ( \33089 , \33087 , \33088 );
xnor \U$24026 ( \33090 , \33089 , \15342 );
and \U$24027 ( \33091 , \19558 , \21005 );
and \U$24028 ( \33092 , \20544 , \20557 );
nor \U$24029 ( \33093 , \33091 , \33092 );
xnor \U$24030 ( \33094 , \33093 , \21011 );
xor \U$24031 ( \33095 , \33090 , \33094 );
and \U$24032 ( \33096 , \18035 , \22542 );
and \U$24033 ( \33097 , \19032 , \22103 );
nor \U$24034 ( \33098 , \33096 , \33097 );
xnor \U$24035 ( \33099 , \33098 , \22548 );
xor \U$24036 ( \33100 , \33095 , \33099 );
and \U$24037 ( \33101 , \29084 , \12790 );
and \U$24038 ( \33102 , \30268 , \12461 );
nor \U$24039 ( \33103 , \33101 , \33102 );
xnor \U$24040 ( \33104 , \33103 , \12780 );
and \U$24041 ( \33105 , \24199 , \16635 );
and \U$24042 ( \33106 , \25272 , \16301 );
nor \U$24043 ( \33107 , \33105 , \33106 );
xnor \U$24044 ( \33108 , \33107 , \16625 );
xor \U$24045 ( \33109 , \33104 , \33108 );
and \U$24046 ( \33110 , \16655 , \24138 );
and \U$24047 ( \33111 , \17627 , \23630 );
nor \U$24048 ( \33112 , \33110 , \33111 );
xnor \U$24049 ( \33113 , \33112 , \24144 );
xor \U$24050 ( \33114 , \33109 , \33113 );
xor \U$24051 ( \33115 , \33100 , \33114 );
and \U$24052 ( \33116 , \22556 , \18090 );
and \U$24053 ( \33117 , \23617 , \17655 );
nor \U$24054 ( \33118 , \33116 , \33117 );
xnor \U$24055 ( \33119 , \33118 , \18046 );
and \U$24056 ( \33120 , \15321 , \25826 );
and \U$24057 ( \33121 , \16267 , \25264 );
nor \U$24058 ( \33122 , \33120 , \33121 );
xnor \U$24059 ( \33123 , \33122 , \25773 );
xor \U$24060 ( \33124 , \33119 , \33123 );
and \U$24061 ( \33125 , \14024 , \27397 );
and \U$24062 ( \33126 , \14950 , \26807 );
nor \U$24063 ( \33127 , \33125 , \33126 );
xnor \U$24064 ( \33128 , \33127 , \27295 );
xor \U$24065 ( \33129 , \33124 , \33128 );
xor \U$24066 ( \33130 , \33115 , \33129 );
xor \U$24067 ( \33131 , \33086 , \33130 );
xor \U$24068 ( \33132 , \33067 , \33131 );
and \U$24069 ( \33133 , \32512 , \32526 );
and \U$24070 ( \33134 , \32526 , \32817 );
and \U$24071 ( \33135 , \32512 , \32817 );
or \U$24072 ( \33136 , \33133 , \33134 , \33135 );
and \U$24073 ( \33137 , \32823 , \32827 );
and \U$24074 ( \33138 , \32827 , \32875 );
and \U$24075 ( \33139 , \32823 , \32875 );
or \U$24076 ( \33140 , \33137 , \33138 , \33139 );
xor \U$24077 ( \33141 , \33136 , \33140 );
and \U$24078 ( \33142 , \32516 , \32520 );
and \U$24079 ( \33143 , \32520 , \32525 );
and \U$24080 ( \33144 , \32516 , \32525 );
or \U$24081 ( \33145 , \33142 , \33143 , \33144 );
and \U$24082 ( \33146 , \27313 , \14054 );
and \U$24083 ( \33147 , \28534 , \13692 );
nor \U$24084 ( \33148 , \33146 , \33147 );
xnor \U$24085 ( \33149 , \33148 , \14035 );
and \U$24086 ( \33150 , \21033 , \19534 );
and \U$24087 ( \33151 , \22090 , \19045 );
nor \U$24088 ( \33152 , \33150 , \33151 );
xnor \U$24089 ( \33153 , \33152 , \19540 );
xor \U$24090 ( \33154 , \33149 , \33153 );
and \U$24091 ( \33155 , \10988 , \32854 );
and \U$24092 ( \33156 , \11270 , \32067 );
nor \U$24093 ( \33157 , \33155 , \33156 );
xnor \U$24094 ( \33158 , \33157 , \32805 );
xor \U$24095 ( \33159 , \33154 , \33158 );
xor \U$24096 ( \33160 , \33145 , \33159 );
and \U$24097 ( \33161 , \32797 , \32806 );
and \U$24098 ( \33162 , \12769 , \29070 );
and \U$24099 ( \33163 , \13679 , \28526 );
nor \U$24100 ( \33164 , \33162 , \33163 );
xnor \U$24101 ( \33165 , \33164 , \29076 );
xor \U$24102 ( \33166 , \33161 , \33165 );
and \U$24103 ( \33167 , \11586 , \30823 );
and \U$24104 ( \33168 , \12448 , \30246 );
nor \U$24105 ( \33169 , \33167 , \33168 );
xnor \U$24106 ( \33170 , \33169 , \30813 );
xor \U$24107 ( \33171 , \33166 , \33170 );
xor \U$24108 ( \33172 , \33160 , \33171 );
xor \U$24109 ( \33173 , \33141 , \33172 );
xor \U$24110 ( \33174 , \33132 , \33173 );
xor \U$24111 ( \33175 , \33037 , \33174 );
xor \U$24112 ( \33176 , \33028 , \33175 );
and \U$24113 ( \33177 , \32878 , \32882 );
and \U$24114 ( \33178 , \32883 , \32886 );
or \U$24115 ( \33179 , \33177 , \33178 );
xor \U$24116 ( \33180 , \33176 , \33179 );
buf g9bae ( \33181_nG9bae , \33180 );
and \U$24117 ( \33182 , \10704 , \33181_nG9bae );
or \U$24118 ( \33183 , \33024 , \33182 );
xor \U$24119 ( \33184 , \10703 , \33183 );
buf \U$24120 ( \33185 , \33184 );
buf \U$24122 ( \33186 , \33185 );
xor \U$24123 ( \33187 , \33023 , \33186 );
buf \U$24124 ( \33188 , \33187 );
xor \U$24125 ( \33189 , \32934 , \33188 );
and \U$24126 ( \33190 , \32429 , \32434 );
and \U$24127 ( \33191 , \32429 , \32440 );
and \U$24128 ( \33192 , \32434 , \32440 );
or \U$24129 ( \33193 , \33190 , \33191 , \33192 );
buf \U$24130 ( \33194 , \33193 );
xor \U$24131 ( \33195 , \33189 , \33194 );
buf \U$24132 ( \33196 , \33195 );
and \U$24133 ( \33197 , \32272 , \32370 );
and \U$24134 ( \33198 , \32272 , \32376 );
and \U$24135 ( \33199 , \32370 , \32376 );
or \U$24136 ( \33200 , \33197 , \33198 , \33199 );
buf \U$24137 ( \33201 , \33200 );
xor \U$24138 ( \33202 , \33196 , \33201 );
and \U$24139 ( \33203 , \32442 , \32895 );
and \U$24140 ( \33204 , \32442 , \32901 );
and \U$24141 ( \33205 , \32895 , \32901 );
or \U$24142 ( \33206 , \33203 , \33204 , \33205 );
buf \U$24143 ( \33207 , \33206 );
and \U$24144 ( \33208 , \32327 , \32333 );
and \U$24145 ( \33209 , \32327 , \32340 );
and \U$24146 ( \33210 , \32333 , \32340 );
or \U$24147 ( \33211 , \33208 , \33209 , \33210 );
buf \U$24148 ( \33212 , \33211 );
and \U$24149 ( \33213 , \32447 , \32453 );
and \U$24150 ( \33214 , \32447 , \32893 );
and \U$24151 ( \33215 , \32453 , \32893 );
or \U$24152 ( \33216 , \33213 , \33214 , \33215 );
buf \U$24153 ( \33217 , \33216 );
xor \U$24154 ( \33218 , \33212 , \33217 );
and \U$24155 ( \33219 , \13370 , \27416_nG9bc3 );
and \U$24156 ( \33220 , \13367 , \28602_nG9bc0 );
or \U$24157 ( \33221 , \33219 , \33220 );
xor \U$24158 ( \33222 , \13366 , \33221 );
buf \U$24159 ( \33223 , \33222 );
buf \U$24161 ( \33224 , \33223 );
and \U$24162 ( \33225 , \12157 , \29179_nG9bbd );
and \U$24163 ( \33226 , \12154 , \30366_nG9bba );
or \U$24164 ( \33227 , \33225 , \33226 );
xor \U$24165 ( \33228 , \12153 , \33227 );
buf \U$24166 ( \33229 , \33228 );
buf \U$24168 ( \33230 , \33229 );
xor \U$24169 ( \33231 , \33224 , \33230 );
and \U$24170 ( \33232 , \10421 , \30940_nG9bb7 );
and \U$24171 ( \33233 , \10418 , \32179_nG9bb4 );
or \U$24172 ( \33234 , \33232 , \33233 );
xor \U$24173 ( \33235 , \10417 , \33234 );
buf \U$24174 ( \33236 , \33235 );
buf \U$24176 ( \33237 , \33236 );
xor \U$24177 ( \33238 , \33231 , \33237 );
buf \U$24178 ( \33239 , \33238 );
xor \U$24179 ( \33240 , \33218 , \33239 );
buf \U$24180 ( \33241 , \33240 );
xor \U$24181 ( \33242 , \33207 , \33241 );
and \U$24182 ( \33243 , \32415 , \32420 );
and \U$24183 ( \33244 , \32415 , \32427 );
and \U$24184 ( \33245 , \32420 , \32427 );
or \U$24185 ( \33246 , \33243 , \33244 , \33245 );
buf \U$24186 ( \33247 , \33246 );
and \U$24187 ( \33248 , \32312 , \32318 );
and \U$24188 ( \33249 , \32312 , \32325 );
and \U$24189 ( \33250 , \32318 , \32325 );
or \U$24190 ( \33251 , \33248 , \33249 , \33250 );
buf \U$24191 ( \33252 , \33251 );
and \U$24192 ( \33253 , \32391 , \32397 );
and \U$24193 ( \33254 , \32391 , \32404 );
and \U$24194 ( \33255 , \32397 , \32404 );
or \U$24195 ( \33256 , \33253 , \33254 , \33255 );
buf \U$24196 ( \33257 , \33256 );
and \U$24197 ( \33258 , \20155 , \19586_nG9be1 );
and \U$24198 ( \33259 , \20152 , \20608_nG9bde );
or \U$24199 ( \33260 , \33258 , \33259 );
xor \U$24200 ( \33261 , \20151 , \33260 );
buf \U$24201 ( \33262 , \33261 );
buf \U$24203 ( \33263 , \33262 );
xor \U$24204 ( \33264 , \33257 , \33263 );
and \U$24205 ( \33265 , \18702 , \21086_nG9bdb );
and \U$24206 ( \33266 , \18699 , \22129_nG9bd8 );
or \U$24207 ( \33267 , \33265 , \33266 );
xor \U$24208 ( \33268 , \18698 , \33267 );
buf \U$24209 ( \33269 , \33268 );
buf \U$24211 ( \33270 , \33269 );
xor \U$24212 ( \33271 , \33264 , \33270 );
buf \U$24213 ( \33272 , \33271 );
xor \U$24214 ( \33273 , \33252 , \33272 );
and \U$24215 ( \33274 , \14631 , \25860_nG9bc9 );
and \U$24216 ( \33275 , \14628 , \26887_nG9bc6 );
or \U$24217 ( \33276 , \33274 , \33275 );
xor \U$24218 ( \33277 , \14627 , \33276 );
buf \U$24219 ( \33278 , \33277 );
buf \U$24221 ( \33279 , \33278 );
xor \U$24222 ( \33280 , \33273 , \33279 );
buf \U$24223 ( \33281 , \33280 );
xor \U$24224 ( \33282 , \33247 , \33281 );
and \U$24225 ( \33283 , \32347 , \32353 );
and \U$24226 ( \33284 , \32347 , \32360 );
and \U$24227 ( \33285 , \32353 , \32360 );
or \U$24228 ( \33286 , \33283 , \33284 , \33285 );
buf \U$24229 ( \33287 , \33286 );
xor \U$24230 ( \33288 , \33282 , \33287 );
buf \U$24231 ( \33289 , \33288 );
xor \U$24232 ( \33290 , \33242 , \33289 );
buf \U$24233 ( \33291 , \33290 );
xor \U$24234 ( \33292 , \33202 , \33291 );
and \U$24235 ( \33293 , \32924 , \33292 );
and \U$24236 ( \33294 , \32928 , \33292 );
or \U$24237 ( \33295 , \32929 , \33293 , \33294 );
and \U$24238 ( \33296 , \32910 , \32914 );
and \U$24239 ( \33297 , \32910 , \32923 );
and \U$24240 ( \33298 , \32914 , \32923 );
or \U$24241 ( \33299 , \33296 , \33297 , \33298 );
xor \U$24242 ( \33300 , \33295 , \33299 );
xor \U$24246 ( \33301 , \33300 , 1'b0 );
and \U$24247 ( \33302 , \33207 , \33241 );
and \U$24248 ( \33303 , \33207 , \33289 );
and \U$24249 ( \33304 , \33241 , \33289 );
or \U$24250 ( \33305 , \33302 , \33303 , \33304 );
buf \U$24251 ( \33306 , \33305 );
and \U$24252 ( \33307 , \32990 , \33004 );
and \U$24253 ( \33308 , \32990 , \33011 );
and \U$24254 ( \33309 , \33004 , \33011 );
or \U$24255 ( \33310 , \33307 , \33308 , \33309 );
buf \U$24256 ( \33311 , \33310 );
and \U$24257 ( \33312 , \32996 , \33002 );
buf \U$24258 ( \33313 , \33312 );
and \U$24259 ( \33314 , \28118 , \13705_nG9bfc );
and \U$24260 ( \33315 , \28115 , \14070_nG9bf9 );
or \U$24261 ( \33316 , \33314 , \33315 );
xor \U$24262 ( \33317 , \28114 , \33316 );
buf \U$24263 ( \33318 , \33317 );
buf \U$24265 ( \33319 , \33318 );
xor \U$24266 ( \33320 , \33313 , \33319 );
and \U$24267 ( \33321 , \26431 , \14984_nG9bf6 );
and \U$24268 ( \33322 , \26428 , \15373_nG9bf3 );
or \U$24269 ( \33323 , \33321 , \33322 );
xor \U$24270 ( \33324 , \26427 , \33323 );
buf \U$24271 ( \33325 , \33324 );
buf \U$24273 ( \33326 , \33325 );
xor \U$24274 ( \33327 , \33320 , \33326 );
buf \U$24275 ( \33328 , \33327 );
xor \U$24276 ( \33329 , \33311 , \33328 );
and \U$24277 ( \33330 , \23201 , \17665_nG9bea );
and \U$24278 ( \33331 , \23198 , \18107_nG9be7 );
or \U$24279 ( \33332 , \33330 , \33331 );
xor \U$24280 ( \33333 , \23197 , \33332 );
buf \U$24281 ( \33334 , \33333 );
buf \U$24283 ( \33335 , \33334 );
xor \U$24284 ( \33336 , \33329 , \33335 );
buf \U$24285 ( \33337 , \33336 );
and \U$24286 ( \33338 , \32941 , \32947 );
and \U$24287 ( \33339 , \32941 , \32954 );
and \U$24288 ( \33340 , \32947 , \32954 );
or \U$24289 ( \33341 , \33338 , \33339 , \33340 );
buf \U$24290 ( \33342 , \33341 );
and \U$24292 ( \33343 , \32916 , \10995_nG9c0b );
or \U$24293 ( \33344 , 1'b0 , \33343 );
xor \U$24294 ( \33345 , 1'b0 , \33344 );
buf \U$24295 ( \33346 , \33345 );
buf \U$24297 ( \33347 , \33346 );
and \U$24298 ( \33348 , \31636 , \11283_nG9c08 );
and \U$24299 ( \33349 , \31633 , \11598_nG9c05 );
or \U$24300 ( \33350 , \33348 , \33349 );
xor \U$24301 ( \33351 , \31632 , \33350 );
buf \U$24302 ( \33352 , \33351 );
buf \U$24304 ( \33353 , \33352 );
xor \U$24305 ( \33354 , \33347 , \33353 );
and \U$24306 ( \33355 , \29853 , \12470_nG9c02 );
and \U$24307 ( \33356 , \29850 , \12801_nG9bff );
or \U$24308 ( \33357 , \33355 , \33356 );
xor \U$24309 ( \33358 , \29849 , \33357 );
buf \U$24310 ( \33359 , \33358 );
buf \U$24312 ( \33360 , \33359 );
xor \U$24313 ( \33361 , \33354 , \33360 );
buf \U$24314 ( \33362 , \33361 );
xor \U$24315 ( \33363 , \33342 , \33362 );
and \U$24316 ( \33364 , \24792 , \16315_nG9bf0 );
and \U$24317 ( \33365 , \24789 , \16680_nG9bed );
or \U$24318 ( \33366 , \33364 , \33365 );
xor \U$24319 ( \33367 , \24788 , \33366 );
buf \U$24320 ( \33368 , \33367 );
buf \U$24322 ( \33369 , \33368 );
xor \U$24323 ( \33370 , \33363 , \33369 );
buf \U$24324 ( \33371 , \33370 );
and \U$24325 ( \33372 , \21658 , \19091_nG9be4 );
and \U$24326 ( \33373 , \21655 , \19586_nG9be1 );
or \U$24327 ( \33374 , \33372 , \33373 );
xor \U$24328 ( \33375 , \21654 , \33374 );
buf \U$24329 ( \33376 , \33375 );
buf \U$24331 ( \33377 , \33376 );
xor \U$24332 ( \33378 , \33371 , \33377 );
and \U$24333 ( \33379 , \20155 , \20608_nG9bde );
and \U$24334 ( \33380 , \20152 , \21086_nG9bdb );
or \U$24335 ( \33381 , \33379 , \33380 );
xor \U$24336 ( \33382 , \20151 , \33381 );
buf \U$24337 ( \33383 , \33382 );
buf \U$24339 ( \33384 , \33383 );
xor \U$24340 ( \33385 , \33378 , \33384 );
buf \U$24341 ( \33386 , \33385 );
xor \U$24342 ( \33387 , \33337 , \33386 );
and \U$24343 ( \33388 , \33257 , \33263 );
and \U$24344 ( \33389 , \33257 , \33270 );
and \U$24345 ( \33390 , \33263 , \33270 );
or \U$24346 ( \33391 , \33388 , \33389 , \33390 );
buf \U$24347 ( \33392 , \33391 );
xor \U$24348 ( \33393 , \33387 , \33392 );
buf \U$24349 ( \33394 , \33393 );
and \U$24350 ( \33395 , \33252 , \33272 );
and \U$24351 ( \33396 , \33252 , \33279 );
and \U$24352 ( \33397 , \33272 , \33279 );
or \U$24353 ( \33398 , \33395 , \33396 , \33397 );
buf \U$24354 ( \33399 , \33398 );
xor \U$24355 ( \33400 , \33394 , \33399 );
and \U$24356 ( \33401 , \15940 , \25298_nG9bcc );
and \U$24357 ( \33402 , \15937 , \25860_nG9bc9 );
or \U$24358 ( \33403 , \33401 , \33402 );
xor \U$24359 ( \33404 , \15936 , \33403 );
buf \U$24360 ( \33405 , \33404 );
buf \U$24362 ( \33406 , \33405 );
and \U$24363 ( \33407 , \14631 , \26887_nG9bc6 );
and \U$24364 ( \33408 , \14628 , \27416_nG9bc3 );
or \U$24365 ( \33409 , \33407 , \33408 );
xor \U$24366 ( \33410 , \14627 , \33409 );
buf \U$24367 ( \33411 , \33410 );
buf \U$24369 ( \33412 , \33411 );
xor \U$24370 ( \33413 , \33406 , \33412 );
and \U$24371 ( \33414 , \12157 , \30366_nG9bba );
and \U$24372 ( \33415 , \12154 , \30940_nG9bb7 );
or \U$24373 ( \33416 , \33414 , \33415 );
xor \U$24374 ( \33417 , \12153 , \33416 );
buf \U$24375 ( \33418 , \33417 );
buf \U$24377 ( \33419 , \33418 );
xor \U$24378 ( \33420 , \33413 , \33419 );
buf \U$24379 ( \33421 , \33420 );
xor \U$24380 ( \33422 , \33400 , \33421 );
buf \U$24381 ( \33423 , \33422 );
and \U$24382 ( \33424 , \33247 , \33281 );
and \U$24383 ( \33425 , \33247 , \33287 );
and \U$24384 ( \33426 , \33281 , \33287 );
or \U$24385 ( \33427 , \33424 , \33425 , \33426 );
buf \U$24386 ( \33428 , \33427 );
xor \U$24387 ( \33429 , \33423 , \33428 );
and \U$24388 ( \33430 , \32956 , \32962 );
and \U$24389 ( \33431 , \32956 , \32969 );
and \U$24390 ( \33432 , \32962 , \32969 );
or \U$24391 ( \33433 , \33430 , \33431 , \33432 );
buf \U$24392 ( \33434 , \33433 );
and \U$24393 ( \33435 , \18702 , \22129_nG9bd8 );
and \U$24394 ( \33436 , \18699 , \22629_nG9bd5 );
or \U$24395 ( \33437 , \33435 , \33436 );
xor \U$24396 ( \33438 , \18698 , \33437 );
buf \U$24397 ( \33439 , \33438 );
buf \U$24399 ( \33440 , \33439 );
xor \U$24400 ( \33441 , \33434 , \33440 );
and \U$24401 ( \33442 , \17297 , \23696_nG9bd2 );
and \U$24402 ( \33443 , \17294 , \24226_nG9bcf );
or \U$24403 ( \33444 , \33442 , \33443 );
xor \U$24404 ( \33445 , \17293 , \33444 );
buf \U$24405 ( \33446 , \33445 );
buf \U$24407 ( \33447 , \33446 );
xor \U$24408 ( \33448 , \33441 , \33447 );
buf \U$24409 ( \33449 , \33448 );
and \U$24410 ( \33450 , \32939 , \32971 );
and \U$24411 ( \33451 , \32939 , \32978 );
and \U$24412 ( \33452 , \32971 , \32978 );
or \U$24413 ( \33453 , \33450 , \33451 , \33452 );
buf \U$24414 ( \33454 , \33453 );
xor \U$24415 ( \33455 , \33449 , \33454 );
and \U$24416 ( \33456 , \10707 , \33181_nG9bae );
and \U$24417 ( \33457 , \33067 , \33131 );
and \U$24418 ( \33458 , \33131 , \33173 );
and \U$24419 ( \33459 , \33067 , \33173 );
or \U$24420 ( \33460 , \33457 , \33458 , \33459 );
and \U$24421 ( \33461 , \33041 , \33045 );
and \U$24422 ( \33462 , \33045 , \33066 );
and \U$24423 ( \33463 , \33041 , \33066 );
or \U$24424 ( \33464 , \33461 , \33462 , \33463 );
and \U$24425 ( \33465 , \33161 , \33165 );
and \U$24426 ( \33466 , \33165 , \33170 );
and \U$24427 ( \33467 , \33161 , \33170 );
or \U$24428 ( \33468 , \33465 , \33466 , \33467 );
and \U$24429 ( \33469 , \33075 , \33079 );
and \U$24430 ( \33470 , \33079 , \33084 );
and \U$24431 ( \33471 , \33075 , \33084 );
or \U$24432 ( \33472 , \33469 , \33470 , \33471 );
xor \U$24433 ( \33473 , \33468 , \33472 );
and \U$24434 ( \33474 , \33050 , \33054 );
and \U$24435 ( \33475 , \33054 , \33065 );
and \U$24436 ( \33476 , \33050 , \33065 );
or \U$24437 ( \33477 , \33474 , \33475 , \33476 );
xor \U$24438 ( \33478 , \33473 , \33477 );
xor \U$24439 ( \33479 , \33464 , \33478 );
and \U$24440 ( \33480 , \33100 , \33114 );
and \U$24441 ( \33481 , \33114 , \33129 );
and \U$24442 ( \33482 , \33100 , \33129 );
or \U$24443 ( \33483 , \33480 , \33481 , \33482 );
and \U$24444 ( \33484 , \33090 , \33094 );
and \U$24445 ( \33485 , \33094 , \33099 );
and \U$24446 ( \33486 , \33090 , \33099 );
or \U$24447 ( \33487 , \33484 , \33485 , \33486 );
and \U$24448 ( \33488 , \33119 , \33123 );
and \U$24449 ( \33489 , \33123 , \33128 );
and \U$24450 ( \33490 , \33119 , \33128 );
or \U$24451 ( \33491 , \33488 , \33489 , \33490 );
xor \U$24452 ( \33492 , \33487 , \33491 );
and \U$24453 ( \33493 , \33149 , \33153 );
and \U$24454 ( \33494 , \33153 , \33158 );
and \U$24455 ( \33495 , \33149 , \33158 );
or \U$24456 ( \33496 , \33493 , \33494 , \33495 );
xor \U$24457 ( \33497 , \33492 , \33496 );
xor \U$24458 ( \33498 , \33483 , \33497 );
and \U$24459 ( \33499 , \33058 , \33062 );
and \U$24460 ( \33500 , \33062 , \33064 );
and \U$24461 ( \33501 , \33058 , \33064 );
or \U$24462 ( \33502 , \33499 , \33500 , \33501 );
xor \U$24463 ( \33503 , \33502 , \10980 );
and \U$24464 ( \33504 , \12448 , \30823 );
and \U$24465 ( \33505 , \12769 , \30246 );
nor \U$24466 ( \33506 , \33504 , \33505 );
xnor \U$24467 ( \33507 , \33506 , \30813 );
xor \U$24468 ( \33508 , \33503 , \33507 );
xor \U$24469 ( \33509 , \33498 , \33508 );
xor \U$24470 ( \33510 , \33479 , \33509 );
xor \U$24471 ( \33511 , \33460 , \33510 );
and \U$24472 ( \33512 , \33071 , \33085 );
and \U$24473 ( \33513 , \33085 , \33130 );
and \U$24474 ( \33514 , \33071 , \33130 );
or \U$24475 ( \33515 , \33512 , \33513 , \33514 );
and \U$24476 ( \33516 , \33136 , \33140 );
and \U$24477 ( \33517 , \33140 , \33172 );
and \U$24478 ( \33518 , \33136 , \33172 );
or \U$24479 ( \33519 , \33516 , \33517 , \33518 );
xor \U$24480 ( \33520 , \33515 , \33519 );
and \U$24481 ( \33521 , \33145 , \33159 );
and \U$24482 ( \33522 , \33159 , \33171 );
and \U$24483 ( \33523 , \33145 , \33171 );
or \U$24484 ( \33524 , \33521 , \33522 , \33523 );
and \U$24485 ( \33525 , \33104 , \33108 );
and \U$24486 ( \33526 , \33108 , \33113 );
and \U$24487 ( \33527 , \33104 , \33113 );
or \U$24488 ( \33528 , \33525 , \33526 , \33527 );
and \U$24489 ( \33529 , \22090 , \19534 );
and \U$24490 ( \33530 , \22556 , \19045 );
nor \U$24491 ( \33531 , \33529 , \33530 );
xnor \U$24492 ( \33532 , \33531 , \19540 );
and \U$24493 ( \33533 , \11270 , \32854 );
and \U$24494 ( \33534 , \11586 , \32067 );
nor \U$24495 ( \33535 , \33533 , \33534 );
xnor \U$24496 ( \33536 , \33535 , \32805 );
xor \U$24497 ( \33537 , \33532 , \33536 );
and \U$24498 ( \33538 , \10988 , \32802 );
xor \U$24499 ( \33539 , \33537 , \33538 );
xor \U$24500 ( \33540 , \33528 , \33539 );
and \U$24501 ( \33541 , \23617 , \18090 );
and \U$24502 ( \33542 , \24199 , \17655 );
nor \U$24503 ( \33543 , \33541 , \33542 );
xnor \U$24504 ( \33544 , \33543 , \18046 );
and \U$24505 ( \33545 , \14950 , \27397 );
and \U$24506 ( \33546 , \15321 , \26807 );
nor \U$24507 ( \33547 , \33545 , \33546 );
xnor \U$24508 ( \33548 , \33547 , \27295 );
xor \U$24509 ( \33549 , \33544 , \33548 );
and \U$24510 ( \33550 , \13679 , \29070 );
and \U$24511 ( \33551 , \14024 , \28526 );
nor \U$24512 ( \33552 , \33550 , \33551 );
xnor \U$24513 ( \33553 , \33552 , \29076 );
xor \U$24514 ( \33554 , \33549 , \33553 );
xor \U$24515 ( \33555 , \33540 , \33554 );
xor \U$24516 ( \33556 , \33524 , \33555 );
and \U$24517 ( \33557 , \32054 , \11574 );
and \U$24518 ( \33558 , \32794 , \11278 );
nor \U$24519 ( \33559 , \33557 , \33558 );
xnor \U$24520 ( \33560 , \33559 , \11580 );
and \U$24521 ( \33561 , \28534 , \14054 );
and \U$24522 ( \33562 , \29084 , \13692 );
nor \U$24523 ( \33563 , \33561 , \33562 );
xnor \U$24524 ( \33564 , \33563 , \14035 );
xor \U$24525 ( \33565 , \33560 , \33564 );
and \U$24526 ( \33566 , \20544 , \21005 );
and \U$24527 ( \33567 , \21033 , \20557 );
nor \U$24528 ( \33568 , \33566 , \33567 );
xnor \U$24529 ( \33569 , \33568 , \21011 );
xor \U$24530 ( \33570 , \33565 , \33569 );
and \U$24531 ( \33571 , \26829 , \15336 );
and \U$24532 ( \33572 , \27313 , \14963 );
nor \U$24533 ( \33573 , \33571 , \33572 );
xnor \U$24534 ( \33574 , \33573 , \15342 );
and \U$24535 ( \33575 , \19032 , \22542 );
and \U$24536 ( \33576 , \19558 , \22103 );
nor \U$24537 ( \33577 , \33575 , \33576 );
xnor \U$24538 ( \33578 , \33577 , \22548 );
xor \U$24539 ( \33579 , \33574 , \33578 );
and \U$24540 ( \33580 , \17627 , \24138 );
and \U$24541 ( \33581 , \18035 , \23630 );
nor \U$24542 ( \33582 , \33580 , \33581 );
xnor \U$24543 ( \33583 , \33582 , \24144 );
xor \U$24544 ( \33584 , \33579 , \33583 );
xor \U$24545 ( \33585 , \33570 , \33584 );
and \U$24546 ( \33586 , \30268 , \12790 );
and \U$24547 ( \33587 , \30802 , \12461 );
nor \U$24548 ( \33588 , \33586 , \33587 );
xnor \U$24549 ( \33589 , \33588 , \12780 );
and \U$24550 ( \33590 , \25272 , \16635 );
and \U$24551 ( \33591 , \25815 , \16301 );
nor \U$24552 ( \33592 , \33590 , \33591 );
xnor \U$24553 ( \33593 , \33592 , \16625 );
xor \U$24554 ( \33594 , \33589 , \33593 );
and \U$24555 ( \33595 , \16267 , \25826 );
and \U$24556 ( \33596 , \16655 , \25264 );
nor \U$24557 ( \33597 , \33595 , \33596 );
xnor \U$24558 ( \33598 , \33597 , \25773 );
xor \U$24559 ( \33599 , \33594 , \33598 );
xor \U$24560 ( \33600 , \33585 , \33599 );
xor \U$24561 ( \33601 , \33556 , \33600 );
xor \U$24562 ( \33602 , \33520 , \33601 );
xor \U$24563 ( \33603 , \33511 , \33602 );
and \U$24564 ( \33604 , \33032 , \33036 );
and \U$24565 ( \33605 , \33036 , \33174 );
and \U$24566 ( \33606 , \33032 , \33174 );
or \U$24567 ( \33607 , \33604 , \33605 , \33606 );
xor \U$24568 ( \33608 , \33603 , \33607 );
and \U$24569 ( \33609 , \33028 , \33175 );
and \U$24570 ( \33610 , \33176 , \33179 );
or \U$24571 ( \33611 , \33609 , \33610 );
xor \U$24572 ( \33612 , \33608 , \33611 );
buf g9bab ( \33613_nG9bab , \33612 );
and \U$24573 ( \33614 , \10704 , \33613_nG9bab );
or \U$24574 ( \33615 , \33456 , \33614 );
xor \U$24575 ( \33616 , \10703 , \33615 );
buf \U$24576 ( \33617 , \33616 );
buf \U$24578 ( \33618 , \33617 );
xor \U$24579 ( \33619 , \33455 , \33618 );
buf \U$24580 ( \33620 , \33619 );
xor \U$24581 ( \33621 , \33429 , \33620 );
buf \U$24582 ( \33622 , \33621 );
xor \U$24583 ( \33623 , \33306 , \33622 );
and \U$24584 ( \33624 , \32934 , \33188 );
and \U$24585 ( \33625 , \32934 , \33194 );
and \U$24586 ( \33626 , \33188 , \33194 );
or \U$24587 ( \33627 , \33624 , \33625 , \33626 );
buf \U$24588 ( \33628 , \33627 );
and \U$24589 ( \33629 , \32980 , \33022 );
and \U$24590 ( \33630 , \32980 , \33186 );
and \U$24591 ( \33631 , \33022 , \33186 );
or \U$24592 ( \33632 , \33629 , \33630 , \33631 );
buf \U$24593 ( \33633 , \33632 );
and \U$24594 ( \33634 , \33224 , \33230 );
and \U$24595 ( \33635 , \33224 , \33237 );
and \U$24596 ( \33636 , \33230 , \33237 );
or \U$24597 ( \33637 , \33634 , \33635 , \33636 );
buf \U$24598 ( \33638 , \33637 );
xor \U$24599 ( \33639 , \33633 , \33638 );
and \U$24600 ( \33640 , \32985 , \33013 );
and \U$24601 ( \33641 , \32985 , \33020 );
and \U$24602 ( \33642 , \33013 , \33020 );
or \U$24603 ( \33643 , \33640 , \33641 , \33642 );
buf \U$24604 ( \33644 , \33643 );
and \U$24605 ( \33645 , \13370 , \28602_nG9bc0 );
and \U$24606 ( \33646 , \13367 , \29179_nG9bbd );
or \U$24607 ( \33647 , \33645 , \33646 );
xor \U$24608 ( \33648 , \13366 , \33647 );
buf \U$24609 ( \33649 , \33648 );
buf \U$24611 ( \33650 , \33649 );
xor \U$24612 ( \33651 , \33644 , \33650 );
and \U$24613 ( \33652 , \10421 , \32179_nG9bb4 );
and \U$24614 ( \33653 , \10418 , \32888_nG9bb1 );
or \U$24615 ( \33654 , \33652 , \33653 );
xor \U$24616 ( \33655 , \10417 , \33654 );
buf \U$24617 ( \33656 , \33655 );
buf \U$24619 ( \33657 , \33656 );
xor \U$24620 ( \33658 , \33651 , \33657 );
buf \U$24621 ( \33659 , \33658 );
xor \U$24622 ( \33660 , \33639 , \33659 );
buf \U$24623 ( \33661 , \33660 );
xor \U$24624 ( \33662 , \33628 , \33661 );
and \U$24625 ( \33663 , \33212 , \33217 );
and \U$24626 ( \33664 , \33212 , \33239 );
and \U$24627 ( \33665 , \33217 , \33239 );
or \U$24628 ( \33666 , \33663 , \33664 , \33665 );
buf \U$24629 ( \33667 , \33666 );
xor \U$24630 ( \33668 , \33662 , \33667 );
buf \U$24631 ( \33669 , \33668 );
xor \U$24632 ( \33670 , \33623 , \33669 );
and \U$24633 ( \33671 , \33301 , \33670 );
and \U$24634 ( \33672 , \33196 , \33201 );
and \U$24635 ( \33673 , \33196 , \33291 );
and \U$24636 ( \33674 , \33201 , \33291 );
or \U$24637 ( \33675 , \33672 , \33673 , \33674 );
and \U$24638 ( \33676 , \33301 , \33675 );
and \U$24639 ( \33677 , \33670 , \33675 );
or \U$24640 ( \33678 , \33671 , \33676 , \33677 );
and \U$24641 ( \33679 , \33295 , \33299 );
or \U$24644 ( \33680 , \33679 , 1'b0 , 1'b0 );
xor \U$24645 ( \33681 , \33678 , \33680 );
xor \U$24659 ( \33682 , \33681 , 1'b0 );
and \U$24660 ( \33683 , \33306 , \33622 );
and \U$24661 ( \33684 , \33306 , \33669 );
and \U$24662 ( \33685 , \33622 , \33669 );
or \U$24663 ( \33686 , \33683 , \33684 , \33685 );
and \U$24664 ( \33687 , \33682 , \33686 );
and \U$24665 ( \33688 , \33423 , \33428 );
and \U$24666 ( \33689 , \33423 , \33620 );
and \U$24667 ( \33690 , \33428 , \33620 );
or \U$24668 ( \33691 , \33688 , \33689 , \33690 );
buf \U$24669 ( \33692 , \33691 );
and \U$24670 ( \33693 , \33449 , \33454 );
and \U$24671 ( \33694 , \33449 , \33618 );
and \U$24672 ( \33695 , \33454 , \33618 );
or \U$24673 ( \33696 , \33693 , \33694 , \33695 );
buf \U$24674 ( \33697 , \33696 );
and \U$24675 ( \33698 , \15940 , \25860_nG9bc9 );
and \U$24676 ( \33699 , \15937 , \26887_nG9bc6 );
or \U$24677 ( \33700 , \33698 , \33699 );
xor \U$24678 ( \33701 , \15936 , \33700 );
buf \U$24679 ( \33702 , \33701 );
buf \U$24681 ( \33703 , \33702 );
and \U$24682 ( \33704 , \13370 , \29179_nG9bbd );
and \U$24683 ( \33705 , \13367 , \30366_nG9bba );
or \U$24684 ( \33706 , \33704 , \33705 );
xor \U$24685 ( \33707 , \13366 , \33706 );
buf \U$24686 ( \33708 , \33707 );
buf \U$24688 ( \33709 , \33708 );
xor \U$24689 ( \33710 , \33703 , \33709 );
and \U$24690 ( \33711 , \12157 , \30940_nG9bb7 );
and \U$24691 ( \33712 , \12154 , \32179_nG9bb4 );
or \U$24692 ( \33713 , \33711 , \33712 );
xor \U$24693 ( \33714 , \12153 , \33713 );
buf \U$24694 ( \33715 , \33714 );
buf \U$24696 ( \33716 , \33715 );
xor \U$24697 ( \33717 , \33710 , \33716 );
buf \U$24698 ( \33718 , \33717 );
xor \U$24699 ( \33719 , \33697 , \33718 );
and \U$24700 ( \33720 , \33311 , \33328 );
and \U$24701 ( \33721 , \33311 , \33335 );
and \U$24702 ( \33722 , \33328 , \33335 );
or \U$24703 ( \33723 , \33720 , \33721 , \33722 );
buf \U$24704 ( \33724 , \33723 );
and \U$24705 ( \33725 , \33313 , \33319 );
and \U$24706 ( \33726 , \33313 , \33326 );
and \U$24707 ( \33727 , \33319 , \33326 );
or \U$24708 ( \33728 , \33725 , \33726 , \33727 );
buf \U$24709 ( \33729 , \33728 );
and \U$24711 ( \33730 , \32916 , \11283_nG9c08 );
or \U$24712 ( \33731 , 1'b0 , \33730 );
xor \U$24713 ( \33732 , 1'b0 , \33731 );
buf \U$24714 ( \33733 , \33732 );
buf \U$24716 ( \33734 , \33733 );
and \U$24717 ( \33735 , \31636 , \11598_nG9c05 );
and \U$24718 ( \33736 , \31633 , \12470_nG9c02 );
or \U$24719 ( \33737 , \33735 , \33736 );
xor \U$24720 ( \33738 , \31632 , \33737 );
buf \U$24721 ( \33739 , \33738 );
buf \U$24723 ( \33740 , \33739 );
xor \U$24724 ( \33741 , \33734 , \33740 );
buf \U$24725 ( \33742 , \33741 );
and \U$24726 ( \33743 , \29853 , \12801_nG9bff );
and \U$24727 ( \33744 , \29850 , \13705_nG9bfc );
or \U$24728 ( \33745 , \33743 , \33744 );
xor \U$24729 ( \33746 , \29849 , \33745 );
buf \U$24730 ( \33747 , \33746 );
buf \U$24732 ( \33748 , \33747 );
xor \U$24733 ( \33749 , \33742 , \33748 );
buf \U$24734 ( \33750 , \33749 );
xor \U$24735 ( \33751 , \33729 , \33750 );
and \U$24736 ( \33752 , \24792 , \16680_nG9bed );
and \U$24737 ( \33753 , \24789 , \17665_nG9bea );
or \U$24738 ( \33754 , \33752 , \33753 );
xor \U$24739 ( \33755 , \24788 , \33754 );
buf \U$24740 ( \33756 , \33755 );
buf \U$24742 ( \33757 , \33756 );
xor \U$24743 ( \33758 , \33751 , \33757 );
buf \U$24744 ( \33759 , \33758 );
xor \U$24745 ( \33760 , \33724 , \33759 );
and \U$24746 ( \33761 , \17297 , \24226_nG9bcf );
and \U$24747 ( \33762 , \17294 , \25298_nG9bcc );
or \U$24748 ( \33763 , \33761 , \33762 );
xor \U$24749 ( \33764 , \17293 , \33763 );
buf \U$24750 ( \33765 , \33764 );
buf \U$24752 ( \33766 , \33765 );
xor \U$24753 ( \33767 , \33760 , \33766 );
buf \U$24754 ( \33768 , \33767 );
and \U$24755 ( \33769 , \33342 , \33362 );
and \U$24756 ( \33770 , \33342 , \33369 );
and \U$24757 ( \33771 , \33362 , \33369 );
or \U$24758 ( \33772 , \33769 , \33770 , \33771 );
buf \U$24759 ( \33773 , \33772 );
and \U$24760 ( \33774 , \33347 , \33353 );
and \U$24761 ( \33775 , \33347 , \33360 );
and \U$24762 ( \33776 , \33353 , \33360 );
or \U$24763 ( \33777 , \33774 , \33775 , \33776 );
buf \U$24764 ( \33778 , \33777 );
and \U$24765 ( \33779 , \28118 , \14070_nG9bf9 );
and \U$24766 ( \33780 , \28115 , \14984_nG9bf6 );
or \U$24767 ( \33781 , \33779 , \33780 );
xor \U$24768 ( \33782 , \28114 , \33781 );
buf \U$24769 ( \33783 , \33782 );
buf \U$24771 ( \33784 , \33783 );
xor \U$24772 ( \33785 , \33778 , \33784 );
and \U$24773 ( \33786 , \26431 , \15373_nG9bf3 );
and \U$24774 ( \33787 , \26428 , \16315_nG9bf0 );
or \U$24775 ( \33788 , \33786 , \33787 );
xor \U$24776 ( \33789 , \26427 , \33788 );
buf \U$24777 ( \33790 , \33789 );
buf \U$24779 ( \33791 , \33790 );
xor \U$24780 ( \33792 , \33785 , \33791 );
buf \U$24781 ( \33793 , \33792 );
xor \U$24782 ( \33794 , \33773 , \33793 );
and \U$24783 ( \33795 , \18702 , \22629_nG9bd5 );
and \U$24784 ( \33796 , \18699 , \23696_nG9bd2 );
or \U$24785 ( \33797 , \33795 , \33796 );
xor \U$24786 ( \33798 , \18698 , \33797 );
buf \U$24787 ( \33799 , \33798 );
buf \U$24789 ( \33800 , \33799 );
xor \U$24790 ( \33801 , \33794 , \33800 );
buf \U$24791 ( \33802 , \33801 );
xor \U$24792 ( \33803 , \33768 , \33802 );
and \U$24793 ( \33804 , \10421 , \32888_nG9bb1 );
and \U$24794 ( \33805 , \10418 , \33181_nG9bae );
or \U$24795 ( \33806 , \33804 , \33805 );
xor \U$24796 ( \33807 , \10417 , \33806 );
buf \U$24797 ( \33808 , \33807 );
buf \U$24799 ( \33809 , \33808 );
xor \U$24800 ( \33810 , \33803 , \33809 );
buf \U$24801 ( \33811 , \33810 );
xor \U$24802 ( \33812 , \33719 , \33811 );
buf \U$24803 ( \33813 , \33812 );
xor \U$24804 ( \33814 , \33692 , \33813 );
and \U$24805 ( \33815 , \33406 , \33412 );
and \U$24806 ( \33816 , \33406 , \33419 );
and \U$24807 ( \33817 , \33412 , \33419 );
or \U$24808 ( \33818 , \33815 , \33816 , \33817 );
buf \U$24809 ( \33819 , \33818 );
and \U$24810 ( \33820 , \33371 , \33377 );
and \U$24811 ( \33821 , \33371 , \33384 );
and \U$24812 ( \33822 , \33377 , \33384 );
or \U$24813 ( \33823 , \33820 , \33821 , \33822 );
buf \U$24814 ( \33824 , \33823 );
and \U$24815 ( \33825 , \23201 , \18107_nG9be7 );
and \U$24816 ( \33826 , \23198 , \19091_nG9be4 );
or \U$24817 ( \33827 , \33825 , \33826 );
xor \U$24818 ( \33828 , \23197 , \33827 );
buf \U$24819 ( \33829 , \33828 );
buf \U$24821 ( \33830 , \33829 );
and \U$24822 ( \33831 , \21658 , \19586_nG9be1 );
and \U$24823 ( \33832 , \21655 , \20608_nG9bde );
or \U$24824 ( \33833 , \33831 , \33832 );
xor \U$24825 ( \33834 , \21654 , \33833 );
buf \U$24826 ( \33835 , \33834 );
buf \U$24828 ( \33836 , \33835 );
xor \U$24829 ( \33837 , \33830 , \33836 );
and \U$24830 ( \33838 , \20155 , \21086_nG9bdb );
and \U$24831 ( \33839 , \20152 , \22129_nG9bd8 );
or \U$24832 ( \33840 , \33838 , \33839 );
xor \U$24833 ( \33841 , \20151 , \33840 );
buf \U$24834 ( \33842 , \33841 );
buf \U$24836 ( \33843 , \33842 );
xor \U$24837 ( \33844 , \33837 , \33843 );
buf \U$24838 ( \33845 , \33844 );
xor \U$24839 ( \33846 , \33824 , \33845 );
and \U$24840 ( \33847 , \14631 , \27416_nG9bc3 );
and \U$24841 ( \33848 , \14628 , \28602_nG9bc0 );
or \U$24842 ( \33849 , \33847 , \33848 );
xor \U$24843 ( \33850 , \14627 , \33849 );
buf \U$24844 ( \33851 , \33850 );
buf \U$24846 ( \33852 , \33851 );
xor \U$24847 ( \33853 , \33846 , \33852 );
buf \U$24848 ( \33854 , \33853 );
xor \U$24849 ( \33855 , \33819 , \33854 );
and \U$24850 ( \33856 , \33644 , \33650 );
and \U$24851 ( \33857 , \33644 , \33657 );
and \U$24852 ( \33858 , \33650 , \33657 );
or \U$24853 ( \33859 , \33856 , \33857 , \33858 );
buf \U$24854 ( \33860 , \33859 );
xor \U$24855 ( \33861 , \33855 , \33860 );
buf \U$24856 ( \33862 , \33861 );
xor \U$24857 ( \33863 , \33814 , \33862 );
buf \U$24858 ( \33864 , \33863 );
and \U$24859 ( \33865 , \33628 , \33661 );
and \U$24860 ( \33866 , \33628 , \33667 );
and \U$24861 ( \33867 , \33661 , \33667 );
or \U$24862 ( \33868 , \33865 , \33866 , \33867 );
buf \U$24863 ( \33869 , \33868 );
xor \U$24864 ( \33870 , \33864 , \33869 );
and \U$24865 ( \33871 , \33337 , \33386 );
and \U$24866 ( \33872 , \33337 , \33392 );
and \U$24867 ( \33873 , \33386 , \33392 );
or \U$24868 ( \33874 , \33871 , \33872 , \33873 );
buf \U$24869 ( \33875 , \33874 );
and \U$24870 ( \33876 , \33434 , \33440 );
and \U$24871 ( \33877 , \33434 , \33447 );
and \U$24872 ( \33878 , \33440 , \33447 );
or \U$24873 ( \33879 , \33876 , \33877 , \33878 );
buf \U$24874 ( \33880 , \33879 );
xor \U$24875 ( \33881 , \33875 , \33880 );
and \U$24876 ( \33882 , \10707 , \33613_nG9bab );
and \U$24877 ( \33883 , \33515 , \33519 );
and \U$24878 ( \33884 , \33519 , \33601 );
and \U$24879 ( \33885 , \33515 , \33601 );
or \U$24880 ( \33886 , \33883 , \33884 , \33885 );
and \U$24881 ( \33887 , \33468 , \33472 );
and \U$24882 ( \33888 , \33472 , \33477 );
and \U$24883 ( \33889 , \33468 , \33477 );
or \U$24884 ( \33890 , \33887 , \33888 , \33889 );
and \U$24885 ( \33891 , \33487 , \33491 );
and \U$24886 ( \33892 , \33491 , \33496 );
and \U$24887 ( \33893 , \33487 , \33496 );
or \U$24888 ( \33894 , \33891 , \33892 , \33893 );
and \U$24889 ( \33895 , \33502 , \10980 );
and \U$24890 ( \33896 , \10980 , \33507 );
and \U$24891 ( \33897 , \33502 , \33507 );
or \U$24892 ( \33898 , \33895 , \33896 , \33897 );
xor \U$24893 ( \33899 , \33894 , \33898 );
and \U$24894 ( \33900 , \33560 , \33564 );
and \U$24895 ( \33901 , \33564 , \33569 );
and \U$24896 ( \33902 , \33560 , \33569 );
or \U$24897 ( \33903 , \33900 , \33901 , \33902 );
and \U$24898 ( \33904 , \33574 , \33578 );
and \U$24899 ( \33905 , \33578 , \33583 );
and \U$24900 ( \33906 , \33574 , \33583 );
or \U$24901 ( \33907 , \33904 , \33905 , \33906 );
xor \U$24902 ( \33908 , \33903 , \33907 );
and \U$24903 ( \33909 , \33589 , \33593 );
and \U$24904 ( \33910 , \33593 , \33598 );
and \U$24905 ( \33911 , \33589 , \33598 );
or \U$24906 ( \33912 , \33909 , \33910 , \33911 );
xor \U$24907 ( \33913 , \33908 , \33912 );
xor \U$24908 ( \33914 , \33899 , \33913 );
xor \U$24909 ( \33915 , \33890 , \33914 );
and \U$24910 ( \33916 , \33528 , \33539 );
and \U$24911 ( \33917 , \33539 , \33554 );
and \U$24912 ( \33918 , \33528 , \33554 );
or \U$24913 ( \33919 , \33916 , \33917 , \33918 );
and \U$24914 ( \33920 , \33570 , \33584 );
and \U$24915 ( \33921 , \33584 , \33599 );
and \U$24916 ( \33922 , \33570 , \33599 );
or \U$24917 ( \33923 , \33920 , \33921 , \33922 );
xor \U$24918 ( \33924 , \33919 , \33923 );
and \U$24919 ( \33925 , \33532 , \33536 );
and \U$24920 ( \33926 , \33536 , \33538 );
and \U$24921 ( \33927 , \33532 , \33538 );
or \U$24922 ( \33928 , \33925 , \33926 , \33927 );
not \U$24923 ( \33929 , \10980 );
buf \U$24924 ( \33930 , \33929 );
xor \U$24925 ( \33931 , \33928 , \33930 );
and \U$24926 ( \33932 , \32794 , \11574 );
not \U$24927 ( \33933 , \33932 );
xnor \U$24928 ( \33934 , \33933 , \11580 );
not \U$24929 ( \33935 , \33934 );
xor \U$24930 ( \33936 , \33931 , \33935 );
xor \U$24931 ( \33937 , \33924 , \33936 );
xor \U$24932 ( \33938 , \33915 , \33937 );
xor \U$24933 ( \33939 , \33886 , \33938 );
and \U$24934 ( \33940 , \33524 , \33555 );
and \U$24935 ( \33941 , \33555 , \33600 );
and \U$24936 ( \33942 , \33524 , \33600 );
or \U$24937 ( \33943 , \33940 , \33941 , \33942 );
and \U$24938 ( \33944 , \33464 , \33478 );
and \U$24939 ( \33945 , \33478 , \33509 );
and \U$24940 ( \33946 , \33464 , \33509 );
or \U$24941 ( \33947 , \33944 , \33945 , \33946 );
xor \U$24942 ( \33948 , \33943 , \33947 );
and \U$24943 ( \33949 , \33483 , \33497 );
and \U$24944 ( \33950 , \33497 , \33508 );
and \U$24945 ( \33951 , \33483 , \33508 );
or \U$24946 ( \33952 , \33949 , \33950 , \33951 );
and \U$24947 ( \33953 , \30802 , \12790 );
and \U$24948 ( \33954 , \32054 , \12461 );
nor \U$24949 ( \33955 , \33953 , \33954 );
xnor \U$24950 ( \33956 , \33955 , \12780 );
and \U$24951 ( \33957 , \27313 , \15336 );
and \U$24952 ( \33958 , \28534 , \14963 );
nor \U$24953 ( \33959 , \33957 , \33958 );
xnor \U$24954 ( \33960 , \33959 , \15342 );
xor \U$24955 ( \33961 , \33956 , \33960 );
and \U$24956 ( \33962 , \11270 , \32802 );
xor \U$24957 ( \33963 , \33961 , \33962 );
and \U$24958 ( \33964 , \24199 , \18090 );
and \U$24959 ( \33965 , \25272 , \17655 );
nor \U$24960 ( \33966 , \33964 , \33965 );
xnor \U$24961 ( \33967 , \33966 , \18046 );
and \U$24962 ( \33968 , \15321 , \27397 );
and \U$24963 ( \33969 , \16267 , \26807 );
nor \U$24964 ( \33970 , \33968 , \33969 );
xnor \U$24965 ( \33971 , \33970 , \27295 );
xor \U$24966 ( \33972 , \33967 , \33971 );
and \U$24967 ( \33973 , \14024 , \29070 );
and \U$24968 ( \33974 , \14950 , \28526 );
nor \U$24969 ( \33975 , \33973 , \33974 );
xnor \U$24970 ( \33976 , \33975 , \29076 );
xor \U$24971 ( \33977 , \33972 , \33976 );
xor \U$24972 ( \33978 , \33963 , \33977 );
and \U$24973 ( \33979 , \29084 , \14054 );
and \U$24974 ( \33980 , \30268 , \13692 );
nor \U$24975 ( \33981 , \33979 , \33980 );
xnor \U$24976 ( \33982 , \33981 , \14035 );
and \U$24977 ( \33983 , \18035 , \24138 );
and \U$24978 ( \33984 , \19032 , \23630 );
nor \U$24979 ( \33985 , \33983 , \33984 );
xnor \U$24980 ( \33986 , \33985 , \24144 );
xor \U$24981 ( \33987 , \33982 , \33986 );
and \U$24982 ( \33988 , \16655 , \25826 );
and \U$24983 ( \33989 , \17627 , \25264 );
nor \U$24984 ( \33990 , \33988 , \33989 );
xnor \U$24985 ( \33991 , \33990 , \25773 );
xor \U$24986 ( \33992 , \33987 , \33991 );
xor \U$24987 ( \33993 , \33978 , \33992 );
xor \U$24988 ( \33994 , \33952 , \33993 );
and \U$24989 ( \33995 , \33544 , \33548 );
and \U$24990 ( \33996 , \33548 , \33553 );
and \U$24991 ( \33997 , \33544 , \33553 );
or \U$24992 ( \33998 , \33995 , \33996 , \33997 );
and \U$24993 ( \33999 , \22556 , \19534 );
and \U$24994 ( \34000 , \23617 , \19045 );
nor \U$24995 ( \34001 , \33999 , \34000 );
xnor \U$24996 ( \34002 , \34001 , \19540 );
and \U$24997 ( \34003 , \12769 , \30823 );
and \U$24998 ( \34004 , \13679 , \30246 );
nor \U$24999 ( \34005 , \34003 , \34004 );
xnor \U$25000 ( \34006 , \34005 , \30813 );
xor \U$25001 ( \34007 , \34002 , \34006 );
and \U$25002 ( \34008 , \11586 , \32854 );
and \U$25003 ( \34009 , \12448 , \32067 );
nor \U$25004 ( \34010 , \34008 , \34009 );
xnor \U$25005 ( \34011 , \34010 , \32805 );
xor \U$25006 ( \34012 , \34007 , \34011 );
xor \U$25007 ( \34013 , \33998 , \34012 );
and \U$25008 ( \34014 , \25815 , \16635 );
and \U$25009 ( \34015 , \26829 , \16301 );
nor \U$25010 ( \34016 , \34014 , \34015 );
xnor \U$25011 ( \34017 , \34016 , \16625 );
and \U$25012 ( \34018 , \21033 , \21005 );
and \U$25013 ( \34019 , \22090 , \20557 );
nor \U$25014 ( \34020 , \34018 , \34019 );
xnor \U$25015 ( \34021 , \34020 , \21011 );
xor \U$25016 ( \34022 , \34017 , \34021 );
and \U$25017 ( \34023 , \19558 , \22542 );
and \U$25018 ( \34024 , \20544 , \22103 );
nor \U$25019 ( \34025 , \34023 , \34024 );
xnor \U$25020 ( \34026 , \34025 , \22548 );
xor \U$25021 ( \34027 , \34022 , \34026 );
xor \U$25022 ( \34028 , \34013 , \34027 );
xor \U$25023 ( \34029 , \33994 , \34028 );
xor \U$25024 ( \34030 , \33948 , \34029 );
xor \U$25025 ( \34031 , \33939 , \34030 );
and \U$25026 ( \34032 , \33460 , \33510 );
and \U$25027 ( \34033 , \33510 , \33602 );
and \U$25028 ( \34034 , \33460 , \33602 );
or \U$25029 ( \34035 , \34032 , \34033 , \34034 );
xor \U$25030 ( \34036 , \34031 , \34035 );
and \U$25031 ( \34037 , \33603 , \33607 );
and \U$25032 ( \34038 , \33608 , \33611 );
or \U$25033 ( \34039 , \34037 , \34038 );
xor \U$25034 ( \34040 , \34036 , \34039 );
buf g9ba8 ( \34041_nG9ba8 , \34040 );
and \U$25035 ( \34042 , \10704 , \34041_nG9ba8 );
or \U$25036 ( \34043 , \33882 , \34042 );
xor \U$25037 ( \34044 , \10703 , \34043 );
buf \U$25038 ( \34045 , \34044 );
buf \U$25040 ( \34046 , \34045 );
xor \U$25041 ( \34047 , \33881 , \34046 );
buf \U$25042 ( \34048 , \34047 );
and \U$25043 ( \34049 , \33394 , \33399 );
and \U$25044 ( \34050 , \33394 , \33421 );
and \U$25045 ( \34051 , \33399 , \33421 );
or \U$25046 ( \34052 , \34049 , \34050 , \34051 );
buf \U$25047 ( \34053 , \34052 );
xor \U$25048 ( \34054 , \34048 , \34053 );
and \U$25049 ( \34055 , \33633 , \33638 );
and \U$25050 ( \34056 , \33633 , \33659 );
and \U$25051 ( \34057 , \33638 , \33659 );
or \U$25052 ( \34058 , \34055 , \34056 , \34057 );
buf \U$25053 ( \34059 , \34058 );
xor \U$25054 ( \34060 , \34054 , \34059 );
buf \U$25055 ( \34061 , \34060 );
xor \U$25056 ( \34062 , \33870 , \34061 );
and \U$25057 ( \34063 , \33682 , \34062 );
and \U$25058 ( \34064 , \33686 , \34062 );
or \U$25059 ( \34065 , \33687 , \34063 , \34064 );
and \U$25060 ( \34066 , \33678 , \33680 );
or \U$25063 ( \34067 , \34066 , 1'b0 , 1'b0 );
xor \U$25064 ( \34068 , \34065 , \34067 );
xor \U$25068 ( \34069 , \34068 , 1'b0 );
xor \U$25075 ( \34070 , \34069 , 1'b0 );
and \U$25076 ( \34071 , \33864 , \33869 );
and \U$25077 ( \34072 , \33864 , \34061 );
and \U$25078 ( \34073 , \33869 , \34061 );
or \U$25079 ( \34074 , \34071 , \34072 , \34073 );
xor \U$25080 ( \34075 , \34070 , \34074 );
and \U$25081 ( \34076 , \33692 , \33813 );
and \U$25082 ( \34077 , \33692 , \33862 );
and \U$25083 ( \34078 , \33813 , \33862 );
or \U$25084 ( \34079 , \34076 , \34077 , \34078 );
buf \U$25085 ( \34080 , \34079 );
and \U$25086 ( \34081 , \33778 , \33784 );
and \U$25087 ( \34082 , \33778 , \33791 );
and \U$25088 ( \34083 , \33784 , \33791 );
or \U$25089 ( \34084 , \34081 , \34082 , \34083 );
buf \U$25090 ( \34085 , \34084 );
and \U$25092 ( \34086 , \32916 , \11598_nG9c05 );
or \U$25093 ( \34087 , 1'b0 , \34086 );
xor \U$25094 ( \34088 , 1'b0 , \34087 );
buf \U$25095 ( \34089 , \34088 );
buf \U$25097 ( \34090 , \34089 );
and \U$25098 ( \34091 , \31636 , \12470_nG9c02 );
and \U$25099 ( \34092 , \31633 , \12801_nG9bff );
or \U$25100 ( \34093 , \34091 , \34092 );
xor \U$25101 ( \34094 , \31632 , \34093 );
buf \U$25102 ( \34095 , \34094 );
buf \U$25104 ( \34096 , \34095 );
xor \U$25105 ( \34097 , \34090 , \34096 );
buf \U$25106 ( \34098 , \34097 );
and \U$25107 ( \34099 , \33734 , \33740 );
buf \U$25108 ( \34100 , \34099 );
xor \U$25109 ( \34101 , \34098 , \34100 );
and \U$25110 ( \34102 , \29853 , \13705_nG9bfc );
and \U$25111 ( \34103 , \29850 , \14070_nG9bf9 );
or \U$25112 ( \34104 , \34102 , \34103 );
xor \U$25113 ( \34105 , \29849 , \34104 );
buf \U$25114 ( \34106 , \34105 );
buf \U$25116 ( \34107 , \34106 );
xor \U$25117 ( \34108 , \34101 , \34107 );
buf \U$25118 ( \34109 , \34108 );
xor \U$25119 ( \34110 , \34085 , \34109 );
and \U$25120 ( \34111 , \24792 , \17665_nG9bea );
and \U$25121 ( \34112 , \24789 , \18107_nG9be7 );
or \U$25122 ( \34113 , \34111 , \34112 );
xor \U$25123 ( \34114 , \24788 , \34113 );
buf \U$25124 ( \34115 , \34114 );
buf \U$25126 ( \34116 , \34115 );
xor \U$25127 ( \34117 , \34110 , \34116 );
buf \U$25128 ( \34118 , \34117 );
and \U$25129 ( \34119 , \33830 , \33836 );
and \U$25130 ( \34120 , \33830 , \33843 );
and \U$25131 ( \34121 , \33836 , \33843 );
or \U$25132 ( \34122 , \34119 , \34120 , \34121 );
buf \U$25133 ( \34123 , \34122 );
xor \U$25134 ( \34124 , \34118 , \34123 );
and \U$25135 ( \34125 , \15940 , \26887_nG9bc6 );
and \U$25136 ( \34126 , \15937 , \27416_nG9bc3 );
or \U$25137 ( \34127 , \34125 , \34126 );
xor \U$25138 ( \34128 , \15936 , \34127 );
buf \U$25139 ( \34129 , \34128 );
buf \U$25141 ( \34130 , \34129 );
xor \U$25142 ( \34131 , \34124 , \34130 );
buf \U$25143 ( \34132 , \34131 );
and \U$25144 ( \34133 , \33824 , \33845 );
and \U$25145 ( \34134 , \33824 , \33852 );
and \U$25146 ( \34135 , \33845 , \33852 );
or \U$25147 ( \34136 , \34133 , \34134 , \34135 );
buf \U$25148 ( \34137 , \34136 );
xor \U$25149 ( \34138 , \34132 , \34137 );
and \U$25150 ( \34139 , \10707 , \34041_nG9ba8 );
and \U$25151 ( \34140 , \33886 , \33938 );
and \U$25152 ( \34141 , \33938 , \34030 );
and \U$25153 ( \34142 , \33886 , \34030 );
or \U$25154 ( \34143 , \34140 , \34141 , \34142 );
and \U$25155 ( \34144 , \33943 , \33947 );
and \U$25156 ( \34145 , \33947 , \34029 );
and \U$25157 ( \34146 , \33943 , \34029 );
or \U$25158 ( \34147 , \34144 , \34145 , \34146 );
and \U$25159 ( \34148 , \33894 , \33898 );
and \U$25160 ( \34149 , \33898 , \33913 );
and \U$25161 ( \34150 , \33894 , \33913 );
or \U$25162 ( \34151 , \34148 , \34149 , \34150 );
and \U$25163 ( \34152 , \33919 , \33923 );
and \U$25164 ( \34153 , \33923 , \33936 );
and \U$25165 ( \34154 , \33919 , \33936 );
or \U$25166 ( \34155 , \34152 , \34153 , \34154 );
xor \U$25167 ( \34156 , \34151 , \34155 );
and \U$25168 ( \34157 , \33963 , \33977 );
and \U$25169 ( \34158 , \33977 , \33992 );
and \U$25170 ( \34159 , \33963 , \33992 );
or \U$25171 ( \34160 , \34157 , \34158 , \34159 );
and \U$25172 ( \34161 , \33998 , \34012 );
and \U$25173 ( \34162 , \34012 , \34027 );
and \U$25174 ( \34163 , \33998 , \34027 );
or \U$25175 ( \34164 , \34161 , \34162 , \34163 );
xor \U$25176 ( \34165 , \34160 , \34164 );
and \U$25177 ( \34166 , \34017 , \34021 );
and \U$25178 ( \34167 , \34021 , \34026 );
and \U$25179 ( \34168 , \34017 , \34026 );
or \U$25180 ( \34169 , \34166 , \34167 , \34168 );
and \U$25181 ( \34170 , \33967 , \33971 );
and \U$25182 ( \34171 , \33971 , \33976 );
and \U$25183 ( \34172 , \33967 , \33976 );
or \U$25184 ( \34173 , \34170 , \34171 , \34172 );
xor \U$25185 ( \34174 , \34169 , \34173 );
and \U$25186 ( \34175 , \33982 , \33986 );
and \U$25187 ( \34176 , \33986 , \33991 );
and \U$25188 ( \34177 , \33982 , \33991 );
or \U$25189 ( \34178 , \34175 , \34176 , \34177 );
xor \U$25190 ( \34179 , \34174 , \34178 );
xor \U$25191 ( \34180 , \34165 , \34179 );
xor \U$25192 ( \34181 , \34156 , \34180 );
xor \U$25193 ( \34182 , \34147 , \34181 );
and \U$25194 ( \34183 , \33952 , \33993 );
and \U$25195 ( \34184 , \33993 , \34028 );
and \U$25196 ( \34185 , \33952 , \34028 );
or \U$25197 ( \34186 , \34183 , \34184 , \34185 );
and \U$25198 ( \34187 , \33890 , \33914 );
and \U$25199 ( \34188 , \33914 , \33937 );
and \U$25200 ( \34189 , \33890 , \33937 );
or \U$25201 ( \34190 , \34187 , \34188 , \34189 );
xor \U$25202 ( \34191 , \34186 , \34190 );
and \U$25203 ( \34192 , \23617 , \19534 );
and \U$25204 ( \34193 , \24199 , \19045 );
nor \U$25205 ( \34194 , \34192 , \34193 );
xnor \U$25206 ( \34195 , \34194 , \19540 );
and \U$25207 ( \34196 , \14950 , \29070 );
and \U$25208 ( \34197 , \15321 , \28526 );
nor \U$25209 ( \34198 , \34196 , \34197 );
xnor \U$25210 ( \34199 , \34198 , \29076 );
xor \U$25211 ( \34200 , \34195 , \34199 );
and \U$25212 ( \34201 , \13679 , \30823 );
and \U$25213 ( \34202 , \14024 , \30246 );
nor \U$25214 ( \34203 , \34201 , \34202 );
xnor \U$25215 ( \34204 , \34203 , \30813 );
xor \U$25216 ( \34205 , \34200 , \34204 );
and \U$25217 ( \34206 , \26829 , \16635 );
and \U$25218 ( \34207 , \27313 , \16301 );
nor \U$25219 ( \34208 , \34206 , \34207 );
xnor \U$25220 ( \34209 , \34208 , \16625 );
and \U$25221 ( \34210 , \19032 , \24138 );
and \U$25222 ( \34211 , \19558 , \23630 );
nor \U$25223 ( \34212 , \34210 , \34211 );
xnor \U$25224 ( \34213 , \34212 , \24144 );
xor \U$25225 ( \34214 , \34209 , \34213 );
and \U$25226 ( \34215 , \17627 , \25826 );
and \U$25227 ( \34216 , \18035 , \25264 );
nor \U$25228 ( \34217 , \34215 , \34216 );
xnor \U$25229 ( \34218 , \34217 , \25773 );
xor \U$25230 ( \34219 , \34214 , \34218 );
xor \U$25231 ( \34220 , \34205 , \34219 );
and \U$25232 ( \34221 , \30268 , \14054 );
and \U$25233 ( \34222 , \30802 , \13692 );
nor \U$25234 ( \34223 , \34221 , \34222 );
xnor \U$25235 ( \34224 , \34223 , \14035 );
and \U$25236 ( \34225 , \25272 , \18090 );
and \U$25237 ( \34226 , \25815 , \17655 );
nor \U$25238 ( \34227 , \34225 , \34226 );
xnor \U$25239 ( \34228 , \34227 , \18046 );
xor \U$25240 ( \34229 , \34224 , \34228 );
and \U$25241 ( \34230 , \16267 , \27397 );
and \U$25242 ( \34231 , \16655 , \26807 );
nor \U$25243 ( \34232 , \34230 , \34231 );
xnor \U$25244 ( \34233 , \34232 , \27295 );
xor \U$25245 ( \34234 , \34229 , \34233 );
xor \U$25246 ( \34235 , \34220 , \34234 );
and \U$25247 ( \34236 , \34002 , \34006 );
and \U$25248 ( \34237 , \34006 , \34011 );
and \U$25249 ( \34238 , \34002 , \34011 );
or \U$25250 ( \34239 , \34236 , \34237 , \34238 );
not \U$25251 ( \34240 , \11580 );
and \U$25252 ( \34241 , \32054 , \12790 );
and \U$25253 ( \34242 , \32794 , \12461 );
nor \U$25254 ( \34243 , \34241 , \34242 );
xnor \U$25255 ( \34244 , \34243 , \12780 );
xor \U$25256 ( \34245 , \34240 , \34244 );
and \U$25257 ( \34246 , \28534 , \15336 );
and \U$25258 ( \34247 , \29084 , \14963 );
nor \U$25259 ( \34248 , \34246 , \34247 );
xnor \U$25260 ( \34249 , \34248 , \15342 );
xor \U$25261 ( \34250 , \34245 , \34249 );
xor \U$25262 ( \34251 , \34239 , \34250 );
and \U$25263 ( \34252 , \22090 , \21005 );
and \U$25264 ( \34253 , \22556 , \20557 );
nor \U$25265 ( \34254 , \34252 , \34253 );
xnor \U$25266 ( \34255 , \34254 , \21011 );
and \U$25267 ( \34256 , \20544 , \22542 );
and \U$25268 ( \34257 , \21033 , \22103 );
nor \U$25269 ( \34258 , \34256 , \34257 );
xnor \U$25270 ( \34259 , \34258 , \22548 );
xor \U$25271 ( \34260 , \34255 , \34259 );
and \U$25272 ( \34261 , \11586 , \32802 );
xor \U$25273 ( \34262 , \34260 , \34261 );
xor \U$25274 ( \34263 , \34251 , \34262 );
xor \U$25275 ( \34264 , \34235 , \34263 );
and \U$25276 ( \34265 , \33903 , \33907 );
and \U$25277 ( \34266 , \33907 , \33912 );
and \U$25278 ( \34267 , \33903 , \33912 );
or \U$25279 ( \34268 , \34265 , \34266 , \34267 );
and \U$25280 ( \34269 , \33928 , \33930 );
and \U$25281 ( \34270 , \33930 , \33935 );
and \U$25282 ( \34271 , \33928 , \33935 );
or \U$25283 ( \34272 , \34269 , \34270 , \34271 );
xor \U$25284 ( \34273 , \34268 , \34272 );
and \U$25285 ( \34274 , \33956 , \33960 );
and \U$25286 ( \34275 , \33960 , \33962 );
and \U$25287 ( \34276 , \33956 , \33962 );
or \U$25288 ( \34277 , \34274 , \34275 , \34276 );
buf \U$25289 ( \34278 , \33934 );
xor \U$25290 ( \34279 , \34277 , \34278 );
and \U$25291 ( \34280 , \12448 , \32854 );
and \U$25292 ( \34281 , \12769 , \32067 );
nor \U$25293 ( \34282 , \34280 , \34281 );
xnor \U$25294 ( \34283 , \34282 , \32805 );
xor \U$25295 ( \34284 , \34279 , \34283 );
xor \U$25296 ( \34285 , \34273 , \34284 );
xor \U$25297 ( \34286 , \34264 , \34285 );
xor \U$25298 ( \34287 , \34191 , \34286 );
xor \U$25299 ( \34288 , \34182 , \34287 );
xor \U$25300 ( \34289 , \34143 , \34288 );
and \U$25301 ( \34290 , \34031 , \34035 );
and \U$25302 ( \34291 , \34036 , \34039 );
or \U$25303 ( \34292 , \34290 , \34291 );
xor \U$25304 ( \34293 , \34289 , \34292 );
buf g9ba5 ( \34294_nG9ba5 , \34293 );
and \U$25305 ( \34295 , \10704 , \34294_nG9ba5 );
or \U$25306 ( \34296 , \34139 , \34295 );
xor \U$25307 ( \34297 , \10703 , \34296 );
buf \U$25308 ( \34298 , \34297 );
buf \U$25310 ( \34299 , \34298 );
xor \U$25311 ( \34300 , \34138 , \34299 );
buf \U$25312 ( \34301 , \34300 );
and \U$25313 ( \34302 , \33819 , \33854 );
and \U$25314 ( \34303 , \33819 , \33860 );
and \U$25315 ( \34304 , \33854 , \33860 );
or \U$25316 ( \34305 , \34302 , \34303 , \34304 );
buf \U$25317 ( \34306 , \34305 );
xor \U$25318 ( \34307 , \34301 , \34306 );
and \U$25319 ( \34308 , \33724 , \33759 );
and \U$25320 ( \34309 , \33724 , \33766 );
and \U$25321 ( \34310 , \33759 , \33766 );
or \U$25322 ( \34311 , \34308 , \34309 , \34310 );
buf \U$25323 ( \34312 , \34311 );
and \U$25324 ( \34313 , \33773 , \33793 );
and \U$25325 ( \34314 , \33773 , \33800 );
and \U$25326 ( \34315 , \33793 , \33800 );
or \U$25327 ( \34316 , \34313 , \34314 , \34315 );
buf \U$25328 ( \34317 , \34316 );
xor \U$25329 ( \34318 , \34312 , \34317 );
and \U$25330 ( \34319 , \13370 , \30366_nG9bba );
and \U$25331 ( \34320 , \13367 , \30940_nG9bb7 );
or \U$25332 ( \34321 , \34319 , \34320 );
xor \U$25333 ( \34322 , \13366 , \34321 );
buf \U$25334 ( \34323 , \34322 );
buf \U$25336 ( \34324 , \34323 );
xor \U$25337 ( \34325 , \34318 , \34324 );
buf \U$25338 ( \34326 , \34325 );
and \U$25339 ( \34327 , \33742 , \33748 );
buf \U$25340 ( \34328 , \34327 );
and \U$25341 ( \34329 , \28118 , \14984_nG9bf6 );
and \U$25342 ( \34330 , \28115 , \15373_nG9bf3 );
or \U$25343 ( \34331 , \34329 , \34330 );
xor \U$25344 ( \34332 , \28114 , \34331 );
buf \U$25345 ( \34333 , \34332 );
buf \U$25347 ( \34334 , \34333 );
xor \U$25348 ( \34335 , \34328 , \34334 );
and \U$25349 ( \34336 , \26431 , \16315_nG9bf0 );
and \U$25350 ( \34337 , \26428 , \16680_nG9bed );
or \U$25351 ( \34338 , \34336 , \34337 );
xor \U$25352 ( \34339 , \26427 , \34338 );
buf \U$25353 ( \34340 , \34339 );
buf \U$25355 ( \34341 , \34340 );
xor \U$25356 ( \34342 , \34335 , \34341 );
buf \U$25357 ( \34343 , \34342 );
and \U$25358 ( \34344 , \23201 , \19091_nG9be4 );
and \U$25359 ( \34345 , \23198 , \19586_nG9be1 );
or \U$25360 ( \34346 , \34344 , \34345 );
xor \U$25361 ( \34347 , \23197 , \34346 );
buf \U$25362 ( \34348 , \34347 );
buf \U$25364 ( \34349 , \34348 );
xor \U$25365 ( \34350 , \34343 , \34349 );
and \U$25366 ( \34351 , \21658 , \20608_nG9bde );
and \U$25367 ( \34352 , \21655 , \21086_nG9bdb );
or \U$25368 ( \34353 , \34351 , \34352 );
xor \U$25369 ( \34354 , \21654 , \34353 );
buf \U$25370 ( \34355 , \34354 );
buf \U$25372 ( \34356 , \34355 );
xor \U$25373 ( \34357 , \34350 , \34356 );
buf \U$25374 ( \34358 , \34357 );
and \U$25375 ( \34359 , \17297 , \25298_nG9bcc );
and \U$25376 ( \34360 , \17294 , \25860_nG9bc9 );
or \U$25377 ( \34361 , \34359 , \34360 );
xor \U$25378 ( \34362 , \17293 , \34361 );
buf \U$25379 ( \34363 , \34362 );
buf \U$25381 ( \34364 , \34363 );
xor \U$25382 ( \34365 , \34358 , \34364 );
and \U$25383 ( \34366 , \14631 , \28602_nG9bc0 );
and \U$25384 ( \34367 , \14628 , \29179_nG9bbd );
or \U$25385 ( \34368 , \34366 , \34367 );
xor \U$25386 ( \34369 , \14627 , \34368 );
buf \U$25387 ( \34370 , \34369 );
buf \U$25389 ( \34371 , \34370 );
xor \U$25390 ( \34372 , \34365 , \34371 );
buf \U$25391 ( \34373 , \34372 );
xor \U$25392 ( \34374 , \34326 , \34373 );
and \U$25393 ( \34375 , \33703 , \33709 );
and \U$25394 ( \34376 , \33703 , \33716 );
and \U$25395 ( \34377 , \33709 , \33716 );
or \U$25396 ( \34378 , \34375 , \34376 , \34377 );
buf \U$25397 ( \34379 , \34378 );
xor \U$25398 ( \34380 , \34374 , \34379 );
buf \U$25399 ( \34381 , \34380 );
xor \U$25400 ( \34382 , \34307 , \34381 );
buf \U$25401 ( \34383 , \34382 );
xor \U$25402 ( \34384 , \34080 , \34383 );
and \U$25403 ( \34385 , \33697 , \33718 );
and \U$25404 ( \34386 , \33697 , \33811 );
and \U$25405 ( \34387 , \33718 , \33811 );
or \U$25406 ( \34388 , \34385 , \34386 , \34387 );
buf \U$25407 ( \34389 , \34388 );
and \U$25408 ( \34390 , \34048 , \34053 );
and \U$25409 ( \34391 , \34048 , \34059 );
and \U$25410 ( \34392 , \34053 , \34059 );
or \U$25411 ( \34393 , \34390 , \34391 , \34392 );
buf \U$25412 ( \34394 , \34393 );
xor \U$25413 ( \34395 , \34389 , \34394 );
and \U$25414 ( \34396 , \33875 , \33880 );
and \U$25415 ( \34397 , \33875 , \34046 );
and \U$25416 ( \34398 , \33880 , \34046 );
or \U$25417 ( \34399 , \34396 , \34397 , \34398 );
buf \U$25418 ( \34400 , \34399 );
and \U$25419 ( \34401 , \33729 , \33750 );
and \U$25420 ( \34402 , \33729 , \33757 );
and \U$25421 ( \34403 , \33750 , \33757 );
or \U$25422 ( \34404 , \34401 , \34402 , \34403 );
buf \U$25423 ( \34405 , \34404 );
and \U$25424 ( \34406 , \20155 , \22129_nG9bd8 );
and \U$25425 ( \34407 , \20152 , \22629_nG9bd5 );
or \U$25426 ( \34408 , \34406 , \34407 );
xor \U$25427 ( \34409 , \20151 , \34408 );
buf \U$25428 ( \34410 , \34409 );
buf \U$25430 ( \34411 , \34410 );
xor \U$25431 ( \34412 , \34405 , \34411 );
and \U$25432 ( \34413 , \18702 , \23696_nG9bd2 );
and \U$25433 ( \34414 , \18699 , \24226_nG9bcf );
or \U$25434 ( \34415 , \34413 , \34414 );
xor \U$25435 ( \34416 , \18698 , \34415 );
buf \U$25436 ( \34417 , \34416 );
buf \U$25438 ( \34418 , \34417 );
xor \U$25439 ( \34419 , \34412 , \34418 );
buf \U$25440 ( \34420 , \34419 );
and \U$25441 ( \34421 , \12157 , \32179_nG9bb4 );
and \U$25442 ( \34422 , \12154 , \32888_nG9bb1 );
or \U$25443 ( \34423 , \34421 , \34422 );
xor \U$25444 ( \34424 , \12153 , \34423 );
buf \U$25445 ( \34425 , \34424 );
buf \U$25447 ( \34426 , \34425 );
xor \U$25448 ( \34427 , \34420 , \34426 );
and \U$25449 ( \34428 , \10421 , \33181_nG9bae );
and \U$25450 ( \34429 , \10418 , \33613_nG9bab );
or \U$25451 ( \34430 , \34428 , \34429 );
xor \U$25452 ( \34431 , \10417 , \34430 );
buf \U$25453 ( \34432 , \34431 );
buf \U$25455 ( \34433 , \34432 );
xor \U$25456 ( \34434 , \34427 , \34433 );
buf \U$25457 ( \34435 , \34434 );
xor \U$25458 ( \34436 , \34400 , \34435 );
and \U$25459 ( \34437 , \33768 , \33802 );
and \U$25460 ( \34438 , \33768 , \33809 );
and \U$25461 ( \34439 , \33802 , \33809 );
or \U$25462 ( \34440 , \34437 , \34438 , \34439 );
buf \U$25463 ( \34441 , \34440 );
xor \U$25464 ( \34442 , \34436 , \34441 );
buf \U$25465 ( \34443 , \34442 );
xor \U$25466 ( \34444 , \34395 , \34443 );
buf \U$25467 ( \34445 , \34444 );
xor \U$25468 ( \34446 , \34384 , \34445 );
and \U$25469 ( \34447 , \34075 , \34446 );
and \U$25471 ( \34448 , \34069 , \34074 );
or \U$25473 ( \34449 , 1'b0 , \34448 , 1'b0 );
xor \U$25474 ( \34450 , \34447 , \34449 );
and \U$25475 ( \34451 , \34065 , \34067 );
or \U$25478 ( \34452 , \34451 , 1'b0 , 1'b0 );
xor \U$25479 ( \34453 , \34450 , \34452 );
xor \U$25486 ( \34454 , \34453 , 1'b0 );
and \U$25487 ( \34455 , \34080 , \34383 );
and \U$25488 ( \34456 , \34080 , \34445 );
and \U$25489 ( \34457 , \34383 , \34445 );
or \U$25490 ( \34458 , \34455 , \34456 , \34457 );
xor \U$25491 ( \34459 , \34454 , \34458 );
and \U$25492 ( \34460 , \34301 , \34306 );
and \U$25493 ( \34461 , \34301 , \34381 );
and \U$25494 ( \34462 , \34306 , \34381 );
or \U$25495 ( \34463 , \34460 , \34461 , \34462 );
buf \U$25496 ( \34464 , \34463 );
and \U$25497 ( \34465 , \34085 , \34109 );
and \U$25498 ( \34466 , \34085 , \34116 );
and \U$25499 ( \34467 , \34109 , \34116 );
or \U$25500 ( \34468 , \34465 , \34466 , \34467 );
buf \U$25501 ( \34469 , \34468 );
and \U$25502 ( \34470 , \20155 , \22629_nG9bd5 );
and \U$25503 ( \34471 , \20152 , \23696_nG9bd2 );
or \U$25504 ( \34472 , \34470 , \34471 );
xor \U$25505 ( \34473 , \20151 , \34472 );
buf \U$25506 ( \34474 , \34473 );
buf \U$25508 ( \34475 , \34474 );
xor \U$25509 ( \34476 , \34469 , \34475 );
and \U$25510 ( \34477 , \18702 , \24226_nG9bcf );
and \U$25511 ( \34478 , \18699 , \25298_nG9bcc );
or \U$25512 ( \34479 , \34477 , \34478 );
xor \U$25513 ( \34480 , \18698 , \34479 );
buf \U$25514 ( \34481 , \34480 );
buf \U$25516 ( \34482 , \34481 );
xor \U$25517 ( \34483 , \34476 , \34482 );
buf \U$25518 ( \34484 , \34483 );
and \U$25519 ( \34485 , \12157 , \32888_nG9bb1 );
and \U$25520 ( \34486 , \12154 , \33181_nG9bae );
or \U$25521 ( \34487 , \34485 , \34486 );
xor \U$25522 ( \34488 , \12153 , \34487 );
buf \U$25523 ( \34489 , \34488 );
buf \U$25525 ( \34490 , \34489 );
xor \U$25526 ( \34491 , \34484 , \34490 );
and \U$25527 ( \34492 , \10707 , \34294_nG9ba5 );
and \U$25528 ( \34493 , \34186 , \34190 );
and \U$25529 ( \34494 , \34190 , \34286 );
and \U$25530 ( \34495 , \34186 , \34286 );
or \U$25531 ( \34496 , \34493 , \34494 , \34495 );
and \U$25532 ( \34497 , \34160 , \34164 );
and \U$25533 ( \34498 , \34164 , \34179 );
and \U$25534 ( \34499 , \34160 , \34179 );
or \U$25535 ( \34500 , \34497 , \34498 , \34499 );
and \U$25536 ( \34501 , \34169 , \34173 );
and \U$25537 ( \34502 , \34173 , \34178 );
and \U$25538 ( \34503 , \34169 , \34178 );
or \U$25539 ( \34504 , \34501 , \34502 , \34503 );
and \U$25540 ( \34505 , \34277 , \34278 );
and \U$25541 ( \34506 , \34278 , \34283 );
and \U$25542 ( \34507 , \34277 , \34283 );
or \U$25543 ( \34508 , \34505 , \34506 , \34507 );
xor \U$25544 ( \34509 , \34504 , \34508 );
and \U$25545 ( \34510 , \32794 , \12790 );
not \U$25546 ( \34511 , \34510 );
xnor \U$25547 ( \34512 , \34511 , \12780 );
not \U$25548 ( \34513 , \34512 );
and \U$25549 ( \34514 , \12769 , \32854 );
and \U$25550 ( \34515 , \13679 , \32067 );
nor \U$25551 ( \34516 , \34514 , \34515 );
xnor \U$25552 ( \34517 , \34516 , \32805 );
xor \U$25553 ( \34518 , \34513 , \34517 );
and \U$25554 ( \34519 , \12448 , \32802 );
xor \U$25555 ( \34520 , \34518 , \34519 );
xor \U$25556 ( \34521 , \34509 , \34520 );
xor \U$25557 ( \34522 , \34500 , \34521 );
and \U$25558 ( \34523 , \34239 , \34250 );
and \U$25559 ( \34524 , \34250 , \34262 );
and \U$25560 ( \34525 , \34239 , \34262 );
or \U$25561 ( \34526 , \34523 , \34524 , \34525 );
and \U$25562 ( \34527 , \34240 , \34244 );
and \U$25563 ( \34528 , \34244 , \34249 );
and \U$25564 ( \34529 , \34240 , \34249 );
or \U$25565 ( \34530 , \34527 , \34528 , \34529 );
and \U$25566 ( \34531 , \34255 , \34259 );
and \U$25567 ( \34532 , \34259 , \34261 );
and \U$25568 ( \34533 , \34255 , \34261 );
or \U$25569 ( \34534 , \34531 , \34532 , \34533 );
xor \U$25570 ( \34535 , \34530 , \34534 );
and \U$25571 ( \34536 , \34209 , \34213 );
and \U$25572 ( \34537 , \34213 , \34218 );
and \U$25573 ( \34538 , \34209 , \34218 );
or \U$25574 ( \34539 , \34536 , \34537 , \34538 );
xor \U$25575 ( \34540 , \34535 , \34539 );
xor \U$25576 ( \34541 , \34526 , \34540 );
and \U$25577 ( \34542 , \34195 , \34199 );
and \U$25578 ( \34543 , \34199 , \34204 );
and \U$25579 ( \34544 , \34195 , \34204 );
or \U$25580 ( \34545 , \34542 , \34543 , \34544 );
and \U$25581 ( \34546 , \34224 , \34228 );
and \U$25582 ( \34547 , \34228 , \34233 );
and \U$25583 ( \34548 , \34224 , \34233 );
or \U$25584 ( \34549 , \34546 , \34547 , \34548 );
xor \U$25585 ( \34550 , \34545 , \34549 );
and \U$25586 ( \34551 , \30802 , \14054 );
and \U$25587 ( \34552 , \32054 , \13692 );
nor \U$25588 ( \34553 , \34551 , \34552 );
xnor \U$25589 ( \34554 , \34553 , \14035 );
and \U$25590 ( \34555 , \27313 , \16635 );
and \U$25591 ( \34556 , \28534 , \16301 );
nor \U$25592 ( \34557 , \34555 , \34556 );
xnor \U$25593 ( \34558 , \34557 , \16625 );
xor \U$25594 ( \34559 , \34554 , \34558 );
and \U$25595 ( \34560 , \21033 , \22542 );
and \U$25596 ( \34561 , \22090 , \22103 );
nor \U$25597 ( \34562 , \34560 , \34561 );
xnor \U$25598 ( \34563 , \34562 , \22548 );
xor \U$25599 ( \34564 , \34559 , \34563 );
xor \U$25600 ( \34565 , \34550 , \34564 );
xor \U$25601 ( \34566 , \34541 , \34565 );
xor \U$25602 ( \34567 , \34522 , \34566 );
xor \U$25603 ( \34568 , \34496 , \34567 );
and \U$25604 ( \34569 , \34151 , \34155 );
and \U$25605 ( \34570 , \34155 , \34180 );
and \U$25606 ( \34571 , \34151 , \34180 );
or \U$25607 ( \34572 , \34569 , \34570 , \34571 );
and \U$25608 ( \34573 , \34235 , \34263 );
and \U$25609 ( \34574 , \34263 , \34285 );
and \U$25610 ( \34575 , \34235 , \34285 );
or \U$25611 ( \34576 , \34573 , \34574 , \34575 );
xor \U$25612 ( \34577 , \34572 , \34576 );
and \U$25613 ( \34578 , \34205 , \34219 );
and \U$25614 ( \34579 , \34219 , \34234 );
and \U$25615 ( \34580 , \34205 , \34234 );
or \U$25616 ( \34581 , \34578 , \34579 , \34580 );
and \U$25617 ( \34582 , \34268 , \34272 );
and \U$25618 ( \34583 , \34272 , \34284 );
and \U$25619 ( \34584 , \34268 , \34284 );
or \U$25620 ( \34585 , \34582 , \34583 , \34584 );
xor \U$25621 ( \34586 , \34581 , \34585 );
and \U$25622 ( \34587 , \22556 , \21005 );
and \U$25623 ( \34588 , \23617 , \20557 );
nor \U$25624 ( \34589 , \34587 , \34588 );
xnor \U$25625 ( \34590 , \34589 , \21011 );
and \U$25626 ( \34591 , \15321 , \29070 );
and \U$25627 ( \34592 , \16267 , \28526 );
nor \U$25628 ( \34593 , \34591 , \34592 );
xnor \U$25629 ( \34594 , \34593 , \29076 );
xor \U$25630 ( \34595 , \34590 , \34594 );
and \U$25631 ( \34596 , \14024 , \30823 );
and \U$25632 ( \34597 , \14950 , \30246 );
nor \U$25633 ( \34598 , \34596 , \34597 );
xnor \U$25634 ( \34599 , \34598 , \30813 );
xor \U$25635 ( \34600 , \34595 , \34599 );
and \U$25636 ( \34601 , \25815 , \18090 );
and \U$25637 ( \34602 , \26829 , \17655 );
nor \U$25638 ( \34603 , \34601 , \34602 );
xnor \U$25639 ( \34604 , \34603 , \18046 );
and \U$25640 ( \34605 , \19558 , \24138 );
and \U$25641 ( \34606 , \20544 , \23630 );
nor \U$25642 ( \34607 , \34605 , \34606 );
xnor \U$25643 ( \34608 , \34607 , \24144 );
xor \U$25644 ( \34609 , \34604 , \34608 );
and \U$25645 ( \34610 , \18035 , \25826 );
and \U$25646 ( \34611 , \19032 , \25264 );
nor \U$25647 ( \34612 , \34610 , \34611 );
xnor \U$25648 ( \34613 , \34612 , \25773 );
xor \U$25649 ( \34614 , \34609 , \34613 );
xor \U$25650 ( \34615 , \34600 , \34614 );
and \U$25651 ( \34616 , \29084 , \15336 );
and \U$25652 ( \34617 , \30268 , \14963 );
nor \U$25653 ( \34618 , \34616 , \34617 );
xnor \U$25654 ( \34619 , \34618 , \15342 );
and \U$25655 ( \34620 , \24199 , \19534 );
and \U$25656 ( \34621 , \25272 , \19045 );
nor \U$25657 ( \34622 , \34620 , \34621 );
xnor \U$25658 ( \34623 , \34622 , \19540 );
xor \U$25659 ( \34624 , \34619 , \34623 );
and \U$25660 ( \34625 , \16655 , \27397 );
and \U$25661 ( \34626 , \17627 , \26807 );
nor \U$25662 ( \34627 , \34625 , \34626 );
xnor \U$25663 ( \34628 , \34627 , \27295 );
xor \U$25664 ( \34629 , \34624 , \34628 );
xor \U$25665 ( \34630 , \34615 , \34629 );
xor \U$25666 ( \34631 , \34586 , \34630 );
xor \U$25667 ( \34632 , \34577 , \34631 );
xor \U$25668 ( \34633 , \34568 , \34632 );
and \U$25669 ( \34634 , \34147 , \34181 );
and \U$25670 ( \34635 , \34181 , \34287 );
and \U$25671 ( \34636 , \34147 , \34287 );
or \U$25672 ( \34637 , \34634 , \34635 , \34636 );
xor \U$25673 ( \34638 , \34633 , \34637 );
and \U$25674 ( \34639 , \34143 , \34288 );
and \U$25675 ( \34640 , \34289 , \34292 );
or \U$25676 ( \34641 , \34639 , \34640 );
xor \U$25677 ( \34642 , \34638 , \34641 );
buf g9ba2 ( \34643_nG9ba2 , \34642 );
and \U$25678 ( \34644 , \10704 , \34643_nG9ba2 );
or \U$25679 ( \34645 , \34492 , \34644 );
xor \U$25680 ( \34646 , \10703 , \34645 );
buf \U$25681 ( \34647 , \34646 );
buf \U$25683 ( \34648 , \34647 );
xor \U$25684 ( \34649 , \34491 , \34648 );
buf \U$25685 ( \34650 , \34649 );
and \U$25686 ( \34651 , \34132 , \34137 );
and \U$25687 ( \34652 , \34132 , \34299 );
and \U$25688 ( \34653 , \34137 , \34299 );
or \U$25689 ( \34654 , \34651 , \34652 , \34653 );
buf \U$25690 ( \34655 , \34654 );
xor \U$25691 ( \34656 , \34650 , \34655 );
and \U$25692 ( \34657 , \34405 , \34411 );
and \U$25693 ( \34658 , \34405 , \34418 );
and \U$25694 ( \34659 , \34411 , \34418 );
or \U$25695 ( \34660 , \34657 , \34658 , \34659 );
buf \U$25696 ( \34661 , \34660 );
and \U$25697 ( \34662 , \13370 , \30940_nG9bb7 );
and \U$25698 ( \34663 , \13367 , \32179_nG9bb4 );
or \U$25699 ( \34664 , \34662 , \34663 );
xor \U$25700 ( \34665 , \13366 , \34664 );
buf \U$25701 ( \34666 , \34665 );
buf \U$25703 ( \34667 , \34666 );
xor \U$25704 ( \34668 , \34661 , \34667 );
and \U$25705 ( \34669 , \10421 , \33613_nG9bab );
and \U$25706 ( \34670 , \10418 , \34041_nG9ba8 );
or \U$25707 ( \34671 , \34669 , \34670 );
xor \U$25708 ( \34672 , \10417 , \34671 );
buf \U$25709 ( \34673 , \34672 );
buf \U$25711 ( \34674 , \34673 );
xor \U$25712 ( \34675 , \34668 , \34674 );
buf \U$25713 ( \34676 , \34675 );
xor \U$25714 ( \34677 , \34656 , \34676 );
buf \U$25715 ( \34678 , \34677 );
xor \U$25716 ( \34679 , \34464 , \34678 );
and \U$25717 ( \34680 , \34400 , \34435 );
and \U$25718 ( \34681 , \34400 , \34441 );
and \U$25719 ( \34682 , \34435 , \34441 );
or \U$25720 ( \34683 , \34680 , \34681 , \34682 );
buf \U$25721 ( \34684 , \34683 );
xor \U$25722 ( \34685 , \34679 , \34684 );
buf \U$25723 ( \34686 , \34685 );
and \U$25724 ( \34687 , \34389 , \34394 );
and \U$25725 ( \34688 , \34389 , \34443 );
and \U$25726 ( \34689 , \34394 , \34443 );
or \U$25727 ( \34690 , \34687 , \34688 , \34689 );
buf \U$25728 ( \34691 , \34690 );
xor \U$25729 ( \34692 , \34686 , \34691 );
and \U$25730 ( \34693 , \34420 , \34426 );
and \U$25731 ( \34694 , \34420 , \34433 );
and \U$25732 ( \34695 , \34426 , \34433 );
or \U$25733 ( \34696 , \34693 , \34694 , \34695 );
buf \U$25734 ( \34697 , \34696 );
and \U$25735 ( \34698 , \34312 , \34317 );
and \U$25736 ( \34699 , \34312 , \34324 );
and \U$25737 ( \34700 , \34317 , \34324 );
or \U$25738 ( \34701 , \34698 , \34699 , \34700 );
buf \U$25739 ( \34702 , \34701 );
xor \U$25740 ( \34703 , \34697 , \34702 );
and \U$25741 ( \34704 , \34358 , \34364 );
and \U$25742 ( \34705 , \34358 , \34371 );
and \U$25743 ( \34706 , \34364 , \34371 );
or \U$25744 ( \34707 , \34704 , \34705 , \34706 );
buf \U$25745 ( \34708 , \34707 );
xor \U$25746 ( \34709 , \34703 , \34708 );
buf \U$25747 ( \34710 , \34709 );
and \U$25748 ( \34711 , \34326 , \34373 );
and \U$25749 ( \34712 , \34326 , \34379 );
and \U$25750 ( \34713 , \34373 , \34379 );
or \U$25751 ( \34714 , \34711 , \34712 , \34713 );
buf \U$25752 ( \34715 , \34714 );
xor \U$25753 ( \34716 , \34710 , \34715 );
and \U$25754 ( \34717 , \34098 , \34100 );
and \U$25755 ( \34718 , \34098 , \34107 );
and \U$25756 ( \34719 , \34100 , \34107 );
or \U$25757 ( \34720 , \34717 , \34718 , \34719 );
buf \U$25758 ( \34721 , \34720 );
and \U$25759 ( \34722 , \28118 , \15373_nG9bf3 );
and \U$25760 ( \34723 , \28115 , \16315_nG9bf0 );
or \U$25761 ( \34724 , \34722 , \34723 );
xor \U$25762 ( \34725 , \28114 , \34724 );
buf \U$25763 ( \34726 , \34725 );
buf \U$25765 ( \34727 , \34726 );
xor \U$25766 ( \34728 , \34721 , \34727 );
and \U$25767 ( \34729 , \26431 , \16680_nG9bed );
and \U$25768 ( \34730 , \26428 , \17665_nG9bea );
or \U$25769 ( \34731 , \34729 , \34730 );
xor \U$25770 ( \34732 , \26427 , \34731 );
buf \U$25771 ( \34733 , \34732 );
buf \U$25773 ( \34734 , \34733 );
xor \U$25774 ( \34735 , \34728 , \34734 );
buf \U$25775 ( \34736 , \34735 );
and \U$25776 ( \34737 , \34328 , \34334 );
and \U$25777 ( \34738 , \34328 , \34341 );
and \U$25778 ( \34739 , \34334 , \34341 );
or \U$25779 ( \34740 , \34737 , \34738 , \34739 );
buf \U$25780 ( \34741 , \34740 );
xor \U$25781 ( \34742 , \34736 , \34741 );
and \U$25782 ( \34743 , \21658 , \21086_nG9bdb );
and \U$25783 ( \34744 , \21655 , \22129_nG9bd8 );
or \U$25784 ( \34745 , \34743 , \34744 );
xor \U$25785 ( \34746 , \21654 , \34745 );
buf \U$25786 ( \34747 , \34746 );
buf \U$25788 ( \34748 , \34747 );
xor \U$25789 ( \34749 , \34742 , \34748 );
buf \U$25790 ( \34750 , \34749 );
and \U$25791 ( \34751 , \17297 , \25860_nG9bc9 );
and \U$25792 ( \34752 , \17294 , \26887_nG9bc6 );
or \U$25793 ( \34753 , \34751 , \34752 );
xor \U$25794 ( \34754 , \17293 , \34753 );
buf \U$25795 ( \34755 , \34754 );
buf \U$25797 ( \34756 , \34755 );
xor \U$25798 ( \34757 , \34750 , \34756 );
and \U$25799 ( \34758 , \14631 , \29179_nG9bbd );
and \U$25800 ( \34759 , \14628 , \30366_nG9bba );
or \U$25801 ( \34760 , \34758 , \34759 );
xor \U$25802 ( \34761 , \14627 , \34760 );
buf \U$25803 ( \34762 , \34761 );
buf \U$25805 ( \34763 , \34762 );
xor \U$25806 ( \34764 , \34757 , \34763 );
buf \U$25807 ( \34765 , \34764 );
and \U$25809 ( \34766 , \32916 , \12470_nG9c02 );
or \U$25810 ( \34767 , 1'b0 , \34766 );
xor \U$25811 ( \34768 , 1'b0 , \34767 );
buf \U$25812 ( \34769 , \34768 );
buf \U$25814 ( \34770 , \34769 );
and \U$25815 ( \34771 , \31636 , \12801_nG9bff );
and \U$25816 ( \34772 , \31633 , \13705_nG9bfc );
or \U$25817 ( \34773 , \34771 , \34772 );
xor \U$25818 ( \34774 , \31632 , \34773 );
buf \U$25819 ( \34775 , \34774 );
buf \U$25821 ( \34776 , \34775 );
xor \U$25822 ( \34777 , \34770 , \34776 );
buf \U$25823 ( \34778 , \34777 );
and \U$25824 ( \34779 , \34090 , \34096 );
buf \U$25825 ( \34780 , \34779 );
xor \U$25826 ( \34781 , \34778 , \34780 );
and \U$25827 ( \34782 , \29853 , \14070_nG9bf9 );
and \U$25828 ( \34783 , \29850 , \14984_nG9bf6 );
or \U$25829 ( \34784 , \34782 , \34783 );
xor \U$25830 ( \34785 , \29849 , \34784 );
buf \U$25831 ( \34786 , \34785 );
buf \U$25833 ( \34787 , \34786 );
xor \U$25834 ( \34788 , \34781 , \34787 );
buf \U$25835 ( \34789 , \34788 );
and \U$25836 ( \34790 , \24792 , \18107_nG9be7 );
and \U$25837 ( \34791 , \24789 , \19091_nG9be4 );
or \U$25838 ( \34792 , \34790 , \34791 );
xor \U$25839 ( \34793 , \24788 , \34792 );
buf \U$25840 ( \34794 , \34793 );
buf \U$25842 ( \34795 , \34794 );
xor \U$25843 ( \34796 , \34789 , \34795 );
and \U$25844 ( \34797 , \23201 , \19586_nG9be1 );
and \U$25845 ( \34798 , \23198 , \20608_nG9bde );
or \U$25846 ( \34799 , \34797 , \34798 );
xor \U$25847 ( \34800 , \23197 , \34799 );
buf \U$25848 ( \34801 , \34800 );
buf \U$25850 ( \34802 , \34801 );
xor \U$25851 ( \34803 , \34796 , \34802 );
buf \U$25852 ( \34804 , \34803 );
and \U$25853 ( \34805 , \34343 , \34349 );
and \U$25854 ( \34806 , \34343 , \34356 );
and \U$25855 ( \34807 , \34349 , \34356 );
or \U$25856 ( \34808 , \34805 , \34806 , \34807 );
buf \U$25857 ( \34809 , \34808 );
xor \U$25858 ( \34810 , \34804 , \34809 );
and \U$25859 ( \34811 , \15940 , \27416_nG9bc3 );
and \U$25860 ( \34812 , \15937 , \28602_nG9bc0 );
or \U$25861 ( \34813 , \34811 , \34812 );
xor \U$25862 ( \34814 , \15936 , \34813 );
buf \U$25863 ( \34815 , \34814 );
buf \U$25865 ( \34816 , \34815 );
xor \U$25866 ( \34817 , \34810 , \34816 );
buf \U$25867 ( \34818 , \34817 );
xor \U$25868 ( \34819 , \34765 , \34818 );
and \U$25869 ( \34820 , \34118 , \34123 );
and \U$25870 ( \34821 , \34118 , \34130 );
and \U$25871 ( \34822 , \34123 , \34130 );
or \U$25872 ( \34823 , \34820 , \34821 , \34822 );
buf \U$25873 ( \34824 , \34823 );
xor \U$25874 ( \34825 , \34819 , \34824 );
buf \U$25875 ( \34826 , \34825 );
xor \U$25876 ( \34827 , \34716 , \34826 );
buf \U$25877 ( \34828 , \34827 );
xor \U$25878 ( \34829 , \34692 , \34828 );
and \U$25879 ( \34830 , \34459 , \34829 );
and \U$25881 ( \34831 , \34453 , \34458 );
or \U$25883 ( \34832 , 1'b0 , \34831 , 1'b0 );
xor \U$25884 ( \34833 , \34830 , \34832 );
and \U$25886 ( \34834 , \34447 , \34452 );
or \U$25888 ( \34835 , 1'b0 , \34834 , 1'b0 );
xor \U$25889 ( \34836 , \34833 , \34835 );
xor \U$25896 ( \34837 , \34836 , 1'b0 );
and \U$25897 ( \34838 , \34686 , \34691 );
and \U$25898 ( \34839 , \34686 , \34828 );
and \U$25899 ( \34840 , \34691 , \34828 );
or \U$25900 ( \34841 , \34838 , \34839 , \34840 );
xor \U$25901 ( \34842 , \34837 , \34841 );
and \U$25902 ( \34843 , \34650 , \34655 );
and \U$25903 ( \34844 , \34650 , \34676 );
and \U$25904 ( \34845 , \34655 , \34676 );
or \U$25905 ( \34846 , \34843 , \34844 , \34845 );
buf \U$25906 ( \34847 , \34846 );
and \U$25907 ( \34848 , \34697 , \34702 );
and \U$25908 ( \34849 , \34697 , \34708 );
and \U$25909 ( \34850 , \34702 , \34708 );
or \U$25910 ( \34851 , \34848 , \34849 , \34850 );
buf \U$25911 ( \34852 , \34851 );
xor \U$25912 ( \34853 , \34847 , \34852 );
and \U$25913 ( \34854 , \34750 , \34756 );
and \U$25914 ( \34855 , \34750 , \34763 );
and \U$25915 ( \34856 , \34756 , \34763 );
or \U$25916 ( \34857 , \34854 , \34855 , \34856 );
buf \U$25917 ( \34858 , \34857 );
and \U$25918 ( \34859 , \34804 , \34809 );
and \U$25919 ( \34860 , \34804 , \34816 );
and \U$25920 ( \34861 , \34809 , \34816 );
or \U$25921 ( \34862 , \34859 , \34860 , \34861 );
buf \U$25922 ( \34863 , \34862 );
xor \U$25923 ( \34864 , \34858 , \34863 );
and \U$25924 ( \34865 , \34736 , \34741 );
and \U$25925 ( \34866 , \34736 , \34748 );
and \U$25926 ( \34867 , \34741 , \34748 );
or \U$25927 ( \34868 , \34865 , \34866 , \34867 );
buf \U$25928 ( \34869 , \34868 );
and \U$25930 ( \34870 , \32916 , \12801_nG9bff );
or \U$25931 ( \34871 , 1'b0 , \34870 );
xor \U$25932 ( \34872 , 1'b0 , \34871 );
buf \U$25933 ( \34873 , \34872 );
buf \U$25935 ( \34874 , \34873 );
and \U$25936 ( \34875 , \31636 , \13705_nG9bfc );
and \U$25937 ( \34876 , \31633 , \14070_nG9bf9 );
or \U$25938 ( \34877 , \34875 , \34876 );
xor \U$25939 ( \34878 , \31632 , \34877 );
buf \U$25940 ( \34879 , \34878 );
buf \U$25942 ( \34880 , \34879 );
xor \U$25943 ( \34881 , \34874 , \34880 );
buf \U$25944 ( \34882 , \34881 );
and \U$25945 ( \34883 , \34770 , \34776 );
buf \U$25946 ( \34884 , \34883 );
xor \U$25947 ( \34885 , \34882 , \34884 );
and \U$25948 ( \34886 , \29853 , \14984_nG9bf6 );
and \U$25949 ( \34887 , \29850 , \15373_nG9bf3 );
or \U$25950 ( \34888 , \34886 , \34887 );
xor \U$25951 ( \34889 , \29849 , \34888 );
buf \U$25952 ( \34890 , \34889 );
buf \U$25954 ( \34891 , \34890 );
xor \U$25955 ( \34892 , \34885 , \34891 );
buf \U$25956 ( \34893 , \34892 );
and \U$25957 ( \34894 , \24792 , \19091_nG9be4 );
and \U$25958 ( \34895 , \24789 , \19586_nG9be1 );
or \U$25959 ( \34896 , \34894 , \34895 );
xor \U$25960 ( \34897 , \24788 , \34896 );
buf \U$25961 ( \34898 , \34897 );
buf \U$25963 ( \34899 , \34898 );
xor \U$25964 ( \34900 , \34893 , \34899 );
and \U$25965 ( \34901 , \23201 , \20608_nG9bde );
and \U$25966 ( \34902 , \23198 , \21086_nG9bdb );
or \U$25967 ( \34903 , \34901 , \34902 );
xor \U$25968 ( \34904 , \23197 , \34903 );
buf \U$25969 ( \34905 , \34904 );
buf \U$25971 ( \34906 , \34905 );
xor \U$25972 ( \34907 , \34900 , \34906 );
buf \U$25973 ( \34908 , \34907 );
xor \U$25974 ( \34909 , \34869 , \34908 );
and \U$25975 ( \34910 , \17297 , \26887_nG9bc6 );
and \U$25976 ( \34911 , \17294 , \27416_nG9bc3 );
or \U$25977 ( \34912 , \34910 , \34911 );
xor \U$25978 ( \34913 , \17293 , \34912 );
buf \U$25979 ( \34914 , \34913 );
buf \U$25981 ( \34915 , \34914 );
xor \U$25982 ( \34916 , \34909 , \34915 );
buf \U$25983 ( \34917 , \34916 );
xor \U$25984 ( \34918 , \34864 , \34917 );
buf \U$25985 ( \34919 , \34918 );
xor \U$25986 ( \34920 , \34853 , \34919 );
buf \U$25987 ( \34921 , \34920 );
and \U$25988 ( \34922 , \34789 , \34795 );
and \U$25989 ( \34923 , \34789 , \34802 );
and \U$25990 ( \34924 , \34795 , \34802 );
or \U$25991 ( \34925 , \34922 , \34923 , \34924 );
buf \U$25992 ( \34926 , \34925 );
and \U$25993 ( \34927 , \20155 , \23696_nG9bd2 );
and \U$25994 ( \34928 , \20152 , \24226_nG9bcf );
or \U$25995 ( \34929 , \34927 , \34928 );
xor \U$25996 ( \34930 , \20151 , \34929 );
buf \U$25997 ( \34931 , \34930 );
buf \U$25999 ( \34932 , \34931 );
xor \U$26000 ( \34933 , \34926 , \34932 );
and \U$26001 ( \34934 , \18702 , \25298_nG9bcc );
and \U$26002 ( \34935 , \18699 , \25860_nG9bc9 );
or \U$26003 ( \34936 , \34934 , \34935 );
xor \U$26004 ( \34937 , \18698 , \34936 );
buf \U$26005 ( \34938 , \34937 );
buf \U$26007 ( \34939 , \34938 );
xor \U$26008 ( \34940 , \34933 , \34939 );
buf \U$26009 ( \34941 , \34940 );
and \U$26010 ( \34942 , \10421 , \34041_nG9ba8 );
and \U$26011 ( \34943 , \10418 , \34294_nG9ba5 );
or \U$26012 ( \34944 , \34942 , \34943 );
xor \U$26013 ( \34945 , \10417 , \34944 );
buf \U$26014 ( \34946 , \34945 );
buf \U$26016 ( \34947 , \34946 );
xor \U$26017 ( \34948 , \34941 , \34947 );
and \U$26018 ( \34949 , \10707 , \34643_nG9ba2 );
and \U$26019 ( \34950 , \34572 , \34576 );
and \U$26020 ( \34951 , \34576 , \34631 );
and \U$26021 ( \34952 , \34572 , \34631 );
or \U$26022 ( \34953 , \34950 , \34951 , \34952 );
and \U$26023 ( \34954 , \34504 , \34508 );
and \U$26024 ( \34955 , \34508 , \34520 );
and \U$26025 ( \34956 , \34504 , \34520 );
or \U$26026 ( \34957 , \34954 , \34955 , \34956 );
and \U$26027 ( \34958 , \34526 , \34540 );
and \U$26028 ( \34959 , \34540 , \34565 );
and \U$26029 ( \34960 , \34526 , \34565 );
or \U$26030 ( \34961 , \34958 , \34959 , \34960 );
xor \U$26031 ( \34962 , \34957 , \34961 );
and \U$26032 ( \34963 , \34545 , \34549 );
and \U$26033 ( \34964 , \34549 , \34564 );
and \U$26034 ( \34965 , \34545 , \34564 );
or \U$26035 ( \34966 , \34963 , \34964 , \34965 );
and \U$26036 ( \34967 , \34554 , \34558 );
and \U$26037 ( \34968 , \34558 , \34563 );
and \U$26038 ( \34969 , \34554 , \34563 );
or \U$26039 ( \34970 , \34967 , \34968 , \34969 );
and \U$26040 ( \34971 , \34604 , \34608 );
and \U$26041 ( \34972 , \34608 , \34613 );
and \U$26042 ( \34973 , \34604 , \34613 );
or \U$26043 ( \34974 , \34971 , \34972 , \34973 );
xor \U$26044 ( \34975 , \34970 , \34974 );
buf \U$26045 ( \34976 , \34512 );
xor \U$26046 ( \34977 , \34975 , \34976 );
xor \U$26047 ( \34978 , \34966 , \34977 );
and \U$26048 ( \34979 , \34590 , \34594 );
and \U$26049 ( \34980 , \34594 , \34599 );
and \U$26050 ( \34981 , \34590 , \34599 );
or \U$26051 ( \34982 , \34979 , \34980 , \34981 );
and \U$26052 ( \34983 , \34619 , \34623 );
and \U$26053 ( \34984 , \34623 , \34628 );
and \U$26054 ( \34985 , \34619 , \34628 );
or \U$26055 ( \34986 , \34983 , \34984 , \34985 );
xor \U$26056 ( \34987 , \34982 , \34986 );
and \U$26057 ( \34988 , \26829 , \18090 );
and \U$26058 ( \34989 , \27313 , \17655 );
nor \U$26059 ( \34990 , \34988 , \34989 );
xnor \U$26060 ( \34991 , \34990 , \18046 );
and \U$26061 ( \34992 , \22090 , \22542 );
and \U$26062 ( \34993 , \22556 , \22103 );
nor \U$26063 ( \34994 , \34992 , \34993 );
xnor \U$26064 ( \34995 , \34994 , \22548 );
xor \U$26065 ( \34996 , \34991 , \34995 );
and \U$26066 ( \34997 , \20544 , \24138 );
and \U$26067 ( \34998 , \21033 , \23630 );
nor \U$26068 ( \34999 , \34997 , \34998 );
xnor \U$26069 ( \35000 , \34999 , \24144 );
xor \U$26070 ( \35001 , \34996 , \35000 );
xor \U$26071 ( \35002 , \34987 , \35001 );
xor \U$26072 ( \35003 , \34978 , \35002 );
xor \U$26073 ( \35004 , \34962 , \35003 );
xor \U$26074 ( \35005 , \34953 , \35004 );
and \U$26075 ( \35006 , \34581 , \34585 );
and \U$26076 ( \35007 , \34585 , \34630 );
and \U$26077 ( \35008 , \34581 , \34630 );
or \U$26078 ( \35009 , \35006 , \35007 , \35008 );
and \U$26079 ( \35010 , \34500 , \34521 );
and \U$26080 ( \35011 , \34521 , \34566 );
and \U$26081 ( \35012 , \34500 , \34566 );
or \U$26082 ( \35013 , \35010 , \35011 , \35012 );
xor \U$26083 ( \35014 , \35009 , \35013 );
and \U$26084 ( \35015 , \34600 , \34614 );
and \U$26085 ( \35016 , \34614 , \34629 );
and \U$26086 ( \35017 , \34600 , \34629 );
or \U$26087 ( \35018 , \35015 , \35016 , \35017 );
not \U$26088 ( \35019 , \12780 );
and \U$26089 ( \35020 , \32054 , \14054 );
and \U$26090 ( \35021 , \32794 , \13692 );
nor \U$26091 ( \35022 , \35020 , \35021 );
xnor \U$26092 ( \35023 , \35022 , \14035 );
xor \U$26093 ( \35024 , \35019 , \35023 );
and \U$26094 ( \35025 , \28534 , \16635 );
and \U$26095 ( \35026 , \29084 , \16301 );
nor \U$26096 ( \35027 , \35025 , \35026 );
xnor \U$26097 ( \35028 , \35027 , \16625 );
xor \U$26098 ( \35029 , \35024 , \35028 );
and \U$26099 ( \35030 , \25272 , \19534 );
and \U$26100 ( \35031 , \25815 , \19045 );
nor \U$26101 ( \35032 , \35030 , \35031 );
xnor \U$26102 ( \35033 , \35032 , \19540 );
and \U$26103 ( \35034 , \16267 , \29070 );
and \U$26104 ( \35035 , \16655 , \28526 );
nor \U$26105 ( \35036 , \35034 , \35035 );
xnor \U$26106 ( \35037 , \35036 , \29076 );
xor \U$26107 ( \35038 , \35033 , \35037 );
and \U$26108 ( \35039 , \14950 , \30823 );
and \U$26109 ( \35040 , \15321 , \30246 );
nor \U$26110 ( \35041 , \35039 , \35040 );
xnor \U$26111 ( \35042 , \35041 , \30813 );
xor \U$26112 ( \35043 , \35038 , \35042 );
xor \U$26113 ( \35044 , \35029 , \35043 );
and \U$26114 ( \35045 , \23617 , \21005 );
and \U$26115 ( \35046 , \24199 , \20557 );
nor \U$26116 ( \35047 , \35045 , \35046 );
xnor \U$26117 ( \35048 , \35047 , \21011 );
and \U$26118 ( \35049 , \13679 , \32854 );
and \U$26119 ( \35050 , \14024 , \32067 );
nor \U$26120 ( \35051 , \35049 , \35050 );
xnor \U$26121 ( \35052 , \35051 , \32805 );
xor \U$26122 ( \35053 , \35048 , \35052 );
and \U$26123 ( \35054 , \12769 , \32802 );
xor \U$26124 ( \35055 , \35053 , \35054 );
xor \U$26125 ( \35056 , \35044 , \35055 );
xor \U$26126 ( \35057 , \35018 , \35056 );
and \U$26127 ( \35058 , \34530 , \34534 );
and \U$26128 ( \35059 , \34534 , \34539 );
and \U$26129 ( \35060 , \34530 , \34539 );
or \U$26130 ( \35061 , \35058 , \35059 , \35060 );
and \U$26131 ( \35062 , \34513 , \34517 );
and \U$26132 ( \35063 , \34517 , \34519 );
and \U$26133 ( \35064 , \34513 , \34519 );
or \U$26134 ( \35065 , \35062 , \35063 , \35064 );
xor \U$26135 ( \35066 , \35061 , \35065 );
and \U$26136 ( \35067 , \30268 , \15336 );
and \U$26137 ( \35068 , \30802 , \14963 );
nor \U$26138 ( \35069 , \35067 , \35068 );
xnor \U$26139 ( \35070 , \35069 , \15342 );
and \U$26140 ( \35071 , \19032 , \25826 );
and \U$26141 ( \35072 , \19558 , \25264 );
nor \U$26142 ( \35073 , \35071 , \35072 );
xnor \U$26143 ( \35074 , \35073 , \25773 );
xor \U$26144 ( \35075 , \35070 , \35074 );
and \U$26145 ( \35076 , \17627 , \27397 );
and \U$26146 ( \35077 , \18035 , \26807 );
nor \U$26147 ( \35078 , \35076 , \35077 );
xnor \U$26148 ( \35079 , \35078 , \27295 );
xor \U$26149 ( \35080 , \35075 , \35079 );
xor \U$26150 ( \35081 , \35066 , \35080 );
xor \U$26151 ( \35082 , \35057 , \35081 );
xor \U$26152 ( \35083 , \35014 , \35082 );
xor \U$26153 ( \35084 , \35005 , \35083 );
and \U$26154 ( \35085 , \34496 , \34567 );
and \U$26155 ( \35086 , \34567 , \34632 );
and \U$26156 ( \35087 , \34496 , \34632 );
or \U$26157 ( \35088 , \35085 , \35086 , \35087 );
xor \U$26158 ( \35089 , \35084 , \35088 );
and \U$26159 ( \35090 , \34633 , \34637 );
and \U$26160 ( \35091 , \34638 , \34641 );
or \U$26161 ( \35092 , \35090 , \35091 );
xor \U$26162 ( \35093 , \35089 , \35092 );
buf g9b9f ( \35094_nG9b9f , \35093 );
and \U$26163 ( \35095 , \10704 , \35094_nG9b9f );
or \U$26164 ( \35096 , \34949 , \35095 );
xor \U$26165 ( \35097 , \10703 , \35096 );
buf \U$26166 ( \35098 , \35097 );
buf \U$26168 ( \35099 , \35098 );
xor \U$26169 ( \35100 , \34948 , \35099 );
buf \U$26170 ( \35101 , \35100 );
and \U$26171 ( \35102 , \34765 , \34818 );
and \U$26172 ( \35103 , \34765 , \34824 );
and \U$26173 ( \35104 , \34818 , \34824 );
or \U$26174 ( \35105 , \35102 , \35103 , \35104 );
buf \U$26175 ( \35106 , \35105 );
xor \U$26176 ( \35107 , \35101 , \35106 );
and \U$26177 ( \35108 , \34469 , \34475 );
and \U$26178 ( \35109 , \34469 , \34482 );
and \U$26179 ( \35110 , \34475 , \34482 );
or \U$26180 ( \35111 , \35108 , \35109 , \35110 );
buf \U$26181 ( \35112 , \35111 );
and \U$26182 ( \35113 , \34721 , \34727 );
and \U$26183 ( \35114 , \34721 , \34734 );
and \U$26184 ( \35115 , \34727 , \34734 );
or \U$26185 ( \35116 , \35113 , \35114 , \35115 );
buf \U$26186 ( \35117 , \35116 );
and \U$26187 ( \35118 , \34778 , \34780 );
and \U$26188 ( \35119 , \34778 , \34787 );
and \U$26189 ( \35120 , \34780 , \34787 );
or \U$26190 ( \35121 , \35118 , \35119 , \35120 );
buf \U$26191 ( \35122 , \35121 );
and \U$26192 ( \35123 , \28118 , \16315_nG9bf0 );
and \U$26193 ( \35124 , \28115 , \16680_nG9bed );
or \U$26194 ( \35125 , \35123 , \35124 );
xor \U$26195 ( \35126 , \28114 , \35125 );
buf \U$26196 ( \35127 , \35126 );
buf \U$26198 ( \35128 , \35127 );
xor \U$26199 ( \35129 , \35122 , \35128 );
and \U$26200 ( \35130 , \26431 , \17665_nG9bea );
and \U$26201 ( \35131 , \26428 , \18107_nG9be7 );
or \U$26202 ( \35132 , \35130 , \35131 );
xor \U$26203 ( \35133 , \26427 , \35132 );
buf \U$26204 ( \35134 , \35133 );
buf \U$26206 ( \35135 , \35134 );
xor \U$26207 ( \35136 , \35129 , \35135 );
buf \U$26208 ( \35137 , \35136 );
xor \U$26209 ( \35138 , \35117 , \35137 );
and \U$26210 ( \35139 , \21658 , \22129_nG9bd8 );
and \U$26211 ( \35140 , \21655 , \22629_nG9bd5 );
or \U$26212 ( \35141 , \35139 , \35140 );
xor \U$26213 ( \35142 , \21654 , \35141 );
buf \U$26214 ( \35143 , \35142 );
buf \U$26216 ( \35144 , \35143 );
xor \U$26217 ( \35145 , \35138 , \35144 );
buf \U$26218 ( \35146 , \35145 );
xor \U$26219 ( \35147 , \35112 , \35146 );
and \U$26220 ( \35148 , \13370 , \32179_nG9bb4 );
and \U$26221 ( \35149 , \13367 , \32888_nG9bb1 );
or \U$26222 ( \35150 , \35148 , \35149 );
xor \U$26223 ( \35151 , \13366 , \35150 );
buf \U$26224 ( \35152 , \35151 );
buf \U$26226 ( \35153 , \35152 );
xor \U$26227 ( \35154 , \35147 , \35153 );
buf \U$26228 ( \35155 , \35154 );
xor \U$26229 ( \35156 , \35107 , \35155 );
buf \U$26230 ( \35157 , \35156 );
xor \U$26231 ( \35158 , \34921 , \35157 );
and \U$26232 ( \35159 , \34484 , \34490 );
and \U$26233 ( \35160 , \34484 , \34648 );
and \U$26234 ( \35161 , \34490 , \34648 );
or \U$26235 ( \35162 , \35159 , \35160 , \35161 );
buf \U$26236 ( \35163 , \35162 );
and \U$26237 ( \35164 , \34661 , \34667 );
and \U$26238 ( \35165 , \34661 , \34674 );
and \U$26239 ( \35166 , \34667 , \34674 );
or \U$26240 ( \35167 , \35164 , \35165 , \35166 );
buf \U$26241 ( \35168 , \35167 );
xor \U$26242 ( \35169 , \35163 , \35168 );
and \U$26243 ( \35170 , \15940 , \28602_nG9bc0 );
and \U$26244 ( \35171 , \15937 , \29179_nG9bbd );
or \U$26245 ( \35172 , \35170 , \35171 );
xor \U$26246 ( \35173 , \15936 , \35172 );
buf \U$26247 ( \35174 , \35173 );
buf \U$26249 ( \35175 , \35174 );
and \U$26250 ( \35176 , \14631 , \30366_nG9bba );
and \U$26251 ( \35177 , \14628 , \30940_nG9bb7 );
or \U$26252 ( \35178 , \35176 , \35177 );
xor \U$26253 ( \35179 , \14627 , \35178 );
buf \U$26254 ( \35180 , \35179 );
buf \U$26256 ( \35181 , \35180 );
xor \U$26257 ( \35182 , \35175 , \35181 );
and \U$26258 ( \35183 , \12157 , \33181_nG9bae );
and \U$26259 ( \35184 , \12154 , \33613_nG9bab );
or \U$26260 ( \35185 , \35183 , \35184 );
xor \U$26261 ( \35186 , \12153 , \35185 );
buf \U$26262 ( \35187 , \35186 );
buf \U$26264 ( \35188 , \35187 );
xor \U$26265 ( \35189 , \35182 , \35188 );
buf \U$26266 ( \35190 , \35189 );
xor \U$26267 ( \35191 , \35169 , \35190 );
buf \U$26268 ( \35192 , \35191 );
xor \U$26269 ( \35193 , \35158 , \35192 );
buf \U$26270 ( \35194 , \35193 );
and \U$26271 ( \35195 , \34464 , \34678 );
and \U$26272 ( \35196 , \34464 , \34684 );
and \U$26273 ( \35197 , \34678 , \34684 );
or \U$26274 ( \35198 , \35195 , \35196 , \35197 );
buf \U$26275 ( \35199 , \35198 );
xor \U$26276 ( \35200 , \35194 , \35199 );
and \U$26277 ( \35201 , \34710 , \34715 );
and \U$26278 ( \35202 , \34710 , \34826 );
and \U$26279 ( \35203 , \34715 , \34826 );
or \U$26280 ( \35204 , \35201 , \35202 , \35203 );
buf \U$26281 ( \35205 , \35204 );
xor \U$26282 ( \35206 , \35200 , \35205 );
and \U$26283 ( \35207 , \34842 , \35206 );
and \U$26285 ( \35208 , \34836 , \34841 );
or \U$26287 ( \35209 , 1'b0 , \35208 , 1'b0 );
xor \U$26288 ( \35210 , \35207 , \35209 );
and \U$26290 ( \35211 , \34830 , \34835 );
and \U$26291 ( \35212 , \34832 , \34835 );
or \U$26292 ( \35213 , 1'b0 , \35211 , \35212 );
xor \U$26293 ( \35214 , \35210 , \35213 );
xor \U$26300 ( \35215 , \35214 , 1'b0 );
and \U$26301 ( \35216 , \35194 , \35199 );
and \U$26302 ( \35217 , \35194 , \35205 );
and \U$26303 ( \35218 , \35199 , \35205 );
or \U$26304 ( \35219 , \35216 , \35217 , \35218 );
xor \U$26305 ( \35220 , \35215 , \35219 );
and \U$26306 ( \35221 , \34921 , \35157 );
and \U$26307 ( \35222 , \34921 , \35192 );
and \U$26308 ( \35223 , \35157 , \35192 );
or \U$26309 ( \35224 , \35221 , \35222 , \35223 );
buf \U$26310 ( \35225 , \35224 );
and \U$26311 ( \35226 , \34941 , \34947 );
and \U$26312 ( \35227 , \34941 , \35099 );
and \U$26313 ( \35228 , \34947 , \35099 );
or \U$26314 ( \35229 , \35226 , \35227 , \35228 );
buf \U$26315 ( \35230 , \35229 );
and \U$26316 ( \35231 , \34858 , \34863 );
and \U$26317 ( \35232 , \34858 , \34917 );
and \U$26318 ( \35233 , \34863 , \34917 );
or \U$26319 ( \35234 , \35231 , \35232 , \35233 );
buf \U$26320 ( \35235 , \35234 );
xor \U$26321 ( \35236 , \35230 , \35235 );
and \U$26322 ( \35237 , \34869 , \34908 );
and \U$26323 ( \35238 , \34869 , \34915 );
and \U$26324 ( \35239 , \34908 , \34915 );
or \U$26325 ( \35240 , \35237 , \35238 , \35239 );
buf \U$26326 ( \35241 , \35240 );
and \U$26327 ( \35242 , \34926 , \34932 );
and \U$26328 ( \35243 , \34926 , \34939 );
and \U$26329 ( \35244 , \34932 , \34939 );
or \U$26330 ( \35245 , \35242 , \35243 , \35244 );
buf \U$26331 ( \35246 , \35245 );
xor \U$26332 ( \35247 , \35241 , \35246 );
and \U$26333 ( \35248 , \34893 , \34899 );
and \U$26334 ( \35249 , \34893 , \34906 );
and \U$26335 ( \35250 , \34899 , \34906 );
or \U$26336 ( \35251 , \35248 , \35249 , \35250 );
buf \U$26337 ( \35252 , \35251 );
and \U$26338 ( \35253 , \34882 , \34884 );
and \U$26339 ( \35254 , \34882 , \34891 );
and \U$26340 ( \35255 , \34884 , \34891 );
or \U$26341 ( \35256 , \35253 , \35254 , \35255 );
buf \U$26342 ( \35257 , \35256 );
and \U$26343 ( \35258 , \28118 , \16680_nG9bed );
and \U$26344 ( \35259 , \28115 , \17665_nG9bea );
or \U$26345 ( \35260 , \35258 , \35259 );
xor \U$26346 ( \35261 , \28114 , \35260 );
buf \U$26347 ( \35262 , \35261 );
buf \U$26349 ( \35263 , \35262 );
xor \U$26350 ( \35264 , \35257 , \35263 );
and \U$26351 ( \35265 , \26431 , \18107_nG9be7 );
and \U$26352 ( \35266 , \26428 , \19091_nG9be4 );
or \U$26353 ( \35267 , \35265 , \35266 );
xor \U$26354 ( \35268 , \26427 , \35267 );
buf \U$26355 ( \35269 , \35268 );
buf \U$26357 ( \35270 , \35269 );
xor \U$26358 ( \35271 , \35264 , \35270 );
buf \U$26359 ( \35272 , \35271 );
xor \U$26360 ( \35273 , \35252 , \35272 );
and \U$26361 ( \35274 , \18702 , \25860_nG9bc9 );
and \U$26362 ( \35275 , \18699 , \26887_nG9bc6 );
or \U$26363 ( \35276 , \35274 , \35275 );
xor \U$26364 ( \35277 , \18698 , \35276 );
buf \U$26365 ( \35278 , \35277 );
buf \U$26367 ( \35279 , \35278 );
xor \U$26368 ( \35280 , \35273 , \35279 );
buf \U$26369 ( \35281 , \35280 );
xor \U$26370 ( \35282 , \35247 , \35281 );
buf \U$26371 ( \35283 , \35282 );
xor \U$26372 ( \35284 , \35236 , \35283 );
buf \U$26373 ( \35285 , \35284 );
and \U$26374 ( \35286 , \35101 , \35106 );
and \U$26375 ( \35287 , \35101 , \35155 );
and \U$26376 ( \35288 , \35106 , \35155 );
or \U$26377 ( \35289 , \35286 , \35287 , \35288 );
buf \U$26378 ( \35290 , \35289 );
xor \U$26379 ( \35291 , \35285 , \35290 );
and \U$26380 ( \35292 , \34847 , \34852 );
and \U$26381 ( \35293 , \34847 , \34919 );
and \U$26382 ( \35294 , \34852 , \34919 );
or \U$26383 ( \35295 , \35292 , \35293 , \35294 );
buf \U$26384 ( \35296 , \35295 );
xor \U$26385 ( \35297 , \35291 , \35296 );
buf \U$26386 ( \35298 , \35297 );
xor \U$26387 ( \35299 , \35225 , \35298 );
and \U$26388 ( \35300 , \35122 , \35128 );
and \U$26389 ( \35301 , \35122 , \35135 );
and \U$26390 ( \35302 , \35128 , \35135 );
or \U$26391 ( \35303 , \35300 , \35301 , \35302 );
buf \U$26392 ( \35304 , \35303 );
and \U$26393 ( \35305 , \21658 , \22629_nG9bd5 );
and \U$26394 ( \35306 , \21655 , \23696_nG9bd2 );
or \U$26395 ( \35307 , \35305 , \35306 );
xor \U$26396 ( \35308 , \21654 , \35307 );
buf \U$26397 ( \35309 , \35308 );
buf \U$26399 ( \35310 , \35309 );
xor \U$26400 ( \35311 , \35304 , \35310 );
and \U$26401 ( \35312 , \20155 , \24226_nG9bcf );
and \U$26402 ( \35313 , \20152 , \25298_nG9bcc );
or \U$26403 ( \35314 , \35312 , \35313 );
xor \U$26404 ( \35315 , \20151 , \35314 );
buf \U$26405 ( \35316 , \35315 );
buf \U$26407 ( \35317 , \35316 );
xor \U$26408 ( \35318 , \35311 , \35317 );
buf \U$26409 ( \35319 , \35318 );
and \U$26410 ( \35320 , \13370 , \32888_nG9bb1 );
and \U$26411 ( \35321 , \13367 , \33181_nG9bae );
or \U$26412 ( \35322 , \35320 , \35321 );
xor \U$26413 ( \35323 , \13366 , \35322 );
buf \U$26414 ( \35324 , \35323 );
buf \U$26416 ( \35325 , \35324 );
xor \U$26417 ( \35326 , \35319 , \35325 );
and \U$26418 ( \35327 , \10421 , \34294_nG9ba5 );
and \U$26419 ( \35328 , \10418 , \34643_nG9ba2 );
or \U$26420 ( \35329 , \35327 , \35328 );
xor \U$26421 ( \35330 , \10417 , \35329 );
buf \U$26422 ( \35331 , \35330 );
buf \U$26424 ( \35332 , \35331 );
xor \U$26425 ( \35333 , \35326 , \35332 );
buf \U$26426 ( \35334 , \35333 );
and \U$26427 ( \35335 , \35112 , \35146 );
and \U$26428 ( \35336 , \35112 , \35153 );
and \U$26429 ( \35337 , \35146 , \35153 );
or \U$26430 ( \35338 , \35335 , \35336 , \35337 );
buf \U$26431 ( \35339 , \35338 );
xor \U$26432 ( \35340 , \35334 , \35339 );
and \U$26433 ( \35341 , \35175 , \35181 );
and \U$26434 ( \35342 , \35175 , \35188 );
and \U$26435 ( \35343 , \35181 , \35188 );
or \U$26436 ( \35344 , \35341 , \35342 , \35343 );
buf \U$26437 ( \35345 , \35344 );
xor \U$26438 ( \35346 , \35340 , \35345 );
buf \U$26439 ( \35347 , \35346 );
and \U$26440 ( \35348 , \35163 , \35168 );
and \U$26441 ( \35349 , \35163 , \35190 );
and \U$26442 ( \35350 , \35168 , \35190 );
or \U$26443 ( \35351 , \35348 , \35349 , \35350 );
buf \U$26444 ( \35352 , \35351 );
xor \U$26445 ( \35353 , \35347 , \35352 );
and \U$26446 ( \35354 , \15940 , \29179_nG9bbd );
and \U$26447 ( \35355 , \15937 , \30366_nG9bba );
or \U$26448 ( \35356 , \35354 , \35355 );
xor \U$26449 ( \35357 , \15936 , \35356 );
buf \U$26450 ( \35358 , \35357 );
buf \U$26452 ( \35359 , \35358 );
and \U$26453 ( \35360 , \14631 , \30940_nG9bb7 );
and \U$26454 ( \35361 , \14628 , \32179_nG9bb4 );
or \U$26455 ( \35362 , \35360 , \35361 );
xor \U$26456 ( \35363 , \14627 , \35362 );
buf \U$26457 ( \35364 , \35363 );
buf \U$26459 ( \35365 , \35364 );
xor \U$26460 ( \35366 , \35359 , \35365 );
and \U$26461 ( \35367 , \12157 , \33613_nG9bab );
and \U$26462 ( \35368 , \12154 , \34041_nG9ba8 );
or \U$26463 ( \35369 , \35367 , \35368 );
xor \U$26464 ( \35370 , \12153 , \35369 );
buf \U$26465 ( \35371 , \35370 );
buf \U$26467 ( \35372 , \35371 );
xor \U$26468 ( \35373 , \35366 , \35372 );
buf \U$26469 ( \35374 , \35373 );
and \U$26470 ( \35375 , \35117 , \35137 );
and \U$26471 ( \35376 , \35117 , \35144 );
and \U$26472 ( \35377 , \35137 , \35144 );
or \U$26473 ( \35378 , \35375 , \35376 , \35377 );
buf \U$26474 ( \35379 , \35378 );
and \U$26476 ( \35380 , \32916 , \13705_nG9bfc );
or \U$26477 ( \35381 , 1'b0 , \35380 );
xor \U$26478 ( \35382 , 1'b0 , \35381 );
buf \U$26479 ( \35383 , \35382 );
buf \U$26481 ( \35384 , \35383 );
and \U$26482 ( \35385 , \31636 , \14070_nG9bf9 );
and \U$26483 ( \35386 , \31633 , \14984_nG9bf6 );
or \U$26484 ( \35387 , \35385 , \35386 );
xor \U$26485 ( \35388 , \31632 , \35387 );
buf \U$26486 ( \35389 , \35388 );
buf \U$26488 ( \35390 , \35389 );
xor \U$26489 ( \35391 , \35384 , \35390 );
buf \U$26490 ( \35392 , \35391 );
and \U$26491 ( \35393 , \34874 , \34880 );
buf \U$26492 ( \35394 , \35393 );
xor \U$26493 ( \35395 , \35392 , \35394 );
and \U$26494 ( \35396 , \29853 , \15373_nG9bf3 );
and \U$26495 ( \35397 , \29850 , \16315_nG9bf0 );
or \U$26496 ( \35398 , \35396 , \35397 );
xor \U$26497 ( \35399 , \29849 , \35398 );
buf \U$26498 ( \35400 , \35399 );
buf \U$26500 ( \35401 , \35400 );
xor \U$26501 ( \35402 , \35395 , \35401 );
buf \U$26502 ( \35403 , \35402 );
and \U$26503 ( \35404 , \24792 , \19586_nG9be1 );
and \U$26504 ( \35405 , \24789 , \20608_nG9bde );
or \U$26505 ( \35406 , \35404 , \35405 );
xor \U$26506 ( \35407 , \24788 , \35406 );
buf \U$26507 ( \35408 , \35407 );
buf \U$26509 ( \35409 , \35408 );
xor \U$26510 ( \35410 , \35403 , \35409 );
and \U$26511 ( \35411 , \23201 , \21086_nG9bdb );
and \U$26512 ( \35412 , \23198 , \22129_nG9bd8 );
or \U$26513 ( \35413 , \35411 , \35412 );
xor \U$26514 ( \35414 , \23197 , \35413 );
buf \U$26515 ( \35415 , \35414 );
buf \U$26517 ( \35416 , \35415 );
xor \U$26518 ( \35417 , \35410 , \35416 );
buf \U$26519 ( \35418 , \35417 );
xor \U$26520 ( \35419 , \35379 , \35418 );
and \U$26521 ( \35420 , \17297 , \27416_nG9bc3 );
and \U$26522 ( \35421 , \17294 , \28602_nG9bc0 );
or \U$26523 ( \35422 , \35420 , \35421 );
xor \U$26524 ( \35423 , \17293 , \35422 );
buf \U$26525 ( \35424 , \35423 );
buf \U$26527 ( \35425 , \35424 );
xor \U$26528 ( \35426 , \35419 , \35425 );
buf \U$26529 ( \35427 , \35426 );
xor \U$26530 ( \35428 , \35374 , \35427 );
and \U$26531 ( \35429 , \10707 , \35094_nG9b9f );
and \U$26532 ( \35430 , \34957 , \34961 );
and \U$26533 ( \35431 , \34961 , \35003 );
and \U$26534 ( \35432 , \34957 , \35003 );
or \U$26535 ( \35433 , \35430 , \35431 , \35432 );
and \U$26536 ( \35434 , \35009 , \35013 );
and \U$26537 ( \35435 , \35013 , \35082 );
and \U$26538 ( \35436 , \35009 , \35082 );
or \U$26539 ( \35437 , \35434 , \35435 , \35436 );
xor \U$26540 ( \35438 , \35433 , \35437 );
and \U$26541 ( \35439 , \35018 , \35056 );
and \U$26542 ( \35440 , \35056 , \35081 );
and \U$26543 ( \35441 , \35018 , \35081 );
or \U$26544 ( \35442 , \35439 , \35440 , \35441 );
and \U$26545 ( \35443 , \35029 , \35043 );
and \U$26546 ( \35444 , \35043 , \35055 );
and \U$26547 ( \35445 , \35029 , \35055 );
or \U$26548 ( \35446 , \35443 , \35444 , \35445 );
and \U$26549 ( \35447 , \35061 , \35065 );
and \U$26550 ( \35448 , \35065 , \35080 );
and \U$26551 ( \35449 , \35061 , \35080 );
or \U$26552 ( \35450 , \35447 , \35448 , \35449 );
xor \U$26553 ( \35451 , \35446 , \35450 );
and \U$26554 ( \35452 , \35048 , \35052 );
and \U$26555 ( \35453 , \35052 , \35054 );
and \U$26556 ( \35454 , \35048 , \35054 );
or \U$26557 ( \35455 , \35452 , \35453 , \35454 );
and \U$26558 ( \35456 , \29084 , \16635 );
and \U$26559 ( \35457 , \30268 , \16301 );
nor \U$26560 ( \35458 , \35456 , \35457 );
xnor \U$26561 ( \35459 , \35458 , \16625 );
and \U$26562 ( \35460 , \14024 , \32854 );
and \U$26563 ( \35461 , \14950 , \32067 );
nor \U$26564 ( \35462 , \35460 , \35461 );
xnor \U$26565 ( \35463 , \35462 , \32805 );
xor \U$26566 ( \35464 , \35459 , \35463 );
and \U$26567 ( \35465 , \13679 , \32802 );
xor \U$26568 ( \35466 , \35464 , \35465 );
xor \U$26569 ( \35467 , \35455 , \35466 );
and \U$26570 ( \35468 , \27313 , \18090 );
and \U$26571 ( \35469 , \28534 , \17655 );
nor \U$26572 ( \35470 , \35468 , \35469 );
xnor \U$26573 ( \35471 , \35470 , \18046 );
and \U$26574 ( \35472 , \21033 , \24138 );
and \U$26575 ( \35473 , \22090 , \23630 );
nor \U$26576 ( \35474 , \35472 , \35473 );
xnor \U$26577 ( \35475 , \35474 , \24144 );
xor \U$26578 ( \35476 , \35471 , \35475 );
and \U$26579 ( \35477 , \19558 , \25826 );
and \U$26580 ( \35478 , \20544 , \25264 );
nor \U$26581 ( \35479 , \35477 , \35478 );
xnor \U$26582 ( \35480 , \35479 , \25773 );
xor \U$26583 ( \35481 , \35476 , \35480 );
xor \U$26584 ( \35482 , \35467 , \35481 );
xor \U$26585 ( \35483 , \35451 , \35482 );
xor \U$26586 ( \35484 , \35442 , \35483 );
and \U$26587 ( \35485 , \34966 , \34977 );
and \U$26588 ( \35486 , \34977 , \35002 );
and \U$26589 ( \35487 , \34966 , \35002 );
or \U$26590 ( \35488 , \35485 , \35486 , \35487 );
and \U$26591 ( \35489 , \32794 , \14054 );
not \U$26592 ( \35490 , \35489 );
xnor \U$26593 ( \35491 , \35490 , \14035 );
and \U$26594 ( \35492 , \24199 , \21005 );
and \U$26595 ( \35493 , \25272 , \20557 );
nor \U$26596 ( \35494 , \35492 , \35493 );
xnor \U$26597 ( \35495 , \35494 , \21011 );
xor \U$26598 ( \35496 , \35491 , \35495 );
and \U$26599 ( \35497 , \15321 , \30823 );
and \U$26600 ( \35498 , \16267 , \30246 );
nor \U$26601 ( \35499 , \35497 , \35498 );
xnor \U$26602 ( \35500 , \35499 , \30813 );
xor \U$26603 ( \35501 , \35496 , \35500 );
and \U$26604 ( \35502 , \25815 , \19534 );
and \U$26605 ( \35503 , \26829 , \19045 );
nor \U$26606 ( \35504 , \35502 , \35503 );
xnor \U$26607 ( \35505 , \35504 , \19540 );
and \U$26608 ( \35506 , \18035 , \27397 );
and \U$26609 ( \35507 , \19032 , \26807 );
nor \U$26610 ( \35508 , \35506 , \35507 );
xnor \U$26611 ( \35509 , \35508 , \27295 );
xor \U$26612 ( \35510 , \35505 , \35509 );
and \U$26613 ( \35511 , \16655 , \29070 );
and \U$26614 ( \35512 , \17627 , \28526 );
nor \U$26615 ( \35513 , \35511 , \35512 );
xnor \U$26616 ( \35514 , \35513 , \29076 );
xor \U$26617 ( \35515 , \35510 , \35514 );
xor \U$26618 ( \35516 , \35501 , \35515 );
and \U$26619 ( \35517 , \35033 , \35037 );
and \U$26620 ( \35518 , \35037 , \35042 );
and \U$26621 ( \35519 , \35033 , \35042 );
or \U$26622 ( \35520 , \35517 , \35518 , \35519 );
and \U$26623 ( \35521 , \30802 , \15336 );
and \U$26624 ( \35522 , \32054 , \14963 );
nor \U$26625 ( \35523 , \35521 , \35522 );
xnor \U$26626 ( \35524 , \35523 , \15342 );
not \U$26627 ( \35525 , \35524 );
xor \U$26628 ( \35526 , \35520 , \35525 );
and \U$26629 ( \35527 , \22556 , \22542 );
and \U$26630 ( \35528 , \23617 , \22103 );
nor \U$26631 ( \35529 , \35527 , \35528 );
xnor \U$26632 ( \35530 , \35529 , \22548 );
xor \U$26633 ( \35531 , \35526 , \35530 );
xor \U$26634 ( \35532 , \35516 , \35531 );
xor \U$26635 ( \35533 , \35488 , \35532 );
and \U$26636 ( \35534 , \34970 , \34974 );
and \U$26637 ( \35535 , \34974 , \34976 );
and \U$26638 ( \35536 , \34970 , \34976 );
or \U$26639 ( \35537 , \35534 , \35535 , \35536 );
and \U$26640 ( \35538 , \34982 , \34986 );
and \U$26641 ( \35539 , \34986 , \35001 );
and \U$26642 ( \35540 , \34982 , \35001 );
or \U$26643 ( \35541 , \35538 , \35539 , \35540 );
xor \U$26644 ( \35542 , \35537 , \35541 );
and \U$26645 ( \35543 , \34991 , \34995 );
and \U$26646 ( \35544 , \34995 , \35000 );
and \U$26647 ( \35545 , \34991 , \35000 );
or \U$26648 ( \35546 , \35543 , \35544 , \35545 );
and \U$26649 ( \35547 , \35070 , \35074 );
and \U$26650 ( \35548 , \35074 , \35079 );
and \U$26651 ( \35549 , \35070 , \35079 );
or \U$26652 ( \35550 , \35547 , \35548 , \35549 );
xor \U$26653 ( \35551 , \35546 , \35550 );
and \U$26654 ( \35552 , \35019 , \35023 );
and \U$26655 ( \35553 , \35023 , \35028 );
and \U$26656 ( \35554 , \35019 , \35028 );
or \U$26657 ( \35555 , \35552 , \35553 , \35554 );
xor \U$26658 ( \35556 , \35551 , \35555 );
xor \U$26659 ( \35557 , \35542 , \35556 );
xor \U$26660 ( \35558 , \35533 , \35557 );
xor \U$26661 ( \35559 , \35484 , \35558 );
xor \U$26662 ( \35560 , \35438 , \35559 );
and \U$26663 ( \35561 , \34953 , \35004 );
and \U$26664 ( \35562 , \35004 , \35083 );
and \U$26665 ( \35563 , \34953 , \35083 );
or \U$26666 ( \35564 , \35561 , \35562 , \35563 );
xor \U$26667 ( \35565 , \35560 , \35564 );
and \U$26668 ( \35566 , \35084 , \35088 );
and \U$26669 ( \35567 , \35089 , \35092 );
or \U$26670 ( \35568 , \35566 , \35567 );
xor \U$26671 ( \35569 , \35565 , \35568 );
buf g9b9c ( \35570_nG9b9c , \35569 );
and \U$26672 ( \35571 , \10704 , \35570_nG9b9c );
or \U$26673 ( \35572 , \35429 , \35571 );
xor \U$26674 ( \35573 , \10703 , \35572 );
buf \U$26675 ( \35574 , \35573 );
buf \U$26677 ( \35575 , \35574 );
xor \U$26678 ( \35576 , \35428 , \35575 );
buf \U$26679 ( \35577 , \35576 );
xor \U$26680 ( \35578 , \35353 , \35577 );
buf \U$26681 ( \35579 , \35578 );
xor \U$26682 ( \35580 , \35299 , \35579 );
and \U$26683 ( \35581 , \35220 , \35580 );
and \U$26685 ( \35582 , \35214 , \35219 );
or \U$26687 ( \35583 , 1'b0 , \35582 , 1'b0 );
xor \U$26688 ( \35584 , \35581 , \35583 );
and \U$26690 ( \35585 , \35207 , \35213 );
and \U$26691 ( \35586 , \35209 , \35213 );
or \U$26692 ( \35587 , 1'b0 , \35585 , \35586 );
xor \U$26693 ( \35588 , \35584 , \35587 );
xor \U$26700 ( \35589 , \35588 , 1'b0 );
and \U$26701 ( \35590 , \35225 , \35298 );
and \U$26702 ( \35591 , \35225 , \35579 );
and \U$26703 ( \35592 , \35298 , \35579 );
or \U$26704 ( \35593 , \35590 , \35591 , \35592 );
xor \U$26705 ( \35594 , \35589 , \35593 );
and \U$26706 ( \35595 , \35347 , \35352 );
and \U$26707 ( \35596 , \35347 , \35577 );
and \U$26708 ( \35597 , \35352 , \35577 );
or \U$26709 ( \35598 , \35595 , \35596 , \35597 );
buf \U$26710 ( \35599 , \35598 );
and \U$26711 ( \35600 , \35319 , \35325 );
and \U$26712 ( \35601 , \35319 , \35332 );
and \U$26713 ( \35602 , \35325 , \35332 );
or \U$26714 ( \35603 , \35600 , \35601 , \35602 );
buf \U$26715 ( \35604 , \35603 );
and \U$26716 ( \35605 , \35304 , \35310 );
and \U$26717 ( \35606 , \35304 , \35317 );
and \U$26718 ( \35607 , \35310 , \35317 );
or \U$26719 ( \35608 , \35605 , \35606 , \35607 );
buf \U$26720 ( \35609 , \35608 );
and \U$26721 ( \35610 , \14631 , \32179_nG9bb4 );
and \U$26722 ( \35611 , \14628 , \32888_nG9bb1 );
or \U$26723 ( \35612 , \35610 , \35611 );
xor \U$26724 ( \35613 , \14627 , \35612 );
buf \U$26725 ( \35614 , \35613 );
buf \U$26727 ( \35615 , \35614 );
xor \U$26728 ( \35616 , \35609 , \35615 );
and \U$26729 ( \35617 , \13370 , \33181_nG9bae );
and \U$26730 ( \35618 , \13367 , \33613_nG9bab );
or \U$26731 ( \35619 , \35617 , \35618 );
xor \U$26732 ( \35620 , \13366 , \35619 );
buf \U$26733 ( \35621 , \35620 );
buf \U$26735 ( \35622 , \35621 );
xor \U$26736 ( \35623 , \35616 , \35622 );
buf \U$26737 ( \35624 , \35623 );
xor \U$26738 ( \35625 , \35604 , \35624 );
and \U$26739 ( \35626 , \35241 , \35246 );
and \U$26740 ( \35627 , \35241 , \35281 );
and \U$26741 ( \35628 , \35246 , \35281 );
or \U$26742 ( \35629 , \35626 , \35627 , \35628 );
buf \U$26743 ( \35630 , \35629 );
xor \U$26744 ( \35631 , \35625 , \35630 );
buf \U$26745 ( \35632 , \35631 );
xor \U$26746 ( \35633 , \35599 , \35632 );
and \U$26747 ( \35634 , \35374 , \35427 );
and \U$26748 ( \35635 , \35374 , \35575 );
and \U$26749 ( \35636 , \35427 , \35575 );
or \U$26750 ( \35637 , \35634 , \35635 , \35636 );
buf \U$26751 ( \35638 , \35637 );
and \U$26752 ( \35639 , \35403 , \35409 );
and \U$26753 ( \35640 , \35403 , \35416 );
and \U$26754 ( \35641 , \35409 , \35416 );
or \U$26755 ( \35642 , \35639 , \35640 , \35641 );
buf \U$26756 ( \35643 , \35642 );
and \U$26757 ( \35644 , \23201 , \22129_nG9bd8 );
and \U$26758 ( \35645 , \23198 , \22629_nG9bd5 );
or \U$26759 ( \35646 , \35644 , \35645 );
xor \U$26760 ( \35647 , \23197 , \35646 );
buf \U$26761 ( \35648 , \35647 );
buf \U$26763 ( \35649 , \35648 );
xor \U$26764 ( \35650 , \35643 , \35649 );
and \U$26765 ( \35651 , \21658 , \23696_nG9bd2 );
and \U$26766 ( \35652 , \21655 , \24226_nG9bcf );
or \U$26767 ( \35653 , \35651 , \35652 );
xor \U$26768 ( \35654 , \21654 , \35653 );
buf \U$26769 ( \35655 , \35654 );
buf \U$26771 ( \35656 , \35655 );
xor \U$26772 ( \35657 , \35650 , \35656 );
buf \U$26773 ( \35658 , \35657 );
and \U$26774 ( \35659 , \10421 , \34643_nG9ba2 );
and \U$26775 ( \35660 , \10418 , \35094_nG9b9f );
or \U$26776 ( \35661 , \35659 , \35660 );
xor \U$26777 ( \35662 , \10417 , \35661 );
buf \U$26778 ( \35663 , \35662 );
buf \U$26780 ( \35664 , \35663 );
xor \U$26781 ( \35665 , \35658 , \35664 );
and \U$26782 ( \35666 , \10707 , \35570_nG9b9c );
and \U$26783 ( \35667 , \35488 , \35532 );
and \U$26784 ( \35668 , \35532 , \35557 );
and \U$26785 ( \35669 , \35488 , \35557 );
or \U$26786 ( \35670 , \35667 , \35668 , \35669 );
and \U$26787 ( \35671 , \35442 , \35483 );
and \U$26788 ( \35672 , \35483 , \35558 );
and \U$26789 ( \35673 , \35442 , \35558 );
or \U$26790 ( \35674 , \35671 , \35672 , \35673 );
xor \U$26791 ( \35675 , \35670 , \35674 );
and \U$26792 ( \35676 , \35446 , \35450 );
and \U$26793 ( \35677 , \35450 , \35482 );
and \U$26794 ( \35678 , \35446 , \35482 );
or \U$26795 ( \35679 , \35676 , \35677 , \35678 );
and \U$26796 ( \35680 , \35501 , \35515 );
and \U$26797 ( \35681 , \35515 , \35531 );
and \U$26798 ( \35682 , \35501 , \35531 );
or \U$26799 ( \35683 , \35680 , \35681 , \35682 );
and \U$26800 ( \35684 , \35537 , \35541 );
and \U$26801 ( \35685 , \35541 , \35556 );
and \U$26802 ( \35686 , \35537 , \35556 );
or \U$26803 ( \35687 , \35684 , \35685 , \35686 );
xor \U$26804 ( \35688 , \35683 , \35687 );
and \U$26805 ( \35689 , \35546 , \35550 );
and \U$26806 ( \35690 , \35550 , \35555 );
and \U$26807 ( \35691 , \35546 , \35555 );
or \U$26808 ( \35692 , \35689 , \35690 , \35691 );
and \U$26809 ( \35693 , \35520 , \35525 );
and \U$26810 ( \35694 , \35525 , \35530 );
and \U$26811 ( \35695 , \35520 , \35530 );
or \U$26812 ( \35696 , \35693 , \35694 , \35695 );
xor \U$26813 ( \35697 , \35692 , \35696 );
and \U$26814 ( \35698 , \35491 , \35495 );
and \U$26815 ( \35699 , \35495 , \35500 );
and \U$26816 ( \35700 , \35491 , \35500 );
or \U$26817 ( \35701 , \35698 , \35699 , \35700 );
and \U$26818 ( \35702 , \35505 , \35509 );
and \U$26819 ( \35703 , \35509 , \35514 );
and \U$26820 ( \35704 , \35505 , \35514 );
or \U$26821 ( \35705 , \35702 , \35703 , \35704 );
xor \U$26822 ( \35706 , \35701 , \35705 );
and \U$26823 ( \35707 , \35471 , \35475 );
and \U$26824 ( \35708 , \35475 , \35480 );
and \U$26825 ( \35709 , \35471 , \35480 );
or \U$26826 ( \35710 , \35707 , \35708 , \35709 );
xor \U$26827 ( \35711 , \35706 , \35710 );
xor \U$26828 ( \35712 , \35697 , \35711 );
xor \U$26829 ( \35713 , \35688 , \35712 );
xor \U$26830 ( \35714 , \35679 , \35713 );
and \U$26831 ( \35715 , \35455 , \35466 );
and \U$26832 ( \35716 , \35466 , \35481 );
and \U$26833 ( \35717 , \35455 , \35481 );
or \U$26834 ( \35718 , \35715 , \35716 , \35717 );
and \U$26835 ( \35719 , \35459 , \35463 );
and \U$26836 ( \35720 , \35463 , \35465 );
and \U$26837 ( \35721 , \35459 , \35465 );
or \U$26838 ( \35722 , \35719 , \35720 , \35721 );
and \U$26839 ( \35723 , \26829 , \19534 );
and \U$26840 ( \35724 , \27313 , \19045 );
nor \U$26841 ( \35725 , \35723 , \35724 );
xnor \U$26842 ( \35726 , \35725 , \19540 );
and \U$26843 ( \35727 , \22090 , \24138 );
and \U$26844 ( \35728 , \22556 , \23630 );
nor \U$26845 ( \35729 , \35727 , \35728 );
xnor \U$26846 ( \35730 , \35729 , \24144 );
xor \U$26847 ( \35731 , \35726 , \35730 );
and \U$26848 ( \35732 , \20544 , \25826 );
and \U$26849 ( \35733 , \21033 , \25264 );
nor \U$26850 ( \35734 , \35732 , \35733 );
xnor \U$26851 ( \35735 , \35734 , \25773 );
xor \U$26852 ( \35736 , \35731 , \35735 );
xor \U$26853 ( \35737 , \35722 , \35736 );
not \U$26854 ( \35738 , \14035 );
and \U$26855 ( \35739 , \32054 , \15336 );
and \U$26856 ( \35740 , \32794 , \14963 );
nor \U$26857 ( \35741 , \35739 , \35740 );
xnor \U$26858 ( \35742 , \35741 , \15342 );
xor \U$26859 ( \35743 , \35738 , \35742 );
and \U$26860 ( \35744 , \28534 , \18090 );
and \U$26861 ( \35745 , \29084 , \17655 );
nor \U$26862 ( \35746 , \35744 , \35745 );
xnor \U$26863 ( \35747 , \35746 , \18046 );
xor \U$26864 ( \35748 , \35743 , \35747 );
xor \U$26865 ( \35749 , \35737 , \35748 );
xor \U$26866 ( \35750 , \35718 , \35749 );
and \U$26867 ( \35751 , \25272 , \21005 );
and \U$26868 ( \35752 , \25815 , \20557 );
nor \U$26869 ( \35753 , \35751 , \35752 );
xnor \U$26870 ( \35754 , \35753 , \21011 );
and \U$26871 ( \35755 , \16267 , \30823 );
and \U$26872 ( \35756 , \16655 , \30246 );
nor \U$26873 ( \35757 , \35755 , \35756 );
xnor \U$26874 ( \35758 , \35757 , \30813 );
xor \U$26875 ( \35759 , \35754 , \35758 );
and \U$26876 ( \35760 , \14950 , \32854 );
and \U$26877 ( \35761 , \15321 , \32067 );
nor \U$26878 ( \35762 , \35760 , \35761 );
xnor \U$26879 ( \35763 , \35762 , \32805 );
xor \U$26880 ( \35764 , \35759 , \35763 );
and \U$26881 ( \35765 , \30268 , \16635 );
and \U$26882 ( \35766 , \30802 , \16301 );
nor \U$26883 ( \35767 , \35765 , \35766 );
xnor \U$26884 ( \35768 , \35767 , \16625 );
and \U$26885 ( \35769 , \19032 , \27397 );
and \U$26886 ( \35770 , \19558 , \26807 );
nor \U$26887 ( \35771 , \35769 , \35770 );
xnor \U$26888 ( \35772 , \35771 , \27295 );
xor \U$26889 ( \35773 , \35768 , \35772 );
and \U$26890 ( \35774 , \17627 , \29070 );
and \U$26891 ( \35775 , \18035 , \28526 );
nor \U$26892 ( \35776 , \35774 , \35775 );
xnor \U$26893 ( \35777 , \35776 , \29076 );
xor \U$26894 ( \35778 , \35773 , \35777 );
xor \U$26895 ( \35779 , \35764 , \35778 );
buf \U$26896 ( \35780 , \35524 );
and \U$26897 ( \35781 , \23617 , \22542 );
and \U$26898 ( \35782 , \24199 , \22103 );
nor \U$26899 ( \35783 , \35781 , \35782 );
xnor \U$26900 ( \35784 , \35783 , \22548 );
xor \U$26901 ( \35785 , \35780 , \35784 );
and \U$26902 ( \35786 , \14024 , \32802 );
xor \U$26903 ( \35787 , \35785 , \35786 );
xor \U$26904 ( \35788 , \35779 , \35787 );
xor \U$26905 ( \35789 , \35750 , \35788 );
xor \U$26906 ( \35790 , \35714 , \35789 );
xor \U$26907 ( \35791 , \35675 , \35790 );
and \U$26908 ( \35792 , \35433 , \35437 );
and \U$26909 ( \35793 , \35437 , \35559 );
and \U$26910 ( \35794 , \35433 , \35559 );
or \U$26911 ( \35795 , \35792 , \35793 , \35794 );
xor \U$26912 ( \35796 , \35791 , \35795 );
and \U$26913 ( \35797 , \35560 , \35564 );
and \U$26914 ( \35798 , \35565 , \35568 );
or \U$26915 ( \35799 , \35797 , \35798 );
xor \U$26916 ( \35800 , \35796 , \35799 );
buf g9b99 ( \35801_nG9b99 , \35800 );
and \U$26917 ( \35802 , \10704 , \35801_nG9b99 );
or \U$26918 ( \35803 , \35666 , \35802 );
xor \U$26919 ( \35804 , \10703 , \35803 );
buf \U$26920 ( \35805 , \35804 );
buf \U$26922 ( \35806 , \35805 );
xor \U$26923 ( \35807 , \35665 , \35806 );
buf \U$26924 ( \35808 , \35807 );
xor \U$26925 ( \35809 , \35638 , \35808 );
and \U$26926 ( \35810 , \35392 , \35394 );
and \U$26927 ( \35811 , \35392 , \35401 );
and \U$26928 ( \35812 , \35394 , \35401 );
or \U$26929 ( \35813 , \35810 , \35811 , \35812 );
buf \U$26930 ( \35814 , \35813 );
and \U$26931 ( \35815 , \28118 , \17665_nG9bea );
and \U$26932 ( \35816 , \28115 , \18107_nG9be7 );
or \U$26933 ( \35817 , \35815 , \35816 );
xor \U$26934 ( \35818 , \28114 , \35817 );
buf \U$26935 ( \35819 , \35818 );
buf \U$26937 ( \35820 , \35819 );
xor \U$26938 ( \35821 , \35814 , \35820 );
and \U$26939 ( \35822 , \24792 , \20608_nG9bde );
and \U$26940 ( \35823 , \24789 , \21086_nG9bdb );
or \U$26941 ( \35824 , \35822 , \35823 );
xor \U$26942 ( \35825 , \24788 , \35824 );
buf \U$26943 ( \35826 , \35825 );
buf \U$26945 ( \35827 , \35826 );
xor \U$26946 ( \35828 , \35821 , \35827 );
buf \U$26947 ( \35829 , \35828 );
and \U$26948 ( \35830 , \20155 , \25298_nG9bcc );
and \U$26949 ( \35831 , \20152 , \25860_nG9bc9 );
or \U$26950 ( \35832 , \35830 , \35831 );
xor \U$26951 ( \35833 , \20151 , \35832 );
buf \U$26952 ( \35834 , \35833 );
buf \U$26954 ( \35835 , \35834 );
xor \U$26955 ( \35836 , \35829 , \35835 );
and \U$26956 ( \35837 , \18702 , \26887_nG9bc6 );
and \U$26957 ( \35838 , \18699 , \27416_nG9bc3 );
or \U$26958 ( \35839 , \35837 , \35838 );
xor \U$26959 ( \35840 , \18698 , \35839 );
buf \U$26960 ( \35841 , \35840 );
buf \U$26962 ( \35842 , \35841 );
xor \U$26963 ( \35843 , \35836 , \35842 );
buf \U$26964 ( \35844 , \35843 );
and \U$26965 ( \35845 , \35252 , \35272 );
and \U$26966 ( \35846 , \35252 , \35279 );
and \U$26967 ( \35847 , \35272 , \35279 );
or \U$26968 ( \35848 , \35845 , \35846 , \35847 );
buf \U$26969 ( \35849 , \35848 );
xor \U$26970 ( \35850 , \35844 , \35849 );
and \U$26971 ( \35851 , \12157 , \34041_nG9ba8 );
and \U$26972 ( \35852 , \12154 , \34294_nG9ba5 );
or \U$26973 ( \35853 , \35851 , \35852 );
xor \U$26974 ( \35854 , \12153 , \35853 );
buf \U$26975 ( \35855 , \35854 );
buf \U$26977 ( \35856 , \35855 );
xor \U$26978 ( \35857 , \35850 , \35856 );
buf \U$26979 ( \35858 , \35857 );
xor \U$26980 ( \35859 , \35809 , \35858 );
buf \U$26981 ( \35860 , \35859 );
xor \U$26982 ( \35861 , \35633 , \35860 );
buf \U$26983 ( \35862 , \35861 );
and \U$26984 ( \35863 , \35285 , \35290 );
and \U$26985 ( \35864 , \35285 , \35296 );
and \U$26986 ( \35865 , \35290 , \35296 );
or \U$26987 ( \35866 , \35863 , \35864 , \35865 );
buf \U$26988 ( \35867 , \35866 );
xor \U$26989 ( \35868 , \35862 , \35867 );
and \U$26990 ( \35869 , \35334 , \35339 );
and \U$26991 ( \35870 , \35334 , \35345 );
and \U$26992 ( \35871 , \35339 , \35345 );
or \U$26993 ( \35872 , \35869 , \35870 , \35871 );
buf \U$26994 ( \35873 , \35872 );
and \U$26995 ( \35874 , \35230 , \35235 );
and \U$26996 ( \35875 , \35230 , \35283 );
and \U$26997 ( \35876 , \35235 , \35283 );
or \U$26998 ( \35877 , \35874 , \35875 , \35876 );
buf \U$26999 ( \35878 , \35877 );
xor \U$27000 ( \35879 , \35873 , \35878 );
and \U$27001 ( \35880 , \35359 , \35365 );
and \U$27002 ( \35881 , \35359 , \35372 );
and \U$27003 ( \35882 , \35365 , \35372 );
or \U$27004 ( \35883 , \35880 , \35881 , \35882 );
buf \U$27005 ( \35884 , \35883 );
and \U$27006 ( \35885 , \35257 , \35263 );
and \U$27007 ( \35886 , \35257 , \35270 );
and \U$27008 ( \35887 , \35263 , \35270 );
or \U$27009 ( \35888 , \35885 , \35886 , \35887 );
buf \U$27010 ( \35889 , \35888 );
and \U$27012 ( \35890 , \32916 , \14070_nG9bf9 );
or \U$27013 ( \35891 , 1'b0 , \35890 );
xor \U$27014 ( \35892 , 1'b0 , \35891 );
buf \U$27015 ( \35893 , \35892 );
buf \U$27017 ( \35894 , \35893 );
and \U$27018 ( \35895 , \31636 , \14984_nG9bf6 );
and \U$27019 ( \35896 , \31633 , \15373_nG9bf3 );
or \U$27020 ( \35897 , \35895 , \35896 );
xor \U$27021 ( \35898 , \31632 , \35897 );
buf \U$27022 ( \35899 , \35898 );
buf \U$27024 ( \35900 , \35899 );
xor \U$27025 ( \35901 , \35894 , \35900 );
buf \U$27026 ( \35902 , \35901 );
and \U$27027 ( \35903 , \35384 , \35390 );
buf \U$27028 ( \35904 , \35903 );
xor \U$27029 ( \35905 , \35902 , \35904 );
and \U$27030 ( \35906 , \29853 , \16315_nG9bf0 );
and \U$27031 ( \35907 , \29850 , \16680_nG9bed );
or \U$27032 ( \35908 , \35906 , \35907 );
xor \U$27033 ( \35909 , \29849 , \35908 );
buf \U$27034 ( \35910 , \35909 );
buf \U$27036 ( \35911 , \35910 );
xor \U$27037 ( \35912 , \35905 , \35911 );
buf \U$27038 ( \35913 , \35912 );
xor \U$27039 ( \35914 , \35889 , \35913 );
and \U$27040 ( \35915 , \26431 , \19091_nG9be4 );
and \U$27041 ( \35916 , \26428 , \19586_nG9be1 );
or \U$27042 ( \35917 , \35915 , \35916 );
xor \U$27043 ( \35918 , \26427 , \35917 );
buf \U$27044 ( \35919 , \35918 );
buf \U$27046 ( \35920 , \35919 );
xor \U$27047 ( \35921 , \35914 , \35920 );
buf \U$27048 ( \35922 , \35921 );
and \U$27049 ( \35923 , \17297 , \28602_nG9bc0 );
and \U$27050 ( \35924 , \17294 , \29179_nG9bbd );
or \U$27051 ( \35925 , \35923 , \35924 );
xor \U$27052 ( \35926 , \17293 , \35925 );
buf \U$27053 ( \35927 , \35926 );
buf \U$27055 ( \35928 , \35927 );
xor \U$27056 ( \35929 , \35922 , \35928 );
and \U$27057 ( \35930 , \15940 , \30366_nG9bba );
and \U$27058 ( \35931 , \15937 , \30940_nG9bb7 );
or \U$27059 ( \35932 , \35930 , \35931 );
xor \U$27060 ( \35933 , \15936 , \35932 );
buf \U$27061 ( \35934 , \35933 );
buf \U$27063 ( \35935 , \35934 );
xor \U$27064 ( \35936 , \35929 , \35935 );
buf \U$27065 ( \35937 , \35936 );
xor \U$27066 ( \35938 , \35884 , \35937 );
and \U$27067 ( \35939 , \35379 , \35418 );
and \U$27068 ( \35940 , \35379 , \35425 );
and \U$27069 ( \35941 , \35418 , \35425 );
or \U$27070 ( \35942 , \35939 , \35940 , \35941 );
buf \U$27071 ( \35943 , \35942 );
xor \U$27072 ( \35944 , \35938 , \35943 );
buf \U$27073 ( \35945 , \35944 );
xor \U$27074 ( \35946 , \35879 , \35945 );
buf \U$27075 ( \35947 , \35946 );
xor \U$27076 ( \35948 , \35868 , \35947 );
and \U$27077 ( \35949 , \35594 , \35948 );
and \U$27079 ( \35950 , \35588 , \35593 );
or \U$27081 ( \35951 , 1'b0 , \35950 , 1'b0 );
xor \U$27082 ( \35952 , \35949 , \35951 );
and \U$27084 ( \35953 , \35581 , \35587 );
and \U$27085 ( \35954 , \35583 , \35587 );
or \U$27086 ( \35955 , 1'b0 , \35953 , \35954 );
xor \U$27087 ( \35956 , \35952 , \35955 );
xor \U$27094 ( \35957 , \35956 , 1'b0 );
and \U$27095 ( \35958 , \35862 , \35867 );
and \U$27096 ( \35959 , \35862 , \35947 );
and \U$27097 ( \35960 , \35867 , \35947 );
or \U$27098 ( \35961 , \35958 , \35959 , \35960 );
xor \U$27099 ( \35962 , \35957 , \35961 );
and \U$27100 ( \35963 , \35873 , \35878 );
and \U$27101 ( \35964 , \35873 , \35945 );
and \U$27102 ( \35965 , \35878 , \35945 );
or \U$27103 ( \35966 , \35963 , \35964 , \35965 );
buf \U$27104 ( \35967 , \35966 );
and \U$27105 ( \35968 , \35638 , \35808 );
and \U$27106 ( \35969 , \35638 , \35858 );
and \U$27107 ( \35970 , \35808 , \35858 );
or \U$27108 ( \35971 , \35968 , \35969 , \35970 );
buf \U$27109 ( \35972 , \35971 );
xor \U$27110 ( \35973 , \35967 , \35972 );
and \U$27111 ( \35974 , \35884 , \35937 );
and \U$27112 ( \35975 , \35884 , \35943 );
and \U$27113 ( \35976 , \35937 , \35943 );
or \U$27114 ( \35977 , \35974 , \35975 , \35976 );
buf \U$27115 ( \35978 , \35977 );
and \U$27116 ( \35979 , \35922 , \35928 );
and \U$27117 ( \35980 , \35922 , \35935 );
and \U$27118 ( \35981 , \35928 , \35935 );
or \U$27119 ( \35982 , \35979 , \35980 , \35981 );
buf \U$27120 ( \35983 , \35982 );
and \U$27121 ( \35984 , \35814 , \35820 );
and \U$27122 ( \35985 , \35814 , \35827 );
and \U$27123 ( \35986 , \35820 , \35827 );
or \U$27124 ( \35987 , \35984 , \35985 , \35986 );
buf \U$27125 ( \35988 , \35987 );
and \U$27126 ( \35989 , \21658 , \24226_nG9bcf );
and \U$27127 ( \35990 , \21655 , \25298_nG9bcc );
or \U$27128 ( \35991 , \35989 , \35990 );
xor \U$27129 ( \35992 , \21654 , \35991 );
buf \U$27130 ( \35993 , \35992 );
buf \U$27132 ( \35994 , \35993 );
xor \U$27133 ( \35995 , \35988 , \35994 );
and \U$27134 ( \35996 , \18702 , \27416_nG9bc3 );
and \U$27135 ( \35997 , \18699 , \28602_nG9bc0 );
or \U$27136 ( \35998 , \35996 , \35997 );
xor \U$27137 ( \35999 , \18698 , \35998 );
buf \U$27138 ( \36000 , \35999 );
buf \U$27140 ( \36001 , \36000 );
xor \U$27141 ( \36002 , \35995 , \36001 );
buf \U$27142 ( \36003 , \36002 );
xor \U$27143 ( \36004 , \35983 , \36003 );
and \U$27144 ( \36005 , \12157 , \34294_nG9ba5 );
and \U$27145 ( \36006 , \12154 , \34643_nG9ba2 );
or \U$27146 ( \36007 , \36005 , \36006 );
xor \U$27147 ( \36008 , \12153 , \36007 );
buf \U$27148 ( \36009 , \36008 );
buf \U$27150 ( \36010 , \36009 );
xor \U$27151 ( \36011 , \36004 , \36010 );
buf \U$27152 ( \36012 , \36011 );
xor \U$27153 ( \36013 , \35978 , \36012 );
and \U$27154 ( \36014 , \35844 , \35849 );
and \U$27155 ( \36015 , \35844 , \35856 );
and \U$27156 ( \36016 , \35849 , \35856 );
or \U$27157 ( \36017 , \36014 , \36015 , \36016 );
buf \U$27158 ( \36018 , \36017 );
xor \U$27159 ( \36019 , \36013 , \36018 );
buf \U$27160 ( \36020 , \36019 );
xor \U$27161 ( \36021 , \35973 , \36020 );
buf \U$27162 ( \36022 , \36021 );
and \U$27163 ( \36023 , \35599 , \35632 );
and \U$27164 ( \36024 , \35599 , \35860 );
and \U$27165 ( \36025 , \35632 , \35860 );
or \U$27166 ( \36026 , \36023 , \36024 , \36025 );
buf \U$27167 ( \36027 , \36026 );
xor \U$27168 ( \36028 , \36022 , \36027 );
and \U$27169 ( \36029 , \35829 , \35835 );
and \U$27170 ( \36030 , \35829 , \35842 );
and \U$27171 ( \36031 , \35835 , \35842 );
or \U$27172 ( \36032 , \36029 , \36030 , \36031 );
buf \U$27173 ( \36033 , \36032 );
and \U$27174 ( \36034 , \10421 , \35094_nG9b9f );
and \U$27175 ( \36035 , \10418 , \35570_nG9b9c );
or \U$27176 ( \36036 , \36034 , \36035 );
xor \U$27177 ( \36037 , \10417 , \36036 );
buf \U$27178 ( \36038 , \36037 );
buf \U$27180 ( \36039 , \36038 );
xor \U$27181 ( \36040 , \36033 , \36039 );
and \U$27182 ( \36041 , \10707 , \35801_nG9b99 );
and \U$27183 ( \36042 , \35679 , \35713 );
and \U$27184 ( \36043 , \35713 , \35789 );
and \U$27185 ( \36044 , \35679 , \35789 );
or \U$27186 ( \36045 , \36042 , \36043 , \36044 );
and \U$27187 ( \36046 , \35692 , \35696 );
and \U$27188 ( \36047 , \35696 , \35711 );
and \U$27189 ( \36048 , \35692 , \35711 );
or \U$27190 ( \36049 , \36046 , \36047 , \36048 );
and \U$27191 ( \36050 , \27313 , \19534 );
and \U$27192 ( \36051 , \28534 , \19045 );
nor \U$27193 ( \36052 , \36050 , \36051 );
xnor \U$27194 ( \36053 , \36052 , \19540 );
and \U$27195 ( \36054 , \21033 , \25826 );
and \U$27196 ( \36055 , \22090 , \25264 );
nor \U$27197 ( \36056 , \36054 , \36055 );
xnor \U$27198 ( \36057 , \36056 , \25773 );
xor \U$27199 ( \36058 , \36053 , \36057 );
and \U$27200 ( \36059 , \19558 , \27397 );
and \U$27201 ( \36060 , \20544 , \26807 );
nor \U$27202 ( \36061 , \36059 , \36060 );
xnor \U$27203 ( \36062 , \36061 , \27295 );
xor \U$27204 ( \36063 , \36058 , \36062 );
and \U$27205 ( \36064 , \32794 , \15336 );
not \U$27206 ( \36065 , \36064 );
xnor \U$27207 ( \36066 , \36065 , \15342 );
and \U$27208 ( \36067 , \24199 , \22542 );
and \U$27209 ( \36068 , \25272 , \22103 );
nor \U$27210 ( \36069 , \36067 , \36068 );
xnor \U$27211 ( \36070 , \36069 , \22548 );
xor \U$27212 ( \36071 , \36066 , \36070 );
and \U$27213 ( \36072 , \15321 , \32854 );
and \U$27214 ( \36073 , \16267 , \32067 );
nor \U$27215 ( \36074 , \36072 , \36073 );
xnor \U$27216 ( \36075 , \36074 , \32805 );
xor \U$27217 ( \36076 , \36071 , \36075 );
xor \U$27218 ( \36077 , \36063 , \36076 );
and \U$27219 ( \36078 , \25815 , \21005 );
and \U$27220 ( \36079 , \26829 , \20557 );
nor \U$27221 ( \36080 , \36078 , \36079 );
xnor \U$27222 ( \36081 , \36080 , \21011 );
and \U$27223 ( \36082 , \18035 , \29070 );
and \U$27224 ( \36083 , \19032 , \28526 );
nor \U$27225 ( \36084 , \36082 , \36083 );
xnor \U$27226 ( \36085 , \36084 , \29076 );
xor \U$27227 ( \36086 , \36081 , \36085 );
and \U$27228 ( \36087 , \16655 , \30823 );
and \U$27229 ( \36088 , \17627 , \30246 );
nor \U$27230 ( \36089 , \36087 , \36088 );
xnor \U$27231 ( \36090 , \36089 , \30813 );
xor \U$27232 ( \36091 , \36086 , \36090 );
xor \U$27233 ( \36092 , \36077 , \36091 );
xor \U$27234 ( \36093 , \36049 , \36092 );
and \U$27235 ( \36094 , \35701 , \35705 );
and \U$27236 ( \36095 , \35705 , \35710 );
and \U$27237 ( \36096 , \35701 , \35710 );
or \U$27238 ( \36097 , \36094 , \36095 , \36096 );
and \U$27239 ( \36098 , \35780 , \35784 );
and \U$27240 ( \36099 , \35784 , \35786 );
and \U$27241 ( \36100 , \35780 , \35786 );
or \U$27242 ( \36101 , \36098 , \36099 , \36100 );
xor \U$27243 ( \36102 , \36097 , \36101 );
and \U$27244 ( \36103 , \35726 , \35730 );
and \U$27245 ( \36104 , \35730 , \35735 );
and \U$27246 ( \36105 , \35726 , \35735 );
or \U$27247 ( \36106 , \36103 , \36104 , \36105 );
and \U$27248 ( \36107 , \35768 , \35772 );
and \U$27249 ( \36108 , \35772 , \35777 );
and \U$27250 ( \36109 , \35768 , \35777 );
or \U$27251 ( \36110 , \36107 , \36108 , \36109 );
xor \U$27252 ( \36111 , \36106 , \36110 );
and \U$27253 ( \36112 , \30802 , \16635 );
and \U$27254 ( \36113 , \32054 , \16301 );
nor \U$27255 ( \36114 , \36112 , \36113 );
xnor \U$27256 ( \36115 , \36114 , \16625 );
not \U$27257 ( \36116 , \36115 );
xor \U$27258 ( \36117 , \36111 , \36116 );
xor \U$27259 ( \36118 , \36102 , \36117 );
xor \U$27260 ( \36119 , \36093 , \36118 );
xor \U$27261 ( \36120 , \36045 , \36119 );
and \U$27262 ( \36121 , \35683 , \35687 );
and \U$27263 ( \36122 , \35687 , \35712 );
and \U$27264 ( \36123 , \35683 , \35712 );
or \U$27265 ( \36124 , \36121 , \36122 , \36123 );
and \U$27266 ( \36125 , \35718 , \35749 );
and \U$27267 ( \36126 , \35749 , \35788 );
and \U$27268 ( \36127 , \35718 , \35788 );
or \U$27269 ( \36128 , \36125 , \36126 , \36127 );
xor \U$27270 ( \36129 , \36124 , \36128 );
and \U$27271 ( \36130 , \35722 , \35736 );
and \U$27272 ( \36131 , \35736 , \35748 );
and \U$27273 ( \36132 , \35722 , \35748 );
or \U$27274 ( \36133 , \36130 , \36131 , \36132 );
and \U$27275 ( \36134 , \35764 , \35778 );
and \U$27276 ( \36135 , \35778 , \35787 );
and \U$27277 ( \36136 , \35764 , \35787 );
or \U$27278 ( \36137 , \36134 , \36135 , \36136 );
xor \U$27279 ( \36138 , \36133 , \36137 );
and \U$27280 ( \36139 , \35738 , \35742 );
and \U$27281 ( \36140 , \35742 , \35747 );
and \U$27282 ( \36141 , \35738 , \35747 );
or \U$27283 ( \36142 , \36139 , \36140 , \36141 );
and \U$27284 ( \36143 , \35754 , \35758 );
and \U$27285 ( \36144 , \35758 , \35763 );
and \U$27286 ( \36145 , \35754 , \35763 );
or \U$27287 ( \36146 , \36143 , \36144 , \36145 );
xor \U$27288 ( \36147 , \36142 , \36146 );
and \U$27289 ( \36148 , \29084 , \18090 );
and \U$27290 ( \36149 , \30268 , \17655 );
nor \U$27291 ( \36150 , \36148 , \36149 );
xnor \U$27292 ( \36151 , \36150 , \18046 );
and \U$27293 ( \36152 , \22556 , \24138 );
and \U$27294 ( \36153 , \23617 , \23630 );
nor \U$27295 ( \36154 , \36152 , \36153 );
xnor \U$27296 ( \36155 , \36154 , \24144 );
xor \U$27297 ( \36156 , \36151 , \36155 );
and \U$27298 ( \36157 , \14950 , \32802 );
xor \U$27299 ( \36158 , \36156 , \36157 );
xor \U$27300 ( \36159 , \36147 , \36158 );
xor \U$27301 ( \36160 , \36138 , \36159 );
xor \U$27302 ( \36161 , \36129 , \36160 );
xor \U$27303 ( \36162 , \36120 , \36161 );
and \U$27304 ( \36163 , \35670 , \35674 );
and \U$27305 ( \36164 , \35674 , \35790 );
and \U$27306 ( \36165 , \35670 , \35790 );
or \U$27307 ( \36166 , \36163 , \36164 , \36165 );
xor \U$27308 ( \36167 , \36162 , \36166 );
and \U$27309 ( \36168 , \35791 , \35795 );
and \U$27310 ( \36169 , \35796 , \35799 );
or \U$27311 ( \36170 , \36168 , \36169 );
xor \U$27312 ( \36171 , \36167 , \36170 );
buf g9b96 ( \36172_nG9b96 , \36171 );
and \U$27313 ( \36173 , \10704 , \36172_nG9b96 );
or \U$27314 ( \36174 , \36041 , \36173 );
xor \U$27315 ( \36175 , \10703 , \36174 );
buf \U$27316 ( \36176 , \36175 );
buf \U$27318 ( \36177 , \36176 );
xor \U$27319 ( \36178 , \36040 , \36177 );
buf \U$27320 ( \36179 , \36178 );
and \U$27321 ( \36180 , \35658 , \35664 );
and \U$27322 ( \36181 , \35658 , \35806 );
and \U$27323 ( \36182 , \35664 , \35806 );
or \U$27324 ( \36183 , \36180 , \36181 , \36182 );
buf \U$27325 ( \36184 , \36183 );
xor \U$27326 ( \36185 , \36179 , \36184 );
and \U$27327 ( \36186 , \35643 , \35649 );
and \U$27328 ( \36187 , \35643 , \35656 );
and \U$27329 ( \36188 , \35649 , \35656 );
or \U$27330 ( \36189 , \36186 , \36187 , \36188 );
buf \U$27331 ( \36190 , \36189 );
and \U$27333 ( \36191 , \32916 , \14984_nG9bf6 );
or \U$27334 ( \36192 , 1'b0 , \36191 );
xor \U$27335 ( \36193 , 1'b0 , \36192 );
buf \U$27336 ( \36194 , \36193 );
buf \U$27338 ( \36195 , \36194 );
and \U$27339 ( \36196 , \31636 , \15373_nG9bf3 );
and \U$27340 ( \36197 , \31633 , \16315_nG9bf0 );
or \U$27341 ( \36198 , \36196 , \36197 );
xor \U$27342 ( \36199 , \31632 , \36198 );
buf \U$27343 ( \36200 , \36199 );
buf \U$27345 ( \36201 , \36200 );
xor \U$27346 ( \36202 , \36195 , \36201 );
buf \U$27347 ( \36203 , \36202 );
and \U$27348 ( \36204 , \35894 , \35900 );
buf \U$27349 ( \36205 , \36204 );
xor \U$27350 ( \36206 , \36203 , \36205 );
and \U$27351 ( \36207 , \29853 , \16680_nG9bed );
and \U$27352 ( \36208 , \29850 , \17665_nG9bea );
or \U$27353 ( \36209 , \36207 , \36208 );
xor \U$27354 ( \36210 , \29849 , \36209 );
buf \U$27355 ( \36211 , \36210 );
buf \U$27357 ( \36212 , \36211 );
xor \U$27358 ( \36213 , \36206 , \36212 );
buf \U$27359 ( \36214 , \36213 );
and \U$27360 ( \36215 , \35902 , \35904 );
and \U$27361 ( \36216 , \35902 , \35911 );
and \U$27362 ( \36217 , \35904 , \35911 );
or \U$27363 ( \36218 , \36215 , \36216 , \36217 );
buf \U$27364 ( \36219 , \36218 );
xor \U$27365 ( \36220 , \36214 , \36219 );
and \U$27366 ( \36221 , \23201 , \22629_nG9bd5 );
and \U$27367 ( \36222 , \23198 , \23696_nG9bd2 );
or \U$27368 ( \36223 , \36221 , \36222 );
xor \U$27369 ( \36224 , \23197 , \36223 );
buf \U$27370 ( \36225 , \36224 );
buf \U$27372 ( \36226 , \36225 );
xor \U$27373 ( \36227 , \36220 , \36226 );
buf \U$27374 ( \36228 , \36227 );
xor \U$27375 ( \36229 , \36190 , \36228 );
and \U$27376 ( \36230 , \13370 , \33613_nG9bab );
and \U$27377 ( \36231 , \13367 , \34041_nG9ba8 );
or \U$27378 ( \36232 , \36230 , \36231 );
xor \U$27379 ( \36233 , \13366 , \36232 );
buf \U$27380 ( \36234 , \36233 );
buf \U$27382 ( \36235 , \36234 );
xor \U$27383 ( \36236 , \36229 , \36235 );
buf \U$27384 ( \36237 , \36236 );
xor \U$27385 ( \36238 , \36185 , \36237 );
buf \U$27386 ( \36239 , \36238 );
and \U$27387 ( \36240 , \35604 , \35624 );
and \U$27388 ( \36241 , \35604 , \35630 );
and \U$27389 ( \36242 , \35624 , \35630 );
or \U$27390 ( \36243 , \36240 , \36241 , \36242 );
buf \U$27391 ( \36244 , \36243 );
xor \U$27392 ( \36245 , \36239 , \36244 );
and \U$27393 ( \36246 , \35889 , \35913 );
and \U$27394 ( \36247 , \35889 , \35920 );
and \U$27395 ( \36248 , \35913 , \35920 );
or \U$27396 ( \36249 , \36246 , \36247 , \36248 );
buf \U$27397 ( \36250 , \36249 );
and \U$27398 ( \36251 , \17297 , \29179_nG9bbd );
and \U$27399 ( \36252 , \17294 , \30366_nG9bba );
or \U$27400 ( \36253 , \36251 , \36252 );
xor \U$27401 ( \36254 , \17293 , \36253 );
buf \U$27402 ( \36255 , \36254 );
buf \U$27404 ( \36256 , \36255 );
xor \U$27405 ( \36257 , \36250 , \36256 );
and \U$27406 ( \36258 , \14631 , \32888_nG9bb1 );
and \U$27407 ( \36259 , \14628 , \33181_nG9bae );
or \U$27408 ( \36260 , \36258 , \36259 );
xor \U$27409 ( \36261 , \14627 , \36260 );
buf \U$27410 ( \36262 , \36261 );
buf \U$27412 ( \36263 , \36262 );
xor \U$27413 ( \36264 , \36257 , \36263 );
buf \U$27414 ( \36265 , \36264 );
and \U$27415 ( \36266 , \35609 , \35615 );
and \U$27416 ( \36267 , \35609 , \35622 );
and \U$27417 ( \36268 , \35615 , \35622 );
or \U$27418 ( \36269 , \36266 , \36267 , \36268 );
buf \U$27419 ( \36270 , \36269 );
xor \U$27420 ( \36271 , \36265 , \36270 );
and \U$27421 ( \36272 , \28118 , \18107_nG9be7 );
and \U$27422 ( \36273 , \28115 , \19091_nG9be4 );
or \U$27423 ( \36274 , \36272 , \36273 );
xor \U$27424 ( \36275 , \28114 , \36274 );
buf \U$27425 ( \36276 , \36275 );
buf \U$27427 ( \36277 , \36276 );
and \U$27428 ( \36278 , \26431 , \19586_nG9be1 );
and \U$27429 ( \36279 , \26428 , \20608_nG9bde );
or \U$27430 ( \36280 , \36278 , \36279 );
xor \U$27431 ( \36281 , \26427 , \36280 );
buf \U$27432 ( \36282 , \36281 );
buf \U$27434 ( \36283 , \36282 );
xor \U$27435 ( \36284 , \36277 , \36283 );
and \U$27436 ( \36285 , \24792 , \21086_nG9bdb );
and \U$27437 ( \36286 , \24789 , \22129_nG9bd8 );
or \U$27438 ( \36287 , \36285 , \36286 );
xor \U$27439 ( \36288 , \24788 , \36287 );
buf \U$27440 ( \36289 , \36288 );
buf \U$27442 ( \36290 , \36289 );
xor \U$27443 ( \36291 , \36284 , \36290 );
buf \U$27444 ( \36292 , \36291 );
and \U$27445 ( \36293 , \20155 , \25860_nG9bc9 );
and \U$27446 ( \36294 , \20152 , \26887_nG9bc6 );
or \U$27447 ( \36295 , \36293 , \36294 );
xor \U$27448 ( \36296 , \20151 , \36295 );
buf \U$27449 ( \36297 , \36296 );
buf \U$27451 ( \36298 , \36297 );
xor \U$27452 ( \36299 , \36292 , \36298 );
and \U$27453 ( \36300 , \15940 , \30940_nG9bb7 );
and \U$27454 ( \36301 , \15937 , \32179_nG9bb4 );
or \U$27455 ( \36302 , \36300 , \36301 );
xor \U$27456 ( \36303 , \15936 , \36302 );
buf \U$27457 ( \36304 , \36303 );
buf \U$27459 ( \36305 , \36304 );
xor \U$27460 ( \36306 , \36299 , \36305 );
buf \U$27461 ( \36307 , \36306 );
xor \U$27462 ( \36308 , \36271 , \36307 );
buf \U$27463 ( \36309 , \36308 );
xor \U$27464 ( \36310 , \36245 , \36309 );
buf \U$27465 ( \36311 , \36310 );
xor \U$27466 ( \36312 , \36028 , \36311 );
and \U$27467 ( \36313 , \35962 , \36312 );
and \U$27469 ( \36314 , \35956 , \35961 );
or \U$27471 ( \36315 , 1'b0 , \36314 , 1'b0 );
xor \U$27472 ( \36316 , \36313 , \36315 );
and \U$27474 ( \36317 , \35949 , \35955 );
and \U$27475 ( \36318 , \35951 , \35955 );
or \U$27476 ( \36319 , 1'b0 , \36317 , \36318 );
xor \U$27477 ( \36320 , \36316 , \36319 );
xor \U$27484 ( \36321 , \36320 , 1'b0 );
and \U$27485 ( \36322 , \36022 , \36027 );
and \U$27486 ( \36323 , \36022 , \36311 );
and \U$27487 ( \36324 , \36027 , \36311 );
or \U$27488 ( \36325 , \36322 , \36323 , \36324 );
xor \U$27489 ( \36326 , \36321 , \36325 );
and \U$27490 ( \36327 , \35967 , \35972 );
and \U$27491 ( \36328 , \35967 , \36020 );
and \U$27492 ( \36329 , \35972 , \36020 );
or \U$27493 ( \36330 , \36327 , \36328 , \36329 );
buf \U$27494 ( \36331 , \36330 );
and \U$27495 ( \36332 , \36239 , \36244 );
and \U$27496 ( \36333 , \36239 , \36309 );
and \U$27497 ( \36334 , \36244 , \36309 );
or \U$27498 ( \36335 , \36332 , \36333 , \36334 );
buf \U$27499 ( \36336 , \36335 );
and \U$27500 ( \36337 , \36214 , \36219 );
and \U$27501 ( \36338 , \36214 , \36226 );
and \U$27502 ( \36339 , \36219 , \36226 );
or \U$27503 ( \36340 , \36337 , \36338 , \36339 );
buf \U$27504 ( \36341 , \36340 );
and \U$27505 ( \36342 , \36203 , \36205 );
and \U$27506 ( \36343 , \36203 , \36212 );
and \U$27507 ( \36344 , \36205 , \36212 );
or \U$27508 ( \36345 , \36342 , \36343 , \36344 );
buf \U$27509 ( \36346 , \36345 );
and \U$27510 ( \36347 , \28118 , \19091_nG9be4 );
and \U$27511 ( \36348 , \28115 , \19586_nG9be1 );
or \U$27512 ( \36349 , \36347 , \36348 );
xor \U$27513 ( \36350 , \28114 , \36349 );
buf \U$27514 ( \36351 , \36350 );
buf \U$27516 ( \36352 , \36351 );
xor \U$27517 ( \36353 , \36346 , \36352 );
and \U$27518 ( \36354 , \26431 , \20608_nG9bde );
and \U$27519 ( \36355 , \26428 , \21086_nG9bdb );
or \U$27520 ( \36356 , \36354 , \36355 );
xor \U$27521 ( \36357 , \26427 , \36356 );
buf \U$27522 ( \36358 , \36357 );
buf \U$27524 ( \36359 , \36358 );
xor \U$27525 ( \36360 , \36353 , \36359 );
buf \U$27526 ( \36361 , \36360 );
xor \U$27527 ( \36362 , \36341 , \36361 );
and \U$27528 ( \36363 , \18702 , \28602_nG9bc0 );
and \U$27529 ( \36364 , \18699 , \29179_nG9bbd );
or \U$27530 ( \36365 , \36363 , \36364 );
xor \U$27531 ( \36366 , \18698 , \36365 );
buf \U$27532 ( \36367 , \36366 );
buf \U$27534 ( \36368 , \36367 );
xor \U$27535 ( \36369 , \36362 , \36368 );
buf \U$27536 ( \36370 , \36369 );
and \U$27537 ( \36371 , \36292 , \36298 );
and \U$27538 ( \36372 , \36292 , \36305 );
and \U$27539 ( \36373 , \36298 , \36305 );
or \U$27540 ( \36374 , \36371 , \36372 , \36373 );
buf \U$27541 ( \36375 , \36374 );
xor \U$27542 ( \36376 , \36370 , \36375 );
and \U$27544 ( \36377 , \32916 , \15373_nG9bf3 );
or \U$27545 ( \36378 , 1'b0 , \36377 );
xor \U$27546 ( \36379 , 1'b0 , \36378 );
buf \U$27547 ( \36380 , \36379 );
buf \U$27549 ( \36381 , \36380 );
and \U$27550 ( \36382 , \31636 , \16315_nG9bf0 );
and \U$27551 ( \36383 , \31633 , \16680_nG9bed );
or \U$27552 ( \36384 , \36382 , \36383 );
xor \U$27553 ( \36385 , \31632 , \36384 );
buf \U$27554 ( \36386 , \36385 );
buf \U$27556 ( \36387 , \36386 );
xor \U$27557 ( \36388 , \36381 , \36387 );
buf \U$27558 ( \36389 , \36388 );
and \U$27559 ( \36390 , \36195 , \36201 );
buf \U$27560 ( \36391 , \36390 );
xor \U$27561 ( \36392 , \36389 , \36391 );
and \U$27562 ( \36393 , \29853 , \17665_nG9bea );
and \U$27563 ( \36394 , \29850 , \18107_nG9be7 );
or \U$27564 ( \36395 , \36393 , \36394 );
xor \U$27565 ( \36396 , \29849 , \36395 );
buf \U$27566 ( \36397 , \36396 );
buf \U$27568 ( \36398 , \36397 );
xor \U$27569 ( \36399 , \36392 , \36398 );
buf \U$27570 ( \36400 , \36399 );
and \U$27571 ( \36401 , \21658 , \25298_nG9bcc );
and \U$27572 ( \36402 , \21655 , \25860_nG9bc9 );
or \U$27573 ( \36403 , \36401 , \36402 );
xor \U$27574 ( \36404 , \21654 , \36403 );
buf \U$27575 ( \36405 , \36404 );
buf \U$27577 ( \36406 , \36405 );
xor \U$27578 ( \36407 , \36400 , \36406 );
and \U$27579 ( \36408 , \20155 , \26887_nG9bc6 );
and \U$27580 ( \36409 , \20152 , \27416_nG9bc3 );
or \U$27581 ( \36410 , \36408 , \36409 );
xor \U$27582 ( \36411 , \20151 , \36410 );
buf \U$27583 ( \36412 , \36411 );
buf \U$27585 ( \36413 , \36412 );
xor \U$27586 ( \36414 , \36407 , \36413 );
buf \U$27587 ( \36415 , \36414 );
xor \U$27588 ( \36416 , \36376 , \36415 );
buf \U$27589 ( \36417 , \36416 );
and \U$27590 ( \36418 , \35983 , \36003 );
and \U$27591 ( \36419 , \35983 , \36010 );
and \U$27592 ( \36420 , \36003 , \36010 );
or \U$27593 ( \36421 , \36418 , \36419 , \36420 );
buf \U$27594 ( \36422 , \36421 );
xor \U$27595 ( \36423 , \36417 , \36422 );
and \U$27596 ( \36424 , \36265 , \36270 );
and \U$27597 ( \36425 , \36265 , \36307 );
and \U$27598 ( \36426 , \36270 , \36307 );
or \U$27599 ( \36427 , \36424 , \36425 , \36426 );
buf \U$27600 ( \36428 , \36427 );
xor \U$27601 ( \36429 , \36423 , \36428 );
buf \U$27602 ( \36430 , \36429 );
xor \U$27603 ( \36431 , \36336 , \36430 );
and \U$27604 ( \36432 , \36033 , \36039 );
and \U$27605 ( \36433 , \36033 , \36177 );
and \U$27606 ( \36434 , \36039 , \36177 );
or \U$27607 ( \36435 , \36432 , \36433 , \36434 );
buf \U$27608 ( \36436 , \36435 );
and \U$27609 ( \36437 , \36277 , \36283 );
and \U$27610 ( \36438 , \36277 , \36290 );
and \U$27611 ( \36439 , \36283 , \36290 );
or \U$27612 ( \36440 , \36437 , \36438 , \36439 );
buf \U$27613 ( \36441 , \36440 );
and \U$27614 ( \36442 , \24792 , \22129_nG9bd8 );
and \U$27615 ( \36443 , \24789 , \22629_nG9bd5 );
or \U$27616 ( \36444 , \36442 , \36443 );
xor \U$27617 ( \36445 , \24788 , \36444 );
buf \U$27618 ( \36446 , \36445 );
buf \U$27620 ( \36447 , \36446 );
xor \U$27621 ( \36448 , \36441 , \36447 );
and \U$27622 ( \36449 , \23201 , \23696_nG9bd2 );
and \U$27623 ( \36450 , \23198 , \24226_nG9bcf );
or \U$27624 ( \36451 , \36449 , \36450 );
xor \U$27625 ( \36452 , \23197 , \36451 );
buf \U$27626 ( \36453 , \36452 );
buf \U$27628 ( \36454 , \36453 );
xor \U$27629 ( \36455 , \36448 , \36454 );
buf \U$27630 ( \36456 , \36455 );
and \U$27631 ( \36457 , \12157 , \34643_nG9ba2 );
and \U$27632 ( \36458 , \12154 , \35094_nG9b9f );
or \U$27633 ( \36459 , \36457 , \36458 );
xor \U$27634 ( \36460 , \12153 , \36459 );
buf \U$27635 ( \36461 , \36460 );
buf \U$27637 ( \36462 , \36461 );
xor \U$27638 ( \36463 , \36456 , \36462 );
and \U$27639 ( \36464 , \10707 , \36172_nG9b96 );
and \U$27640 ( \36465 , \36124 , \36128 );
and \U$27641 ( \36466 , \36128 , \36160 );
and \U$27642 ( \36467 , \36124 , \36160 );
or \U$27643 ( \36468 , \36465 , \36466 , \36467 );
and \U$27644 ( \36469 , \36097 , \36101 );
and \U$27645 ( \36470 , \36101 , \36117 );
and \U$27646 ( \36471 , \36097 , \36117 );
or \U$27647 ( \36472 , \36469 , \36470 , \36471 );
and \U$27648 ( \36473 , \26829 , \21005 );
and \U$27649 ( \36474 , \27313 , \20557 );
nor \U$27650 ( \36475 , \36473 , \36474 );
xnor \U$27651 ( \36476 , \36475 , \21011 );
and \U$27652 ( \36477 , \22090 , \25826 );
and \U$27653 ( \36478 , \22556 , \25264 );
nor \U$27654 ( \36479 , \36477 , \36478 );
xnor \U$27655 ( \36480 , \36479 , \25773 );
xor \U$27656 ( \36481 , \36476 , \36480 );
and \U$27657 ( \36482 , \20544 , \27397 );
and \U$27658 ( \36483 , \21033 , \26807 );
nor \U$27659 ( \36484 , \36482 , \36483 );
xnor \U$27660 ( \36485 , \36484 , \27295 );
xor \U$27661 ( \36486 , \36481 , \36485 );
not \U$27662 ( \36487 , \15342 );
and \U$27663 ( \36488 , \32054 , \16635 );
and \U$27664 ( \36489 , \32794 , \16301 );
nor \U$27665 ( \36490 , \36488 , \36489 );
xnor \U$27666 ( \36491 , \36490 , \16625 );
xor \U$27667 ( \36492 , \36487 , \36491 );
and \U$27668 ( \36493 , \28534 , \19534 );
and \U$27669 ( \36494 , \29084 , \19045 );
nor \U$27670 ( \36495 , \36493 , \36494 );
xnor \U$27671 ( \36496 , \36495 , \19540 );
xor \U$27672 ( \36497 , \36492 , \36496 );
xor \U$27673 ( \36498 , \36486 , \36497 );
and \U$27674 ( \36499 , \30268 , \18090 );
and \U$27675 ( \36500 , \30802 , \17655 );
nor \U$27676 ( \36501 , \36499 , \36500 );
xnor \U$27677 ( \36502 , \36501 , \18046 );
and \U$27678 ( \36503 , \19032 , \29070 );
and \U$27679 ( \36504 , \19558 , \28526 );
nor \U$27680 ( \36505 , \36503 , \36504 );
xnor \U$27681 ( \36506 , \36505 , \29076 );
xor \U$27682 ( \36507 , \36502 , \36506 );
and \U$27683 ( \36508 , \17627 , \30823 );
and \U$27684 ( \36509 , \18035 , \30246 );
nor \U$27685 ( \36510 , \36508 , \36509 );
xnor \U$27686 ( \36511 , \36510 , \30813 );
xor \U$27687 ( \36512 , \36507 , \36511 );
xor \U$27688 ( \36513 , \36498 , \36512 );
xor \U$27689 ( \36514 , \36472 , \36513 );
and \U$27690 ( \36515 , \36106 , \36110 );
and \U$27691 ( \36516 , \36110 , \36116 );
and \U$27692 ( \36517 , \36106 , \36116 );
or \U$27693 ( \36518 , \36515 , \36516 , \36517 );
and \U$27694 ( \36519 , \25272 , \22542 );
and \U$27695 ( \36520 , \25815 , \22103 );
nor \U$27696 ( \36521 , \36519 , \36520 );
xnor \U$27697 ( \36522 , \36521 , \22548 );
and \U$27698 ( \36523 , \16267 , \32854 );
and \U$27699 ( \36524 , \16655 , \32067 );
nor \U$27700 ( \36525 , \36523 , \36524 );
xnor \U$27701 ( \36526 , \36525 , \32805 );
xor \U$27702 ( \36527 , \36522 , \36526 );
and \U$27703 ( \36528 , \15321 , \32802 );
xor \U$27704 ( \36529 , \36527 , \36528 );
xor \U$27705 ( \36530 , \36518 , \36529 );
and \U$27706 ( \36531 , \36081 , \36085 );
and \U$27707 ( \36532 , \36085 , \36090 );
and \U$27708 ( \36533 , \36081 , \36090 );
or \U$27709 ( \36534 , \36531 , \36532 , \36533 );
buf \U$27710 ( \36535 , \36115 );
xor \U$27711 ( \36536 , \36534 , \36535 );
and \U$27712 ( \36537 , \23617 , \24138 );
and \U$27713 ( \36538 , \24199 , \23630 );
nor \U$27714 ( \36539 , \36537 , \36538 );
xnor \U$27715 ( \36540 , \36539 , \24144 );
xor \U$27716 ( \36541 , \36536 , \36540 );
xor \U$27717 ( \36542 , \36530 , \36541 );
xor \U$27718 ( \36543 , \36514 , \36542 );
xor \U$27719 ( \36544 , \36468 , \36543 );
and \U$27720 ( \36545 , \36133 , \36137 );
and \U$27721 ( \36546 , \36137 , \36159 );
and \U$27722 ( \36547 , \36133 , \36159 );
or \U$27723 ( \36548 , \36545 , \36546 , \36547 );
and \U$27724 ( \36549 , \36049 , \36092 );
and \U$27725 ( \36550 , \36092 , \36118 );
and \U$27726 ( \36551 , \36049 , \36118 );
or \U$27727 ( \36552 , \36549 , \36550 , \36551 );
xor \U$27728 ( \36553 , \36548 , \36552 );
and \U$27729 ( \36554 , \36142 , \36146 );
and \U$27730 ( \36555 , \36146 , \36158 );
and \U$27731 ( \36556 , \36142 , \36158 );
or \U$27732 ( \36557 , \36554 , \36555 , \36556 );
and \U$27733 ( \36558 , \36063 , \36076 );
and \U$27734 ( \36559 , \36076 , \36091 );
and \U$27735 ( \36560 , \36063 , \36091 );
or \U$27736 ( \36561 , \36558 , \36559 , \36560 );
xor \U$27737 ( \36562 , \36557 , \36561 );
and \U$27738 ( \36563 , \36151 , \36155 );
and \U$27739 ( \36564 , \36155 , \36157 );
and \U$27740 ( \36565 , \36151 , \36157 );
or \U$27741 ( \36566 , \36563 , \36564 , \36565 );
and \U$27742 ( \36567 , \36053 , \36057 );
and \U$27743 ( \36568 , \36057 , \36062 );
and \U$27744 ( \36569 , \36053 , \36062 );
or \U$27745 ( \36570 , \36567 , \36568 , \36569 );
xor \U$27746 ( \36571 , \36566 , \36570 );
and \U$27747 ( \36572 , \36066 , \36070 );
and \U$27748 ( \36573 , \36070 , \36075 );
and \U$27749 ( \36574 , \36066 , \36075 );
or \U$27750 ( \36575 , \36572 , \36573 , \36574 );
xor \U$27751 ( \36576 , \36571 , \36575 );
xor \U$27752 ( \36577 , \36562 , \36576 );
xor \U$27753 ( \36578 , \36553 , \36577 );
xor \U$27754 ( \36579 , \36544 , \36578 );
and \U$27755 ( \36580 , \36045 , \36119 );
and \U$27756 ( \36581 , \36119 , \36161 );
and \U$27757 ( \36582 , \36045 , \36161 );
or \U$27758 ( \36583 , \36580 , \36581 , \36582 );
xor \U$27759 ( \36584 , \36579 , \36583 );
and \U$27760 ( \36585 , \36162 , \36166 );
and \U$27761 ( \36586 , \36167 , \36170 );
or \U$27762 ( \36587 , \36585 , \36586 );
xor \U$27763 ( \36588 , \36584 , \36587 );
buf g9b93 ( \36589_nG9b93 , \36588 );
and \U$27764 ( \36590 , \10704 , \36589_nG9b93 );
or \U$27765 ( \36591 , \36464 , \36590 );
xor \U$27766 ( \36592 , \10703 , \36591 );
buf \U$27767 ( \36593 , \36592 );
buf \U$27769 ( \36594 , \36593 );
xor \U$27770 ( \36595 , \36463 , \36594 );
buf \U$27771 ( \36596 , \36595 );
xor \U$27772 ( \36597 , \36436 , \36596 );
and \U$27773 ( \36598 , \35988 , \35994 );
and \U$27774 ( \36599 , \35988 , \36001 );
and \U$27775 ( \36600 , \35994 , \36001 );
or \U$27776 ( \36601 , \36598 , \36599 , \36600 );
buf \U$27777 ( \36602 , \36601 );
and \U$27778 ( \36603 , \13370 , \34041_nG9ba8 );
and \U$27779 ( \36604 , \13367 , \34294_nG9ba5 );
or \U$27780 ( \36605 , \36603 , \36604 );
xor \U$27781 ( \36606 , \13366 , \36605 );
buf \U$27782 ( \36607 , \36606 );
buf \U$27784 ( \36608 , \36607 );
xor \U$27785 ( \36609 , \36602 , \36608 );
and \U$27786 ( \36610 , \10421 , \35570_nG9b9c );
and \U$27787 ( \36611 , \10418 , \35801_nG9b99 );
or \U$27788 ( \36612 , \36610 , \36611 );
xor \U$27789 ( \36613 , \10417 , \36612 );
buf \U$27790 ( \36614 , \36613 );
buf \U$27792 ( \36615 , \36614 );
xor \U$27793 ( \36616 , \36609 , \36615 );
buf \U$27794 ( \36617 , \36616 );
xor \U$27795 ( \36618 , \36597 , \36617 );
buf \U$27796 ( \36619 , \36618 );
xor \U$27797 ( \36620 , \36431 , \36619 );
buf \U$27798 ( \36621 , \36620 );
xor \U$27799 ( \36622 , \36331 , \36621 );
and \U$27800 ( \36623 , \35978 , \36012 );
and \U$27801 ( \36624 , \35978 , \36018 );
and \U$27802 ( \36625 , \36012 , \36018 );
or \U$27803 ( \36626 , \36623 , \36624 , \36625 );
buf \U$27804 ( \36627 , \36626 );
and \U$27805 ( \36628 , \36179 , \36184 );
and \U$27806 ( \36629 , \36179 , \36237 );
and \U$27807 ( \36630 , \36184 , \36237 );
or \U$27808 ( \36631 , \36628 , \36629 , \36630 );
buf \U$27809 ( \36632 , \36631 );
xor \U$27810 ( \36633 , \36627 , \36632 );
and \U$27811 ( \36634 , \17297 , \30366_nG9bba );
and \U$27812 ( \36635 , \17294 , \30940_nG9bb7 );
or \U$27813 ( \36636 , \36634 , \36635 );
xor \U$27814 ( \36637 , \17293 , \36636 );
buf \U$27815 ( \36638 , \36637 );
buf \U$27817 ( \36639 , \36638 );
and \U$27818 ( \36640 , \15940 , \32179_nG9bb4 );
and \U$27819 ( \36641 , \15937 , \32888_nG9bb1 );
or \U$27820 ( \36642 , \36640 , \36641 );
xor \U$27821 ( \36643 , \15936 , \36642 );
buf \U$27822 ( \36644 , \36643 );
buf \U$27824 ( \36645 , \36644 );
xor \U$27825 ( \36646 , \36639 , \36645 );
and \U$27826 ( \36647 , \14631 , \33181_nG9bae );
and \U$27827 ( \36648 , \14628 , \33613_nG9bab );
or \U$27828 ( \36649 , \36647 , \36648 );
xor \U$27829 ( \36650 , \14627 , \36649 );
buf \U$27830 ( \36651 , \36650 );
buf \U$27832 ( \36652 , \36651 );
xor \U$27833 ( \36653 , \36646 , \36652 );
buf \U$27834 ( \36654 , \36653 );
and \U$27835 ( \36655 , \36190 , \36228 );
and \U$27836 ( \36656 , \36190 , \36235 );
and \U$27837 ( \36657 , \36228 , \36235 );
or \U$27838 ( \36658 , \36655 , \36656 , \36657 );
buf \U$27839 ( \36659 , \36658 );
xor \U$27840 ( \36660 , \36654 , \36659 );
and \U$27841 ( \36661 , \36250 , \36256 );
and \U$27842 ( \36662 , \36250 , \36263 );
and \U$27843 ( \36663 , \36256 , \36263 );
or \U$27844 ( \36664 , \36661 , \36662 , \36663 );
buf \U$27845 ( \36665 , \36664 );
xor \U$27846 ( \36666 , \36660 , \36665 );
buf \U$27847 ( \36667 , \36666 );
xor \U$27848 ( \36668 , \36633 , \36667 );
buf \U$27849 ( \36669 , \36668 );
xor \U$27850 ( \36670 , \36622 , \36669 );
and \U$27851 ( \36671 , \36326 , \36670 );
and \U$27853 ( \36672 , \36320 , \36325 );
or \U$27855 ( \36673 , 1'b0 , \36672 , 1'b0 );
xor \U$27856 ( \36674 , \36671 , \36673 );
and \U$27858 ( \36675 , \36313 , \36319 );
and \U$27859 ( \36676 , \36315 , \36319 );
or \U$27860 ( \36677 , 1'b0 , \36675 , \36676 );
xor \U$27861 ( \36678 , \36674 , \36677 );
xor \U$27868 ( \36679 , \36678 , 1'b0 );
and \U$27869 ( \36680 , \36331 , \36621 );
and \U$27870 ( \36681 , \36331 , \36669 );
and \U$27871 ( \36682 , \36621 , \36669 );
or \U$27872 ( \36683 , \36680 , \36681 , \36682 );
xor \U$27873 ( \36684 , \36679 , \36683 );
and \U$27874 ( \36685 , \36336 , \36430 );
and \U$27875 ( \36686 , \36336 , \36619 );
and \U$27876 ( \36687 , \36430 , \36619 );
or \U$27877 ( \36688 , \36685 , \36686 , \36687 );
buf \U$27878 ( \36689 , \36688 );
and \U$27879 ( \36690 , \36417 , \36422 );
and \U$27880 ( \36691 , \36417 , \36428 );
and \U$27881 ( \36692 , \36422 , \36428 );
or \U$27882 ( \36693 , \36690 , \36691 , \36692 );
buf \U$27883 ( \36694 , \36693 );
and \U$27884 ( \36695 , \36436 , \36596 );
and \U$27885 ( \36696 , \36436 , \36617 );
and \U$27886 ( \36697 , \36596 , \36617 );
or \U$27887 ( \36698 , \36695 , \36696 , \36697 );
buf \U$27888 ( \36699 , \36698 );
xor \U$27889 ( \36700 , \36694 , \36699 );
and \U$27890 ( \36701 , \36441 , \36447 );
and \U$27891 ( \36702 , \36441 , \36454 );
and \U$27892 ( \36703 , \36447 , \36454 );
or \U$27893 ( \36704 , \36701 , \36702 , \36703 );
buf \U$27894 ( \36705 , \36704 );
and \U$27895 ( \36706 , \15940 , \32888_nG9bb1 );
and \U$27896 ( \36707 , \15937 , \33181_nG9bae );
or \U$27897 ( \36708 , \36706 , \36707 );
xor \U$27898 ( \36709 , \15936 , \36708 );
buf \U$27899 ( \36710 , \36709 );
buf \U$27901 ( \36711 , \36710 );
xor \U$27902 ( \36712 , \36705 , \36711 );
and \U$27903 ( \36713 , \14631 , \33613_nG9bab );
and \U$27904 ( \36714 , \14628 , \34041_nG9ba8 );
or \U$27905 ( \36715 , \36713 , \36714 );
xor \U$27906 ( \36716 , \14627 , \36715 );
buf \U$27907 ( \36717 , \36716 );
buf \U$27909 ( \36718 , \36717 );
xor \U$27910 ( \36719 , \36712 , \36718 );
buf \U$27911 ( \36720 , \36719 );
and \U$27912 ( \36721 , \36389 , \36391 );
and \U$27913 ( \36722 , \36389 , \36398 );
and \U$27914 ( \36723 , \36391 , \36398 );
or \U$27915 ( \36724 , \36721 , \36722 , \36723 );
buf \U$27916 ( \36725 , \36724 );
and \U$27917 ( \36726 , \28118 , \19586_nG9be1 );
and \U$27918 ( \36727 , \28115 , \20608_nG9bde );
or \U$27919 ( \36728 , \36726 , \36727 );
xor \U$27920 ( \36729 , \28114 , \36728 );
buf \U$27921 ( \36730 , \36729 );
buf \U$27923 ( \36731 , \36730 );
xor \U$27924 ( \36732 , \36725 , \36731 );
and \U$27925 ( \36733 , \26431 , \21086_nG9bdb );
and \U$27926 ( \36734 , \26428 , \22129_nG9bd8 );
or \U$27927 ( \36735 , \36733 , \36734 );
xor \U$27928 ( \36736 , \26427 , \36735 );
buf \U$27929 ( \36737 , \36736 );
buf \U$27931 ( \36738 , \36737 );
xor \U$27932 ( \36739 , \36732 , \36738 );
buf \U$27933 ( \36740 , \36739 );
and \U$27934 ( \36741 , \18702 , \29179_nG9bbd );
and \U$27935 ( \36742 , \18699 , \30366_nG9bba );
or \U$27936 ( \36743 , \36741 , \36742 );
xor \U$27937 ( \36744 , \18698 , \36743 );
buf \U$27938 ( \36745 , \36744 );
buf \U$27940 ( \36746 , \36745 );
xor \U$27941 ( \36747 , \36740 , \36746 );
and \U$27942 ( \36748 , \17297 , \30940_nG9bb7 );
and \U$27943 ( \36749 , \17294 , \32179_nG9bb4 );
or \U$27944 ( \36750 , \36748 , \36749 );
xor \U$27945 ( \36751 , \17293 , \36750 );
buf \U$27946 ( \36752 , \36751 );
buf \U$27948 ( \36753 , \36752 );
xor \U$27949 ( \36754 , \36747 , \36753 );
buf \U$27950 ( \36755 , \36754 );
xor \U$27951 ( \36756 , \36720 , \36755 );
and \U$27952 ( \36757 , \36602 , \36608 );
and \U$27953 ( \36758 , \36602 , \36615 );
and \U$27954 ( \36759 , \36608 , \36615 );
or \U$27955 ( \36760 , \36757 , \36758 , \36759 );
buf \U$27956 ( \36761 , \36760 );
xor \U$27957 ( \36762 , \36756 , \36761 );
buf \U$27958 ( \36763 , \36762 );
xor \U$27959 ( \36764 , \36700 , \36763 );
buf \U$27960 ( \36765 , \36764 );
xor \U$27961 ( \36766 , \36689 , \36765 );
and \U$27962 ( \36767 , \36627 , \36632 );
and \U$27963 ( \36768 , \36627 , \36667 );
and \U$27964 ( \36769 , \36632 , \36667 );
or \U$27965 ( \36770 , \36767 , \36768 , \36769 );
buf \U$27966 ( \36771 , \36770 );
and \U$27967 ( \36772 , \36654 , \36659 );
and \U$27968 ( \36773 , \36654 , \36665 );
and \U$27969 ( \36774 , \36659 , \36665 );
or \U$27970 ( \36775 , \36772 , \36773 , \36774 );
buf \U$27971 ( \36776 , \36775 );
and \U$27972 ( \36777 , \36639 , \36645 );
and \U$27973 ( \36778 , \36639 , \36652 );
and \U$27974 ( \36779 , \36645 , \36652 );
or \U$27975 ( \36780 , \36777 , \36778 , \36779 );
buf \U$27976 ( \36781 , \36780 );
and \U$27977 ( \36782 , \36341 , \36361 );
and \U$27978 ( \36783 , \36341 , \36368 );
and \U$27979 ( \36784 , \36361 , \36368 );
or \U$27980 ( \36785 , \36782 , \36783 , \36784 );
buf \U$27981 ( \36786 , \36785 );
xor \U$27982 ( \36787 , \36781 , \36786 );
and \U$27983 ( \36788 , \36346 , \36352 );
and \U$27984 ( \36789 , \36346 , \36359 );
and \U$27985 ( \36790 , \36352 , \36359 );
or \U$27986 ( \36791 , \36788 , \36789 , \36790 );
buf \U$27987 ( \36792 , \36791 );
and \U$27988 ( \36793 , \21658 , \25860_nG9bc9 );
and \U$27989 ( \36794 , \21655 , \26887_nG9bc6 );
or \U$27990 ( \36795 , \36793 , \36794 );
xor \U$27991 ( \36796 , \21654 , \36795 );
buf \U$27992 ( \36797 , \36796 );
buf \U$27994 ( \36798 , \36797 );
xor \U$27995 ( \36799 , \36792 , \36798 );
and \U$27996 ( \36800 , \20155 , \27416_nG9bc3 );
and \U$27997 ( \36801 , \20152 , \28602_nG9bc0 );
or \U$27998 ( \36802 , \36800 , \36801 );
xor \U$27999 ( \36803 , \20151 , \36802 );
buf \U$28000 ( \36804 , \36803 );
buf \U$28002 ( \36805 , \36804 );
xor \U$28003 ( \36806 , \36799 , \36805 );
buf \U$28004 ( \36807 , \36806 );
xor \U$28005 ( \36808 , \36787 , \36807 );
buf \U$28006 ( \36809 , \36808 );
xor \U$28007 ( \36810 , \36776 , \36809 );
and \U$28008 ( \36811 , \36370 , \36375 );
and \U$28009 ( \36812 , \36370 , \36415 );
and \U$28010 ( \36813 , \36375 , \36415 );
or \U$28011 ( \36814 , \36811 , \36812 , \36813 );
buf \U$28012 ( \36815 , \36814 );
xor \U$28013 ( \36816 , \36810 , \36815 );
buf \U$28014 ( \36817 , \36816 );
xor \U$28015 ( \36818 , \36771 , \36817 );
and \U$28017 ( \36819 , \32916 , \16315_nG9bf0 );
or \U$28018 ( \36820 , 1'b0 , \36819 );
xor \U$28019 ( \36821 , 1'b0 , \36820 );
buf \U$28020 ( \36822 , \36821 );
buf \U$28022 ( \36823 , \36822 );
and \U$28023 ( \36824 , \31636 , \16680_nG9bed );
and \U$28024 ( \36825 , \31633 , \17665_nG9bea );
or \U$28025 ( \36826 , \36824 , \36825 );
xor \U$28026 ( \36827 , \31632 , \36826 );
buf \U$28027 ( \36828 , \36827 );
buf \U$28029 ( \36829 , \36828 );
xor \U$28030 ( \36830 , \36823 , \36829 );
buf \U$28031 ( \36831 , \36830 );
and \U$28032 ( \36832 , \36381 , \36387 );
buf \U$28033 ( \36833 , \36832 );
xor \U$28034 ( \36834 , \36831 , \36833 );
and \U$28035 ( \36835 , \29853 , \18107_nG9be7 );
and \U$28036 ( \36836 , \29850 , \19091_nG9be4 );
or \U$28037 ( \36837 , \36835 , \36836 );
xor \U$28038 ( \36838 , \29849 , \36837 );
buf \U$28039 ( \36839 , \36838 );
buf \U$28041 ( \36840 , \36839 );
xor \U$28042 ( \36841 , \36834 , \36840 );
buf \U$28043 ( \36842 , \36841 );
and \U$28044 ( \36843 , \24792 , \22629_nG9bd5 );
and \U$28045 ( \36844 , \24789 , \23696_nG9bd2 );
or \U$28046 ( \36845 , \36843 , \36844 );
xor \U$28047 ( \36846 , \24788 , \36845 );
buf \U$28048 ( \36847 , \36846 );
buf \U$28050 ( \36848 , \36847 );
xor \U$28051 ( \36849 , \36842 , \36848 );
and \U$28052 ( \36850 , \23201 , \24226_nG9bcf );
and \U$28053 ( \36851 , \23198 , \25298_nG9bcc );
or \U$28054 ( \36852 , \36850 , \36851 );
xor \U$28055 ( \36853 , \23197 , \36852 );
buf \U$28056 ( \36854 , \36853 );
buf \U$28058 ( \36855 , \36854 );
xor \U$28059 ( \36856 , \36849 , \36855 );
buf \U$28060 ( \36857 , \36856 );
and \U$28061 ( \36858 , \12157 , \35094_nG9b9f );
and \U$28062 ( \36859 , \12154 , \35570_nG9b9c );
or \U$28063 ( \36860 , \36858 , \36859 );
xor \U$28064 ( \36861 , \12153 , \36860 );
buf \U$28065 ( \36862 , \36861 );
buf \U$28067 ( \36863 , \36862 );
xor \U$28068 ( \36864 , \36857 , \36863 );
and \U$28069 ( \36865 , \10707 , \36589_nG9b93 );
and \U$28070 ( \36866 , \36548 , \36552 );
and \U$28071 ( \36867 , \36552 , \36577 );
and \U$28072 ( \36868 , \36548 , \36577 );
or \U$28073 ( \36869 , \36866 , \36867 , \36868 );
and \U$28074 ( \36870 , \36518 , \36529 );
and \U$28075 ( \36871 , \36529 , \36541 );
and \U$28076 ( \36872 , \36518 , \36541 );
or \U$28077 ( \36873 , \36870 , \36871 , \36872 );
and \U$28078 ( \36874 , \36476 , \36480 );
and \U$28079 ( \36875 , \36480 , \36485 );
and \U$28080 ( \36876 , \36476 , \36485 );
or \U$28081 ( \36877 , \36874 , \36875 , \36876 );
and \U$28082 ( \36878 , \32794 , \16635 );
not \U$28083 ( \36879 , \36878 );
xnor \U$28084 ( \36880 , \36879 , \16625 );
and \U$28085 ( \36881 , \29084 , \19534 );
and \U$28086 ( \36882 , \30268 , \19045 );
nor \U$28087 ( \36883 , \36881 , \36882 );
xnor \U$28088 ( \36884 , \36883 , \19540 );
xor \U$28089 ( \36885 , \36880 , \36884 );
and \U$28090 ( \36886 , \16267 , \32802 );
xor \U$28091 ( \36887 , \36885 , \36886 );
xor \U$28092 ( \36888 , \36877 , \36887 );
and \U$28093 ( \36889 , \27313 , \21005 );
and \U$28094 ( \36890 , \28534 , \20557 );
nor \U$28095 ( \36891 , \36889 , \36890 );
xnor \U$28096 ( \36892 , \36891 , \21011 );
and \U$28097 ( \36893 , \21033 , \27397 );
and \U$28098 ( \36894 , \22090 , \26807 );
nor \U$28099 ( \36895 , \36893 , \36894 );
xnor \U$28100 ( \36896 , \36895 , \27295 );
xor \U$28101 ( \36897 , \36892 , \36896 );
and \U$28102 ( \36898 , \19558 , \29070 );
and \U$28103 ( \36899 , \20544 , \28526 );
nor \U$28104 ( \36900 , \36898 , \36899 );
xnor \U$28105 ( \36901 , \36900 , \29076 );
xor \U$28106 ( \36902 , \36897 , \36901 );
xor \U$28107 ( \36903 , \36888 , \36902 );
xor \U$28108 ( \36904 , \36873 , \36903 );
and \U$28109 ( \36905 , \36566 , \36570 );
and \U$28110 ( \36906 , \36570 , \36575 );
and \U$28111 ( \36907 , \36566 , \36575 );
or \U$28112 ( \36908 , \36905 , \36906 , \36907 );
and \U$28113 ( \36909 , \25815 , \22542 );
and \U$28114 ( \36910 , \26829 , \22103 );
nor \U$28115 ( \36911 , \36909 , \36910 );
xnor \U$28116 ( \36912 , \36911 , \22548 );
and \U$28117 ( \36913 , \18035 , \30823 );
and \U$28118 ( \36914 , \19032 , \30246 );
nor \U$28119 ( \36915 , \36913 , \36914 );
xnor \U$28120 ( \36916 , \36915 , \30813 );
xor \U$28121 ( \36917 , \36912 , \36916 );
and \U$28122 ( \36918 , \16655 , \32854 );
and \U$28123 ( \36919 , \17627 , \32067 );
nor \U$28124 ( \36920 , \36918 , \36919 );
xnor \U$28125 ( \36921 , \36920 , \32805 );
xor \U$28126 ( \36922 , \36917 , \36921 );
xor \U$28127 ( \36923 , \36908 , \36922 );
and \U$28128 ( \36924 , \30802 , \18090 );
and \U$28129 ( \36925 , \32054 , \17655 );
nor \U$28130 ( \36926 , \36924 , \36925 );
xnor \U$28131 ( \36927 , \36926 , \18046 );
not \U$28132 ( \36928 , \36927 );
and \U$28133 ( \36929 , \24199 , \24138 );
and \U$28134 ( \36930 , \25272 , \23630 );
nor \U$28135 ( \36931 , \36929 , \36930 );
xnor \U$28136 ( \36932 , \36931 , \24144 );
xor \U$28137 ( \36933 , \36928 , \36932 );
and \U$28138 ( \36934 , \22556 , \25826 );
and \U$28139 ( \36935 , \23617 , \25264 );
nor \U$28140 ( \36936 , \36934 , \36935 );
xnor \U$28141 ( \36937 , \36936 , \25773 );
xor \U$28142 ( \36938 , \36933 , \36937 );
xor \U$28143 ( \36939 , \36923 , \36938 );
xor \U$28144 ( \36940 , \36904 , \36939 );
xor \U$28145 ( \36941 , \36869 , \36940 );
and \U$28146 ( \36942 , \36557 , \36561 );
and \U$28147 ( \36943 , \36561 , \36576 );
and \U$28148 ( \36944 , \36557 , \36576 );
or \U$28149 ( \36945 , \36942 , \36943 , \36944 );
and \U$28150 ( \36946 , \36472 , \36513 );
and \U$28151 ( \36947 , \36513 , \36542 );
and \U$28152 ( \36948 , \36472 , \36542 );
or \U$28153 ( \36949 , \36946 , \36947 , \36948 );
xor \U$28154 ( \36950 , \36945 , \36949 );
and \U$28155 ( \36951 , \36534 , \36535 );
and \U$28156 ( \36952 , \36535 , \36540 );
and \U$28157 ( \36953 , \36534 , \36540 );
or \U$28158 ( \36954 , \36951 , \36952 , \36953 );
and \U$28159 ( \36955 , \36486 , \36497 );
and \U$28160 ( \36956 , \36497 , \36512 );
and \U$28161 ( \36957 , \36486 , \36512 );
or \U$28162 ( \36958 , \36955 , \36956 , \36957 );
xor \U$28163 ( \36959 , \36954 , \36958 );
and \U$28164 ( \36960 , \36522 , \36526 );
and \U$28165 ( \36961 , \36526 , \36528 );
and \U$28166 ( \36962 , \36522 , \36528 );
or \U$28167 ( \36963 , \36960 , \36961 , \36962 );
and \U$28168 ( \36964 , \36487 , \36491 );
and \U$28169 ( \36965 , \36491 , \36496 );
and \U$28170 ( \36966 , \36487 , \36496 );
or \U$28171 ( \36967 , \36964 , \36965 , \36966 );
xor \U$28172 ( \36968 , \36963 , \36967 );
and \U$28173 ( \36969 , \36502 , \36506 );
and \U$28174 ( \36970 , \36506 , \36511 );
and \U$28175 ( \36971 , \36502 , \36511 );
or \U$28176 ( \36972 , \36969 , \36970 , \36971 );
xor \U$28177 ( \36973 , \36968 , \36972 );
xor \U$28178 ( \36974 , \36959 , \36973 );
xor \U$28179 ( \36975 , \36950 , \36974 );
xor \U$28180 ( \36976 , \36941 , \36975 );
and \U$28181 ( \36977 , \36468 , \36543 );
and \U$28182 ( \36978 , \36543 , \36578 );
and \U$28183 ( \36979 , \36468 , \36578 );
or \U$28184 ( \36980 , \36977 , \36978 , \36979 );
xor \U$28185 ( \36981 , \36976 , \36980 );
and \U$28186 ( \36982 , \36579 , \36583 );
and \U$28187 ( \36983 , \36584 , \36587 );
or \U$28188 ( \36984 , \36982 , \36983 );
xor \U$28189 ( \36985 , \36981 , \36984 );
buf g9b90 ( \36986_nG9b90 , \36985 );
and \U$28190 ( \36987 , \10704 , \36986_nG9b90 );
or \U$28191 ( \36988 , \36865 , \36987 );
xor \U$28192 ( \36989 , \10703 , \36988 );
buf \U$28193 ( \36990 , \36989 );
buf \U$28195 ( \36991 , \36990 );
xor \U$28196 ( \36992 , \36864 , \36991 );
buf \U$28197 ( \36993 , \36992 );
and \U$28198 ( \36994 , \36400 , \36406 );
and \U$28199 ( \36995 , \36400 , \36413 );
and \U$28200 ( \36996 , \36406 , \36413 );
or \U$28201 ( \36997 , \36994 , \36995 , \36996 );
buf \U$28202 ( \36998 , \36997 );
and \U$28203 ( \36999 , \13370 , \34294_nG9ba5 );
and \U$28204 ( \37000 , \13367 , \34643_nG9ba2 );
or \U$28205 ( \37001 , \36999 , \37000 );
xor \U$28206 ( \37002 , \13366 , \37001 );
buf \U$28207 ( \37003 , \37002 );
buf \U$28209 ( \37004 , \37003 );
xor \U$28210 ( \37005 , \36998 , \37004 );
and \U$28211 ( \37006 , \10421 , \35801_nG9b99 );
and \U$28212 ( \37007 , \10418 , \36172_nG9b96 );
or \U$28213 ( \37008 , \37006 , \37007 );
xor \U$28214 ( \37009 , \10417 , \37008 );
buf \U$28215 ( \37010 , \37009 );
buf \U$28217 ( \37011 , \37010 );
xor \U$28218 ( \37012 , \37005 , \37011 );
buf \U$28219 ( \37013 , \37012 );
xor \U$28220 ( \37014 , \36993 , \37013 );
and \U$28221 ( \37015 , \36456 , \36462 );
and \U$28222 ( \37016 , \36456 , \36594 );
and \U$28223 ( \37017 , \36462 , \36594 );
or \U$28224 ( \37018 , \37015 , \37016 , \37017 );
buf \U$28225 ( \37019 , \37018 );
xor \U$28226 ( \37020 , \37014 , \37019 );
buf \U$28227 ( \37021 , \37020 );
xor \U$28228 ( \37022 , \36818 , \37021 );
buf \U$28229 ( \37023 , \37022 );
xor \U$28230 ( \37024 , \36766 , \37023 );
and \U$28231 ( \37025 , \36684 , \37024 );
and \U$28233 ( \37026 , \36678 , \36683 );
or \U$28235 ( \37027 , 1'b0 , \37026 , 1'b0 );
xor \U$28236 ( \37028 , \37025 , \37027 );
and \U$28238 ( \37029 , \36671 , \36677 );
and \U$28239 ( \37030 , \36673 , \36677 );
or \U$28240 ( \37031 , 1'b0 , \37029 , \37030 );
xor \U$28241 ( \37032 , \37028 , \37031 );
xor \U$28248 ( \37033 , \37032 , 1'b0 );
and \U$28249 ( \37034 , \36689 , \36765 );
and \U$28250 ( \37035 , \36689 , \37023 );
and \U$28251 ( \37036 , \36765 , \37023 );
or \U$28252 ( \37037 , \37034 , \37035 , \37036 );
xor \U$28253 ( \37038 , \37033 , \37037 );
and \U$28254 ( \37039 , \36771 , \36817 );
and \U$28255 ( \37040 , \36771 , \37021 );
and \U$28256 ( \37041 , \36817 , \37021 );
or \U$28257 ( \37042 , \37039 , \37040 , \37041 );
buf \U$28258 ( \37043 , \37042 );
and \U$28259 ( \37044 , \36781 , \36786 );
and \U$28260 ( \37045 , \36781 , \36807 );
and \U$28261 ( \37046 , \36786 , \36807 );
or \U$28262 ( \37047 , \37044 , \37045 , \37046 );
buf \U$28263 ( \37048 , \37047 );
and \U$28264 ( \37049 , \36725 , \36731 );
and \U$28265 ( \37050 , \36725 , \36738 );
and \U$28266 ( \37051 , \36731 , \36738 );
or \U$28267 ( \37052 , \37049 , \37050 , \37051 );
buf \U$28268 ( \37053 , \37052 );
and \U$28269 ( \37054 , \36823 , \36829 );
buf \U$28270 ( \37055 , \37054 );
and \U$28271 ( \37056 , \29853 , \19091_nG9be4 );
and \U$28272 ( \37057 , \29850 , \19586_nG9be1 );
or \U$28273 ( \37058 , \37056 , \37057 );
xor \U$28274 ( \37059 , \29849 , \37058 );
buf \U$28275 ( \37060 , \37059 );
buf \U$28277 ( \37061 , \37060 );
xor \U$28278 ( \37062 , \37055 , \37061 );
and \U$28279 ( \37063 , \28118 , \20608_nG9bde );
and \U$28280 ( \37064 , \28115 , \21086_nG9bdb );
or \U$28281 ( \37065 , \37063 , \37064 );
xor \U$28282 ( \37066 , \28114 , \37065 );
buf \U$28283 ( \37067 , \37066 );
buf \U$28285 ( \37068 , \37067 );
xor \U$28286 ( \37069 , \37062 , \37068 );
buf \U$28287 ( \37070 , \37069 );
xor \U$28288 ( \37071 , \37053 , \37070 );
and \U$28289 ( \37072 , \18702 , \30366_nG9bba );
and \U$28290 ( \37073 , \18699 , \30940_nG9bb7 );
or \U$28291 ( \37074 , \37072 , \37073 );
xor \U$28292 ( \37075 , \18698 , \37074 );
buf \U$28293 ( \37076 , \37075 );
buf \U$28295 ( \37077 , \37076 );
xor \U$28296 ( \37078 , \37071 , \37077 );
buf \U$28297 ( \37079 , \37078 );
and \U$28298 ( \37080 , \24792 , \23696_nG9bd2 );
and \U$28299 ( \37081 , \24789 , \24226_nG9bcf );
or \U$28300 ( \37082 , \37080 , \37081 );
xor \U$28301 ( \37083 , \24788 , \37082 );
buf \U$28302 ( \37084 , \37083 );
buf \U$28304 ( \37085 , \37084 );
and \U$28305 ( \37086 , \23201 , \25298_nG9bcc );
and \U$28306 ( \37087 , \23198 , \25860_nG9bc9 );
or \U$28307 ( \37088 , \37086 , \37087 );
xor \U$28308 ( \37089 , \23197 , \37088 );
buf \U$28309 ( \37090 , \37089 );
buf \U$28311 ( \37091 , \37090 );
xor \U$28312 ( \37092 , \37085 , \37091 );
and \U$28313 ( \37093 , \21658 , \26887_nG9bc6 );
and \U$28314 ( \37094 , \21655 , \27416_nG9bc3 );
or \U$28315 ( \37095 , \37093 , \37094 );
xor \U$28316 ( \37096 , \21654 , \37095 );
buf \U$28317 ( \37097 , \37096 );
buf \U$28319 ( \37098 , \37097 );
xor \U$28320 ( \37099 , \37092 , \37098 );
buf \U$28321 ( \37100 , \37099 );
xor \U$28322 ( \37101 , \37079 , \37100 );
and \U$28323 ( \37102 , \36705 , \36711 );
and \U$28324 ( \37103 , \36705 , \36718 );
and \U$28325 ( \37104 , \36711 , \36718 );
or \U$28326 ( \37105 , \37102 , \37103 , \37104 );
buf \U$28327 ( \37106 , \37105 );
xor \U$28328 ( \37107 , \37101 , \37106 );
buf \U$28329 ( \37108 , \37107 );
xor \U$28330 ( \37109 , \37048 , \37108 );
and \U$28331 ( \37110 , \36720 , \36755 );
and \U$28332 ( \37111 , \36720 , \36761 );
and \U$28333 ( \37112 , \36755 , \36761 );
or \U$28334 ( \37113 , \37110 , \37111 , \37112 );
buf \U$28335 ( \37114 , \37113 );
xor \U$28336 ( \37115 , \37109 , \37114 );
buf \U$28337 ( \37116 , \37115 );
and \U$28338 ( \37117 , \36776 , \36809 );
and \U$28339 ( \37118 , \36776 , \36815 );
and \U$28340 ( \37119 , \36809 , \36815 );
or \U$28341 ( \37120 , \37117 , \37118 , \37119 );
buf \U$28342 ( \37121 , \37120 );
xor \U$28343 ( \37122 , \37116 , \37121 );
and \U$28344 ( \37123 , \36740 , \36746 );
and \U$28345 ( \37124 , \36740 , \36753 );
and \U$28346 ( \37125 , \36746 , \36753 );
or \U$28347 ( \37126 , \37123 , \37124 , \37125 );
buf \U$28348 ( \37127 , \37126 );
and \U$28349 ( \37128 , \10421 , \36172_nG9b96 );
and \U$28350 ( \37129 , \10418 , \36589_nG9b93 );
or \U$28351 ( \37130 , \37128 , \37129 );
xor \U$28352 ( \37131 , \10417 , \37130 );
buf \U$28353 ( \37132 , \37131 );
buf \U$28355 ( \37133 , \37132 );
xor \U$28356 ( \37134 , \37127 , \37133 );
and \U$28357 ( \37135 , \10707 , \36986_nG9b90 );
and \U$28358 ( \37136 , \36945 , \36949 );
and \U$28359 ( \37137 , \36949 , \36974 );
and \U$28360 ( \37138 , \36945 , \36974 );
or \U$28361 ( \37139 , \37136 , \37137 , \37138 );
and \U$28362 ( \37140 , \36908 , \36922 );
and \U$28363 ( \37141 , \36922 , \36938 );
and \U$28364 ( \37142 , \36908 , \36938 );
or \U$28365 ( \37143 , \37140 , \37141 , \37142 );
and \U$28366 ( \37144 , \36928 , \36932 );
and \U$28367 ( \37145 , \36932 , \36937 );
and \U$28368 ( \37146 , \36928 , \36937 );
or \U$28369 ( \37147 , \37144 , \37145 , \37146 );
not \U$28370 ( \37148 , \16625 );
and \U$28371 ( \37149 , \32054 , \18090 );
and \U$28372 ( \37150 , \32794 , \17655 );
nor \U$28373 ( \37151 , \37149 , \37150 );
xnor \U$28374 ( \37152 , \37151 , \18046 );
xor \U$28375 ( \37153 , \37148 , \37152 );
and \U$28376 ( \37154 , \28534 , \21005 );
and \U$28377 ( \37155 , \29084 , \20557 );
nor \U$28378 ( \37156 , \37154 , \37155 );
xnor \U$28379 ( \37157 , \37156 , \21011 );
xor \U$28380 ( \37158 , \37153 , \37157 );
xor \U$28381 ( \37159 , \37147 , \37158 );
and \U$28382 ( \37160 , \26829 , \22542 );
and \U$28383 ( \37161 , \27313 , \22103 );
nor \U$28384 ( \37162 , \37160 , \37161 );
xnor \U$28385 ( \37163 , \37162 , \22548 );
and \U$28386 ( \37164 , \22090 , \27397 );
and \U$28387 ( \37165 , \22556 , \26807 );
nor \U$28388 ( \37166 , \37164 , \37165 );
xnor \U$28389 ( \37167 , \37166 , \27295 );
xor \U$28390 ( \37168 , \37163 , \37167 );
and \U$28391 ( \37169 , \20544 , \29070 );
and \U$28392 ( \37170 , \21033 , \28526 );
nor \U$28393 ( \37171 , \37169 , \37170 );
xnor \U$28394 ( \37172 , \37171 , \29076 );
xor \U$28395 ( \37173 , \37168 , \37172 );
xor \U$28396 ( \37174 , \37159 , \37173 );
xor \U$28397 ( \37175 , \37143 , \37174 );
and \U$28398 ( \37176 , \36912 , \36916 );
and \U$28399 ( \37177 , \36916 , \36921 );
and \U$28400 ( \37178 , \36912 , \36921 );
or \U$28401 ( \37179 , \37176 , \37177 , \37178 );
and \U$28402 ( \37180 , \30268 , \19534 );
and \U$28403 ( \37181 , \30802 , \19045 );
nor \U$28404 ( \37182 , \37180 , \37181 );
xnor \U$28405 ( \37183 , \37182 , \19540 );
and \U$28406 ( \37184 , \19032 , \30823 );
and \U$28407 ( \37185 , \19558 , \30246 );
nor \U$28408 ( \37186 , \37184 , \37185 );
xnor \U$28409 ( \37187 , \37186 , \30813 );
xor \U$28410 ( \37188 , \37183 , \37187 );
and \U$28411 ( \37189 , \17627 , \32854 );
and \U$28412 ( \37190 , \18035 , \32067 );
nor \U$28413 ( \37191 , \37189 , \37190 );
xnor \U$28414 ( \37192 , \37191 , \32805 );
xor \U$28415 ( \37193 , \37188 , \37192 );
xor \U$28416 ( \37194 , \37179 , \37193 );
and \U$28417 ( \37195 , \25272 , \24138 );
and \U$28418 ( \37196 , \25815 , \23630 );
nor \U$28419 ( \37197 , \37195 , \37196 );
xnor \U$28420 ( \37198 , \37197 , \24144 );
and \U$28421 ( \37199 , \23617 , \25826 );
and \U$28422 ( \37200 , \24199 , \25264 );
nor \U$28423 ( \37201 , \37199 , \37200 );
xnor \U$28424 ( \37202 , \37201 , \25773 );
xor \U$28425 ( \37203 , \37198 , \37202 );
and \U$28426 ( \37204 , \16655 , \32802 );
xor \U$28427 ( \37205 , \37203 , \37204 );
xor \U$28428 ( \37206 , \37194 , \37205 );
xor \U$28429 ( \37207 , \37175 , \37206 );
xor \U$28430 ( \37208 , \37139 , \37207 );
and \U$28431 ( \37209 , \36954 , \36958 );
and \U$28432 ( \37210 , \36958 , \36973 );
and \U$28433 ( \37211 , \36954 , \36973 );
or \U$28434 ( \37212 , \37209 , \37210 , \37211 );
and \U$28435 ( \37213 , \36873 , \36903 );
and \U$28436 ( \37214 , \36903 , \36939 );
and \U$28437 ( \37215 , \36873 , \36939 );
or \U$28438 ( \37216 , \37213 , \37214 , \37215 );
xor \U$28439 ( \37217 , \37212 , \37216 );
and \U$28440 ( \37218 , \36963 , \36967 );
and \U$28441 ( \37219 , \36967 , \36972 );
and \U$28442 ( \37220 , \36963 , \36972 );
or \U$28443 ( \37221 , \37218 , \37219 , \37220 );
and \U$28444 ( \37222 , \36877 , \36887 );
and \U$28445 ( \37223 , \36887 , \36902 );
and \U$28446 ( \37224 , \36877 , \36902 );
or \U$28447 ( \37225 , \37222 , \37223 , \37224 );
xor \U$28448 ( \37226 , \37221 , \37225 );
and \U$28449 ( \37227 , \36880 , \36884 );
and \U$28450 ( \37228 , \36884 , \36886 );
and \U$28451 ( \37229 , \36880 , \36886 );
or \U$28452 ( \37230 , \37227 , \37228 , \37229 );
and \U$28453 ( \37231 , \36892 , \36896 );
and \U$28454 ( \37232 , \36896 , \36901 );
and \U$28455 ( \37233 , \36892 , \36901 );
or \U$28456 ( \37234 , \37231 , \37232 , \37233 );
xor \U$28457 ( \37235 , \37230 , \37234 );
buf \U$28458 ( \37236 , \36927 );
xor \U$28459 ( \37237 , \37235 , \37236 );
xor \U$28460 ( \37238 , \37226 , \37237 );
xor \U$28461 ( \37239 , \37217 , \37238 );
xor \U$28462 ( \37240 , \37208 , \37239 );
and \U$28463 ( \37241 , \36869 , \36940 );
and \U$28464 ( \37242 , \36940 , \36975 );
and \U$28465 ( \37243 , \36869 , \36975 );
or \U$28466 ( \37244 , \37241 , \37242 , \37243 );
xor \U$28467 ( \37245 , \37240 , \37244 );
and \U$28468 ( \37246 , \36976 , \36980 );
and \U$28469 ( \37247 , \36981 , \36984 );
or \U$28470 ( \37248 , \37246 , \37247 );
xor \U$28471 ( \37249 , \37245 , \37248 );
buf g9b8d ( \37250_nG9b8d , \37249 );
and \U$28472 ( \37251 , \10704 , \37250_nG9b8d );
or \U$28473 ( \37252 , \37135 , \37251 );
xor \U$28474 ( \37253 , \10703 , \37252 );
buf \U$28475 ( \37254 , \37253 );
buf \U$28477 ( \37255 , \37254 );
xor \U$28478 ( \37256 , \37134 , \37255 );
buf \U$28479 ( \37257 , \37256 );
and \U$28480 ( \37258 , \36857 , \36863 );
and \U$28481 ( \37259 , \36857 , \36991 );
and \U$28482 ( \37260 , \36863 , \36991 );
or \U$28483 ( \37261 , \37258 , \37259 , \37260 );
buf \U$28484 ( \37262 , \37261 );
xor \U$28485 ( \37263 , \37257 , \37262 );
and \U$28486 ( \37264 , \36792 , \36798 );
and \U$28487 ( \37265 , \36792 , \36805 );
and \U$28488 ( \37266 , \36798 , \36805 );
or \U$28489 ( \37267 , \37264 , \37265 , \37266 );
buf \U$28490 ( \37268 , \37267 );
and \U$28491 ( \37269 , \14631 , \34041_nG9ba8 );
and \U$28492 ( \37270 , \14628 , \34294_nG9ba5 );
or \U$28493 ( \37271 , \37269 , \37270 );
xor \U$28494 ( \37272 , \14627 , \37271 );
buf \U$28495 ( \37273 , \37272 );
buf \U$28497 ( \37274 , \37273 );
xor \U$28498 ( \37275 , \37268 , \37274 );
and \U$28499 ( \37276 , \12157 , \35570_nG9b9c );
and \U$28500 ( \37277 , \12154 , \35801_nG9b99 );
or \U$28501 ( \37278 , \37276 , \37277 );
xor \U$28502 ( \37279 , \12153 , \37278 );
buf \U$28503 ( \37280 , \37279 );
buf \U$28505 ( \37281 , \37280 );
xor \U$28506 ( \37282 , \37275 , \37281 );
buf \U$28507 ( \37283 , \37282 );
xor \U$28508 ( \37284 , \37263 , \37283 );
buf \U$28509 ( \37285 , \37284 );
and \U$28510 ( \37286 , \36998 , \37004 );
and \U$28511 ( \37287 , \36998 , \37011 );
and \U$28512 ( \37288 , \37004 , \37011 );
or \U$28513 ( \37289 , \37286 , \37287 , \37288 );
buf \U$28514 ( \37290 , \37289 );
and \U$28515 ( \37291 , \36831 , \36833 );
and \U$28516 ( \37292 , \36831 , \36840 );
and \U$28517 ( \37293 , \36833 , \36840 );
or \U$28518 ( \37294 , \37291 , \37292 , \37293 );
buf \U$28519 ( \37295 , \37294 );
and \U$28521 ( \37296 , \32916 , \16680_nG9bed );
or \U$28522 ( \37297 , 1'b0 , \37296 );
xor \U$28523 ( \37298 , 1'b0 , \37297 );
buf \U$28524 ( \37299 , \37298 );
buf \U$28526 ( \37300 , \37299 );
and \U$28527 ( \37301 , \31636 , \17665_nG9bea );
and \U$28528 ( \37302 , \31633 , \18107_nG9be7 );
or \U$28529 ( \37303 , \37301 , \37302 );
xor \U$28530 ( \37304 , \31632 , \37303 );
buf \U$28531 ( \37305 , \37304 );
buf \U$28533 ( \37306 , \37305 );
xor \U$28534 ( \37307 , \37300 , \37306 );
buf \U$28535 ( \37308 , \37307 );
xor \U$28536 ( \37309 , \37295 , \37308 );
and \U$28537 ( \37310 , \26431 , \22129_nG9bd8 );
and \U$28538 ( \37311 , \26428 , \22629_nG9bd5 );
or \U$28539 ( \37312 , \37310 , \37311 );
xor \U$28540 ( \37313 , \26427 , \37312 );
buf \U$28541 ( \37314 , \37313 );
buf \U$28543 ( \37315 , \37314 );
xor \U$28544 ( \37316 , \37309 , \37315 );
buf \U$28545 ( \37317 , \37316 );
and \U$28546 ( \37318 , \17297 , \32179_nG9bb4 );
and \U$28547 ( \37319 , \17294 , \32888_nG9bb1 );
or \U$28548 ( \37320 , \37318 , \37319 );
xor \U$28549 ( \37321 , \17293 , \37320 );
buf \U$28550 ( \37322 , \37321 );
buf \U$28552 ( \37323 , \37322 );
xor \U$28553 ( \37324 , \37317 , \37323 );
and \U$28554 ( \37325 , \13370 , \34643_nG9ba2 );
and \U$28555 ( \37326 , \13367 , \35094_nG9b9f );
or \U$28556 ( \37327 , \37325 , \37326 );
xor \U$28557 ( \37328 , \13366 , \37327 );
buf \U$28558 ( \37329 , \37328 );
buf \U$28560 ( \37330 , \37329 );
xor \U$28561 ( \37331 , \37324 , \37330 );
buf \U$28562 ( \37332 , \37331 );
xor \U$28563 ( \37333 , \37290 , \37332 );
and \U$28564 ( \37334 , \36842 , \36848 );
and \U$28565 ( \37335 , \36842 , \36855 );
and \U$28566 ( \37336 , \36848 , \36855 );
or \U$28567 ( \37337 , \37334 , \37335 , \37336 );
buf \U$28568 ( \37338 , \37337 );
and \U$28569 ( \37339 , \20155 , \28602_nG9bc0 );
and \U$28570 ( \37340 , \20152 , \29179_nG9bbd );
or \U$28571 ( \37341 , \37339 , \37340 );
xor \U$28572 ( \37342 , \20151 , \37341 );
buf \U$28573 ( \37343 , \37342 );
buf \U$28575 ( \37344 , \37343 );
xor \U$28576 ( \37345 , \37338 , \37344 );
and \U$28577 ( \37346 , \15940 , \33181_nG9bae );
and \U$28578 ( \37347 , \15937 , \33613_nG9bab );
or \U$28579 ( \37348 , \37346 , \37347 );
xor \U$28580 ( \37349 , \15936 , \37348 );
buf \U$28581 ( \37350 , \37349 );
buf \U$28583 ( \37351 , \37350 );
xor \U$28584 ( \37352 , \37345 , \37351 );
buf \U$28585 ( \37353 , \37352 );
xor \U$28586 ( \37354 , \37333 , \37353 );
buf \U$28587 ( \37355 , \37354 );
xor \U$28588 ( \37356 , \37285 , \37355 );
and \U$28589 ( \37357 , \36993 , \37013 );
and \U$28590 ( \37358 , \36993 , \37019 );
and \U$28591 ( \37359 , \37013 , \37019 );
or \U$28592 ( \37360 , \37357 , \37358 , \37359 );
buf \U$28593 ( \37361 , \37360 );
xor \U$28594 ( \37362 , \37356 , \37361 );
buf \U$28595 ( \37363 , \37362 );
xor \U$28596 ( \37364 , \37122 , \37363 );
buf \U$28597 ( \37365 , \37364 );
xor \U$28598 ( \37366 , \37043 , \37365 );
and \U$28599 ( \37367 , \36694 , \36699 );
and \U$28600 ( \37368 , \36694 , \36763 );
and \U$28601 ( \37369 , \36699 , \36763 );
or \U$28602 ( \37370 , \37367 , \37368 , \37369 );
buf \U$28603 ( \37371 , \37370 );
xor \U$28604 ( \37372 , \37366 , \37371 );
and \U$28605 ( \37373 , \37038 , \37372 );
and \U$28607 ( \37374 , \37032 , \37037 );
or \U$28609 ( \37375 , 1'b0 , \37374 , 1'b0 );
xor \U$28610 ( \37376 , \37373 , \37375 );
and \U$28612 ( \37377 , \37025 , \37031 );
and \U$28613 ( \37378 , \37027 , \37031 );
or \U$28614 ( \37379 , 1'b0 , \37377 , \37378 );
xor \U$28615 ( \37380 , \37376 , \37379 );
xor \U$28622 ( \37381 , \37380 , 1'b0 );
and \U$28623 ( \37382 , \37043 , \37365 );
and \U$28624 ( \37383 , \37043 , \37371 );
and \U$28625 ( \37384 , \37365 , \37371 );
or \U$28626 ( \37385 , \37382 , \37383 , \37384 );
xor \U$28627 ( \37386 , \37381 , \37385 );
and \U$28628 ( \37387 , \37285 , \37355 );
and \U$28629 ( \37388 , \37285 , \37361 );
and \U$28630 ( \37389 , \37355 , \37361 );
or \U$28631 ( \37390 , \37387 , \37388 , \37389 );
buf \U$28632 ( \37391 , \37390 );
and \U$28633 ( \37392 , \37290 , \37332 );
and \U$28634 ( \37393 , \37290 , \37353 );
and \U$28635 ( \37394 , \37332 , \37353 );
or \U$28636 ( \37395 , \37392 , \37393 , \37394 );
buf \U$28637 ( \37396 , \37395 );
and \U$28638 ( \37397 , \37338 , \37344 );
and \U$28639 ( \37398 , \37338 , \37351 );
and \U$28640 ( \37399 , \37344 , \37351 );
or \U$28641 ( \37400 , \37397 , \37398 , \37399 );
buf \U$28642 ( \37401 , \37400 );
and \U$28643 ( \37402 , \37300 , \37306 );
buf \U$28644 ( \37403 , \37402 );
and \U$28645 ( \37404 , \29853 , \19586_nG9be1 );
and \U$28646 ( \37405 , \29850 , \20608_nG9bde );
or \U$28647 ( \37406 , \37404 , \37405 );
xor \U$28648 ( \37407 , \29849 , \37406 );
buf \U$28649 ( \37408 , \37407 );
buf \U$28651 ( \37409 , \37408 );
xor \U$28652 ( \37410 , \37403 , \37409 );
and \U$28653 ( \37411 , \28118 , \21086_nG9bdb );
and \U$28654 ( \37412 , \28115 , \22129_nG9bd8 );
or \U$28655 ( \37413 , \37411 , \37412 );
xor \U$28656 ( \37414 , \28114 , \37413 );
buf \U$28657 ( \37415 , \37414 );
buf \U$28659 ( \37416 , \37415 );
xor \U$28660 ( \37417 , \37410 , \37416 );
buf \U$28661 ( \37418 , \37417 );
and \U$28662 ( \37419 , \20155 , \29179_nG9bbd );
and \U$28663 ( \37420 , \20152 , \30366_nG9bba );
or \U$28664 ( \37421 , \37419 , \37420 );
xor \U$28665 ( \37422 , \20151 , \37421 );
buf \U$28666 ( \37423 , \37422 );
buf \U$28668 ( \37424 , \37423 );
xor \U$28669 ( \37425 , \37418 , \37424 );
and \U$28670 ( \37426 , \18702 , \30940_nG9bb7 );
and \U$28671 ( \37427 , \18699 , \32179_nG9bb4 );
or \U$28672 ( \37428 , \37426 , \37427 );
xor \U$28673 ( \37429 , \18698 , \37428 );
buf \U$28674 ( \37430 , \37429 );
buf \U$28676 ( \37431 , \37430 );
xor \U$28677 ( \37432 , \37425 , \37431 );
buf \U$28678 ( \37433 , \37432 );
xor \U$28679 ( \37434 , \37401 , \37433 );
and \U$28680 ( \37435 , \37317 , \37323 );
and \U$28681 ( \37436 , \37317 , \37330 );
and \U$28682 ( \37437 , \37323 , \37330 );
or \U$28683 ( \37438 , \37435 , \37436 , \37437 );
buf \U$28684 ( \37439 , \37438 );
xor \U$28685 ( \37440 , \37434 , \37439 );
buf \U$28686 ( \37441 , \37440 );
xor \U$28687 ( \37442 , \37396 , \37441 );
and \U$28688 ( \37443 , \37079 , \37100 );
and \U$28689 ( \37444 , \37079 , \37106 );
and \U$28690 ( \37445 , \37100 , \37106 );
or \U$28691 ( \37446 , \37443 , \37444 , \37445 );
buf \U$28692 ( \37447 , \37446 );
xor \U$28693 ( \37448 , \37442 , \37447 );
buf \U$28694 ( \37449 , \37448 );
xor \U$28695 ( \37450 , \37391 , \37449 );
and \U$28696 ( \37451 , \37048 , \37108 );
and \U$28697 ( \37452 , \37048 , \37114 );
and \U$28698 ( \37453 , \37108 , \37114 );
or \U$28699 ( \37454 , \37451 , \37452 , \37453 );
buf \U$28700 ( \37455 , \37454 );
xor \U$28701 ( \37456 , \37450 , \37455 );
buf \U$28702 ( \37457 , \37456 );
and \U$28703 ( \37458 , \37257 , \37262 );
and \U$28704 ( \37459 , \37257 , \37283 );
and \U$28705 ( \37460 , \37262 , \37283 );
or \U$28706 ( \37461 , \37458 , \37459 , \37460 );
buf \U$28707 ( \37462 , \37461 );
and \U$28708 ( \37463 , \37127 , \37133 );
and \U$28709 ( \37464 , \37127 , \37255 );
and \U$28710 ( \37465 , \37133 , \37255 );
or \U$28711 ( \37466 , \37463 , \37464 , \37465 );
buf \U$28712 ( \37467 , \37466 );
and \U$28713 ( \37468 , \24792 , \24226_nG9bcf );
and \U$28714 ( \37469 , \24789 , \25298_nG9bcc );
or \U$28715 ( \37470 , \37468 , \37469 );
xor \U$28716 ( \37471 , \24788 , \37470 );
buf \U$28717 ( \37472 , \37471 );
buf \U$28719 ( \37473 , \37472 );
and \U$28720 ( \37474 , \23201 , \25860_nG9bc9 );
and \U$28721 ( \37475 , \23198 , \26887_nG9bc6 );
or \U$28722 ( \37476 , \37474 , \37475 );
xor \U$28723 ( \37477 , \23197 , \37476 );
buf \U$28724 ( \37478 , \37477 );
buf \U$28726 ( \37479 , \37478 );
xor \U$28727 ( \37480 , \37473 , \37479 );
and \U$28728 ( \37481 , \21658 , \27416_nG9bc3 );
and \U$28729 ( \37482 , \21655 , \28602_nG9bc0 );
or \U$28730 ( \37483 , \37481 , \37482 );
xor \U$28731 ( \37484 , \21654 , \37483 );
buf \U$28732 ( \37485 , \37484 );
buf \U$28734 ( \37486 , \37485 );
xor \U$28735 ( \37487 , \37480 , \37486 );
buf \U$28736 ( \37488 , \37487 );
and \U$28737 ( \37489 , \10421 , \36589_nG9b93 );
and \U$28738 ( \37490 , \10418 , \36986_nG9b90 );
or \U$28739 ( \37491 , \37489 , \37490 );
xor \U$28740 ( \37492 , \10417 , \37491 );
buf \U$28741 ( \37493 , \37492 );
buf \U$28743 ( \37494 , \37493 );
xor \U$28744 ( \37495 , \37488 , \37494 );
and \U$28745 ( \37496 , \10707 , \37250_nG9b8d );
and \U$28746 ( \37497 , \37212 , \37216 );
and \U$28747 ( \37498 , \37216 , \37238 );
and \U$28748 ( \37499 , \37212 , \37238 );
or \U$28749 ( \37500 , \37497 , \37498 , \37499 );
and \U$28750 ( \37501 , \37147 , \37158 );
and \U$28751 ( \37502 , \37158 , \37173 );
and \U$28752 ( \37503 , \37147 , \37173 );
or \U$28753 ( \37504 , \37501 , \37502 , \37503 );
and \U$28754 ( \37505 , \37179 , \37193 );
and \U$28755 ( \37506 , \37193 , \37205 );
and \U$28756 ( \37507 , \37179 , \37205 );
or \U$28757 ( \37508 , \37505 , \37506 , \37507 );
xor \U$28758 ( \37509 , \37504 , \37508 );
and \U$28759 ( \37510 , \27313 , \22542 );
and \U$28760 ( \37511 , \28534 , \22103 );
nor \U$28761 ( \37512 , \37510 , \37511 );
xnor \U$28762 ( \37513 , \37512 , \22548 );
and \U$28763 ( \37514 , \21033 , \29070 );
and \U$28764 ( \37515 , \22090 , \28526 );
nor \U$28765 ( \37516 , \37514 , \37515 );
xnor \U$28766 ( \37517 , \37516 , \29076 );
xor \U$28767 ( \37518 , \37513 , \37517 );
and \U$28768 ( \37519 , \19558 , \30823 );
and \U$28769 ( \37520 , \20544 , \30246 );
nor \U$28770 ( \37521 , \37519 , \37520 );
xnor \U$28771 ( \37522 , \37521 , \30813 );
xor \U$28772 ( \37523 , \37518 , \37522 );
and \U$28773 ( \37524 , \25815 , \24138 );
and \U$28774 ( \37525 , \26829 , \23630 );
nor \U$28775 ( \37526 , \37524 , \37525 );
xnor \U$28776 ( \37527 , \37526 , \24144 );
and \U$28777 ( \37528 , \18035 , \32854 );
and \U$28778 ( \37529 , \19032 , \32067 );
nor \U$28779 ( \37530 , \37528 , \37529 );
xnor \U$28780 ( \37531 , \37530 , \32805 );
xor \U$28781 ( \37532 , \37527 , \37531 );
and \U$28782 ( \37533 , \17627 , \32802 );
xor \U$28783 ( \37534 , \37532 , \37533 );
xor \U$28784 ( \37535 , \37523 , \37534 );
and \U$28785 ( \37536 , \32794 , \18090 );
not \U$28786 ( \37537 , \37536 );
xnor \U$28787 ( \37538 , \37537 , \18046 );
and \U$28788 ( \37539 , \29084 , \21005 );
and \U$28789 ( \37540 , \30268 , \20557 );
nor \U$28790 ( \37541 , \37539 , \37540 );
xnor \U$28791 ( \37542 , \37541 , \21011 );
xor \U$28792 ( \37543 , \37538 , \37542 );
and \U$28793 ( \37544 , \24199 , \25826 );
and \U$28794 ( \37545 , \25272 , \25264 );
nor \U$28795 ( \37546 , \37544 , \37545 );
xnor \U$28796 ( \37547 , \37546 , \25773 );
xor \U$28797 ( \37548 , \37543 , \37547 );
xor \U$28798 ( \37549 , \37535 , \37548 );
xor \U$28799 ( \37550 , \37509 , \37549 );
xor \U$28800 ( \37551 , \37500 , \37550 );
and \U$28801 ( \37552 , \37221 , \37225 );
and \U$28802 ( \37553 , \37225 , \37237 );
and \U$28803 ( \37554 , \37221 , \37237 );
or \U$28804 ( \37555 , \37552 , \37553 , \37554 );
and \U$28805 ( \37556 , \37143 , \37174 );
and \U$28806 ( \37557 , \37174 , \37206 );
and \U$28807 ( \37558 , \37143 , \37206 );
or \U$28808 ( \37559 , \37556 , \37557 , \37558 );
xor \U$28809 ( \37560 , \37555 , \37559 );
and \U$28810 ( \37561 , \37230 , \37234 );
and \U$28811 ( \37562 , \37234 , \37236 );
and \U$28812 ( \37563 , \37230 , \37236 );
or \U$28813 ( \37564 , \37561 , \37562 , \37563 );
and \U$28814 ( \37565 , \37198 , \37202 );
and \U$28815 ( \37566 , \37202 , \37204 );
and \U$28816 ( \37567 , \37198 , \37204 );
or \U$28817 ( \37568 , \37565 , \37566 , \37567 );
and \U$28818 ( \37569 , \37148 , \37152 );
and \U$28819 ( \37570 , \37152 , \37157 );
and \U$28820 ( \37571 , \37148 , \37157 );
or \U$28821 ( \37572 , \37569 , \37570 , \37571 );
xor \U$28822 ( \37573 , \37568 , \37572 );
and \U$28823 ( \37574 , \37163 , \37167 );
and \U$28824 ( \37575 , \37167 , \37172 );
and \U$28825 ( \37576 , \37163 , \37172 );
or \U$28826 ( \37577 , \37574 , \37575 , \37576 );
xor \U$28827 ( \37578 , \37573 , \37577 );
xor \U$28828 ( \37579 , \37564 , \37578 );
and \U$28829 ( \37580 , \37183 , \37187 );
and \U$28830 ( \37581 , \37187 , \37192 );
and \U$28831 ( \37582 , \37183 , \37192 );
or \U$28832 ( \37583 , \37580 , \37581 , \37582 );
and \U$28833 ( \37584 , \30802 , \19534 );
and \U$28834 ( \37585 , \32054 , \19045 );
nor \U$28835 ( \37586 , \37584 , \37585 );
xnor \U$28836 ( \37587 , \37586 , \19540 );
not \U$28837 ( \37588 , \37587 );
xor \U$28838 ( \37589 , \37583 , \37588 );
and \U$28839 ( \37590 , \22556 , \27397 );
and \U$28840 ( \37591 , \23617 , \26807 );
nor \U$28841 ( \37592 , \37590 , \37591 );
xnor \U$28842 ( \37593 , \37592 , \27295 );
xor \U$28843 ( \37594 , \37589 , \37593 );
xor \U$28844 ( \37595 , \37579 , \37594 );
xor \U$28845 ( \37596 , \37560 , \37595 );
xor \U$28846 ( \37597 , \37551 , \37596 );
and \U$28847 ( \37598 , \37139 , \37207 );
and \U$28848 ( \37599 , \37207 , \37239 );
and \U$28849 ( \37600 , \37139 , \37239 );
or \U$28850 ( \37601 , \37598 , \37599 , \37600 );
xor \U$28851 ( \37602 , \37597 , \37601 );
and \U$28852 ( \37603 , \37240 , \37244 );
and \U$28853 ( \37604 , \37245 , \37248 );
or \U$28854 ( \37605 , \37603 , \37604 );
xor \U$28855 ( \37606 , \37602 , \37605 );
buf g9b8a ( \37607_nG9b8a , \37606 );
and \U$28856 ( \37608 , \10704 , \37607_nG9b8a );
or \U$28857 ( \37609 , \37496 , \37608 );
xor \U$28858 ( \37610 , \10703 , \37609 );
buf \U$28859 ( \37611 , \37610 );
buf \U$28861 ( \37612 , \37611 );
xor \U$28862 ( \37613 , \37495 , \37612 );
buf \U$28863 ( \37614 , \37613 );
xor \U$28864 ( \37615 , \37467 , \37614 );
and \U$28865 ( \37616 , \37053 , \37070 );
and \U$28866 ( \37617 , \37053 , \37077 );
and \U$28867 ( \37618 , \37070 , \37077 );
or \U$28868 ( \37619 , \37616 , \37617 , \37618 );
buf \U$28869 ( \37620 , \37619 );
and \U$28870 ( \37621 , \37085 , \37091 );
and \U$28871 ( \37622 , \37085 , \37098 );
and \U$28872 ( \37623 , \37091 , \37098 );
or \U$28873 ( \37624 , \37621 , \37622 , \37623 );
buf \U$28874 ( \37625 , \37624 );
xor \U$28875 ( \37626 , \37620 , \37625 );
and \U$28876 ( \37627 , \12157 , \35801_nG9b99 );
and \U$28877 ( \37628 , \12154 , \36172_nG9b96 );
or \U$28878 ( \37629 , \37627 , \37628 );
xor \U$28879 ( \37630 , \12153 , \37629 );
buf \U$28880 ( \37631 , \37630 );
buf \U$28882 ( \37632 , \37631 );
xor \U$28883 ( \37633 , \37626 , \37632 );
buf \U$28884 ( \37634 , \37633 );
xor \U$28885 ( \37635 , \37615 , \37634 );
buf \U$28886 ( \37636 , \37635 );
xor \U$28887 ( \37637 , \37462 , \37636 );
and \U$28888 ( \37638 , \37268 , \37274 );
and \U$28889 ( \37639 , \37268 , \37281 );
and \U$28890 ( \37640 , \37274 , \37281 );
or \U$28891 ( \37641 , \37638 , \37639 , \37640 );
buf \U$28892 ( \37642 , \37641 );
and \U$28893 ( \37643 , \37295 , \37308 );
and \U$28894 ( \37644 , \37295 , \37315 );
and \U$28895 ( \37645 , \37308 , \37315 );
or \U$28896 ( \37646 , \37643 , \37644 , \37645 );
buf \U$28897 ( \37647 , \37646 );
and \U$28898 ( \37648 , \17297 , \32888_nG9bb1 );
and \U$28899 ( \37649 , \17294 , \33181_nG9bae );
or \U$28900 ( \37650 , \37648 , \37649 );
xor \U$28901 ( \37651 , \17293 , \37650 );
buf \U$28902 ( \37652 , \37651 );
buf \U$28904 ( \37653 , \37652 );
xor \U$28905 ( \37654 , \37647 , \37653 );
and \U$28906 ( \37655 , \15940 , \33613_nG9bab );
and \U$28907 ( \37656 , \15937 , \34041_nG9ba8 );
or \U$28908 ( \37657 , \37655 , \37656 );
xor \U$28909 ( \37658 , \15936 , \37657 );
buf \U$28910 ( \37659 , \37658 );
buf \U$28912 ( \37660 , \37659 );
xor \U$28913 ( \37661 , \37654 , \37660 );
buf \U$28914 ( \37662 , \37661 );
xor \U$28915 ( \37663 , \37642 , \37662 );
and \U$28916 ( \37664 , \37055 , \37061 );
and \U$28917 ( \37665 , \37055 , \37068 );
and \U$28918 ( \37666 , \37061 , \37068 );
or \U$28919 ( \37667 , \37664 , \37665 , \37666 );
buf \U$28920 ( \37668 , \37667 );
and \U$28922 ( \37669 , \32916 , \17665_nG9bea );
or \U$28923 ( \37670 , 1'b0 , \37669 );
xor \U$28924 ( \37671 , 1'b0 , \37670 );
buf \U$28925 ( \37672 , \37671 );
buf \U$28927 ( \37673 , \37672 );
and \U$28928 ( \37674 , \31636 , \18107_nG9be7 );
and \U$28929 ( \37675 , \31633 , \19091_nG9be4 );
or \U$28930 ( \37676 , \37674 , \37675 );
xor \U$28931 ( \37677 , \31632 , \37676 );
buf \U$28932 ( \37678 , \37677 );
buf \U$28934 ( \37679 , \37678 );
xor \U$28935 ( \37680 , \37673 , \37679 );
buf \U$28936 ( \37681 , \37680 );
xor \U$28937 ( \37682 , \37668 , \37681 );
and \U$28938 ( \37683 , \26431 , \22629_nG9bd5 );
and \U$28939 ( \37684 , \26428 , \23696_nG9bd2 );
or \U$28940 ( \37685 , \37683 , \37684 );
xor \U$28941 ( \37686 , \26427 , \37685 );
buf \U$28942 ( \37687 , \37686 );
buf \U$28944 ( \37688 , \37687 );
xor \U$28945 ( \37689 , \37682 , \37688 );
buf \U$28946 ( \37690 , \37689 );
and \U$28947 ( \37691 , \14631 , \34294_nG9ba5 );
and \U$28948 ( \37692 , \14628 , \34643_nG9ba2 );
or \U$28949 ( \37693 , \37691 , \37692 );
xor \U$28950 ( \37694 , \14627 , \37693 );
buf \U$28951 ( \37695 , \37694 );
buf \U$28953 ( \37696 , \37695 );
xor \U$28954 ( \37697 , \37690 , \37696 );
and \U$28955 ( \37698 , \13370 , \35094_nG9b9f );
and \U$28956 ( \37699 , \13367 , \35570_nG9b9c );
or \U$28957 ( \37700 , \37698 , \37699 );
xor \U$28958 ( \37701 , \13366 , \37700 );
buf \U$28959 ( \37702 , \37701 );
buf \U$28961 ( \37703 , \37702 );
xor \U$28962 ( \37704 , \37697 , \37703 );
buf \U$28963 ( \37705 , \37704 );
xor \U$28964 ( \37706 , \37663 , \37705 );
buf \U$28965 ( \37707 , \37706 );
xor \U$28966 ( \37708 , \37637 , \37707 );
buf \U$28967 ( \37709 , \37708 );
xor \U$28968 ( \37710 , \37457 , \37709 );
and \U$28969 ( \37711 , \37116 , \37121 );
and \U$28970 ( \37712 , \37116 , \37363 );
and \U$28971 ( \37713 , \37121 , \37363 );
or \U$28972 ( \37714 , \37711 , \37712 , \37713 );
buf \U$28973 ( \37715 , \37714 );
xor \U$28974 ( \37716 , \37710 , \37715 );
and \U$28975 ( \37717 , \37386 , \37716 );
and \U$28977 ( \37718 , \37380 , \37385 );
or \U$28979 ( \37719 , 1'b0 , \37718 , 1'b0 );
xor \U$28980 ( \37720 , \37717 , \37719 );
and \U$28982 ( \37721 , \37373 , \37379 );
and \U$28983 ( \37722 , \37375 , \37379 );
or \U$28984 ( \37723 , 1'b0 , \37721 , \37722 );
xor \U$28985 ( \37724 , \37720 , \37723 );
xor \U$28992 ( \37725 , \37724 , 1'b0 );
and \U$28993 ( \37726 , \37457 , \37709 );
and \U$28994 ( \37727 , \37457 , \37715 );
and \U$28995 ( \37728 , \37709 , \37715 );
or \U$28996 ( \37729 , \37726 , \37727 , \37728 );
xor \U$28997 ( \37730 , \37725 , \37729 );
and \U$28998 ( \37731 , \37391 , \37449 );
and \U$28999 ( \37732 , \37391 , \37455 );
and \U$29000 ( \37733 , \37449 , \37455 );
or \U$29001 ( \37734 , \37731 , \37732 , \37733 );
buf \U$29002 ( \37735 , \37734 );
and \U$29003 ( \37736 , \37396 , \37441 );
and \U$29004 ( \37737 , \37396 , \37447 );
and \U$29005 ( \37738 , \37441 , \37447 );
or \U$29006 ( \37739 , \37736 , \37737 , \37738 );
buf \U$29007 ( \37740 , \37739 );
and \U$29008 ( \37741 , \37462 , \37636 );
and \U$29009 ( \37742 , \37462 , \37707 );
and \U$29010 ( \37743 , \37636 , \37707 );
or \U$29011 ( \37744 , \37741 , \37742 , \37743 );
buf \U$29012 ( \37745 , \37744 );
xor \U$29013 ( \37746 , \37740 , \37745 );
and \U$29014 ( \37747 , \37401 , \37433 );
and \U$29015 ( \37748 , \37401 , \37439 );
and \U$29016 ( \37749 , \37433 , \37439 );
or \U$29017 ( \37750 , \37747 , \37748 , \37749 );
buf \U$29018 ( \37751 , \37750 );
and \U$29019 ( \37752 , \37642 , \37662 );
and \U$29020 ( \37753 , \37642 , \37705 );
and \U$29021 ( \37754 , \37662 , \37705 );
or \U$29022 ( \37755 , \37752 , \37753 , \37754 );
buf \U$29023 ( \37756 , \37755 );
xor \U$29024 ( \37757 , \37751 , \37756 );
and \U$29026 ( \37758 , \32916 , \18107_nG9be7 );
or \U$29027 ( \37759 , 1'b0 , \37758 );
xor \U$29028 ( \37760 , 1'b0 , \37759 );
buf \U$29029 ( \37761 , \37760 );
buf \U$29031 ( \37762 , \37761 );
and \U$29032 ( \37763 , \29853 , \20608_nG9bde );
and \U$29033 ( \37764 , \29850 , \21086_nG9bdb );
or \U$29034 ( \37765 , \37763 , \37764 );
xor \U$29035 ( \37766 , \29849 , \37765 );
buf \U$29036 ( \37767 , \37766 );
buf \U$29038 ( \37768 , \37767 );
xor \U$29039 ( \37769 , \37762 , \37768 );
buf \U$29040 ( \37770 , \37769 );
and \U$29041 ( \37771 , \37673 , \37679 );
buf \U$29042 ( \37772 , \37771 );
xor \U$29043 ( \37773 , \37770 , \37772 );
and \U$29044 ( \37774 , \31636 , \19091_nG9be4 );
and \U$29045 ( \37775 , \31633 , \19586_nG9be1 );
or \U$29046 ( \37776 , \37774 , \37775 );
xor \U$29047 ( \37777 , \31632 , \37776 );
buf \U$29048 ( \37778 , \37777 );
buf \U$29050 ( \37779 , \37778 );
xor \U$29051 ( \37780 , \37773 , \37779 );
buf \U$29052 ( \37781 , \37780 );
and \U$29053 ( \37782 , \21658 , \28602_nG9bc0 );
and \U$29054 ( \37783 , \21655 , \29179_nG9bbd );
or \U$29055 ( \37784 , \37782 , \37783 );
xor \U$29056 ( \37785 , \21654 , \37784 );
buf \U$29057 ( \37786 , \37785 );
buf \U$29059 ( \37787 , \37786 );
xor \U$29060 ( \37788 , \37781 , \37787 );
and \U$29061 ( \37789 , \18702 , \32179_nG9bb4 );
and \U$29062 ( \37790 , \18699 , \32888_nG9bb1 );
or \U$29063 ( \37791 , \37789 , \37790 );
xor \U$29064 ( \37792 , \18698 , \37791 );
buf \U$29065 ( \37793 , \37792 );
buf \U$29067 ( \37794 , \37793 );
xor \U$29068 ( \37795 , \37788 , \37794 );
buf \U$29069 ( \37796 , \37795 );
and \U$29070 ( \37797 , \37690 , \37696 );
and \U$29071 ( \37798 , \37690 , \37703 );
and \U$29072 ( \37799 , \37696 , \37703 );
or \U$29073 ( \37800 , \37797 , \37798 , \37799 );
buf \U$29074 ( \37801 , \37800 );
xor \U$29075 ( \37802 , \37796 , \37801 );
and \U$29076 ( \37803 , \37647 , \37653 );
and \U$29077 ( \37804 , \37647 , \37660 );
and \U$29078 ( \37805 , \37653 , \37660 );
or \U$29079 ( \37806 , \37803 , \37804 , \37805 );
buf \U$29080 ( \37807 , \37806 );
xor \U$29081 ( \37808 , \37802 , \37807 );
buf \U$29082 ( \37809 , \37808 );
xor \U$29083 ( \37810 , \37757 , \37809 );
buf \U$29084 ( \37811 , \37810 );
xor \U$29085 ( \37812 , \37746 , \37811 );
buf \U$29086 ( \37813 , \37812 );
xor \U$29087 ( \37814 , \37735 , \37813 );
and \U$29088 ( \37815 , \37418 , \37424 );
and \U$29089 ( \37816 , \37418 , \37431 );
and \U$29090 ( \37817 , \37424 , \37431 );
or \U$29091 ( \37818 , \37815 , \37816 , \37817 );
buf \U$29092 ( \37819 , \37818 );
and \U$29093 ( \37820 , \24792 , \25298_nG9bcc );
and \U$29094 ( \37821 , \24789 , \25860_nG9bc9 );
or \U$29095 ( \37822 , \37820 , \37821 );
xor \U$29096 ( \37823 , \24788 , \37822 );
buf \U$29097 ( \37824 , \37823 );
buf \U$29099 ( \37825 , \37824 );
and \U$29100 ( \37826 , \23201 , \26887_nG9bc6 );
and \U$29101 ( \37827 , \23198 , \27416_nG9bc3 );
or \U$29102 ( \37828 , \37826 , \37827 );
xor \U$29103 ( \37829 , \23197 , \37828 );
buf \U$29104 ( \37830 , \37829 );
buf \U$29106 ( \37831 , \37830 );
xor \U$29107 ( \37832 , \37825 , \37831 );
and \U$29108 ( \37833 , \20155 , \30366_nG9bba );
and \U$29109 ( \37834 , \20152 , \30940_nG9bb7 );
or \U$29110 ( \37835 , \37833 , \37834 );
xor \U$29111 ( \37836 , \20151 , \37835 );
buf \U$29112 ( \37837 , \37836 );
buf \U$29114 ( \37838 , \37837 );
xor \U$29115 ( \37839 , \37832 , \37838 );
buf \U$29116 ( \37840 , \37839 );
xor \U$29117 ( \37841 , \37819 , \37840 );
and \U$29118 ( \37842 , \12157 , \36172_nG9b96 );
and \U$29119 ( \37843 , \12154 , \36589_nG9b93 );
or \U$29120 ( \37844 , \37842 , \37843 );
xor \U$29121 ( \37845 , \12153 , \37844 );
buf \U$29122 ( \37846 , \37845 );
buf \U$29124 ( \37847 , \37846 );
xor \U$29125 ( \37848 , \37841 , \37847 );
buf \U$29126 ( \37849 , \37848 );
and \U$29127 ( \37850 , \37488 , \37494 );
and \U$29128 ( \37851 , \37488 , \37612 );
and \U$29129 ( \37852 , \37494 , \37612 );
or \U$29130 ( \37853 , \37850 , \37851 , \37852 );
buf \U$29131 ( \37854 , \37853 );
xor \U$29132 ( \37855 , \37849 , \37854 );
and \U$29133 ( \37856 , \15940 , \34041_nG9ba8 );
and \U$29134 ( \37857 , \15937 , \34294_nG9ba5 );
or \U$29135 ( \37858 , \37856 , \37857 );
xor \U$29136 ( \37859 , \15936 , \37858 );
buf \U$29137 ( \37860 , \37859 );
buf \U$29139 ( \37861 , \37860 );
and \U$29140 ( \37862 , \10421 , \36986_nG9b90 );
and \U$29141 ( \37863 , \10418 , \37250_nG9b8d );
or \U$29142 ( \37864 , \37862 , \37863 );
xor \U$29143 ( \37865 , \10417 , \37864 );
buf \U$29144 ( \37866 , \37865 );
buf \U$29146 ( \37867 , \37866 );
xor \U$29147 ( \37868 , \37861 , \37867 );
and \U$29148 ( \37869 , \10707 , \37607_nG9b8a );
and \U$29149 ( \37870 , \37504 , \37508 );
and \U$29150 ( \37871 , \37508 , \37549 );
and \U$29151 ( \37872 , \37504 , \37549 );
or \U$29152 ( \37873 , \37870 , \37871 , \37872 );
and \U$29153 ( \37874 , \37555 , \37559 );
and \U$29154 ( \37875 , \37559 , \37595 );
and \U$29155 ( \37876 , \37555 , \37595 );
or \U$29156 ( \37877 , \37874 , \37875 , \37876 );
xor \U$29157 ( \37878 , \37873 , \37877 );
and \U$29158 ( \37879 , \37564 , \37578 );
and \U$29159 ( \37880 , \37578 , \37594 );
and \U$29160 ( \37881 , \37564 , \37594 );
or \U$29161 ( \37882 , \37879 , \37880 , \37881 );
and \U$29162 ( \37883 , \37568 , \37572 );
and \U$29163 ( \37884 , \37572 , \37577 );
and \U$29164 ( \37885 , \37568 , \37577 );
or \U$29165 ( \37886 , \37883 , \37884 , \37885 );
and \U$29166 ( \37887 , \37583 , \37588 );
and \U$29167 ( \37888 , \37588 , \37593 );
and \U$29168 ( \37889 , \37583 , \37593 );
or \U$29169 ( \37890 , \37887 , \37888 , \37889 );
xor \U$29170 ( \37891 , \37886 , \37890 );
buf \U$29171 ( \37892 , \37587 );
and \U$29172 ( \37893 , \25272 , \25826 );
and \U$29173 ( \37894 , \25815 , \25264 );
nor \U$29174 ( \37895 , \37893 , \37894 );
xnor \U$29175 ( \37896 , \37895 , \25773 );
xor \U$29176 ( \37897 , \37892 , \37896 );
and \U$29177 ( \37898 , \23617 , \27397 );
and \U$29178 ( \37899 , \24199 , \26807 );
nor \U$29179 ( \37900 , \37898 , \37899 );
xnor \U$29180 ( \37901 , \37900 , \27295 );
xor \U$29181 ( \37902 , \37897 , \37901 );
xor \U$29182 ( \37903 , \37891 , \37902 );
xor \U$29183 ( \37904 , \37882 , \37903 );
and \U$29184 ( \37905 , \37523 , \37534 );
and \U$29185 ( \37906 , \37534 , \37548 );
and \U$29186 ( \37907 , \37523 , \37548 );
or \U$29187 ( \37908 , \37905 , \37906 , \37907 );
and \U$29188 ( \37909 , \37513 , \37517 );
and \U$29189 ( \37910 , \37517 , \37522 );
and \U$29190 ( \37911 , \37513 , \37522 );
or \U$29191 ( \37912 , \37909 , \37910 , \37911 );
and \U$29192 ( \37913 , \37527 , \37531 );
and \U$29193 ( \37914 , \37531 , \37533 );
and \U$29194 ( \37915 , \37527 , \37533 );
or \U$29195 ( \37916 , \37913 , \37914 , \37915 );
xor \U$29196 ( \37917 , \37912 , \37916 );
and \U$29197 ( \37918 , \37538 , \37542 );
and \U$29198 ( \37919 , \37542 , \37547 );
and \U$29199 ( \37920 , \37538 , \37547 );
or \U$29200 ( \37921 , \37918 , \37919 , \37920 );
xor \U$29201 ( \37922 , \37917 , \37921 );
xor \U$29202 ( \37923 , \37908 , \37922 );
and \U$29203 ( \37924 , \30268 , \21005 );
and \U$29204 ( \37925 , \30802 , \20557 );
nor \U$29205 ( \37926 , \37924 , \37925 );
xnor \U$29206 ( \37927 , \37926 , \21011 );
and \U$29207 ( \37928 , \19032 , \32854 );
and \U$29208 ( \37929 , \19558 , \32067 );
nor \U$29209 ( \37930 , \37928 , \37929 );
xnor \U$29210 ( \37931 , \37930 , \32805 );
xor \U$29211 ( \37932 , \37927 , \37931 );
and \U$29212 ( \37933 , \18035 , \32802 );
xor \U$29213 ( \37934 , \37932 , \37933 );
and \U$29214 ( \37935 , \26829 , \24138 );
and \U$29215 ( \37936 , \27313 , \23630 );
nor \U$29216 ( \37937 , \37935 , \37936 );
xnor \U$29217 ( \37938 , \37937 , \24144 );
and \U$29218 ( \37939 , \22090 , \29070 );
and \U$29219 ( \37940 , \22556 , \28526 );
nor \U$29220 ( \37941 , \37939 , \37940 );
xnor \U$29221 ( \37942 , \37941 , \29076 );
xor \U$29222 ( \37943 , \37938 , \37942 );
and \U$29223 ( \37944 , \20544 , \30823 );
and \U$29224 ( \37945 , \21033 , \30246 );
nor \U$29225 ( \37946 , \37944 , \37945 );
xnor \U$29226 ( \37947 , \37946 , \30813 );
xor \U$29227 ( \37948 , \37943 , \37947 );
xor \U$29228 ( \37949 , \37934 , \37948 );
not \U$29229 ( \37950 , \18046 );
and \U$29230 ( \37951 , \32054 , \19534 );
and \U$29231 ( \37952 , \32794 , \19045 );
nor \U$29232 ( \37953 , \37951 , \37952 );
xnor \U$29233 ( \37954 , \37953 , \19540 );
xor \U$29234 ( \37955 , \37950 , \37954 );
and \U$29235 ( \37956 , \28534 , \22542 );
and \U$29236 ( \37957 , \29084 , \22103 );
nor \U$29237 ( \37958 , \37956 , \37957 );
xnor \U$29238 ( \37959 , \37958 , \22548 );
xor \U$29239 ( \37960 , \37955 , \37959 );
xor \U$29240 ( \37961 , \37949 , \37960 );
xor \U$29241 ( \37962 , \37923 , \37961 );
xor \U$29242 ( \37963 , \37904 , \37962 );
xor \U$29243 ( \37964 , \37878 , \37963 );
and \U$29244 ( \37965 , \37500 , \37550 );
and \U$29245 ( \37966 , \37550 , \37596 );
and \U$29246 ( \37967 , \37500 , \37596 );
or \U$29247 ( \37968 , \37965 , \37966 , \37967 );
xor \U$29248 ( \37969 , \37964 , \37968 );
and \U$29249 ( \37970 , \37597 , \37601 );
and \U$29250 ( \37971 , \37602 , \37605 );
or \U$29251 ( \37972 , \37970 , \37971 );
xor \U$29252 ( \37973 , \37969 , \37972 );
buf g9b87 ( \37974_nG9b87 , \37973 );
and \U$29253 ( \37975 , \10704 , \37974_nG9b87 );
or \U$29254 ( \37976 , \37869 , \37975 );
xor \U$29255 ( \37977 , \10703 , \37976 );
buf \U$29256 ( \37978 , \37977 );
buf \U$29258 ( \37979 , \37978 );
xor \U$29259 ( \37980 , \37868 , \37979 );
buf \U$29260 ( \37981 , \37980 );
xor \U$29261 ( \37982 , \37855 , \37981 );
buf \U$29262 ( \37983 , \37982 );
and \U$29263 ( \37984 , \37620 , \37625 );
and \U$29264 ( \37985 , \37620 , \37632 );
and \U$29265 ( \37986 , \37625 , \37632 );
or \U$29266 ( \37987 , \37984 , \37985 , \37986 );
buf \U$29267 ( \37988 , \37987 );
and \U$29268 ( \37989 , \37668 , \37681 );
and \U$29269 ( \37990 , \37668 , \37688 );
and \U$29270 ( \37991 , \37681 , \37688 );
or \U$29271 ( \37992 , \37989 , \37990 , \37991 );
buf \U$29272 ( \37993 , \37992 );
and \U$29273 ( \37994 , \17297 , \33181_nG9bae );
and \U$29274 ( \37995 , \17294 , \33613_nG9bab );
or \U$29275 ( \37996 , \37994 , \37995 );
xor \U$29276 ( \37997 , \17293 , \37996 );
buf \U$29277 ( \37998 , \37997 );
buf \U$29279 ( \37999 , \37998 );
xor \U$29280 ( \38000 , \37993 , \37999 );
and \U$29281 ( \38001 , \14631 , \34643_nG9ba2 );
and \U$29282 ( \38002 , \14628 , \35094_nG9b9f );
or \U$29283 ( \38003 , \38001 , \38002 );
xor \U$29284 ( \38004 , \14627 , \38003 );
buf \U$29285 ( \38005 , \38004 );
buf \U$29287 ( \38006 , \38005 );
xor \U$29288 ( \38007 , \38000 , \38006 );
buf \U$29289 ( \38008 , \38007 );
xor \U$29290 ( \38009 , \37988 , \38008 );
and \U$29291 ( \38010 , \37473 , \37479 );
and \U$29292 ( \38011 , \37473 , \37486 );
and \U$29293 ( \38012 , \37479 , \37486 );
or \U$29294 ( \38013 , \38010 , \38011 , \38012 );
buf \U$29295 ( \38014 , \38013 );
and \U$29296 ( \38015 , \37403 , \37409 );
and \U$29297 ( \38016 , \37403 , \37416 );
and \U$29298 ( \38017 , \37409 , \37416 );
or \U$29299 ( \38018 , \38015 , \38016 , \38017 );
buf \U$29300 ( \38019 , \38018 );
and \U$29301 ( \38020 , \28118 , \22129_nG9bd8 );
and \U$29302 ( \38021 , \28115 , \22629_nG9bd5 );
or \U$29303 ( \38022 , \38020 , \38021 );
xor \U$29304 ( \38023 , \28114 , \38022 );
buf \U$29305 ( \38024 , \38023 );
buf \U$29307 ( \38025 , \38024 );
xor \U$29308 ( \38026 , \38019 , \38025 );
and \U$29309 ( \38027 , \26431 , \23696_nG9bd2 );
and \U$29310 ( \38028 , \26428 , \24226_nG9bcf );
or \U$29311 ( \38029 , \38027 , \38028 );
xor \U$29312 ( \38030 , \26427 , \38029 );
buf \U$29313 ( \38031 , \38030 );
buf \U$29315 ( \38032 , \38031 );
xor \U$29316 ( \38033 , \38026 , \38032 );
buf \U$29317 ( \38034 , \38033 );
xor \U$29318 ( \38035 , \38014 , \38034 );
and \U$29319 ( \38036 , \13370 , \35570_nG9b9c );
and \U$29320 ( \38037 , \13367 , \35801_nG9b99 );
or \U$29321 ( \38038 , \38036 , \38037 );
xor \U$29322 ( \38039 , \13366 , \38038 );
buf \U$29323 ( \38040 , \38039 );
buf \U$29325 ( \38041 , \38040 );
xor \U$29326 ( \38042 , \38035 , \38041 );
buf \U$29327 ( \38043 , \38042 );
xor \U$29328 ( \38044 , \38009 , \38043 );
buf \U$29329 ( \38045 , \38044 );
xor \U$29330 ( \38046 , \37983 , \38045 );
and \U$29331 ( \38047 , \37467 , \37614 );
and \U$29332 ( \38048 , \37467 , \37634 );
and \U$29333 ( \38049 , \37614 , \37634 );
or \U$29334 ( \38050 , \38047 , \38048 , \38049 );
buf \U$29335 ( \38051 , \38050 );
xor \U$29336 ( \38052 , \38046 , \38051 );
buf \U$29337 ( \38053 , \38052 );
xor \U$29338 ( \38054 , \37814 , \38053 );
and \U$29339 ( \38055 , \37730 , \38054 );
and \U$29341 ( \38056 , \37724 , \37729 );
or \U$29343 ( \38057 , 1'b0 , \38056 , 1'b0 );
xor \U$29344 ( \38058 , \38055 , \38057 );
and \U$29346 ( \38059 , \37717 , \37723 );
and \U$29347 ( \38060 , \37719 , \37723 );
or \U$29348 ( \38061 , 1'b0 , \38059 , \38060 );
xor \U$29349 ( \38062 , \38058 , \38061 );
xor \U$29356 ( \38063 , \38062 , 1'b0 );
and \U$29357 ( \38064 , \37735 , \37813 );
and \U$29358 ( \38065 , \37735 , \38053 );
and \U$29359 ( \38066 , \37813 , \38053 );
or \U$29360 ( \38067 , \38064 , \38065 , \38066 );
xor \U$29361 ( \38068 , \38063 , \38067 );
and \U$29362 ( \38069 , \37983 , \38045 );
and \U$29363 ( \38070 , \37983 , \38051 );
and \U$29364 ( \38071 , \38045 , \38051 );
or \U$29365 ( \38072 , \38069 , \38070 , \38071 );
buf \U$29366 ( \38073 , \38072 );
and \U$29367 ( \38074 , \37796 , \37801 );
and \U$29368 ( \38075 , \37796 , \37807 );
and \U$29369 ( \38076 , \37801 , \37807 );
or \U$29370 ( \38077 , \38074 , \38075 , \38076 );
buf \U$29371 ( \38078 , \38077 );
and \U$29372 ( \38079 , \21658 , \29179_nG9bbd );
and \U$29373 ( \38080 , \21655 , \30366_nG9bba );
or \U$29374 ( \38081 , \38079 , \38080 );
xor \U$29375 ( \38082 , \21654 , \38081 );
buf \U$29376 ( \38083 , \38082 );
buf \U$29378 ( \38084 , \38083 );
and \U$29379 ( \38085 , \18702 , \32888_nG9bb1 );
and \U$29380 ( \38086 , \18699 , \33181_nG9bae );
or \U$29381 ( \38087 , \38085 , \38086 );
xor \U$29382 ( \38088 , \18698 , \38087 );
buf \U$29383 ( \38089 , \38088 );
buf \U$29385 ( \38090 , \38089 );
xor \U$29386 ( \38091 , \38084 , \38090 );
and \U$29387 ( \38092 , \17297 , \33613_nG9bab );
and \U$29388 ( \38093 , \17294 , \34041_nG9ba8 );
or \U$29389 ( \38094 , \38092 , \38093 );
xor \U$29390 ( \38095 , \17293 , \38094 );
buf \U$29391 ( \38096 , \38095 );
buf \U$29393 ( \38097 , \38096 );
xor \U$29394 ( \38098 , \38091 , \38097 );
buf \U$29395 ( \38099 , \38098 );
and \U$29396 ( \38100 , \38014 , \38034 );
and \U$29397 ( \38101 , \38014 , \38041 );
and \U$29398 ( \38102 , \38034 , \38041 );
or \U$29399 ( \38103 , \38100 , \38101 , \38102 );
buf \U$29400 ( \38104 , \38103 );
xor \U$29401 ( \38105 , \38099 , \38104 );
and \U$29402 ( \38106 , \37993 , \37999 );
and \U$29403 ( \38107 , \37993 , \38006 );
and \U$29404 ( \38108 , \37999 , \38006 );
or \U$29405 ( \38109 , \38106 , \38107 , \38108 );
buf \U$29406 ( \38110 , \38109 );
xor \U$29407 ( \38111 , \38105 , \38110 );
buf \U$29408 ( \38112 , \38111 );
xor \U$29409 ( \38113 , \38078 , \38112 );
and \U$29410 ( \38114 , \37988 , \38008 );
and \U$29411 ( \38115 , \37988 , \38043 );
and \U$29412 ( \38116 , \38008 , \38043 );
or \U$29413 ( \38117 , \38114 , \38115 , \38116 );
buf \U$29414 ( \38118 , \38117 );
xor \U$29415 ( \38119 , \38113 , \38118 );
buf \U$29416 ( \38120 , \38119 );
xor \U$29417 ( \38121 , \38073 , \38120 );
and \U$29418 ( \38122 , \37751 , \37756 );
and \U$29419 ( \38123 , \37751 , \37809 );
and \U$29420 ( \38124 , \37756 , \37809 );
or \U$29421 ( \38125 , \38122 , \38123 , \38124 );
buf \U$29422 ( \38126 , \38125 );
xor \U$29423 ( \38127 , \38121 , \38126 );
buf \U$29424 ( \38128 , \38127 );
and \U$29425 ( \38129 , \37740 , \37745 );
and \U$29426 ( \38130 , \37740 , \37811 );
and \U$29427 ( \38131 , \37745 , \37811 );
or \U$29428 ( \38132 , \38129 , \38130 , \38131 );
buf \U$29429 ( \38133 , \38132 );
xor \U$29430 ( \38134 , \38128 , \38133 );
and \U$29431 ( \38135 , \37849 , \37854 );
and \U$29432 ( \38136 , \37849 , \37981 );
and \U$29433 ( \38137 , \37854 , \37981 );
or \U$29434 ( \38138 , \38135 , \38136 , \38137 );
buf \U$29435 ( \38139 , \38138 );
and \U$29436 ( \38140 , \37861 , \37867 );
and \U$29437 ( \38141 , \37861 , \37979 );
and \U$29438 ( \38142 , \37867 , \37979 );
or \U$29439 ( \38143 , \38140 , \38141 , \38142 );
buf \U$29440 ( \38144 , \38143 );
and \U$29441 ( \38145 , \28118 , \22629_nG9bd5 );
and \U$29442 ( \38146 , \28115 , \23696_nG9bd2 );
or \U$29443 ( \38147 , \38145 , \38146 );
xor \U$29444 ( \38148 , \28114 , \38147 );
buf \U$29445 ( \38149 , \38148 );
buf \U$29447 ( \38150 , \38149 );
and \U$29448 ( \38151 , \26431 , \24226_nG9bcf );
and \U$29449 ( \38152 , \26428 , \25298_nG9bcc );
or \U$29450 ( \38153 , \38151 , \38152 );
xor \U$29451 ( \38154 , \26427 , \38153 );
buf \U$29452 ( \38155 , \38154 );
buf \U$29454 ( \38156 , \38155 );
xor \U$29455 ( \38157 , \38150 , \38156 );
and \U$29456 ( \38158 , \24792 , \25860_nG9bc9 );
and \U$29457 ( \38159 , \24789 , \26887_nG9bc6 );
or \U$29458 ( \38160 , \38158 , \38159 );
xor \U$29459 ( \38161 , \24788 , \38160 );
buf \U$29460 ( \38162 , \38161 );
buf \U$29462 ( \38163 , \38162 );
xor \U$29463 ( \38164 , \38157 , \38163 );
buf \U$29464 ( \38165 , \38164 );
and \U$29465 ( \38166 , \15940 , \34294_nG9ba5 );
and \U$29466 ( \38167 , \15937 , \34643_nG9ba2 );
or \U$29467 ( \38168 , \38166 , \38167 );
xor \U$29468 ( \38169 , \15936 , \38168 );
buf \U$29469 ( \38170 , \38169 );
buf \U$29471 ( \38171 , \38170 );
xor \U$29472 ( \38172 , \38165 , \38171 );
and \U$29473 ( \38173 , \13370 , \35801_nG9b99 );
and \U$29474 ( \38174 , \13367 , \36172_nG9b96 );
or \U$29475 ( \38175 , \38173 , \38174 );
xor \U$29476 ( \38176 , \13366 , \38175 );
buf \U$29477 ( \38177 , \38176 );
buf \U$29479 ( \38178 , \38177 );
xor \U$29480 ( \38179 , \38172 , \38178 );
buf \U$29481 ( \38180 , \38179 );
xor \U$29482 ( \38181 , \38144 , \38180 );
and \U$29483 ( \38182 , \37819 , \37840 );
and \U$29484 ( \38183 , \37819 , \37847 );
and \U$29485 ( \38184 , \37840 , \37847 );
or \U$29486 ( \38185 , \38182 , \38183 , \38184 );
buf \U$29487 ( \38186 , \38185 );
xor \U$29488 ( \38187 , \38181 , \38186 );
buf \U$29489 ( \38188 , \38187 );
xor \U$29490 ( \38189 , \38139 , \38188 );
and \U$29491 ( \38190 , \37781 , \37787 );
and \U$29492 ( \38191 , \37781 , \37794 );
and \U$29493 ( \38192 , \37787 , \37794 );
or \U$29494 ( \38193 , \38190 , \38191 , \38192 );
buf \U$29495 ( \38194 , \38193 );
and \U$29496 ( \38195 , \37770 , \37772 );
and \U$29497 ( \38196 , \37770 , \37779 );
and \U$29498 ( \38197 , \37772 , \37779 );
or \U$29499 ( \38198 , \38195 , \38196 , \38197 );
buf \U$29500 ( \38199 , \38198 );
and \U$29501 ( \38200 , \23201 , \27416_nG9bc3 );
and \U$29502 ( \38201 , \23198 , \28602_nG9bc0 );
or \U$29503 ( \38202 , \38200 , \38201 );
xor \U$29504 ( \38203 , \23197 , \38202 );
buf \U$29505 ( \38204 , \38203 );
buf \U$29507 ( \38205 , \38204 );
xor \U$29508 ( \38206 , \38199 , \38205 );
and \U$29509 ( \38207 , \20155 , \30940_nG9bb7 );
and \U$29510 ( \38208 , \20152 , \32179_nG9bb4 );
or \U$29511 ( \38209 , \38207 , \38208 );
xor \U$29512 ( \38210 , \20151 , \38209 );
buf \U$29513 ( \38211 , \38210 );
buf \U$29515 ( \38212 , \38211 );
xor \U$29516 ( \38213 , \38206 , \38212 );
buf \U$29517 ( \38214 , \38213 );
xor \U$29518 ( \38215 , \38194 , \38214 );
and \U$29519 ( \38216 , \12157 , \36589_nG9b93 );
and \U$29520 ( \38217 , \12154 , \36986_nG9b90 );
or \U$29521 ( \38218 , \38216 , \38217 );
xor \U$29522 ( \38219 , \12153 , \38218 );
buf \U$29523 ( \38220 , \38219 );
buf \U$29525 ( \38221 , \38220 );
xor \U$29526 ( \38222 , \38215 , \38221 );
buf \U$29527 ( \38223 , \38222 );
and \U$29528 ( \38224 , \37825 , \37831 );
and \U$29529 ( \38225 , \37825 , \37838 );
and \U$29530 ( \38226 , \37831 , \37838 );
or \U$29531 ( \38227 , \38224 , \38225 , \38226 );
buf \U$29532 ( \38228 , \38227 );
and \U$29533 ( \38229 , \10421 , \37250_nG9b8d );
and \U$29534 ( \38230 , \10418 , \37607_nG9b8a );
or \U$29535 ( \38231 , \38229 , \38230 );
xor \U$29536 ( \38232 , \10417 , \38231 );
buf \U$29537 ( \38233 , \38232 );
buf \U$29539 ( \38234 , \38233 );
xor \U$29540 ( \38235 , \38228 , \38234 );
and \U$29541 ( \38236 , \10707 , \37974_nG9b87 );
and \U$29542 ( \38237 , \37882 , \37903 );
and \U$29543 ( \38238 , \37903 , \37962 );
and \U$29544 ( \38239 , \37882 , \37962 );
or \U$29545 ( \38240 , \38237 , \38238 , \38239 );
and \U$29546 ( \38241 , \37934 , \37948 );
and \U$29547 ( \38242 , \37948 , \37960 );
and \U$29548 ( \38243 , \37934 , \37960 );
or \U$29549 ( \38244 , \38241 , \38242 , \38243 );
and \U$29550 ( \38245 , \37938 , \37942 );
and \U$29551 ( \38246 , \37942 , \37947 );
and \U$29552 ( \38247 , \37938 , \37947 );
or \U$29553 ( \38248 , \38245 , \38246 , \38247 );
and \U$29554 ( \38249 , \37950 , \37954 );
and \U$29555 ( \38250 , \37954 , \37959 );
and \U$29556 ( \38251 , \37950 , \37959 );
or \U$29557 ( \38252 , \38249 , \38250 , \38251 );
xor \U$29558 ( \38253 , \38248 , \38252 );
and \U$29559 ( \38254 , \32794 , \19534 );
not \U$29560 ( \38255 , \38254 );
xnor \U$29561 ( \38256 , \38255 , \19540 );
not \U$29562 ( \38257 , \38256 );
xor \U$29563 ( \38258 , \38253 , \38257 );
xor \U$29564 ( \38259 , \38244 , \38258 );
and \U$29565 ( \38260 , \37927 , \37931 );
and \U$29566 ( \38261 , \37931 , \37933 );
and \U$29567 ( \38262 , \37927 , \37933 );
or \U$29568 ( \38263 , \38260 , \38261 , \38262 );
and \U$29569 ( \38264 , \30802 , \21005 );
and \U$29570 ( \38265 , \32054 , \20557 );
nor \U$29571 ( \38266 , \38264 , \38265 );
xnor \U$29572 ( \38267 , \38266 , \21011 );
and \U$29573 ( \38268 , \25815 , \25826 );
and \U$29574 ( \38269 , \26829 , \25264 );
nor \U$29575 ( \38270 , \38268 , \38269 );
xnor \U$29576 ( \38271 , \38270 , \25773 );
xor \U$29577 ( \38272 , \38267 , \38271 );
and \U$29578 ( \38273 , \19032 , \32802 );
xor \U$29579 ( \38274 , \38272 , \38273 );
xor \U$29580 ( \38275 , \38263 , \38274 );
and \U$29581 ( \38276 , \27313 , \24138 );
and \U$29582 ( \38277 , \28534 , \23630 );
nor \U$29583 ( \38278 , \38276 , \38277 );
xnor \U$29584 ( \38279 , \38278 , \24144 );
and \U$29585 ( \38280 , \21033 , \30823 );
and \U$29586 ( \38281 , \22090 , \30246 );
nor \U$29587 ( \38282 , \38280 , \38281 );
xnor \U$29588 ( \38283 , \38282 , \30813 );
xor \U$29589 ( \38284 , \38279 , \38283 );
and \U$29590 ( \38285 , \19558 , \32854 );
and \U$29591 ( \38286 , \20544 , \32067 );
nor \U$29592 ( \38287 , \38285 , \38286 );
xnor \U$29593 ( \38288 , \38287 , \32805 );
xor \U$29594 ( \38289 , \38284 , \38288 );
xor \U$29595 ( \38290 , \38275 , \38289 );
xor \U$29596 ( \38291 , \38259 , \38290 );
xor \U$29597 ( \38292 , \38240 , \38291 );
and \U$29598 ( \38293 , \37886 , \37890 );
and \U$29599 ( \38294 , \37890 , \37902 );
and \U$29600 ( \38295 , \37886 , \37902 );
or \U$29601 ( \38296 , \38293 , \38294 , \38295 );
and \U$29602 ( \38297 , \37908 , \37922 );
and \U$29603 ( \38298 , \37922 , \37961 );
and \U$29604 ( \38299 , \37908 , \37961 );
or \U$29605 ( \38300 , \38297 , \38298 , \38299 );
xor \U$29606 ( \38301 , \38296 , \38300 );
and \U$29607 ( \38302 , \37912 , \37916 );
and \U$29608 ( \38303 , \37916 , \37921 );
and \U$29609 ( \38304 , \37912 , \37921 );
or \U$29610 ( \38305 , \38302 , \38303 , \38304 );
and \U$29611 ( \38306 , \37892 , \37896 );
and \U$29612 ( \38307 , \37896 , \37901 );
and \U$29613 ( \38308 , \37892 , \37901 );
or \U$29614 ( \38309 , \38306 , \38307 , \38308 );
xor \U$29615 ( \38310 , \38305 , \38309 );
and \U$29616 ( \38311 , \29084 , \22542 );
and \U$29617 ( \38312 , \30268 , \22103 );
nor \U$29618 ( \38313 , \38311 , \38312 );
xnor \U$29619 ( \38314 , \38313 , \22548 );
and \U$29620 ( \38315 , \24199 , \27397 );
and \U$29621 ( \38316 , \25272 , \26807 );
nor \U$29622 ( \38317 , \38315 , \38316 );
xnor \U$29623 ( \38318 , \38317 , \27295 );
xor \U$29624 ( \38319 , \38314 , \38318 );
and \U$29625 ( \38320 , \22556 , \29070 );
and \U$29626 ( \38321 , \23617 , \28526 );
nor \U$29627 ( \38322 , \38320 , \38321 );
xnor \U$29628 ( \38323 , \38322 , \29076 );
xor \U$29629 ( \38324 , \38319 , \38323 );
xor \U$29630 ( \38325 , \38310 , \38324 );
xor \U$29631 ( \38326 , \38301 , \38325 );
xor \U$29632 ( \38327 , \38292 , \38326 );
and \U$29633 ( \38328 , \37873 , \37877 );
and \U$29634 ( \38329 , \37877 , \37963 );
and \U$29635 ( \38330 , \37873 , \37963 );
or \U$29636 ( \38331 , \38328 , \38329 , \38330 );
xor \U$29637 ( \38332 , \38327 , \38331 );
and \U$29638 ( \38333 , \37964 , \37968 );
and \U$29639 ( \38334 , \37969 , \37972 );
or \U$29640 ( \38335 , \38333 , \38334 );
xor \U$29641 ( \38336 , \38332 , \38335 );
buf g9b84 ( \38337_nG9b84 , \38336 );
and \U$29642 ( \38338 , \10704 , \38337_nG9b84 );
or \U$29643 ( \38339 , \38236 , \38338 );
xor \U$29644 ( \38340 , \10703 , \38339 );
buf \U$29645 ( \38341 , \38340 );
buf \U$29647 ( \38342 , \38341 );
xor \U$29648 ( \38343 , \38235 , \38342 );
buf \U$29649 ( \38344 , \38343 );
xor \U$29650 ( \38345 , \38223 , \38344 );
and \U$29651 ( \38346 , \38019 , \38025 );
and \U$29652 ( \38347 , \38019 , \38032 );
and \U$29653 ( \38348 , \38025 , \38032 );
or \U$29654 ( \38349 , \38346 , \38347 , \38348 );
buf \U$29655 ( \38350 , \38349 );
and \U$29657 ( \38351 , \32916 , \19091_nG9be4 );
or \U$29658 ( \38352 , 1'b0 , \38351 );
xor \U$29659 ( \38353 , 1'b0 , \38352 );
buf \U$29660 ( \38354 , \38353 );
buf \U$29662 ( \38355 , \38354 );
and \U$29663 ( \38356 , \29853 , \21086_nG9bdb );
and \U$29664 ( \38357 , \29850 , \22129_nG9bd8 );
or \U$29665 ( \38358 , \38356 , \38357 );
xor \U$29666 ( \38359 , \29849 , \38358 );
buf \U$29667 ( \38360 , \38359 );
buf \U$29669 ( \38361 , \38360 );
xor \U$29670 ( \38362 , \38355 , \38361 );
buf \U$29671 ( \38363 , \38362 );
and \U$29672 ( \38364 , \37762 , \37768 );
buf \U$29673 ( \38365 , \38364 );
xor \U$29674 ( \38366 , \38363 , \38365 );
and \U$29675 ( \38367 , \31636 , \19586_nG9be1 );
and \U$29676 ( \38368 , \31633 , \20608_nG9bde );
or \U$29677 ( \38369 , \38367 , \38368 );
xor \U$29678 ( \38370 , \31632 , \38369 );
buf \U$29679 ( \38371 , \38370 );
buf \U$29681 ( \38372 , \38371 );
xor \U$29682 ( \38373 , \38366 , \38372 );
buf \U$29683 ( \38374 , \38373 );
xor \U$29684 ( \38375 , \38350 , \38374 );
and \U$29685 ( \38376 , \14631 , \35094_nG9b9f );
and \U$29686 ( \38377 , \14628 , \35570_nG9b9c );
or \U$29687 ( \38378 , \38376 , \38377 );
xor \U$29688 ( \38379 , \14627 , \38378 );
buf \U$29689 ( \38380 , \38379 );
buf \U$29691 ( \38381 , \38380 );
xor \U$29692 ( \38382 , \38375 , \38381 );
buf \U$29693 ( \38383 , \38382 );
xor \U$29694 ( \38384 , \38345 , \38383 );
buf \U$29695 ( \38385 , \38384 );
xor \U$29696 ( \38386 , \38189 , \38385 );
buf \U$29697 ( \38387 , \38386 );
xor \U$29698 ( \38388 , \38134 , \38387 );
and \U$29699 ( \38389 , \38068 , \38388 );
and \U$29701 ( \38390 , \38062 , \38067 );
or \U$29703 ( \38391 , 1'b0 , \38390 , 1'b0 );
xor \U$29704 ( \38392 , \38389 , \38391 );
and \U$29706 ( \38393 , \38055 , \38061 );
and \U$29707 ( \38394 , \38057 , \38061 );
or \U$29708 ( \38395 , 1'b0 , \38393 , \38394 );
xor \U$29709 ( \38396 , \38392 , \38395 );
xor \U$29716 ( \38397 , \38396 , 1'b0 );
and \U$29717 ( \38398 , \38165 , \38171 );
and \U$29718 ( \38399 , \38165 , \38178 );
and \U$29719 ( \38400 , \38171 , \38178 );
or \U$29720 ( \38401 , \38398 , \38399 , \38400 );
buf \U$29721 ( \38402 , \38401 );
and \U$29722 ( \38403 , \38350 , \38374 );
and \U$29723 ( \38404 , \38350 , \38381 );
and \U$29724 ( \38405 , \38374 , \38381 );
or \U$29725 ( \38406 , \38403 , \38404 , \38405 );
buf \U$29726 ( \38407 , \38406 );
xor \U$29727 ( \38408 , \38402 , \38407 );
and \U$29729 ( \38409 , \32916 , \19586_nG9be1 );
or \U$29730 ( \38410 , 1'b0 , \38409 );
xor \U$29731 ( \38411 , 1'b0 , \38410 );
buf \U$29732 ( \38412 , \38411 );
buf \U$29734 ( \38413 , \38412 );
and \U$29735 ( \38414 , \31636 , \20608_nG9bde );
and \U$29736 ( \38415 , \31633 , \21086_nG9bdb );
or \U$29737 ( \38416 , \38414 , \38415 );
xor \U$29738 ( \38417 , \31632 , \38416 );
buf \U$29739 ( \38418 , \38417 );
buf \U$29741 ( \38419 , \38418 );
xor \U$29742 ( \38420 , \38413 , \38419 );
buf \U$29743 ( \38421 , \38420 );
and \U$29744 ( \38422 , \38355 , \38361 );
buf \U$29745 ( \38423 , \38422 );
xor \U$29746 ( \38424 , \38421 , \38423 );
and \U$29747 ( \38425 , \29853 , \22129_nG9bd8 );
and \U$29748 ( \38426 , \29850 , \22629_nG9bd5 );
or \U$29749 ( \38427 , \38425 , \38426 );
xor \U$29750 ( \38428 , \29849 , \38427 );
buf \U$29751 ( \38429 , \38428 );
buf \U$29753 ( \38430 , \38429 );
xor \U$29754 ( \38431 , \38424 , \38430 );
buf \U$29755 ( \38432 , \38431 );
and \U$29756 ( \38433 , \20155 , \32179_nG9bb4 );
and \U$29757 ( \38434 , \20152 , \32888_nG9bb1 );
or \U$29758 ( \38435 , \38433 , \38434 );
xor \U$29759 ( \38436 , \20151 , \38435 );
buf \U$29760 ( \38437 , \38436 );
buf \U$29762 ( \38438 , \38437 );
xor \U$29763 ( \38439 , \38432 , \38438 );
and \U$29764 ( \38440 , \18702 , \33181_nG9bae );
and \U$29765 ( \38441 , \18699 , \33613_nG9bab );
or \U$29766 ( \38442 , \38440 , \38441 );
xor \U$29767 ( \38443 , \18698 , \38442 );
buf \U$29768 ( \38444 , \38443 );
buf \U$29770 ( \38445 , \38444 );
xor \U$29771 ( \38446 , \38439 , \38445 );
buf \U$29772 ( \38447 , \38446 );
xor \U$29773 ( \38448 , \38408 , \38447 );
buf \U$29774 ( \38449 , \38448 );
and \U$29775 ( \38450 , \38144 , \38180 );
and \U$29776 ( \38451 , \38144 , \38186 );
and \U$29777 ( \38452 , \38180 , \38186 );
or \U$29778 ( \38453 , \38450 , \38451 , \38452 );
buf \U$29779 ( \38454 , \38453 );
xor \U$29780 ( \38455 , \38449 , \38454 );
and \U$29781 ( \38456 , \38099 , \38104 );
and \U$29782 ( \38457 , \38099 , \38110 );
and \U$29783 ( \38458 , \38104 , \38110 );
or \U$29784 ( \38459 , \38456 , \38457 , \38458 );
buf \U$29785 ( \38460 , \38459 );
xor \U$29786 ( \38461 , \38455 , \38460 );
buf \U$29787 ( \38462 , \38461 );
and \U$29788 ( \38463 , \38078 , \38112 );
and \U$29789 ( \38464 , \38078 , \38118 );
and \U$29790 ( \38465 , \38112 , \38118 );
or \U$29791 ( \38466 , \38463 , \38464 , \38465 );
buf \U$29792 ( \38467 , \38466 );
xor \U$29793 ( \38468 , \38462 , \38467 );
and \U$29794 ( \38469 , \38139 , \38188 );
and \U$29795 ( \38470 , \38139 , \38385 );
and \U$29796 ( \38471 , \38188 , \38385 );
or \U$29797 ( \38472 , \38469 , \38470 , \38471 );
buf \U$29798 ( \38473 , \38472 );
xor \U$29799 ( \38474 , \38468 , \38473 );
buf \U$29800 ( \38475 , \38474 );
and \U$29801 ( \38476 , \38073 , \38120 );
and \U$29802 ( \38477 , \38073 , \38126 );
and \U$29803 ( \38478 , \38120 , \38126 );
or \U$29804 ( \38479 , \38476 , \38477 , \38478 );
buf \U$29805 ( \38480 , \38479 );
xor \U$29806 ( \38481 , \38475 , \38480 );
and \U$29807 ( \38482 , \38223 , \38344 );
and \U$29808 ( \38483 , \38223 , \38383 );
and \U$29809 ( \38484 , \38344 , \38383 );
or \U$29810 ( \38485 , \38482 , \38483 , \38484 );
buf \U$29811 ( \38486 , \38485 );
and \U$29812 ( \38487 , \38194 , \38214 );
and \U$29813 ( \38488 , \38194 , \38221 );
and \U$29814 ( \38489 , \38214 , \38221 );
or \U$29815 ( \38490 , \38487 , \38488 , \38489 );
buf \U$29816 ( \38491 , \38490 );
and \U$29817 ( \38492 , \38228 , \38234 );
and \U$29818 ( \38493 , \38228 , \38342 );
and \U$29819 ( \38494 , \38234 , \38342 );
or \U$29820 ( \38495 , \38492 , \38493 , \38494 );
buf \U$29821 ( \38496 , \38495 );
xor \U$29822 ( \38497 , \38491 , \38496 );
and \U$29823 ( \38498 , \38150 , \38156 );
and \U$29824 ( \38499 , \38150 , \38163 );
and \U$29825 ( \38500 , \38156 , \38163 );
or \U$29826 ( \38501 , \38498 , \38499 , \38500 );
buf \U$29827 ( \38502 , \38501 );
and \U$29828 ( \38503 , \15940 , \34643_nG9ba2 );
and \U$29829 ( \38504 , \15937 , \35094_nG9b9f );
or \U$29830 ( \38505 , \38503 , \38504 );
xor \U$29831 ( \38506 , \15936 , \38505 );
buf \U$29832 ( \38507 , \38506 );
buf \U$29834 ( \38508 , \38507 );
xor \U$29835 ( \38509 , \38502 , \38508 );
and \U$29836 ( \38510 , \14631 , \35570_nG9b9c );
and \U$29837 ( \38511 , \14628 , \35801_nG9b99 );
or \U$29838 ( \38512 , \38510 , \38511 );
xor \U$29839 ( \38513 , \14627 , \38512 );
buf \U$29840 ( \38514 , \38513 );
buf \U$29842 ( \38515 , \38514 );
xor \U$29843 ( \38516 , \38509 , \38515 );
buf \U$29844 ( \38517 , \38516 );
xor \U$29845 ( \38518 , \38497 , \38517 );
buf \U$29846 ( \38519 , \38518 );
xor \U$29847 ( \38520 , \38486 , \38519 );
and \U$29848 ( \38521 , \38084 , \38090 );
and \U$29849 ( \38522 , \38084 , \38097 );
and \U$29850 ( \38523 , \38090 , \38097 );
or \U$29851 ( \38524 , \38521 , \38522 , \38523 );
buf \U$29852 ( \38525 , \38524 );
and \U$29853 ( \38526 , \38363 , \38365 );
and \U$29854 ( \38527 , \38363 , \38372 );
and \U$29855 ( \38528 , \38365 , \38372 );
or \U$29856 ( \38529 , \38526 , \38527 , \38528 );
buf \U$29857 ( \38530 , \38529 );
and \U$29858 ( \38531 , \23201 , \28602_nG9bc0 );
and \U$29859 ( \38532 , \23198 , \29179_nG9bbd );
or \U$29860 ( \38533 , \38531 , \38532 );
xor \U$29861 ( \38534 , \23197 , \38533 );
buf \U$29862 ( \38535 , \38534 );
buf \U$29864 ( \38536 , \38535 );
xor \U$29865 ( \38537 , \38530 , \38536 );
and \U$29866 ( \38538 , \21658 , \30366_nG9bba );
and \U$29867 ( \38539 , \21655 , \30940_nG9bb7 );
or \U$29868 ( \38540 , \38538 , \38539 );
xor \U$29869 ( \38541 , \21654 , \38540 );
buf \U$29870 ( \38542 , \38541 );
buf \U$29872 ( \38543 , \38542 );
xor \U$29873 ( \38544 , \38537 , \38543 );
buf \U$29874 ( \38545 , \38544 );
xor \U$29875 ( \38546 , \38525 , \38545 );
and \U$29876 ( \38547 , \12157 , \36986_nG9b90 );
and \U$29877 ( \38548 , \12154 , \37250_nG9b8d );
or \U$29878 ( \38549 , \38547 , \38548 );
xor \U$29879 ( \38550 , \12153 , \38549 );
buf \U$29880 ( \38551 , \38550 );
buf \U$29882 ( \38552 , \38551 );
xor \U$29883 ( \38553 , \38546 , \38552 );
buf \U$29884 ( \38554 , \38553 );
and \U$29885 ( \38555 , \17297 , \34041_nG9ba8 );
and \U$29886 ( \38556 , \17294 , \34294_nG9ba5 );
or \U$29887 ( \38557 , \38555 , \38556 );
xor \U$29888 ( \38558 , \17293 , \38557 );
buf \U$29889 ( \38559 , \38558 );
buf \U$29891 ( \38560 , \38559 );
and \U$29892 ( \38561 , \13370 , \36172_nG9b96 );
and \U$29893 ( \38562 , \13367 , \36589_nG9b93 );
or \U$29894 ( \38563 , \38561 , \38562 );
xor \U$29895 ( \38564 , \13366 , \38563 );
buf \U$29896 ( \38565 , \38564 );
buf \U$29898 ( \38566 , \38565 );
xor \U$29899 ( \38567 , \38560 , \38566 );
and \U$29900 ( \38568 , \10707 , \38337_nG9b84 );
and \U$29901 ( \38569 , \38296 , \38300 );
and \U$29902 ( \38570 , \38300 , \38325 );
and \U$29903 ( \38571 , \38296 , \38325 );
or \U$29904 ( \38572 , \38569 , \38570 , \38571 );
and \U$29905 ( \38573 , \38248 , \38252 );
and \U$29906 ( \38574 , \38252 , \38257 );
and \U$29907 ( \38575 , \38248 , \38257 );
or \U$29908 ( \38576 , \38573 , \38574 , \38575 );
and \U$29909 ( \38577 , \38263 , \38274 );
and \U$29910 ( \38578 , \38274 , \38289 );
and \U$29911 ( \38579 , \38263 , \38289 );
or \U$29912 ( \38580 , \38577 , \38578 , \38579 );
xor \U$29913 ( \38581 , \38576 , \38580 );
and \U$29914 ( \38582 , \38267 , \38271 );
and \U$29915 ( \38583 , \38271 , \38273 );
and \U$29916 ( \38584 , \38267 , \38273 );
or \U$29917 ( \38585 , \38582 , \38583 , \38584 );
and \U$29918 ( \38586 , \38314 , \38318 );
and \U$29919 ( \38587 , \38318 , \38323 );
and \U$29920 ( \38588 , \38314 , \38323 );
or \U$29921 ( \38589 , \38586 , \38587 , \38588 );
xor \U$29922 ( \38590 , \38585 , \38589 );
and \U$29923 ( \38591 , \30268 , \22542 );
and \U$29924 ( \38592 , \30802 , \22103 );
nor \U$29925 ( \38593 , \38591 , \38592 );
xnor \U$29926 ( \38594 , \38593 , \22548 );
and \U$29927 ( \38595 , \25272 , \27397 );
and \U$29928 ( \38596 , \25815 , \26807 );
nor \U$29929 ( \38597 , \38595 , \38596 );
xnor \U$29930 ( \38598 , \38597 , \27295 );
xor \U$29931 ( \38599 , \38594 , \38598 );
and \U$29932 ( \38600 , \19558 , \32802 );
xor \U$29933 ( \38601 , \38599 , \38600 );
xor \U$29934 ( \38602 , \38590 , \38601 );
xor \U$29935 ( \38603 , \38581 , \38602 );
xor \U$29936 ( \38604 , \38572 , \38603 );
and \U$29937 ( \38605 , \38305 , \38309 );
and \U$29938 ( \38606 , \38309 , \38324 );
and \U$29939 ( \38607 , \38305 , \38324 );
or \U$29940 ( \38608 , \38605 , \38606 , \38607 );
and \U$29941 ( \38609 , \38244 , \38258 );
and \U$29942 ( \38610 , \38258 , \38290 );
and \U$29943 ( \38611 , \38244 , \38290 );
or \U$29944 ( \38612 , \38609 , \38610 , \38611 );
xor \U$29945 ( \38613 , \38608 , \38612 );
not \U$29946 ( \38614 , \19540 );
and \U$29947 ( \38615 , \32054 , \21005 );
and \U$29948 ( \38616 , \32794 , \20557 );
nor \U$29949 ( \38617 , \38615 , \38616 );
xnor \U$29950 ( \38618 , \38617 , \21011 );
xor \U$29951 ( \38619 , \38614 , \38618 );
and \U$29952 ( \38620 , \28534 , \24138 );
and \U$29953 ( \38621 , \29084 , \23630 );
nor \U$29954 ( \38622 , \38620 , \38621 );
xnor \U$29955 ( \38623 , \38622 , \24144 );
xor \U$29956 ( \38624 , \38619 , \38623 );
and \U$29957 ( \38625 , \26829 , \25826 );
and \U$29958 ( \38626 , \27313 , \25264 );
nor \U$29959 ( \38627 , \38625 , \38626 );
xnor \U$29960 ( \38628 , \38627 , \25773 );
and \U$29961 ( \38629 , \22090 , \30823 );
and \U$29962 ( \38630 , \22556 , \30246 );
nor \U$29963 ( \38631 , \38629 , \38630 );
xnor \U$29964 ( \38632 , \38631 , \30813 );
xor \U$29965 ( \38633 , \38628 , \38632 );
and \U$29966 ( \38634 , \20544 , \32854 );
and \U$29967 ( \38635 , \21033 , \32067 );
nor \U$29968 ( \38636 , \38634 , \38635 );
xnor \U$29969 ( \38637 , \38636 , \32805 );
xor \U$29970 ( \38638 , \38633 , \38637 );
xor \U$29971 ( \38639 , \38624 , \38638 );
and \U$29972 ( \38640 , \38279 , \38283 );
and \U$29973 ( \38641 , \38283 , \38288 );
and \U$29974 ( \38642 , \38279 , \38288 );
or \U$29975 ( \38643 , \38640 , \38641 , \38642 );
buf \U$29976 ( \38644 , \38256 );
xor \U$29977 ( \38645 , \38643 , \38644 );
and \U$29978 ( \38646 , \23617 , \29070 );
and \U$29979 ( \38647 , \24199 , \28526 );
nor \U$29980 ( \38648 , \38646 , \38647 );
xnor \U$29981 ( \38649 , \38648 , \29076 );
xor \U$29982 ( \38650 , \38645 , \38649 );
xor \U$29983 ( \38651 , \38639 , \38650 );
xor \U$29984 ( \38652 , \38613 , \38651 );
xor \U$29985 ( \38653 , \38604 , \38652 );
and \U$29986 ( \38654 , \38240 , \38291 );
and \U$29987 ( \38655 , \38291 , \38326 );
and \U$29988 ( \38656 , \38240 , \38326 );
or \U$29989 ( \38657 , \38654 , \38655 , \38656 );
xor \U$29990 ( \38658 , \38653 , \38657 );
and \U$29991 ( \38659 , \38327 , \38331 );
and \U$29992 ( \38660 , \38332 , \38335 );
or \U$29993 ( \38661 , \38659 , \38660 );
xor \U$29994 ( \38662 , \38658 , \38661 );
buf g9b81 ( \38663_nG9b81 , \38662 );
and \U$29995 ( \38664 , \10704 , \38663_nG9b81 );
or \U$29996 ( \38665 , \38568 , \38664 );
xor \U$29997 ( \38666 , \10703 , \38665 );
buf \U$29998 ( \38667 , \38666 );
buf \U$30000 ( \38668 , \38667 );
xor \U$30001 ( \38669 , \38567 , \38668 );
buf \U$30002 ( \38670 , \38669 );
xor \U$30003 ( \38671 , \38554 , \38670 );
and \U$30004 ( \38672 , \38199 , \38205 );
and \U$30005 ( \38673 , \38199 , \38212 );
and \U$30006 ( \38674 , \38205 , \38212 );
or \U$30007 ( \38675 , \38672 , \38673 , \38674 );
buf \U$30008 ( \38676 , \38675 );
and \U$30009 ( \38677 , \28118 , \23696_nG9bd2 );
and \U$30010 ( \38678 , \28115 , \24226_nG9bcf );
or \U$30011 ( \38679 , \38677 , \38678 );
xor \U$30012 ( \38680 , \28114 , \38679 );
buf \U$30013 ( \38681 , \38680 );
buf \U$30015 ( \38682 , \38681 );
and \U$30016 ( \38683 , \26431 , \25298_nG9bcc );
and \U$30017 ( \38684 , \26428 , \25860_nG9bc9 );
or \U$30018 ( \38685 , \38683 , \38684 );
xor \U$30019 ( \38686 , \26427 , \38685 );
buf \U$30020 ( \38687 , \38686 );
buf \U$30022 ( \38688 , \38687 );
xor \U$30023 ( \38689 , \38682 , \38688 );
and \U$30024 ( \38690 , \24792 , \26887_nG9bc6 );
and \U$30025 ( \38691 , \24789 , \27416_nG9bc3 );
or \U$30026 ( \38692 , \38690 , \38691 );
xor \U$30027 ( \38693 , \24788 , \38692 );
buf \U$30028 ( \38694 , \38693 );
buf \U$30030 ( \38695 , \38694 );
xor \U$30031 ( \38696 , \38689 , \38695 );
buf \U$30032 ( \38697 , \38696 );
xor \U$30033 ( \38698 , \38676 , \38697 );
and \U$30034 ( \38699 , \10421 , \37607_nG9b8a );
and \U$30035 ( \38700 , \10418 , \37974_nG9b87 );
or \U$30036 ( \38701 , \38699 , \38700 );
xor \U$30037 ( \38702 , \10417 , \38701 );
buf \U$30038 ( \38703 , \38702 );
buf \U$30040 ( \38704 , \38703 );
xor \U$30041 ( \38705 , \38698 , \38704 );
buf \U$30042 ( \38706 , \38705 );
xor \U$30043 ( \38707 , \38671 , \38706 );
buf \U$30044 ( \38708 , \38707 );
xor \U$30045 ( \38709 , \38520 , \38708 );
buf \U$30046 ( \38710 , \38709 );
xor \U$30047 ( \38711 , \38481 , \38710 );
xor \U$30048 ( \38712 , \38397 , \38711 );
and \U$30049 ( \38713 , \38128 , \38133 );
and \U$30050 ( \38714 , \38128 , \38387 );
and \U$30051 ( \38715 , \38133 , \38387 );
or \U$30052 ( \38716 , \38713 , \38714 , \38715 );
and \U$30053 ( \38717 , \38712 , \38716 );
and \U$30055 ( \38718 , \38396 , \38711 );
or \U$30057 ( \38719 , 1'b0 , \38718 , 1'b0 );
xor \U$30058 ( \38720 , \38717 , \38719 );
and \U$30060 ( \38721 , \38389 , \38395 );
and \U$30061 ( \38722 , \38391 , \38395 );
or \U$30062 ( \38723 , 1'b0 , \38721 , \38722 );
xor \U$30063 ( \38724 , \38720 , \38723 );
xor \U$30070 ( \38725 , \38724 , 1'b0 );
and \U$30071 ( \38726 , \38475 , \38480 );
and \U$30072 ( \38727 , \38475 , \38710 );
and \U$30073 ( \38728 , \38480 , \38710 );
or \U$30074 ( \38729 , \38726 , \38727 , \38728 );
xor \U$30075 ( \38730 , \38725 , \38729 );
and \U$30076 ( \38731 , \38486 , \38519 );
and \U$30077 ( \38732 , \38486 , \38708 );
and \U$30078 ( \38733 , \38519 , \38708 );
or \U$30079 ( \38734 , \38731 , \38732 , \38733 );
buf \U$30080 ( \38735 , \38734 );
and \U$30081 ( \38736 , \38491 , \38496 );
and \U$30082 ( \38737 , \38491 , \38517 );
and \U$30083 ( \38738 , \38496 , \38517 );
or \U$30084 ( \38739 , \38736 , \38737 , \38738 );
buf \U$30085 ( \38740 , \38739 );
and \U$30086 ( \38741 , \38682 , \38688 );
and \U$30087 ( \38742 , \38682 , \38695 );
and \U$30088 ( \38743 , \38688 , \38695 );
or \U$30089 ( \38744 , \38741 , \38742 , \38743 );
buf \U$30090 ( \38745 , \38744 );
and \U$30091 ( \38746 , \15940 , \35094_nG9b9f );
and \U$30092 ( \38747 , \15937 , \35570_nG9b9c );
or \U$30093 ( \38748 , \38746 , \38747 );
xor \U$30094 ( \38749 , \15936 , \38748 );
buf \U$30095 ( \38750 , \38749 );
buf \U$30097 ( \38751 , \38750 );
xor \U$30098 ( \38752 , \38745 , \38751 );
and \U$30099 ( \38753 , \14631 , \35801_nG9b99 );
and \U$30100 ( \38754 , \14628 , \36172_nG9b96 );
or \U$30101 ( \38755 , \38753 , \38754 );
xor \U$30102 ( \38756 , \14627 , \38755 );
buf \U$30103 ( \38757 , \38756 );
buf \U$30105 ( \38758 , \38757 );
xor \U$30106 ( \38759 , \38752 , \38758 );
buf \U$30107 ( \38760 , \38759 );
and \U$30109 ( \38761 , \32916 , \20608_nG9bde );
or \U$30110 ( \38762 , 1'b0 , \38761 );
xor \U$30111 ( \38763 , 1'b0 , \38762 );
buf \U$30112 ( \38764 , \38763 );
buf \U$30114 ( \38765 , \38764 );
and \U$30115 ( \38766 , \31636 , \21086_nG9bdb );
and \U$30116 ( \38767 , \31633 , \22129_nG9bd8 );
or \U$30117 ( \38768 , \38766 , \38767 );
xor \U$30118 ( \38769 , \31632 , \38768 );
buf \U$30119 ( \38770 , \38769 );
buf \U$30121 ( \38771 , \38770 );
xor \U$30122 ( \38772 , \38765 , \38771 );
buf \U$30123 ( \38773 , \38772 );
and \U$30124 ( \38774 , \38413 , \38419 );
buf \U$30125 ( \38775 , \38774 );
xor \U$30126 ( \38776 , \38773 , \38775 );
and \U$30127 ( \38777 , \29853 , \22629_nG9bd5 );
and \U$30128 ( \38778 , \29850 , \23696_nG9bd2 );
or \U$30129 ( \38779 , \38777 , \38778 );
xor \U$30130 ( \38780 , \29849 , \38779 );
buf \U$30131 ( \38781 , \38780 );
buf \U$30133 ( \38782 , \38781 );
xor \U$30134 ( \38783 , \38776 , \38782 );
buf \U$30135 ( \38784 , \38783 );
and \U$30136 ( \38785 , \20155 , \32888_nG9bb1 );
and \U$30137 ( \38786 , \20152 , \33181_nG9bae );
or \U$30138 ( \38787 , \38785 , \38786 );
xor \U$30139 ( \38788 , \20151 , \38787 );
buf \U$30140 ( \38789 , \38788 );
buf \U$30142 ( \38790 , \38789 );
xor \U$30143 ( \38791 , \38784 , \38790 );
and \U$30144 ( \38792 , \18702 , \33613_nG9bab );
and \U$30145 ( \38793 , \18699 , \34041_nG9ba8 );
or \U$30146 ( \38794 , \38792 , \38793 );
xor \U$30147 ( \38795 , \18698 , \38794 );
buf \U$30148 ( \38796 , \38795 );
buf \U$30150 ( \38797 , \38796 );
xor \U$30151 ( \38798 , \38791 , \38797 );
buf \U$30152 ( \38799 , \38798 );
xor \U$30153 ( \38800 , \38760 , \38799 );
and \U$30154 ( \38801 , \38502 , \38508 );
and \U$30155 ( \38802 , \38502 , \38515 );
and \U$30156 ( \38803 , \38508 , \38515 );
or \U$30157 ( \38804 , \38801 , \38802 , \38803 );
buf \U$30158 ( \38805 , \38804 );
xor \U$30159 ( \38806 , \38800 , \38805 );
buf \U$30160 ( \38807 , \38806 );
xor \U$30161 ( \38808 , \38740 , \38807 );
and \U$30162 ( \38809 , \38402 , \38407 );
and \U$30163 ( \38810 , \38402 , \38447 );
and \U$30164 ( \38811 , \38407 , \38447 );
or \U$30165 ( \38812 , \38809 , \38810 , \38811 );
buf \U$30166 ( \38813 , \38812 );
xor \U$30167 ( \38814 , \38808 , \38813 );
buf \U$30168 ( \38815 , \38814 );
xor \U$30169 ( \38816 , \38735 , \38815 );
and \U$30170 ( \38817 , \38449 , \38454 );
and \U$30171 ( \38818 , \38449 , \38460 );
and \U$30172 ( \38819 , \38454 , \38460 );
or \U$30173 ( \38820 , \38817 , \38818 , \38819 );
buf \U$30174 ( \38821 , \38820 );
xor \U$30175 ( \38822 , \38816 , \38821 );
buf \U$30176 ( \38823 , \38822 );
and \U$30177 ( \38824 , \38462 , \38467 );
and \U$30178 ( \38825 , \38462 , \38473 );
and \U$30179 ( \38826 , \38467 , \38473 );
or \U$30180 ( \38827 , \38824 , \38825 , \38826 );
buf \U$30181 ( \38828 , \38827 );
xor \U$30182 ( \38829 , \38823 , \38828 );
and \U$30183 ( \38830 , \38432 , \38438 );
and \U$30184 ( \38831 , \38432 , \38445 );
and \U$30185 ( \38832 , \38438 , \38445 );
or \U$30186 ( \38833 , \38830 , \38831 , \38832 );
buf \U$30187 ( \38834 , \38833 );
and \U$30188 ( \38835 , \38421 , \38423 );
and \U$30189 ( \38836 , \38421 , \38430 );
and \U$30190 ( \38837 , \38423 , \38430 );
or \U$30191 ( \38838 , \38835 , \38836 , \38837 );
buf \U$30192 ( \38839 , \38838 );
and \U$30193 ( \38840 , \23201 , \29179_nG9bbd );
and \U$30194 ( \38841 , \23198 , \30366_nG9bba );
or \U$30195 ( \38842 , \38840 , \38841 );
xor \U$30196 ( \38843 , \23197 , \38842 );
buf \U$30197 ( \38844 , \38843 );
buf \U$30199 ( \38845 , \38844 );
xor \U$30200 ( \38846 , \38839 , \38845 );
and \U$30201 ( \38847 , \21658 , \30940_nG9bb7 );
and \U$30202 ( \38848 , \21655 , \32179_nG9bb4 );
or \U$30203 ( \38849 , \38847 , \38848 );
xor \U$30204 ( \38850 , \21654 , \38849 );
buf \U$30205 ( \38851 , \38850 );
buf \U$30207 ( \38852 , \38851 );
xor \U$30208 ( \38853 , \38846 , \38852 );
buf \U$30209 ( \38854 , \38853 );
xor \U$30210 ( \38855 , \38834 , \38854 );
and \U$30211 ( \38856 , \12157 , \37250_nG9b8d );
and \U$30212 ( \38857 , \12154 , \37607_nG9b8a );
or \U$30213 ( \38858 , \38856 , \38857 );
xor \U$30214 ( \38859 , \12153 , \38858 );
buf \U$30215 ( \38860 , \38859 );
buf \U$30217 ( \38861 , \38860 );
xor \U$30218 ( \38862 , \38855 , \38861 );
buf \U$30219 ( \38863 , \38862 );
and \U$30220 ( \38864 , \17297 , \34294_nG9ba5 );
and \U$30221 ( \38865 , \17294 , \34643_nG9ba2 );
or \U$30222 ( \38866 , \38864 , \38865 );
xor \U$30223 ( \38867 , \17293 , \38866 );
buf \U$30224 ( \38868 , \38867 );
buf \U$30226 ( \38869 , \38868 );
and \U$30227 ( \38870 , \13370 , \36589_nG9b93 );
and \U$30228 ( \38871 , \13367 , \36986_nG9b90 );
or \U$30229 ( \38872 , \38870 , \38871 );
xor \U$30230 ( \38873 , \13366 , \38872 );
buf \U$30231 ( \38874 , \38873 );
buf \U$30233 ( \38875 , \38874 );
xor \U$30234 ( \38876 , \38869 , \38875 );
and \U$30235 ( \38877 , \10707 , \38663_nG9b81 );
and \U$30236 ( \38878 , \38608 , \38612 );
and \U$30237 ( \38879 , \38612 , \38651 );
and \U$30238 ( \38880 , \38608 , \38651 );
or \U$30239 ( \38881 , \38878 , \38879 , \38880 );
and \U$30240 ( \38882 , \38643 , \38644 );
and \U$30241 ( \38883 , \38644 , \38649 );
and \U$30242 ( \38884 , \38643 , \38649 );
or \U$30243 ( \38885 , \38882 , \38883 , \38884 );
and \U$30244 ( \38886 , \38585 , \38589 );
and \U$30245 ( \38887 , \38589 , \38601 );
and \U$30246 ( \38888 , \38585 , \38601 );
or \U$30247 ( \38889 , \38886 , \38887 , \38888 );
xor \U$30248 ( \38890 , \38885 , \38889 );
and \U$30249 ( \38891 , \38594 , \38598 );
and \U$30250 ( \38892 , \38598 , \38600 );
and \U$30251 ( \38893 , \38594 , \38600 );
or \U$30252 ( \38894 , \38891 , \38892 , \38893 );
and \U$30253 ( \38895 , \38614 , \38618 );
and \U$30254 ( \38896 , \38618 , \38623 );
and \U$30255 ( \38897 , \38614 , \38623 );
or \U$30256 ( \38898 , \38895 , \38896 , \38897 );
xor \U$30257 ( \38899 , \38894 , \38898 );
and \U$30258 ( \38900 , \38628 , \38632 );
and \U$30259 ( \38901 , \38632 , \38637 );
and \U$30260 ( \38902 , \38628 , \38637 );
or \U$30261 ( \38903 , \38900 , \38901 , \38902 );
xor \U$30262 ( \38904 , \38899 , \38903 );
xor \U$30263 ( \38905 , \38890 , \38904 );
xor \U$30264 ( \38906 , \38881 , \38905 );
and \U$30265 ( \38907 , \38624 , \38638 );
and \U$30266 ( \38908 , \38638 , \38650 );
and \U$30267 ( \38909 , \38624 , \38650 );
or \U$30268 ( \38910 , \38907 , \38908 , \38909 );
and \U$30269 ( \38911 , \38576 , \38580 );
and \U$30270 ( \38912 , \38580 , \38602 );
and \U$30271 ( \38913 , \38576 , \38602 );
or \U$30272 ( \38914 , \38911 , \38912 , \38913 );
xor \U$30273 ( \38915 , \38910 , \38914 );
and \U$30274 ( \38916 , \30802 , \22542 );
and \U$30275 ( \38917 , \32054 , \22103 );
nor \U$30276 ( \38918 , \38916 , \38917 );
xnor \U$30277 ( \38919 , \38918 , \22548 );
and \U$30278 ( \38920 , \29084 , \24138 );
and \U$30279 ( \38921 , \30268 , \23630 );
nor \U$30280 ( \38922 , \38920 , \38921 );
xnor \U$30281 ( \38923 , \38922 , \24144 );
xor \U$30282 ( \38924 , \38919 , \38923 );
and \U$30283 ( \38925 , \25815 , \27397 );
and \U$30284 ( \38926 , \26829 , \26807 );
nor \U$30285 ( \38927 , \38925 , \38926 );
xnor \U$30286 ( \38928 , \38927 , \27295 );
xor \U$30287 ( \38929 , \38924 , \38928 );
and \U$30288 ( \38930 , \27313 , \25826 );
and \U$30289 ( \38931 , \28534 , \25264 );
nor \U$30290 ( \38932 , \38930 , \38931 );
xnor \U$30291 ( \38933 , \38932 , \25773 );
and \U$30292 ( \38934 , \21033 , \32854 );
and \U$30293 ( \38935 , \22090 , \32067 );
nor \U$30294 ( \38936 , \38934 , \38935 );
xnor \U$30295 ( \38937 , \38936 , \32805 );
xor \U$30296 ( \38938 , \38933 , \38937 );
and \U$30297 ( \38939 , \20544 , \32802 );
xor \U$30298 ( \38940 , \38938 , \38939 );
xor \U$30299 ( \38941 , \38929 , \38940 );
and \U$30300 ( \38942 , \32794 , \21005 );
not \U$30301 ( \38943 , \38942 );
xnor \U$30302 ( \38944 , \38943 , \21011 );
not \U$30303 ( \38945 , \38944 );
and \U$30304 ( \38946 , \24199 , \29070 );
and \U$30305 ( \38947 , \25272 , \28526 );
nor \U$30306 ( \38948 , \38946 , \38947 );
xnor \U$30307 ( \38949 , \38948 , \29076 );
xor \U$30308 ( \38950 , \38945 , \38949 );
and \U$30309 ( \38951 , \22556 , \30823 );
and \U$30310 ( \38952 , \23617 , \30246 );
nor \U$30311 ( \38953 , \38951 , \38952 );
xnor \U$30312 ( \38954 , \38953 , \30813 );
xor \U$30313 ( \38955 , \38950 , \38954 );
xor \U$30314 ( \38956 , \38941 , \38955 );
xor \U$30315 ( \38957 , \38915 , \38956 );
xor \U$30316 ( \38958 , \38906 , \38957 );
and \U$30317 ( \38959 , \38572 , \38603 );
and \U$30318 ( \38960 , \38603 , \38652 );
and \U$30319 ( \38961 , \38572 , \38652 );
or \U$30320 ( \38962 , \38959 , \38960 , \38961 );
xor \U$30321 ( \38963 , \38958 , \38962 );
and \U$30322 ( \38964 , \38653 , \38657 );
and \U$30323 ( \38965 , \38658 , \38661 );
or \U$30324 ( \38966 , \38964 , \38965 );
xor \U$30325 ( \38967 , \38963 , \38966 );
buf g9b7e ( \38968_nG9b7e , \38967 );
and \U$30326 ( \38969 , \10704 , \38968_nG9b7e );
or \U$30327 ( \38970 , \38877 , \38969 );
xor \U$30328 ( \38971 , \10703 , \38970 );
buf \U$30329 ( \38972 , \38971 );
buf \U$30331 ( \38973 , \38972 );
xor \U$30332 ( \38974 , \38876 , \38973 );
buf \U$30333 ( \38975 , \38974 );
xor \U$30334 ( \38976 , \38863 , \38975 );
and \U$30335 ( \38977 , \38530 , \38536 );
and \U$30336 ( \38978 , \38530 , \38543 );
and \U$30337 ( \38979 , \38536 , \38543 );
or \U$30338 ( \38980 , \38977 , \38978 , \38979 );
buf \U$30339 ( \38981 , \38980 );
and \U$30340 ( \38982 , \28118 , \24226_nG9bcf );
and \U$30341 ( \38983 , \28115 , \25298_nG9bcc );
or \U$30342 ( \38984 , \38982 , \38983 );
xor \U$30343 ( \38985 , \28114 , \38984 );
buf \U$30344 ( \38986 , \38985 );
buf \U$30346 ( \38987 , \38986 );
and \U$30347 ( \38988 , \26431 , \25860_nG9bc9 );
and \U$30348 ( \38989 , \26428 , \26887_nG9bc6 );
or \U$30349 ( \38990 , \38988 , \38989 );
xor \U$30350 ( \38991 , \26427 , \38990 );
buf \U$30351 ( \38992 , \38991 );
buf \U$30353 ( \38993 , \38992 );
xor \U$30354 ( \38994 , \38987 , \38993 );
and \U$30355 ( \38995 , \24792 , \27416_nG9bc3 );
and \U$30356 ( \38996 , \24789 , \28602_nG9bc0 );
or \U$30357 ( \38997 , \38995 , \38996 );
xor \U$30358 ( \38998 , \24788 , \38997 );
buf \U$30359 ( \38999 , \38998 );
buf \U$30361 ( \39000 , \38999 );
xor \U$30362 ( \39001 , \38994 , \39000 );
buf \U$30363 ( \39002 , \39001 );
xor \U$30364 ( \39003 , \38981 , \39002 );
and \U$30365 ( \39004 , \10421 , \37974_nG9b87 );
and \U$30366 ( \39005 , \10418 , \38337_nG9b84 );
or \U$30367 ( \39006 , \39004 , \39005 );
xor \U$30368 ( \39007 , \10417 , \39006 );
buf \U$30369 ( \39008 , \39007 );
buf \U$30371 ( \39009 , \39008 );
xor \U$30372 ( \39010 , \39003 , \39009 );
buf \U$30373 ( \39011 , \39010 );
xor \U$30374 ( \39012 , \38976 , \39011 );
buf \U$30375 ( \39013 , \39012 );
and \U$30376 ( \39014 , \38525 , \38545 );
and \U$30377 ( \39015 , \38525 , \38552 );
and \U$30378 ( \39016 , \38545 , \38552 );
or \U$30379 ( \39017 , \39014 , \39015 , \39016 );
buf \U$30380 ( \39018 , \39017 );
and \U$30381 ( \39019 , \38560 , \38566 );
and \U$30382 ( \39020 , \38560 , \38668 );
and \U$30383 ( \39021 , \38566 , \38668 );
or \U$30384 ( \39022 , \39019 , \39020 , \39021 );
buf \U$30385 ( \39023 , \39022 );
xor \U$30386 ( \39024 , \39018 , \39023 );
and \U$30387 ( \39025 , \38676 , \38697 );
and \U$30388 ( \39026 , \38676 , \38704 );
and \U$30389 ( \39027 , \38697 , \38704 );
or \U$30390 ( \39028 , \39025 , \39026 , \39027 );
buf \U$30391 ( \39029 , \39028 );
xor \U$30392 ( \39030 , \39024 , \39029 );
buf \U$30393 ( \39031 , \39030 );
xor \U$30394 ( \39032 , \39013 , \39031 );
and \U$30395 ( \39033 , \38554 , \38670 );
and \U$30396 ( \39034 , \38554 , \38706 );
and \U$30397 ( \39035 , \38670 , \38706 );
or \U$30398 ( \39036 , \39033 , \39034 , \39035 );
buf \U$30399 ( \39037 , \39036 );
xor \U$30400 ( \39038 , \39032 , \39037 );
buf \U$30401 ( \39039 , \39038 );
xor \U$30402 ( \39040 , \38829 , \39039 );
and \U$30403 ( \39041 , \38730 , \39040 );
and \U$30405 ( \39042 , \38724 , \38729 );
or \U$30407 ( \39043 , 1'b0 , \39042 , 1'b0 );
xor \U$30408 ( \39044 , \39041 , \39043 );
and \U$30410 ( \39045 , \38717 , \38723 );
and \U$30411 ( \39046 , \38719 , \38723 );
or \U$30412 ( \39047 , 1'b0 , \39045 , \39046 );
xor \U$30413 ( \39048 , \39044 , \39047 );
xor \U$30420 ( \39049 , \39048 , 1'b0 );
and \U$30421 ( \39050 , \38823 , \38828 );
and \U$30422 ( \39051 , \38823 , \39039 );
and \U$30423 ( \39052 , \38828 , \39039 );
or \U$30424 ( \39053 , \39050 , \39051 , \39052 );
xor \U$30425 ( \39054 , \39049 , \39053 );
and \U$30426 ( \39055 , \38760 , \38799 );
and \U$30427 ( \39056 , \38760 , \38805 );
and \U$30428 ( \39057 , \38799 , \38805 );
or \U$30429 ( \39058 , \39055 , \39056 , \39057 );
buf \U$30430 ( \39059 , \39058 );
and \U$30431 ( \39060 , \38839 , \38845 );
and \U$30432 ( \39061 , \38839 , \38852 );
and \U$30433 ( \39062 , \38845 , \38852 );
or \U$30434 ( \39063 , \39060 , \39061 , \39062 );
buf \U$30435 ( \39064 , \39063 );
and \U$30436 ( \39065 , \38773 , \38775 );
and \U$30437 ( \39066 , \38773 , \38782 );
and \U$30438 ( \39067 , \38775 , \38782 );
or \U$30439 ( \39068 , \39065 , \39066 , \39067 );
buf \U$30440 ( \39069 , \39068 );
and \U$30441 ( \39070 , \28118 , \25298_nG9bcc );
and \U$30442 ( \39071 , \28115 , \25860_nG9bc9 );
or \U$30443 ( \39072 , \39070 , \39071 );
xor \U$30444 ( \39073 , \28114 , \39072 );
buf \U$30445 ( \39074 , \39073 );
buf \U$30447 ( \39075 , \39074 );
xor \U$30448 ( \39076 , \39069 , \39075 );
and \U$30449 ( \39077 , \26431 , \26887_nG9bc6 );
and \U$30450 ( \39078 , \26428 , \27416_nG9bc3 );
or \U$30451 ( \39079 , \39077 , \39078 );
xor \U$30452 ( \39080 , \26427 , \39079 );
buf \U$30453 ( \39081 , \39080 );
buf \U$30455 ( \39082 , \39081 );
xor \U$30456 ( \39083 , \39076 , \39082 );
buf \U$30457 ( \39084 , \39083 );
xor \U$30458 ( \39085 , \39064 , \39084 );
and \U$30459 ( \39086 , \12157 , \37607_nG9b8a );
and \U$30460 ( \39087 , \12154 , \37974_nG9b87 );
or \U$30461 ( \39088 , \39086 , \39087 );
xor \U$30462 ( \39089 , \12153 , \39088 );
buf \U$30463 ( \39090 , \39089 );
buf \U$30465 ( \39091 , \39090 );
xor \U$30466 ( \39092 , \39085 , \39091 );
buf \U$30467 ( \39093 , \39092 );
and \U$30468 ( \39094 , \38981 , \39002 );
and \U$30469 ( \39095 , \38981 , \39009 );
and \U$30470 ( \39096 , \39002 , \39009 );
or \U$30471 ( \39097 , \39094 , \39095 , \39096 );
buf \U$30472 ( \39098 , \39097 );
xor \U$30473 ( \39099 , \39093 , \39098 );
and \U$30474 ( \39100 , \38987 , \38993 );
and \U$30475 ( \39101 , \38987 , \39000 );
and \U$30476 ( \39102 , \38993 , \39000 );
or \U$30477 ( \39103 , \39100 , \39101 , \39102 );
buf \U$30478 ( \39104 , \39103 );
and \U$30479 ( \39105 , \21658 , \32179_nG9bb4 );
and \U$30480 ( \39106 , \21655 , \32888_nG9bb1 );
or \U$30481 ( \39107 , \39105 , \39106 );
xor \U$30482 ( \39108 , \21654 , \39107 );
buf \U$30483 ( \39109 , \39108 );
buf \U$30485 ( \39110 , \39109 );
xor \U$30486 ( \39111 , \39104 , \39110 );
and \U$30487 ( \39112 , \18702 , \34041_nG9ba8 );
and \U$30488 ( \39113 , \18699 , \34294_nG9ba5 );
or \U$30489 ( \39114 , \39112 , \39113 );
xor \U$30490 ( \39115 , \18698 , \39114 );
buf \U$30491 ( \39116 , \39115 );
buf \U$30493 ( \39117 , \39116 );
xor \U$30494 ( \39118 , \39111 , \39117 );
buf \U$30495 ( \39119 , \39118 );
xor \U$30496 ( \39120 , \39099 , \39119 );
buf \U$30497 ( \39121 , \39120 );
xor \U$30498 ( \39122 , \39059 , \39121 );
and \U$30500 ( \39123 , \32916 , \21086_nG9bdb );
or \U$30501 ( \39124 , 1'b0 , \39123 );
xor \U$30502 ( \39125 , 1'b0 , \39124 );
buf \U$30503 ( \39126 , \39125 );
buf \U$30505 ( \39127 , \39126 );
and \U$30506 ( \39128 , \31636 , \22129_nG9bd8 );
and \U$30507 ( \39129 , \31633 , \22629_nG9bd5 );
or \U$30508 ( \39130 , \39128 , \39129 );
xor \U$30509 ( \39131 , \31632 , \39130 );
buf \U$30510 ( \39132 , \39131 );
buf \U$30512 ( \39133 , \39132 );
xor \U$30513 ( \39134 , \39127 , \39133 );
buf \U$30514 ( \39135 , \39134 );
and \U$30515 ( \39136 , \38765 , \38771 );
buf \U$30516 ( \39137 , \39136 );
xor \U$30517 ( \39138 , \39135 , \39137 );
and \U$30518 ( \39139 , \29853 , \23696_nG9bd2 );
and \U$30519 ( \39140 , \29850 , \24226_nG9bcf );
or \U$30520 ( \39141 , \39139 , \39140 );
xor \U$30521 ( \39142 , \29849 , \39141 );
buf \U$30522 ( \39143 , \39142 );
buf \U$30524 ( \39144 , \39143 );
xor \U$30525 ( \39145 , \39138 , \39144 );
buf \U$30526 ( \39146 , \39145 );
and \U$30527 ( \39147 , \17297 , \34643_nG9ba2 );
and \U$30528 ( \39148 , \17294 , \35094_nG9b9f );
or \U$30529 ( \39149 , \39147 , \39148 );
xor \U$30530 ( \39150 , \17293 , \39149 );
buf \U$30531 ( \39151 , \39150 );
buf \U$30533 ( \39152 , \39151 );
xor \U$30534 ( \39153 , \39146 , \39152 );
and \U$30535 ( \39154 , \15940 , \35570_nG9b9c );
and \U$30536 ( \39155 , \15937 , \35801_nG9b99 );
or \U$30537 ( \39156 , \39154 , \39155 );
xor \U$30538 ( \39157 , \15936 , \39156 );
buf \U$30539 ( \39158 , \39157 );
buf \U$30541 ( \39159 , \39158 );
xor \U$30542 ( \39160 , \39153 , \39159 );
buf \U$30543 ( \39161 , \39160 );
and \U$30544 ( \39162 , \38745 , \38751 );
and \U$30545 ( \39163 , \38745 , \38758 );
and \U$30546 ( \39164 , \38751 , \38758 );
or \U$30547 ( \39165 , \39162 , \39163 , \39164 );
buf \U$30548 ( \39166 , \39165 );
xor \U$30549 ( \39167 , \39161 , \39166 );
and \U$30550 ( \39168 , \38869 , \38875 );
and \U$30551 ( \39169 , \38869 , \38973 );
and \U$30552 ( \39170 , \38875 , \38973 );
or \U$30553 ( \39171 , \39168 , \39169 , \39170 );
buf \U$30554 ( \39172 , \39171 );
xor \U$30555 ( \39173 , \39167 , \39172 );
buf \U$30556 ( \39174 , \39173 );
xor \U$30557 ( \39175 , \39122 , \39174 );
buf \U$30558 ( \39176 , \39175 );
and \U$30559 ( \39177 , \39013 , \39031 );
and \U$30560 ( \39178 , \39013 , \39037 );
and \U$30561 ( \39179 , \39031 , \39037 );
or \U$30562 ( \39180 , \39177 , \39178 , \39179 );
buf \U$30563 ( \39181 , \39180 );
xor \U$30564 ( \39182 , \39176 , \39181 );
and \U$30565 ( \39183 , \38740 , \38807 );
and \U$30566 ( \39184 , \38740 , \38813 );
and \U$30567 ( \39185 , \38807 , \38813 );
or \U$30568 ( \39186 , \39183 , \39184 , \39185 );
buf \U$30569 ( \39187 , \39186 );
xor \U$30570 ( \39188 , \39182 , \39187 );
buf \U$30571 ( \39189 , \39188 );
and \U$30572 ( \39190 , \38735 , \38815 );
and \U$30573 ( \39191 , \38735 , \38821 );
and \U$30574 ( \39192 , \38815 , \38821 );
or \U$30575 ( \39193 , \39190 , \39191 , \39192 );
buf \U$30576 ( \39194 , \39193 );
xor \U$30577 ( \39195 , \39189 , \39194 );
and \U$30578 ( \39196 , \38863 , \38975 );
and \U$30579 ( \39197 , \38863 , \39011 );
and \U$30580 ( \39198 , \38975 , \39011 );
or \U$30581 ( \39199 , \39196 , \39197 , \39198 );
buf \U$30582 ( \39200 , \39199 );
and \U$30583 ( \39201 , \14631 , \36172_nG9b96 );
and \U$30584 ( \39202 , \14628 , \36589_nG9b93 );
or \U$30585 ( \39203 , \39201 , \39202 );
xor \U$30586 ( \39204 , \14627 , \39203 );
buf \U$30587 ( \39205 , \39204 );
buf \U$30589 ( \39206 , \39205 );
and \U$30590 ( \39207 , \13370 , \36986_nG9b90 );
and \U$30591 ( \39208 , \13367 , \37250_nG9b8d );
or \U$30592 ( \39209 , \39207 , \39208 );
xor \U$30593 ( \39210 , \13366 , \39209 );
buf \U$30594 ( \39211 , \39210 );
buf \U$30596 ( \39212 , \39211 );
xor \U$30597 ( \39213 , \39206 , \39212 );
and \U$30598 ( \39214 , \10421 , \38337_nG9b84 );
and \U$30599 ( \39215 , \10418 , \38663_nG9b81 );
or \U$30600 ( \39216 , \39214 , \39215 );
xor \U$30601 ( \39217 , \10417 , \39216 );
buf \U$30602 ( \39218 , \39217 );
buf \U$30604 ( \39219 , \39218 );
xor \U$30605 ( \39220 , \39213 , \39219 );
buf \U$30606 ( \39221 , \39220 );
and \U$30607 ( \39222 , \38784 , \38790 );
and \U$30608 ( \39223 , \38784 , \38797 );
and \U$30609 ( \39224 , \38790 , \38797 );
or \U$30610 ( \39225 , \39222 , \39223 , \39224 );
buf \U$30611 ( \39226 , \39225 );
and \U$30612 ( \39227 , \24792 , \28602_nG9bc0 );
and \U$30613 ( \39228 , \24789 , \29179_nG9bbd );
or \U$30614 ( \39229 , \39227 , \39228 );
xor \U$30615 ( \39230 , \24788 , \39229 );
buf \U$30616 ( \39231 , \39230 );
buf \U$30618 ( \39232 , \39231 );
and \U$30619 ( \39233 , \23201 , \30366_nG9bba );
and \U$30620 ( \39234 , \23198 , \30940_nG9bb7 );
or \U$30621 ( \39235 , \39233 , \39234 );
xor \U$30622 ( \39236 , \23197 , \39235 );
buf \U$30623 ( \39237 , \39236 );
buf \U$30625 ( \39238 , \39237 );
xor \U$30626 ( \39239 , \39232 , \39238 );
and \U$30627 ( \39240 , \20155 , \33181_nG9bae );
and \U$30628 ( \39241 , \20152 , \33613_nG9bab );
or \U$30629 ( \39242 , \39240 , \39241 );
xor \U$30630 ( \39243 , \20151 , \39242 );
buf \U$30631 ( \39244 , \39243 );
buf \U$30633 ( \39245 , \39244 );
xor \U$30634 ( \39246 , \39239 , \39245 );
buf \U$30635 ( \39247 , \39246 );
xor \U$30636 ( \39248 , \39226 , \39247 );
and \U$30637 ( \39249 , \10707 , \38968_nG9b7e );
and \U$30638 ( \39250 , \38910 , \38914 );
and \U$30639 ( \39251 , \38914 , \38956 );
and \U$30640 ( \39252 , \38910 , \38956 );
or \U$30641 ( \39253 , \39250 , \39251 , \39252 );
and \U$30642 ( \39254 , \38894 , \38898 );
and \U$30643 ( \39255 , \38898 , \38903 );
and \U$30644 ( \39256 , \38894 , \38903 );
or \U$30645 ( \39257 , \39254 , \39255 , \39256 );
and \U$30646 ( \39258 , \38945 , \38949 );
and \U$30647 ( \39259 , \38949 , \38954 );
and \U$30648 ( \39260 , \38945 , \38954 );
or \U$30649 ( \39261 , \39258 , \39259 , \39260 );
xor \U$30650 ( \39262 , \39257 , \39261 );
and \U$30651 ( \39263 , \38919 , \38923 );
and \U$30652 ( \39264 , \38923 , \38928 );
and \U$30653 ( \39265 , \38919 , \38928 );
or \U$30654 ( \39266 , \39263 , \39264 , \39265 );
and \U$30655 ( \39267 , \38933 , \38937 );
and \U$30656 ( \39268 , \38937 , \38939 );
and \U$30657 ( \39269 , \38933 , \38939 );
or \U$30658 ( \39270 , \39267 , \39268 , \39269 );
xor \U$30659 ( \39271 , \39266 , \39270 );
buf \U$30660 ( \39272 , \38944 );
xor \U$30661 ( \39273 , \39271 , \39272 );
xor \U$30662 ( \39274 , \39262 , \39273 );
xor \U$30663 ( \39275 , \39253 , \39274 );
and \U$30664 ( \39276 , \38929 , \38940 );
and \U$30665 ( \39277 , \38940 , \38955 );
and \U$30666 ( \39278 , \38929 , \38955 );
or \U$30667 ( \39279 , \39276 , \39277 , \39278 );
and \U$30668 ( \39280 , \38885 , \38889 );
and \U$30669 ( \39281 , \38889 , \38904 );
and \U$30670 ( \39282 , \38885 , \38904 );
or \U$30671 ( \39283 , \39280 , \39281 , \39282 );
xor \U$30672 ( \39284 , \39279 , \39283 );
and \U$30673 ( \39285 , \26829 , \27397 );
and \U$30674 ( \39286 , \27313 , \26807 );
nor \U$30675 ( \39287 , \39285 , \39286 );
xnor \U$30676 ( \39288 , \39287 , \27295 );
and \U$30677 ( \39289 , \22090 , \32854 );
and \U$30678 ( \39290 , \22556 , \32067 );
nor \U$30679 ( \39291 , \39289 , \39290 );
xnor \U$30680 ( \39292 , \39291 , \32805 );
xor \U$30681 ( \39293 , \39288 , \39292 );
and \U$30682 ( \39294 , \21033 , \32802 );
xor \U$30683 ( \39295 , \39293 , \39294 );
not \U$30684 ( \39296 , \21011 );
and \U$30685 ( \39297 , \32054 , \22542 );
and \U$30686 ( \39298 , \32794 , \22103 );
nor \U$30687 ( \39299 , \39297 , \39298 );
xnor \U$30688 ( \39300 , \39299 , \22548 );
xor \U$30689 ( \39301 , \39296 , \39300 );
and \U$30690 ( \39302 , \28534 , \25826 );
and \U$30691 ( \39303 , \29084 , \25264 );
nor \U$30692 ( \39304 , \39302 , \39303 );
xnor \U$30693 ( \39305 , \39304 , \25773 );
xor \U$30694 ( \39306 , \39301 , \39305 );
xor \U$30695 ( \39307 , \39295 , \39306 );
and \U$30696 ( \39308 , \30268 , \24138 );
and \U$30697 ( \39309 , \30802 , \23630 );
nor \U$30698 ( \39310 , \39308 , \39309 );
xnor \U$30699 ( \39311 , \39310 , \24144 );
and \U$30700 ( \39312 , \25272 , \29070 );
and \U$30701 ( \39313 , \25815 , \28526 );
nor \U$30702 ( \39314 , \39312 , \39313 );
xnor \U$30703 ( \39315 , \39314 , \29076 );
xor \U$30704 ( \39316 , \39311 , \39315 );
and \U$30705 ( \39317 , \23617 , \30823 );
and \U$30706 ( \39318 , \24199 , \30246 );
nor \U$30707 ( \39319 , \39317 , \39318 );
xnor \U$30708 ( \39320 , \39319 , \30813 );
xor \U$30709 ( \39321 , \39316 , \39320 );
xor \U$30710 ( \39322 , \39307 , \39321 );
xor \U$30711 ( \39323 , \39284 , \39322 );
xor \U$30712 ( \39324 , \39275 , \39323 );
and \U$30713 ( \39325 , \38881 , \38905 );
and \U$30714 ( \39326 , \38905 , \38957 );
and \U$30715 ( \39327 , \38881 , \38957 );
or \U$30716 ( \39328 , \39325 , \39326 , \39327 );
xor \U$30717 ( \39329 , \39324 , \39328 );
and \U$30718 ( \39330 , \38958 , \38962 );
and \U$30719 ( \39331 , \38963 , \38966 );
or \U$30720 ( \39332 , \39330 , \39331 );
xor \U$30721 ( \39333 , \39329 , \39332 );
buf g9b7b ( \39334_nG9b7b , \39333 );
and \U$30722 ( \39335 , \10704 , \39334_nG9b7b );
or \U$30723 ( \39336 , \39249 , \39335 );
xor \U$30724 ( \39337 , \10703 , \39336 );
buf \U$30725 ( \39338 , \39337 );
buf \U$30727 ( \39339 , \39338 );
xor \U$30728 ( \39340 , \39248 , \39339 );
buf \U$30729 ( \39341 , \39340 );
xor \U$30730 ( \39342 , \39221 , \39341 );
and \U$30731 ( \39343 , \38834 , \38854 );
and \U$30732 ( \39344 , \38834 , \38861 );
and \U$30733 ( \39345 , \38854 , \38861 );
or \U$30734 ( \39346 , \39343 , \39344 , \39345 );
buf \U$30735 ( \39347 , \39346 );
xor \U$30736 ( \39348 , \39342 , \39347 );
buf \U$30737 ( \39349 , \39348 );
xor \U$30738 ( \39350 , \39200 , \39349 );
and \U$30739 ( \39351 , \39018 , \39023 );
and \U$30740 ( \39352 , \39018 , \39029 );
and \U$30741 ( \39353 , \39023 , \39029 );
or \U$30742 ( \39354 , \39351 , \39352 , \39353 );
buf \U$30743 ( \39355 , \39354 );
xor \U$30744 ( \39356 , \39350 , \39355 );
buf \U$30745 ( \39357 , \39356 );
xor \U$30746 ( \39358 , \39195 , \39357 );
and \U$30747 ( \39359 , \39054 , \39358 );
and \U$30749 ( \39360 , \39048 , \39053 );
or \U$30751 ( \39361 , 1'b0 , \39360 , 1'b0 );
xor \U$30752 ( \39362 , \39359 , \39361 );
and \U$30754 ( \39363 , \39041 , \39047 );
and \U$30755 ( \39364 , \39043 , \39047 );
or \U$30756 ( \39365 , 1'b0 , \39363 , \39364 );
xor \U$30757 ( \39366 , \39362 , \39365 );
xor \U$30764 ( \39367 , \39366 , 1'b0 );
and \U$30765 ( \39368 , \39189 , \39194 );
and \U$30766 ( \39369 , \39189 , \39357 );
and \U$30767 ( \39370 , \39194 , \39357 );
or \U$30768 ( \39371 , \39368 , \39369 , \39370 );
xor \U$30769 ( \39372 , \39367 , \39371 );
and \U$30770 ( \39373 , \39200 , \39349 );
and \U$30771 ( \39374 , \39200 , \39355 );
and \U$30772 ( \39375 , \39349 , \39355 );
or \U$30773 ( \39376 , \39373 , \39374 , \39375 );
buf \U$30774 ( \39377 , \39376 );
and \U$30775 ( \39378 , \39161 , \39166 );
and \U$30776 ( \39379 , \39161 , \39172 );
and \U$30777 ( \39380 , \39166 , \39172 );
or \U$30778 ( \39381 , \39378 , \39379 , \39380 );
buf \U$30779 ( \39382 , \39381 );
and \U$30780 ( \39383 , \39093 , \39098 );
and \U$30781 ( \39384 , \39093 , \39119 );
and \U$30782 ( \39385 , \39098 , \39119 );
or \U$30783 ( \39386 , \39383 , \39384 , \39385 );
buf \U$30784 ( \39387 , \39386 );
xor \U$30785 ( \39388 , \39382 , \39387 );
and \U$30786 ( \39389 , \39064 , \39084 );
and \U$30787 ( \39390 , \39064 , \39091 );
and \U$30788 ( \39391 , \39084 , \39091 );
or \U$30789 ( \39392 , \39389 , \39390 , \39391 );
buf \U$30790 ( \39393 , \39392 );
and \U$30791 ( \39394 , \39135 , \39137 );
and \U$30792 ( \39395 , \39135 , \39144 );
and \U$30793 ( \39396 , \39137 , \39144 );
or \U$30794 ( \39397 , \39394 , \39395 , \39396 );
buf \U$30795 ( \39398 , \39397 );
and \U$30796 ( \39399 , \18702 , \34294_nG9ba5 );
and \U$30797 ( \39400 , \18699 , \34643_nG9ba2 );
or \U$30798 ( \39401 , \39399 , \39400 );
xor \U$30799 ( \39402 , \18698 , \39401 );
buf \U$30800 ( \39403 , \39402 );
buf \U$30802 ( \39404 , \39403 );
xor \U$30803 ( \39405 , \39398 , \39404 );
and \U$30804 ( \39406 , \15940 , \35801_nG9b99 );
and \U$30805 ( \39407 , \15937 , \36172_nG9b96 );
or \U$30806 ( \39408 , \39406 , \39407 );
xor \U$30807 ( \39409 , \15936 , \39408 );
buf \U$30808 ( \39410 , \39409 );
buf \U$30810 ( \39411 , \39410 );
xor \U$30811 ( \39412 , \39405 , \39411 );
buf \U$30812 ( \39413 , \39412 );
xor \U$30813 ( \39414 , \39393 , \39413 );
and \U$30814 ( \39415 , \23201 , \30940_nG9bb7 );
and \U$30815 ( \39416 , \23198 , \32179_nG9bb4 );
or \U$30816 ( \39417 , \39415 , \39416 );
xor \U$30817 ( \39418 , \23197 , \39417 );
buf \U$30818 ( \39419 , \39418 );
buf \U$30820 ( \39420 , \39419 );
and \U$30821 ( \39421 , \21658 , \32888_nG9bb1 );
and \U$30822 ( \39422 , \21655 , \33181_nG9bae );
or \U$30823 ( \39423 , \39421 , \39422 );
xor \U$30824 ( \39424 , \21654 , \39423 );
buf \U$30825 ( \39425 , \39424 );
buf \U$30827 ( \39426 , \39425 );
xor \U$30828 ( \39427 , \39420 , \39426 );
and \U$30829 ( \39428 , \20155 , \33613_nG9bab );
and \U$30830 ( \39429 , \20152 , \34041_nG9ba8 );
or \U$30831 ( \39430 , \39428 , \39429 );
xor \U$30832 ( \39431 , \20151 , \39430 );
buf \U$30833 ( \39432 , \39431 );
buf \U$30835 ( \39433 , \39432 );
xor \U$30836 ( \39434 , \39427 , \39433 );
buf \U$30837 ( \39435 , \39434 );
xor \U$30838 ( \39436 , \39414 , \39435 );
buf \U$30839 ( \39437 , \39436 );
xor \U$30840 ( \39438 , \39388 , \39437 );
buf \U$30841 ( \39439 , \39438 );
xor \U$30842 ( \39440 , \39377 , \39439 );
and \U$30843 ( \39441 , \39059 , \39121 );
and \U$30844 ( \39442 , \39059 , \39174 );
and \U$30845 ( \39443 , \39121 , \39174 );
or \U$30846 ( \39444 , \39441 , \39442 , \39443 );
buf \U$30847 ( \39445 , \39444 );
xor \U$30848 ( \39446 , \39440 , \39445 );
buf \U$30849 ( \39447 , \39446 );
and \U$30850 ( \39448 , \39176 , \39181 );
and \U$30851 ( \39449 , \39176 , \39187 );
and \U$30852 ( \39450 , \39181 , \39187 );
or \U$30853 ( \39451 , \39448 , \39449 , \39450 );
buf \U$30854 ( \39452 , \39451 );
xor \U$30855 ( \39453 , \39447 , \39452 );
and \U$30856 ( \39454 , \39221 , \39341 );
and \U$30857 ( \39455 , \39221 , \39347 );
and \U$30858 ( \39456 , \39341 , \39347 );
or \U$30859 ( \39457 , \39454 , \39455 , \39456 );
buf \U$30860 ( \39458 , \39457 );
and \U$30861 ( \39459 , \39226 , \39247 );
and \U$30862 ( \39460 , \39226 , \39339 );
and \U$30863 ( \39461 , \39247 , \39339 );
or \U$30864 ( \39462 , \39459 , \39460 , \39461 );
buf \U$30865 ( \39463 , \39462 );
and \U$30866 ( \39464 , \28118 , \25860_nG9bc9 );
and \U$30867 ( \39465 , \28115 , \26887_nG9bc6 );
or \U$30868 ( \39466 , \39464 , \39465 );
xor \U$30869 ( \39467 , \28114 , \39466 );
buf \U$30870 ( \39468 , \39467 );
buf \U$30872 ( \39469 , \39468 );
and \U$30873 ( \39470 , \26431 , \27416_nG9bc3 );
and \U$30874 ( \39471 , \26428 , \28602_nG9bc0 );
or \U$30875 ( \39472 , \39470 , \39471 );
xor \U$30876 ( \39473 , \26427 , \39472 );
buf \U$30877 ( \39474 , \39473 );
buf \U$30879 ( \39475 , \39474 );
xor \U$30880 ( \39476 , \39469 , \39475 );
and \U$30881 ( \39477 , \24792 , \29179_nG9bbd );
and \U$30882 ( \39478 , \24789 , \30366_nG9bba );
or \U$30883 ( \39479 , \39477 , \39478 );
xor \U$30884 ( \39480 , \24788 , \39479 );
buf \U$30885 ( \39481 , \39480 );
buf \U$30887 ( \39482 , \39481 );
xor \U$30888 ( \39483 , \39476 , \39482 );
buf \U$30889 ( \39484 , \39483 );
and \U$30891 ( \39485 , \32916 , \22129_nG9bd8 );
or \U$30892 ( \39486 , 1'b0 , \39485 );
xor \U$30893 ( \39487 , 1'b0 , \39486 );
buf \U$30894 ( \39488 , \39487 );
buf \U$30896 ( \39489 , \39488 );
and \U$30897 ( \39490 , \31636 , \22629_nG9bd5 );
and \U$30898 ( \39491 , \31633 , \23696_nG9bd2 );
or \U$30899 ( \39492 , \39490 , \39491 );
xor \U$30900 ( \39493 , \31632 , \39492 );
buf \U$30901 ( \39494 , \39493 );
buf \U$30903 ( \39495 , \39494 );
xor \U$30904 ( \39496 , \39489 , \39495 );
buf \U$30905 ( \39497 , \39496 );
and \U$30906 ( \39498 , \39127 , \39133 );
buf \U$30907 ( \39499 , \39498 );
xor \U$30908 ( \39500 , \39497 , \39499 );
and \U$30909 ( \39501 , \29853 , \24226_nG9bcf );
and \U$30910 ( \39502 , \29850 , \25298_nG9bcc );
or \U$30911 ( \39503 , \39501 , \39502 );
xor \U$30912 ( \39504 , \29849 , \39503 );
buf \U$30913 ( \39505 , \39504 );
buf \U$30915 ( \39506 , \39505 );
xor \U$30916 ( \39507 , \39500 , \39506 );
buf \U$30917 ( \39508 , \39507 );
xor \U$30918 ( \39509 , \39484 , \39508 );
and \U$30919 ( \39510 , \10707 , \39334_nG9b7b );
and \U$30920 ( \39511 , \39257 , \39261 );
and \U$30921 ( \39512 , \39261 , \39273 );
and \U$30922 ( \39513 , \39257 , \39273 );
or \U$30923 ( \39514 , \39511 , \39512 , \39513 );
and \U$30924 ( \39515 , \39279 , \39283 );
and \U$30925 ( \39516 , \39283 , \39322 );
and \U$30926 ( \39517 , \39279 , \39322 );
or \U$30927 ( \39518 , \39515 , \39516 , \39517 );
xor \U$30928 ( \39519 , \39514 , \39518 );
and \U$30929 ( \39520 , \39295 , \39306 );
and \U$30930 ( \39521 , \39306 , \39321 );
and \U$30931 ( \39522 , \39295 , \39321 );
or \U$30932 ( \39523 , \39520 , \39521 , \39522 );
and \U$30933 ( \39524 , \39288 , \39292 );
and \U$30934 ( \39525 , \39292 , \39294 );
and \U$30935 ( \39526 , \39288 , \39294 );
or \U$30936 ( \39527 , \39524 , \39525 , \39526 );
and \U$30937 ( \39528 , \39311 , \39315 );
and \U$30938 ( \39529 , \39315 , \39320 );
and \U$30939 ( \39530 , \39311 , \39320 );
or \U$30940 ( \39531 , \39528 , \39529 , \39530 );
xor \U$30941 ( \39532 , \39527 , \39531 );
and \U$30942 ( \39533 , \29084 , \25826 );
and \U$30943 ( \39534 , \30268 , \25264 );
nor \U$30944 ( \39535 , \39533 , \39534 );
xnor \U$30945 ( \39536 , \39535 , \25773 );
and \U$30946 ( \39537 , \25815 , \29070 );
and \U$30947 ( \39538 , \26829 , \28526 );
nor \U$30948 ( \39539 , \39537 , \39538 );
xnor \U$30949 ( \39540 , \39539 , \29076 );
xor \U$30950 ( \39541 , \39536 , \39540 );
and \U$30951 ( \39542 , \24199 , \30823 );
and \U$30952 ( \39543 , \25272 , \30246 );
nor \U$30953 ( \39544 , \39542 , \39543 );
xnor \U$30954 ( \39545 , \39544 , \30813 );
xor \U$30955 ( \39546 , \39541 , \39545 );
xor \U$30956 ( \39547 , \39532 , \39546 );
xor \U$30957 ( \39548 , \39523 , \39547 );
and \U$30958 ( \39549 , \39266 , \39270 );
and \U$30959 ( \39550 , \39270 , \39272 );
and \U$30960 ( \39551 , \39266 , \39272 );
or \U$30961 ( \39552 , \39549 , \39550 , \39551 );
and \U$30962 ( \39553 , \30802 , \24138 );
and \U$30963 ( \39554 , \32054 , \23630 );
nor \U$30964 ( \39555 , \39553 , \39554 );
xnor \U$30965 ( \39556 , \39555 , \24144 );
and \U$30966 ( \39557 , \27313 , \27397 );
and \U$30967 ( \39558 , \28534 , \26807 );
nor \U$30968 ( \39559 , \39557 , \39558 );
xnor \U$30969 ( \39560 , \39559 , \27295 );
xor \U$30970 ( \39561 , \39556 , \39560 );
and \U$30971 ( \39562 , \22090 , \32802 );
xor \U$30972 ( \39563 , \39561 , \39562 );
xor \U$30973 ( \39564 , \39552 , \39563 );
and \U$30974 ( \39565 , \39296 , \39300 );
and \U$30975 ( \39566 , \39300 , \39305 );
and \U$30976 ( \39567 , \39296 , \39305 );
or \U$30977 ( \39568 , \39565 , \39566 , \39567 );
and \U$30978 ( \39569 , \32794 , \22542 );
not \U$30979 ( \39570 , \39569 );
xnor \U$30980 ( \39571 , \39570 , \22548 );
not \U$30981 ( \39572 , \39571 );
xor \U$30982 ( \39573 , \39568 , \39572 );
and \U$30983 ( \39574 , \22556 , \32854 );
and \U$30984 ( \39575 , \23617 , \32067 );
nor \U$30985 ( \39576 , \39574 , \39575 );
xnor \U$30986 ( \39577 , \39576 , \32805 );
xor \U$30987 ( \39578 , \39573 , \39577 );
xor \U$30988 ( \39579 , \39564 , \39578 );
xor \U$30989 ( \39580 , \39548 , \39579 );
xor \U$30990 ( \39581 , \39519 , \39580 );
and \U$30991 ( \39582 , \39253 , \39274 );
and \U$30992 ( \39583 , \39274 , \39323 );
and \U$30993 ( \39584 , \39253 , \39323 );
or \U$30994 ( \39585 , \39582 , \39583 , \39584 );
xor \U$30995 ( \39586 , \39581 , \39585 );
and \U$30996 ( \39587 , \39324 , \39328 );
and \U$30997 ( \39588 , \39329 , \39332 );
or \U$30998 ( \39589 , \39587 , \39588 );
xor \U$30999 ( \39590 , \39586 , \39589 );
buf g9b78 ( \39591_nG9b78 , \39590 );
and \U$31000 ( \39592 , \10704 , \39591_nG9b78 );
or \U$31001 ( \39593 , \39510 , \39592 );
xor \U$31002 ( \39594 , \10703 , \39593 );
buf \U$31003 ( \39595 , \39594 );
buf \U$31005 ( \39596 , \39595 );
xor \U$31006 ( \39597 , \39509 , \39596 );
buf \U$31007 ( \39598 , \39597 );
xor \U$31008 ( \39599 , \39463 , \39598 );
and \U$31009 ( \39600 , \39206 , \39212 );
and \U$31010 ( \39601 , \39206 , \39219 );
and \U$31011 ( \39602 , \39212 , \39219 );
or \U$31012 ( \39603 , \39600 , \39601 , \39602 );
buf \U$31013 ( \39604 , \39603 );
xor \U$31014 ( \39605 , \39599 , \39604 );
buf \U$31015 ( \39606 , \39605 );
xor \U$31016 ( \39607 , \39458 , \39606 );
and \U$31017 ( \39608 , \39146 , \39152 );
and \U$31018 ( \39609 , \39146 , \39159 );
and \U$31019 ( \39610 , \39152 , \39159 );
or \U$31020 ( \39611 , \39608 , \39609 , \39610 );
buf \U$31021 ( \39612 , \39611 );
and \U$31022 ( \39613 , \39104 , \39110 );
and \U$31023 ( \39614 , \39104 , \39117 );
and \U$31024 ( \39615 , \39110 , \39117 );
or \U$31025 ( \39616 , \39613 , \39614 , \39615 );
buf \U$31026 ( \39617 , \39616 );
xor \U$31027 ( \39618 , \39612 , \39617 );
and \U$31028 ( \39619 , \39232 , \39238 );
and \U$31029 ( \39620 , \39232 , \39245 );
and \U$31030 ( \39621 , \39238 , \39245 );
or \U$31031 ( \39622 , \39619 , \39620 , \39621 );
buf \U$31032 ( \39623 , \39622 );
xor \U$31033 ( \39624 , \39618 , \39623 );
buf \U$31034 ( \39625 , \39624 );
and \U$31035 ( \39626 , \17297 , \35094_nG9b9f );
and \U$31036 ( \39627 , \17294 , \35570_nG9b9c );
or \U$31037 ( \39628 , \39626 , \39627 );
xor \U$31038 ( \39629 , \17293 , \39628 );
buf \U$31039 ( \39630 , \39629 );
buf \U$31041 ( \39631 , \39630 );
and \U$31042 ( \39632 , \13370 , \37250_nG9b8d );
and \U$31043 ( \39633 , \13367 , \37607_nG9b8a );
or \U$31044 ( \39634 , \39632 , \39633 );
xor \U$31045 ( \39635 , \13366 , \39634 );
buf \U$31046 ( \39636 , \39635 );
buf \U$31048 ( \39637 , \39636 );
xor \U$31049 ( \39638 , \39631 , \39637 );
and \U$31050 ( \39639 , \10421 , \38663_nG9b81 );
and \U$31051 ( \39640 , \10418 , \38968_nG9b7e );
or \U$31052 ( \39641 , \39639 , \39640 );
xor \U$31053 ( \39642 , \10417 , \39641 );
buf \U$31054 ( \39643 , \39642 );
buf \U$31056 ( \39644 , \39643 );
xor \U$31057 ( \39645 , \39638 , \39644 );
buf \U$31058 ( \39646 , \39645 );
xor \U$31059 ( \39647 , \39625 , \39646 );
and \U$31060 ( \39648 , \39069 , \39075 );
and \U$31061 ( \39649 , \39069 , \39082 );
and \U$31062 ( \39650 , \39075 , \39082 );
or \U$31063 ( \39651 , \39648 , \39649 , \39650 );
buf \U$31064 ( \39652 , \39651 );
and \U$31065 ( \39653 , \14631 , \36589_nG9b93 );
and \U$31066 ( \39654 , \14628 , \36986_nG9b90 );
or \U$31067 ( \39655 , \39653 , \39654 );
xor \U$31068 ( \39656 , \14627 , \39655 );
buf \U$31069 ( \39657 , \39656 );
buf \U$31071 ( \39658 , \39657 );
xor \U$31072 ( \39659 , \39652 , \39658 );
and \U$31073 ( \39660 , \12157 , \37974_nG9b87 );
and \U$31074 ( \39661 , \12154 , \38337_nG9b84 );
or \U$31075 ( \39662 , \39660 , \39661 );
xor \U$31076 ( \39663 , \12153 , \39662 );
buf \U$31077 ( \39664 , \39663 );
buf \U$31079 ( \39665 , \39664 );
xor \U$31080 ( \39666 , \39659 , \39665 );
buf \U$31081 ( \39667 , \39666 );
xor \U$31082 ( \39668 , \39647 , \39667 );
buf \U$31083 ( \39669 , \39668 );
xor \U$31084 ( \39670 , \39607 , \39669 );
buf \U$31085 ( \39671 , \39670 );
xor \U$31086 ( \39672 , \39453 , \39671 );
and \U$31087 ( \39673 , \39372 , \39672 );
and \U$31089 ( \39674 , \39366 , \39371 );
or \U$31091 ( \39675 , 1'b0 , \39674 , 1'b0 );
xor \U$31092 ( \39676 , \39673 , \39675 );
and \U$31094 ( \39677 , \39359 , \39365 );
and \U$31095 ( \39678 , \39361 , \39365 );
or \U$31096 ( \39679 , 1'b0 , \39677 , \39678 );
xor \U$31097 ( \39680 , \39676 , \39679 );
xor \U$31104 ( \39681 , \39680 , 1'b0 );
and \U$31105 ( \39682 , \39458 , \39606 );
and \U$31106 ( \39683 , \39458 , \39669 );
and \U$31107 ( \39684 , \39606 , \39669 );
or \U$31108 ( \39685 , \39682 , \39683 , \39684 );
buf \U$31109 ( \39686 , \39685 );
and \U$31110 ( \39687 , \39463 , \39598 );
and \U$31111 ( \39688 , \39463 , \39604 );
and \U$31112 ( \39689 , \39598 , \39604 );
or \U$31113 ( \39690 , \39687 , \39688 , \39689 );
buf \U$31114 ( \39691 , \39690 );
and \U$31115 ( \39692 , \39484 , \39508 );
and \U$31116 ( \39693 , \39484 , \39596 );
and \U$31117 ( \39694 , \39508 , \39596 );
or \U$31118 ( \39695 , \39692 , \39693 , \39694 );
buf \U$31119 ( \39696 , \39695 );
and \U$31120 ( \39697 , \39631 , \39637 );
and \U$31121 ( \39698 , \39631 , \39644 );
and \U$31122 ( \39699 , \39637 , \39644 );
or \U$31123 ( \39700 , \39697 , \39698 , \39699 );
buf \U$31124 ( \39701 , \39700 );
xor \U$31125 ( \39702 , \39696 , \39701 );
and \U$31126 ( \39703 , \39652 , \39658 );
and \U$31127 ( \39704 , \39652 , \39665 );
and \U$31128 ( \39705 , \39658 , \39665 );
or \U$31129 ( \39706 , \39703 , \39704 , \39705 );
buf \U$31130 ( \39707 , \39706 );
xor \U$31131 ( \39708 , \39702 , \39707 );
buf \U$31132 ( \39709 , \39708 );
xor \U$31133 ( \39710 , \39691 , \39709 );
and \U$31134 ( \39711 , \39393 , \39413 );
and \U$31135 ( \39712 , \39393 , \39435 );
and \U$31136 ( \39713 , \39413 , \39435 );
or \U$31137 ( \39714 , \39711 , \39712 , \39713 );
buf \U$31138 ( \39715 , \39714 );
xor \U$31139 ( \39716 , \39710 , \39715 );
buf \U$31140 ( \39717 , \39716 );
xor \U$31141 ( \39718 , \39686 , \39717 );
and \U$31142 ( \39719 , \39382 , \39387 );
and \U$31143 ( \39720 , \39382 , \39437 );
and \U$31144 ( \39721 , \39387 , \39437 );
or \U$31145 ( \39722 , \39719 , \39720 , \39721 );
buf \U$31146 ( \39723 , \39722 );
xor \U$31147 ( \39724 , \39718 , \39723 );
buf \U$31148 ( \39725 , \39724 );
and \U$31149 ( \39726 , \39377 , \39439 );
and \U$31150 ( \39727 , \39377 , \39445 );
and \U$31151 ( \39728 , \39439 , \39445 );
or \U$31152 ( \39729 , \39726 , \39727 , \39728 );
buf \U$31153 ( \39730 , \39729 );
xor \U$31154 ( \39731 , \39725 , \39730 );
and \U$31155 ( \39732 , \39625 , \39646 );
and \U$31156 ( \39733 , \39625 , \39667 );
and \U$31157 ( \39734 , \39646 , \39667 );
or \U$31158 ( \39735 , \39732 , \39733 , \39734 );
buf \U$31159 ( \39736 , \39735 );
and \U$31160 ( \39737 , \39489 , \39495 );
buf \U$31161 ( \39738 , \39737 );
and \U$31162 ( \39739 , \29853 , \25298_nG9bcc );
and \U$31163 ( \39740 , \29850 , \25860_nG9bc9 );
or \U$31164 ( \39741 , \39739 , \39740 );
xor \U$31165 ( \39742 , \29849 , \39741 );
buf \U$31166 ( \39743 , \39742 );
buf \U$31168 ( \39744 , \39743 );
xor \U$31169 ( \39745 , \39738 , \39744 );
and \U$31170 ( \39746 , \28118 , \26887_nG9bc6 );
and \U$31171 ( \39747 , \28115 , \27416_nG9bc3 );
or \U$31172 ( \39748 , \39746 , \39747 );
xor \U$31173 ( \39749 , \28114 , \39748 );
buf \U$31174 ( \39750 , \39749 );
buf \U$31176 ( \39751 , \39750 );
xor \U$31177 ( \39752 , \39745 , \39751 );
buf \U$31178 ( \39753 , \39752 );
and \U$31179 ( \39754 , \39420 , \39426 );
and \U$31180 ( \39755 , \39420 , \39433 );
and \U$31181 ( \39756 , \39426 , \39433 );
or \U$31182 ( \39757 , \39754 , \39755 , \39756 );
buf \U$31183 ( \39758 , \39757 );
xor \U$31184 ( \39759 , \39753 , \39758 );
and \U$31185 ( \39760 , \12157 , \38337_nG9b84 );
and \U$31186 ( \39761 , \12154 , \38663_nG9b81 );
or \U$31187 ( \39762 , \39760 , \39761 );
xor \U$31188 ( \39763 , \12153 , \39762 );
buf \U$31189 ( \39764 , \39763 );
buf \U$31191 ( \39765 , \39764 );
xor \U$31192 ( \39766 , \39759 , \39765 );
buf \U$31193 ( \39767 , \39766 );
and \U$31194 ( \39768 , \14631 , \36986_nG9b90 );
and \U$31195 ( \39769 , \14628 , \37250_nG9b8d );
or \U$31196 ( \39770 , \39768 , \39769 );
xor \U$31197 ( \39771 , \14627 , \39770 );
buf \U$31198 ( \39772 , \39771 );
buf \U$31200 ( \39773 , \39772 );
and \U$31201 ( \39774 , \13370 , \37607_nG9b8a );
and \U$31202 ( \39775 , \13367 , \37974_nG9b87 );
or \U$31203 ( \39776 , \39774 , \39775 );
xor \U$31204 ( \39777 , \13366 , \39776 );
buf \U$31205 ( \39778 , \39777 );
buf \U$31207 ( \39779 , \39778 );
xor \U$31208 ( \39780 , \39773 , \39779 );
and \U$31209 ( \39781 , \10421 , \38968_nG9b7e );
and \U$31210 ( \39782 , \10418 , \39334_nG9b7b );
or \U$31211 ( \39783 , \39781 , \39782 );
xor \U$31212 ( \39784 , \10417 , \39783 );
buf \U$31213 ( \39785 , \39784 );
buf \U$31215 ( \39786 , \39785 );
xor \U$31216 ( \39787 , \39780 , \39786 );
buf \U$31217 ( \39788 , \39787 );
xor \U$31218 ( \39789 , \39767 , \39788 );
and \U$31219 ( \39790 , \39497 , \39499 );
and \U$31220 ( \39791 , \39497 , \39506 );
and \U$31221 ( \39792 , \39499 , \39506 );
or \U$31222 ( \39793 , \39790 , \39791 , \39792 );
buf \U$31223 ( \39794 , \39793 );
and \U$31224 ( \39795 , \18702 , \34643_nG9ba2 );
and \U$31225 ( \39796 , \18699 , \35094_nG9b9f );
or \U$31226 ( \39797 , \39795 , \39796 );
xor \U$31227 ( \39798 , \18698 , \39797 );
buf \U$31228 ( \39799 , \39798 );
buf \U$31230 ( \39800 , \39799 );
xor \U$31231 ( \39801 , \39794 , \39800 );
and \U$31232 ( \39802 , \17297 , \35570_nG9b9c );
and \U$31233 ( \39803 , \17294 , \35801_nG9b99 );
or \U$31234 ( \39804 , \39802 , \39803 );
xor \U$31235 ( \39805 , \17293 , \39804 );
buf \U$31236 ( \39806 , \39805 );
buf \U$31238 ( \39807 , \39806 );
xor \U$31239 ( \39808 , \39801 , \39807 );
buf \U$31240 ( \39809 , \39808 );
xor \U$31241 ( \39810 , \39789 , \39809 );
buf \U$31242 ( \39811 , \39810 );
xor \U$31243 ( \39812 , \39736 , \39811 );
and \U$31244 ( \39813 , \39398 , \39404 );
and \U$31245 ( \39814 , \39398 , \39411 );
and \U$31246 ( \39815 , \39404 , \39411 );
or \U$31247 ( \39816 , \39813 , \39814 , \39815 );
buf \U$31248 ( \39817 , \39816 );
and \U$31249 ( \39818 , \23201 , \32179_nG9bb4 );
and \U$31250 ( \39819 , \23198 , \32888_nG9bb1 );
or \U$31251 ( \39820 , \39818 , \39819 );
xor \U$31252 ( \39821 , \23197 , \39820 );
buf \U$31253 ( \39822 , \39821 );
buf \U$31255 ( \39823 , \39822 );
and \U$31256 ( \39824 , \21658 , \33181_nG9bae );
and \U$31257 ( \39825 , \21655 , \33613_nG9bab );
or \U$31258 ( \39826 , \39824 , \39825 );
xor \U$31259 ( \39827 , \21654 , \39826 );
buf \U$31260 ( \39828 , \39827 );
buf \U$31262 ( \39829 , \39828 );
xor \U$31263 ( \39830 , \39823 , \39829 );
and \U$31264 ( \39831 , \20155 , \34041_nG9ba8 );
and \U$31265 ( \39832 , \20152 , \34294_nG9ba5 );
or \U$31266 ( \39833 , \39831 , \39832 );
xor \U$31267 ( \39834 , \20151 , \39833 );
buf \U$31268 ( \39835 , \39834 );
buf \U$31270 ( \39836 , \39835 );
xor \U$31271 ( \39837 , \39830 , \39836 );
buf \U$31272 ( \39838 , \39837 );
xor \U$31273 ( \39839 , \39817 , \39838 );
and \U$31275 ( \39840 , \32916 , \22629_nG9bd5 );
or \U$31276 ( \39841 , 1'b0 , \39840 );
xor \U$31277 ( \39842 , 1'b0 , \39841 );
buf \U$31278 ( \39843 , \39842 );
buf \U$31280 ( \39844 , \39843 );
and \U$31281 ( \39845 , \31636 , \23696_nG9bd2 );
and \U$31282 ( \39846 , \31633 , \24226_nG9bcf );
or \U$31283 ( \39847 , \39845 , \39846 );
xor \U$31284 ( \39848 , \31632 , \39847 );
buf \U$31285 ( \39849 , \39848 );
buf \U$31287 ( \39850 , \39849 );
xor \U$31288 ( \39851 , \39844 , \39850 );
buf \U$31289 ( \39852 , \39851 );
and \U$31290 ( \39853 , \26431 , \28602_nG9bc0 );
and \U$31291 ( \39854 , \26428 , \29179_nG9bbd );
or \U$31292 ( \39855 , \39853 , \39854 );
xor \U$31293 ( \39856 , \26427 , \39855 );
buf \U$31294 ( \39857 , \39856 );
buf \U$31296 ( \39858 , \39857 );
xor \U$31297 ( \39859 , \39852 , \39858 );
and \U$31298 ( \39860 , \24792 , \30366_nG9bba );
and \U$31299 ( \39861 , \24789 , \30940_nG9bb7 );
or \U$31300 ( \39862 , \39860 , \39861 );
xor \U$31301 ( \39863 , \24788 , \39862 );
buf \U$31302 ( \39864 , \39863 );
buf \U$31304 ( \39865 , \39864 );
xor \U$31305 ( \39866 , \39859 , \39865 );
buf \U$31306 ( \39867 , \39866 );
xor \U$31307 ( \39868 , \39839 , \39867 );
buf \U$31308 ( \39869 , \39868 );
and \U$31309 ( \39870 , \39612 , \39617 );
and \U$31310 ( \39871 , \39612 , \39623 );
and \U$31311 ( \39872 , \39617 , \39623 );
or \U$31312 ( \39873 , \39870 , \39871 , \39872 );
buf \U$31313 ( \39874 , \39873 );
xor \U$31314 ( \39875 , \39869 , \39874 );
and \U$31315 ( \39876 , \39469 , \39475 );
and \U$31316 ( \39877 , \39469 , \39482 );
and \U$31317 ( \39878 , \39475 , \39482 );
or \U$31318 ( \39879 , \39876 , \39877 , \39878 );
buf \U$31319 ( \39880 , \39879 );
and \U$31320 ( \39881 , \15940 , \36172_nG9b96 );
and \U$31321 ( \39882 , \15937 , \36589_nG9b93 );
or \U$31322 ( \39883 , \39881 , \39882 );
xor \U$31323 ( \39884 , \15936 , \39883 );
buf \U$31324 ( \39885 , \39884 );
buf \U$31326 ( \39886 , \39885 );
xor \U$31327 ( \39887 , \39880 , \39886 );
and \U$31328 ( \39888 , \10707 , \39591_nG9b78 );
and \U$31329 ( \39889 , \39523 , \39547 );
and \U$31330 ( \39890 , \39547 , \39579 );
and \U$31331 ( \39891 , \39523 , \39579 );
or \U$31332 ( \39892 , \39889 , \39890 , \39891 );
and \U$31333 ( \39893 , \39568 , \39572 );
and \U$31334 ( \39894 , \39572 , \39577 );
and \U$31335 ( \39895 , \39568 , \39577 );
or \U$31336 ( \39896 , \39893 , \39894 , \39895 );
and \U$31337 ( \39897 , \30268 , \25826 );
and \U$31338 ( \39898 , \30802 , \25264 );
nor \U$31339 ( \39899 , \39897 , \39898 );
xnor \U$31340 ( \39900 , \39899 , \25773 );
and \U$31341 ( \39901 , \26829 , \29070 );
and \U$31342 ( \39902 , \27313 , \28526 );
nor \U$31343 ( \39903 , \39901 , \39902 );
xnor \U$31344 ( \39904 , \39903 , \29076 );
xor \U$31345 ( \39905 , \39900 , \39904 );
and \U$31346 ( \39906 , \22556 , \32802 );
xor \U$31347 ( \39907 , \39905 , \39906 );
xor \U$31348 ( \39908 , \39896 , \39907 );
buf \U$31349 ( \39909 , \39571 );
and \U$31350 ( \39910 , \25272 , \30823 );
and \U$31351 ( \39911 , \25815 , \30246 );
nor \U$31352 ( \39912 , \39910 , \39911 );
xnor \U$31353 ( \39913 , \39912 , \30813 );
xor \U$31354 ( \39914 , \39909 , \39913 );
and \U$31355 ( \39915 , \23617 , \32854 );
and \U$31356 ( \39916 , \24199 , \32067 );
nor \U$31357 ( \39917 , \39915 , \39916 );
xnor \U$31358 ( \39918 , \39917 , \32805 );
xor \U$31359 ( \39919 , \39914 , \39918 );
xor \U$31360 ( \39920 , \39908 , \39919 );
xor \U$31361 ( \39921 , \39892 , \39920 );
and \U$31362 ( \39922 , \39527 , \39531 );
and \U$31363 ( \39923 , \39531 , \39546 );
and \U$31364 ( \39924 , \39527 , \39546 );
or \U$31365 ( \39925 , \39922 , \39923 , \39924 );
and \U$31366 ( \39926 , \39552 , \39563 );
and \U$31367 ( \39927 , \39563 , \39578 );
and \U$31368 ( \39928 , \39552 , \39578 );
or \U$31369 ( \39929 , \39926 , \39927 , \39928 );
xor \U$31370 ( \39930 , \39925 , \39929 );
and \U$31371 ( \39931 , \39536 , \39540 );
and \U$31372 ( \39932 , \39540 , \39545 );
and \U$31373 ( \39933 , \39536 , \39545 );
or \U$31374 ( \39934 , \39931 , \39932 , \39933 );
and \U$31375 ( \39935 , \39556 , \39560 );
and \U$31376 ( \39936 , \39560 , \39562 );
and \U$31377 ( \39937 , \39556 , \39562 );
or \U$31378 ( \39938 , \39935 , \39936 , \39937 );
xor \U$31379 ( \39939 , \39934 , \39938 );
not \U$31380 ( \39940 , \22548 );
and \U$31381 ( \39941 , \32054 , \24138 );
and \U$31382 ( \39942 , \32794 , \23630 );
nor \U$31383 ( \39943 , \39941 , \39942 );
xnor \U$31384 ( \39944 , \39943 , \24144 );
xor \U$31385 ( \39945 , \39940 , \39944 );
and \U$31386 ( \39946 , \28534 , \27397 );
and \U$31387 ( \39947 , \29084 , \26807 );
nor \U$31388 ( \39948 , \39946 , \39947 );
xnor \U$31389 ( \39949 , \39948 , \27295 );
xor \U$31390 ( \39950 , \39945 , \39949 );
xor \U$31391 ( \39951 , \39939 , \39950 );
xor \U$31392 ( \39952 , \39930 , \39951 );
xor \U$31393 ( \39953 , \39921 , \39952 );
and \U$31394 ( \39954 , \39514 , \39518 );
and \U$31395 ( \39955 , \39518 , \39580 );
and \U$31396 ( \39956 , \39514 , \39580 );
or \U$31397 ( \39957 , \39954 , \39955 , \39956 );
xor \U$31398 ( \39958 , \39953 , \39957 );
and \U$31399 ( \39959 , \39581 , \39585 );
and \U$31400 ( \39960 , \39586 , \39589 );
or \U$31401 ( \39961 , \39959 , \39960 );
xor \U$31402 ( \39962 , \39958 , \39961 );
buf g9b75 ( \39963_nG9b75 , \39962 );
and \U$31403 ( \39964 , \10704 , \39963_nG9b75 );
or \U$31404 ( \39965 , \39888 , \39964 );
xor \U$31405 ( \39966 , \10703 , \39965 );
buf \U$31406 ( \39967 , \39966 );
buf \U$31408 ( \39968 , \39967 );
xor \U$31409 ( \39969 , \39887 , \39968 );
buf \U$31410 ( \39970 , \39969 );
xor \U$31411 ( \39971 , \39875 , \39970 );
buf \U$31412 ( \39972 , \39971 );
xor \U$31413 ( \39973 , \39812 , \39972 );
buf \U$31414 ( \39974 , \39973 );
xor \U$31415 ( \39975 , \39731 , \39974 );
xor \U$31416 ( \39976 , \39681 , \39975 );
and \U$31417 ( \39977 , \39447 , \39452 );
and \U$31418 ( \39978 , \39447 , \39671 );
and \U$31419 ( \39979 , \39452 , \39671 );
or \U$31420 ( \39980 , \39977 , \39978 , \39979 );
and \U$31421 ( \39981 , \39976 , \39980 );
and \U$31423 ( \39982 , \39680 , \39975 );
or \U$31425 ( \39983 , 1'b0 , \39982 , 1'b0 );
xor \U$31426 ( \39984 , \39981 , \39983 );
and \U$31428 ( \39985 , \39673 , \39679 );
and \U$31429 ( \39986 , \39675 , \39679 );
or \U$31430 ( \39987 , 1'b0 , \39985 , \39986 );
xor \U$31431 ( \39988 , \39984 , \39987 );
xor \U$31438 ( \39989 , \39988 , 1'b0 );
and \U$31439 ( \39990 , \39725 , \39730 );
and \U$31440 ( \39991 , \39725 , \39974 );
and \U$31441 ( \39992 , \39730 , \39974 );
or \U$31442 ( \39993 , \39990 , \39991 , \39992 );
xor \U$31443 ( \39994 , \39989 , \39993 );
and \U$31444 ( \39995 , \39736 , \39811 );
and \U$31445 ( \39996 , \39736 , \39972 );
and \U$31446 ( \39997 , \39811 , \39972 );
or \U$31447 ( \39998 , \39995 , \39996 , \39997 );
buf \U$31448 ( \39999 , \39998 );
and \U$31449 ( \40000 , \39691 , \39709 );
and \U$31450 ( \40001 , \39691 , \39715 );
and \U$31451 ( \40002 , \39709 , \39715 );
or \U$31452 ( \40003 , \40000 , \40001 , \40002 );
buf \U$31453 ( \40004 , \40003 );
xor \U$31454 ( \40005 , \39999 , \40004 );
and \U$31455 ( \40006 , \39696 , \39701 );
and \U$31456 ( \40007 , \39696 , \39707 );
and \U$31457 ( \40008 , \39701 , \39707 );
or \U$31458 ( \40009 , \40006 , \40007 , \40008 );
buf \U$31459 ( \40010 , \40009 );
and \U$31460 ( \40011 , \39767 , \39788 );
and \U$31461 ( \40012 , \39767 , \39809 );
and \U$31462 ( \40013 , \39788 , \39809 );
or \U$31463 ( \40014 , \40011 , \40012 , \40013 );
buf \U$31464 ( \40015 , \40014 );
xor \U$31465 ( \40016 , \40010 , \40015 );
and \U$31466 ( \40017 , \39880 , \39886 );
and \U$31467 ( \40018 , \39880 , \39968 );
and \U$31468 ( \40019 , \39886 , \39968 );
or \U$31469 ( \40020 , \40017 , \40018 , \40019 );
buf \U$31470 ( \40021 , \40020 );
and \U$31471 ( \40022 , \39773 , \39779 );
and \U$31472 ( \40023 , \39773 , \39786 );
and \U$31473 ( \40024 , \39779 , \39786 );
or \U$31474 ( \40025 , \40022 , \40023 , \40024 );
buf \U$31475 ( \40026 , \40025 );
xor \U$31476 ( \40027 , \40021 , \40026 );
and \U$31477 ( \40028 , \39738 , \39744 );
and \U$31478 ( \40029 , \39738 , \39751 );
and \U$31479 ( \40030 , \39744 , \39751 );
or \U$31480 ( \40031 , \40028 , \40029 , \40030 );
buf \U$31481 ( \40032 , \40031 );
and \U$31482 ( \40033 , \18702 , \35094_nG9b9f );
and \U$31483 ( \40034 , \18699 , \35570_nG9b9c );
or \U$31484 ( \40035 , \40033 , \40034 );
xor \U$31485 ( \40036 , \18698 , \40035 );
buf \U$31486 ( \40037 , \40036 );
buf \U$31488 ( \40038 , \40037 );
xor \U$31489 ( \40039 , \40032 , \40038 );
and \U$31490 ( \40040 , \17297 , \35801_nG9b99 );
and \U$31491 ( \40041 , \17294 , \36172_nG9b96 );
or \U$31492 ( \40042 , \40040 , \40041 );
xor \U$31493 ( \40043 , \17293 , \40042 );
buf \U$31494 ( \40044 , \40043 );
buf \U$31496 ( \40045 , \40044 );
xor \U$31497 ( \40046 , \40039 , \40045 );
buf \U$31498 ( \40047 , \40046 );
xor \U$31499 ( \40048 , \40027 , \40047 );
buf \U$31500 ( \40049 , \40048 );
xor \U$31501 ( \40050 , \40016 , \40049 );
buf \U$31502 ( \40051 , \40050 );
xor \U$31503 ( \40052 , \40005 , \40051 );
buf \U$31504 ( \40053 , \40052 );
and \U$31505 ( \40054 , \39686 , \39717 );
and \U$31506 ( \40055 , \39686 , \39723 );
and \U$31507 ( \40056 , \39717 , \39723 );
or \U$31508 ( \40057 , \40054 , \40055 , \40056 );
buf \U$31509 ( \40058 , \40057 );
xor \U$31510 ( \40059 , \40053 , \40058 );
and \U$31512 ( \40060 , \32916 , \23696_nG9bd2 );
or \U$31513 ( \40061 , 1'b0 , \40060 );
xor \U$31514 ( \40062 , 1'b0 , \40061 );
buf \U$31515 ( \40063 , \40062 );
buf \U$31517 ( \40064 , \40063 );
and \U$31518 ( \40065 , \31636 , \24226_nG9bcf );
and \U$31519 ( \40066 , \31633 , \25298_nG9bcc );
or \U$31520 ( \40067 , \40065 , \40066 );
xor \U$31521 ( \40068 , \31632 , \40067 );
buf \U$31522 ( \40069 , \40068 );
buf \U$31524 ( \40070 , \40069 );
xor \U$31525 ( \40071 , \40064 , \40070 );
buf \U$31526 ( \40072 , \40071 );
and \U$31527 ( \40073 , \26431 , \29179_nG9bbd );
and \U$31528 ( \40074 , \26428 , \30366_nG9bba );
or \U$31529 ( \40075 , \40073 , \40074 );
xor \U$31530 ( \40076 , \26427 , \40075 );
buf \U$31531 ( \40077 , \40076 );
buf \U$31533 ( \40078 , \40077 );
xor \U$31534 ( \40079 , \40072 , \40078 );
and \U$31535 ( \40080 , \24792 , \30940_nG9bb7 );
and \U$31536 ( \40081 , \24789 , \32179_nG9bb4 );
or \U$31537 ( \40082 , \40080 , \40081 );
xor \U$31538 ( \40083 , \24788 , \40082 );
buf \U$31539 ( \40084 , \40083 );
buf \U$31541 ( \40085 , \40084 );
xor \U$31542 ( \40086 , \40079 , \40085 );
buf \U$31543 ( \40087 , \40086 );
and \U$31544 ( \40088 , \13370 , \37974_nG9b87 );
and \U$31545 ( \40089 , \13367 , \38337_nG9b84 );
or \U$31546 ( \40090 , \40088 , \40089 );
xor \U$31547 ( \40091 , \13366 , \40090 );
buf \U$31548 ( \40092 , \40091 );
buf \U$31550 ( \40093 , \40092 );
xor \U$31551 ( \40094 , \40087 , \40093 );
and \U$31552 ( \40095 , \12157 , \38663_nG9b81 );
and \U$31553 ( \40096 , \12154 , \38968_nG9b7e );
or \U$31554 ( \40097 , \40095 , \40096 );
xor \U$31555 ( \40098 , \12153 , \40097 );
buf \U$31556 ( \40099 , \40098 );
buf \U$31558 ( \40100 , \40099 );
xor \U$31559 ( \40101 , \40094 , \40100 );
buf \U$31560 ( \40102 , \40101 );
and \U$31561 ( \40103 , \39753 , \39758 );
and \U$31562 ( \40104 , \39753 , \39765 );
and \U$31563 ( \40105 , \39758 , \39765 );
or \U$31564 ( \40106 , \40103 , \40104 , \40105 );
buf \U$31565 ( \40107 , \40106 );
xor \U$31566 ( \40108 , \40102 , \40107 );
and \U$31567 ( \40109 , \39844 , \39850 );
buf \U$31568 ( \40110 , \40109 );
and \U$31569 ( \40111 , \29853 , \25860_nG9bc9 );
and \U$31570 ( \40112 , \29850 , \26887_nG9bc6 );
or \U$31571 ( \40113 , \40111 , \40112 );
xor \U$31572 ( \40114 , \29849 , \40113 );
buf \U$31573 ( \40115 , \40114 );
buf \U$31575 ( \40116 , \40115 );
xor \U$31576 ( \40117 , \40110 , \40116 );
and \U$31577 ( \40118 , \28118 , \27416_nG9bc3 );
and \U$31578 ( \40119 , \28115 , \28602_nG9bc0 );
or \U$31579 ( \40120 , \40118 , \40119 );
xor \U$31580 ( \40121 , \28114 , \40120 );
buf \U$31581 ( \40122 , \40121 );
buf \U$31583 ( \40123 , \40122 );
xor \U$31584 ( \40124 , \40117 , \40123 );
buf \U$31585 ( \40125 , \40124 );
and \U$31586 ( \40126 , \15940 , \36589_nG9b93 );
and \U$31587 ( \40127 , \15937 , \36986_nG9b90 );
or \U$31588 ( \40128 , \40126 , \40127 );
xor \U$31589 ( \40129 , \15936 , \40128 );
buf \U$31590 ( \40130 , \40129 );
buf \U$31592 ( \40131 , \40130 );
xor \U$31593 ( \40132 , \40125 , \40131 );
and \U$31594 ( \40133 , \10707 , \39963_nG9b75 );
and \U$31595 ( \40134 , \39892 , \39920 );
and \U$31596 ( \40135 , \39920 , \39952 );
and \U$31597 ( \40136 , \39892 , \39952 );
or \U$31598 ( \40137 , \40134 , \40135 , \40136 );
and \U$31599 ( \40138 , \39896 , \39907 );
and \U$31600 ( \40139 , \39907 , \39919 );
and \U$31601 ( \40140 , \39896 , \39919 );
or \U$31602 ( \40141 , \40138 , \40139 , \40140 );
and \U$31603 ( \40142 , \39925 , \39929 );
and \U$31604 ( \40143 , \39929 , \39951 );
and \U$31605 ( \40144 , \39925 , \39951 );
or \U$31606 ( \40145 , \40142 , \40143 , \40144 );
xor \U$31607 ( \40146 , \40141 , \40145 );
and \U$31608 ( \40147 , \39934 , \39938 );
and \U$31609 ( \40148 , \39938 , \39950 );
and \U$31610 ( \40149 , \39934 , \39950 );
or \U$31611 ( \40150 , \40147 , \40148 , \40149 );
and \U$31612 ( \40151 , \39900 , \39904 );
and \U$31613 ( \40152 , \39904 , \39906 );
and \U$31614 ( \40153 , \39900 , \39906 );
or \U$31615 ( \40154 , \40151 , \40152 , \40153 );
and \U$31616 ( \40155 , \39940 , \39944 );
and \U$31617 ( \40156 , \39944 , \39949 );
and \U$31618 ( \40157 , \39940 , \39949 );
or \U$31619 ( \40158 , \40155 , \40156 , \40157 );
xor \U$31620 ( \40159 , \40154 , \40158 );
and \U$31621 ( \40160 , \32794 , \24138 );
not \U$31622 ( \40161 , \40160 );
xnor \U$31623 ( \40162 , \40161 , \24144 );
not \U$31624 ( \40163 , \40162 );
xor \U$31625 ( \40164 , \40159 , \40163 );
xor \U$31626 ( \40165 , \40150 , \40164 );
and \U$31627 ( \40166 , \39909 , \39913 );
and \U$31628 ( \40167 , \39913 , \39918 );
and \U$31629 ( \40168 , \39909 , \39918 );
or \U$31630 ( \40169 , \40166 , \40167 , \40168 );
and \U$31631 ( \40170 , \30802 , \25826 );
and \U$31632 ( \40171 , \32054 , \25264 );
nor \U$31633 ( \40172 , \40170 , \40171 );
xnor \U$31634 ( \40173 , \40172 , \25773 );
and \U$31635 ( \40174 , \27313 , \29070 );
and \U$31636 ( \40175 , \28534 , \28526 );
nor \U$31637 ( \40176 , \40174 , \40175 );
xnor \U$31638 ( \40177 , \40176 , \29076 );
xor \U$31639 ( \40178 , \40173 , \40177 );
and \U$31640 ( \40179 , \25815 , \30823 );
and \U$31641 ( \40180 , \26829 , \30246 );
nor \U$31642 ( \40181 , \40179 , \40180 );
xnor \U$31643 ( \40182 , \40181 , \30813 );
xor \U$31644 ( \40183 , \40178 , \40182 );
xor \U$31645 ( \40184 , \40169 , \40183 );
and \U$31646 ( \40185 , \29084 , \27397 );
and \U$31647 ( \40186 , \30268 , \26807 );
nor \U$31648 ( \40187 , \40185 , \40186 );
xnor \U$31649 ( \40188 , \40187 , \27295 );
and \U$31650 ( \40189 , \24199 , \32854 );
and \U$31651 ( \40190 , \25272 , \32067 );
nor \U$31652 ( \40191 , \40189 , \40190 );
xnor \U$31653 ( \40192 , \40191 , \32805 );
xor \U$31654 ( \40193 , \40188 , \40192 );
and \U$31655 ( \40194 , \23617 , \32802 );
xor \U$31656 ( \40195 , \40193 , \40194 );
xor \U$31657 ( \40196 , \40184 , \40195 );
xor \U$31658 ( \40197 , \40165 , \40196 );
xor \U$31659 ( \40198 , \40146 , \40197 );
xor \U$31660 ( \40199 , \40137 , \40198 );
and \U$31661 ( \40200 , \39953 , \39957 );
and \U$31662 ( \40201 , \39958 , \39961 );
or \U$31663 ( \40202 , \40200 , \40201 );
xor \U$31664 ( \40203 , \40199 , \40202 );
buf g9b72 ( \40204_nG9b72 , \40203 );
and \U$31665 ( \40205 , \10704 , \40204_nG9b72 );
or \U$31666 ( \40206 , \40133 , \40205 );
xor \U$31667 ( \40207 , \10703 , \40206 );
buf \U$31668 ( \40208 , \40207 );
buf \U$31670 ( \40209 , \40208 );
xor \U$31671 ( \40210 , \40132 , \40209 );
buf \U$31672 ( \40211 , \40210 );
xor \U$31673 ( \40212 , \40108 , \40211 );
buf \U$31674 ( \40213 , \40212 );
and \U$31675 ( \40214 , \39869 , \39874 );
and \U$31676 ( \40215 , \39869 , \39970 );
and \U$31677 ( \40216 , \39874 , \39970 );
or \U$31678 ( \40217 , \40214 , \40215 , \40216 );
buf \U$31679 ( \40218 , \40217 );
xor \U$31680 ( \40219 , \40213 , \40218 );
and \U$31681 ( \40220 , \39794 , \39800 );
and \U$31682 ( \40221 , \39794 , \39807 );
and \U$31683 ( \40222 , \39800 , \39807 );
or \U$31684 ( \40223 , \40220 , \40221 , \40222 );
buf \U$31685 ( \40224 , \40223 );
and \U$31686 ( \40225 , \39823 , \39829 );
and \U$31687 ( \40226 , \39823 , \39836 );
and \U$31688 ( \40227 , \39829 , \39836 );
or \U$31689 ( \40228 , \40225 , \40226 , \40227 );
buf \U$31690 ( \40229 , \40228 );
xor \U$31691 ( \40230 , \40224 , \40229 );
and \U$31692 ( \40231 , \23201 , \32888_nG9bb1 );
and \U$31693 ( \40232 , \23198 , \33181_nG9bae );
or \U$31694 ( \40233 , \40231 , \40232 );
xor \U$31695 ( \40234 , \23197 , \40233 );
buf \U$31696 ( \40235 , \40234 );
buf \U$31698 ( \40236 , \40235 );
and \U$31699 ( \40237 , \21658 , \33613_nG9bab );
and \U$31700 ( \40238 , \21655 , \34041_nG9ba8 );
or \U$31701 ( \40239 , \40237 , \40238 );
xor \U$31702 ( \40240 , \21654 , \40239 );
buf \U$31703 ( \40241 , \40240 );
buf \U$31705 ( \40242 , \40241 );
xor \U$31706 ( \40243 , \40236 , \40242 );
and \U$31707 ( \40244 , \20155 , \34294_nG9ba5 );
and \U$31708 ( \40245 , \20152 , \34643_nG9ba2 );
or \U$31709 ( \40246 , \40244 , \40245 );
xor \U$31710 ( \40247 , \20151 , \40246 );
buf \U$31711 ( \40248 , \40247 );
buf \U$31713 ( \40249 , \40248 );
xor \U$31714 ( \40250 , \40243 , \40249 );
buf \U$31715 ( \40251 , \40250 );
xor \U$31716 ( \40252 , \40230 , \40251 );
buf \U$31717 ( \40253 , \40252 );
and \U$31718 ( \40254 , \39852 , \39858 );
and \U$31719 ( \40255 , \39852 , \39865 );
and \U$31720 ( \40256 , \39858 , \39865 );
or \U$31721 ( \40257 , \40254 , \40255 , \40256 );
buf \U$31722 ( \40258 , \40257 );
and \U$31723 ( \40259 , \14631 , \37250_nG9b8d );
and \U$31724 ( \40260 , \14628 , \37607_nG9b8a );
or \U$31725 ( \40261 , \40259 , \40260 );
xor \U$31726 ( \40262 , \14627 , \40261 );
buf \U$31727 ( \40263 , \40262 );
buf \U$31729 ( \40264 , \40263 );
xor \U$31730 ( \40265 , \40258 , \40264 );
and \U$31731 ( \40266 , \10421 , \39334_nG9b7b );
and \U$31732 ( \40267 , \10418 , \39591_nG9b78 );
or \U$31733 ( \40268 , \40266 , \40267 );
xor \U$31734 ( \40269 , \10417 , \40268 );
buf \U$31735 ( \40270 , \40269 );
buf \U$31737 ( \40271 , \40270 );
xor \U$31738 ( \40272 , \40265 , \40271 );
buf \U$31739 ( \40273 , \40272 );
xor \U$31740 ( \40274 , \40253 , \40273 );
and \U$31741 ( \40275 , \39817 , \39838 );
and \U$31742 ( \40276 , \39817 , \39867 );
and \U$31743 ( \40277 , \39838 , \39867 );
or \U$31744 ( \40278 , \40275 , \40276 , \40277 );
buf \U$31745 ( \40279 , \40278 );
xor \U$31746 ( \40280 , \40274 , \40279 );
buf \U$31747 ( \40281 , \40280 );
xor \U$31748 ( \40282 , \40219 , \40281 );
buf \U$31749 ( \40283 , \40282 );
xor \U$31750 ( \40284 , \40059 , \40283 );
and \U$31751 ( \40285 , \39994 , \40284 );
and \U$31753 ( \40286 , \39988 , \39993 );
or \U$31755 ( \40287 , 1'b0 , \40286 , 1'b0 );
xor \U$31756 ( \40288 , \40285 , \40287 );
and \U$31758 ( \40289 , \39981 , \39987 );
and \U$31759 ( \40290 , \39983 , \39987 );
or \U$31760 ( \40291 , 1'b0 , \40289 , \40290 );
xor \U$31761 ( \40292 , \40288 , \40291 );
xor \U$31768 ( \40293 , \40292 , 1'b0 );
and \U$31769 ( \40294 , \40053 , \40058 );
and \U$31770 ( \40295 , \40053 , \40283 );
and \U$31771 ( \40296 , \40058 , \40283 );
or \U$31772 ( \40297 , \40294 , \40295 , \40296 );
xor \U$31773 ( \40298 , \40293 , \40297 );
and \U$31774 ( \40299 , \39999 , \40004 );
and \U$31775 ( \40300 , \39999 , \40051 );
and \U$31776 ( \40301 , \40004 , \40051 );
or \U$31777 ( \40302 , \40299 , \40300 , \40301 );
buf \U$31778 ( \40303 , \40302 );
and \U$31779 ( \40304 , \40021 , \40026 );
and \U$31780 ( \40305 , \40021 , \40047 );
and \U$31781 ( \40306 , \40026 , \40047 );
or \U$31782 ( \40307 , \40304 , \40305 , \40306 );
buf \U$31783 ( \40308 , \40307 );
and \U$31784 ( \40309 , \40064 , \40070 );
buf \U$31785 ( \40310 , \40309 );
and \U$31786 ( \40311 , \31636 , \25298_nG9bcc );
and \U$31787 ( \40312 , \31633 , \25860_nG9bc9 );
or \U$31788 ( \40313 , \40311 , \40312 );
xor \U$31789 ( \40314 , \31632 , \40313 );
buf \U$31790 ( \40315 , \40314 );
buf \U$31792 ( \40316 , \40315 );
xor \U$31793 ( \40317 , \40310 , \40316 );
and \U$31794 ( \40318 , \26431 , \30366_nG9bba );
and \U$31795 ( \40319 , \26428 , \30940_nG9bb7 );
or \U$31796 ( \40320 , \40318 , \40319 );
xor \U$31797 ( \40321 , \26427 , \40320 );
buf \U$31798 ( \40322 , \40321 );
buf \U$31800 ( \40323 , \40322 );
xor \U$31801 ( \40324 , \40317 , \40323 );
buf \U$31802 ( \40325 , \40324 );
and \U$31803 ( \40326 , \40236 , \40242 );
and \U$31804 ( \40327 , \40236 , \40249 );
and \U$31805 ( \40328 , \40242 , \40249 );
or \U$31806 ( \40329 , \40326 , \40327 , \40328 );
buf \U$31807 ( \40330 , \40329 );
xor \U$31808 ( \40331 , \40325 , \40330 );
and \U$31809 ( \40332 , \17297 , \36172_nG9b96 );
and \U$31810 ( \40333 , \17294 , \36589_nG9b93 );
or \U$31811 ( \40334 , \40332 , \40333 );
xor \U$31812 ( \40335 , \17293 , \40334 );
buf \U$31813 ( \40336 , \40335 );
buf \U$31815 ( \40337 , \40336 );
xor \U$31816 ( \40338 , \40331 , \40337 );
buf \U$31817 ( \40339 , \40338 );
xor \U$31818 ( \40340 , \40308 , \40339 );
and \U$31819 ( \40341 , \40224 , \40229 );
and \U$31820 ( \40342 , \40224 , \40251 );
and \U$31821 ( \40343 , \40229 , \40251 );
or \U$31822 ( \40344 , \40341 , \40342 , \40343 );
buf \U$31823 ( \40345 , \40344 );
xor \U$31824 ( \40346 , \40340 , \40345 );
buf \U$31825 ( \40347 , \40346 );
and \U$31826 ( \40348 , \40253 , \40273 );
and \U$31827 ( \40349 , \40253 , \40279 );
and \U$31828 ( \40350 , \40273 , \40279 );
or \U$31829 ( \40351 , \40348 , \40349 , \40350 );
buf \U$31830 ( \40352 , \40351 );
xor \U$31831 ( \40353 , \40347 , \40352 );
and \U$31832 ( \40354 , \40072 , \40078 );
and \U$31833 ( \40355 , \40072 , \40085 );
and \U$31834 ( \40356 , \40078 , \40085 );
or \U$31835 ( \40357 , \40354 , \40355 , \40356 );
buf \U$31836 ( \40358 , \40357 );
and \U$31837 ( \40359 , \15940 , \36986_nG9b90 );
and \U$31838 ( \40360 , \15937 , \37250_nG9b8d );
or \U$31839 ( \40361 , \40359 , \40360 );
xor \U$31840 ( \40362 , \15936 , \40361 );
buf \U$31841 ( \40363 , \40362 );
buf \U$31843 ( \40364 , \40363 );
xor \U$31844 ( \40365 , \40358 , \40364 );
and \U$31845 ( \40366 , \12157 , \38968_nG9b7e );
and \U$31846 ( \40367 , \12154 , \39334_nG9b7b );
or \U$31847 ( \40368 , \40366 , \40367 );
xor \U$31848 ( \40369 , \12153 , \40368 );
buf \U$31849 ( \40370 , \40369 );
buf \U$31851 ( \40371 , \40370 );
xor \U$31852 ( \40372 , \40365 , \40371 );
buf \U$31853 ( \40373 , \40372 );
and \U$31854 ( \40374 , \21658 , \34041_nG9ba8 );
and \U$31855 ( \40375 , \21655 , \34294_nG9ba5 );
or \U$31856 ( \40376 , \40374 , \40375 );
xor \U$31857 ( \40377 , \21654 , \40376 );
buf \U$31858 ( \40378 , \40377 );
buf \U$31860 ( \40379 , \40378 );
and \U$31861 ( \40380 , \13370 , \38337_nG9b84 );
and \U$31862 ( \40381 , \13367 , \38663_nG9b81 );
or \U$31863 ( \40382 , \40380 , \40381 );
xor \U$31864 ( \40383 , \13366 , \40382 );
buf \U$31865 ( \40384 , \40383 );
buf \U$31867 ( \40385 , \40384 );
xor \U$31868 ( \40386 , \40379 , \40385 );
and \U$31869 ( \40387 , \10707 , \40204_nG9b72 );
and \U$31870 ( \40388 , \40150 , \40164 );
and \U$31871 ( \40389 , \40164 , \40196 );
and \U$31872 ( \40390 , \40150 , \40196 );
or \U$31873 ( \40391 , \40388 , \40389 , \40390 );
and \U$31874 ( \40392 , \40188 , \40192 );
and \U$31875 ( \40393 , \40192 , \40194 );
and \U$31876 ( \40394 , \40188 , \40194 );
or \U$31877 ( \40395 , \40392 , \40393 , \40394 );
not \U$31878 ( \40396 , \24144 );
and \U$31879 ( \40397 , \32054 , \25826 );
and \U$31880 ( \40398 , \32794 , \25264 );
nor \U$31881 ( \40399 , \40397 , \40398 );
xnor \U$31882 ( \40400 , \40399 , \25773 );
xor \U$31883 ( \40401 , \40396 , \40400 );
and \U$31884 ( \40402 , \28534 , \29070 );
and \U$31885 ( \40403 , \29084 , \28526 );
nor \U$31886 ( \40404 , \40402 , \40403 );
xnor \U$31887 ( \40405 , \40404 , \29076 );
xor \U$31888 ( \40406 , \40401 , \40405 );
xor \U$31889 ( \40407 , \40395 , \40406 );
and \U$31890 ( \40408 , \30268 , \27397 );
and \U$31891 ( \40409 , \30802 , \26807 );
nor \U$31892 ( \40410 , \40408 , \40409 );
xnor \U$31893 ( \40411 , \40410 , \27295 );
and \U$31894 ( \40412 , \26829 , \30823 );
and \U$31895 ( \40413 , \27313 , \30246 );
nor \U$31896 ( \40414 , \40412 , \40413 );
xnor \U$31897 ( \40415 , \40414 , \30813 );
xor \U$31898 ( \40416 , \40411 , \40415 );
and \U$31899 ( \40417 , \25272 , \32854 );
and \U$31900 ( \40418 , \25815 , \32067 );
nor \U$31901 ( \40419 , \40417 , \40418 );
xnor \U$31902 ( \40420 , \40419 , \32805 );
xor \U$31903 ( \40421 , \40416 , \40420 );
xor \U$31904 ( \40422 , \40407 , \40421 );
xor \U$31905 ( \40423 , \40391 , \40422 );
and \U$31906 ( \40424 , \40154 , \40158 );
and \U$31907 ( \40425 , \40158 , \40163 );
and \U$31908 ( \40426 , \40154 , \40163 );
or \U$31909 ( \40427 , \40424 , \40425 , \40426 );
and \U$31910 ( \40428 , \40169 , \40183 );
and \U$31911 ( \40429 , \40183 , \40195 );
and \U$31912 ( \40430 , \40169 , \40195 );
or \U$31913 ( \40431 , \40428 , \40429 , \40430 );
xor \U$31914 ( \40432 , \40427 , \40431 );
and \U$31915 ( \40433 , \40173 , \40177 );
and \U$31916 ( \40434 , \40177 , \40182 );
and \U$31917 ( \40435 , \40173 , \40182 );
or \U$31918 ( \40436 , \40433 , \40434 , \40435 );
buf \U$31919 ( \40437 , \40162 );
xor \U$31920 ( \40438 , \40436 , \40437 );
and \U$31921 ( \40439 , \24199 , \32802 );
xor \U$31922 ( \40440 , \40438 , \40439 );
xor \U$31923 ( \40441 , \40432 , \40440 );
xor \U$31924 ( \40442 , \40423 , \40441 );
and \U$31925 ( \40443 , \40141 , \40145 );
and \U$31926 ( \40444 , \40145 , \40197 );
and \U$31927 ( \40445 , \40141 , \40197 );
or \U$31928 ( \40446 , \40443 , \40444 , \40445 );
xor \U$31929 ( \40447 , \40442 , \40446 );
and \U$31930 ( \40448 , \40137 , \40198 );
and \U$31931 ( \40449 , \40199 , \40202 );
or \U$31932 ( \40450 , \40448 , \40449 );
xor \U$31933 ( \40451 , \40447 , \40450 );
buf g9b6f ( \40452_nG9b6f , \40451 );
and \U$31934 ( \40453 , \10704 , \40452_nG9b6f );
or \U$31935 ( \40454 , \40387 , \40453 );
xor \U$31936 ( \40455 , \10703 , \40454 );
buf \U$31937 ( \40456 , \40455 );
buf \U$31939 ( \40457 , \40456 );
xor \U$31940 ( \40458 , \40386 , \40457 );
buf \U$31941 ( \40459 , \40458 );
xor \U$31942 ( \40460 , \40373 , \40459 );
and \U$31943 ( \40461 , \40110 , \40116 );
and \U$31944 ( \40462 , \40110 , \40123 );
and \U$31945 ( \40463 , \40116 , \40123 );
or \U$31946 ( \40464 , \40461 , \40462 , \40463 );
buf \U$31947 ( \40465 , \40464 );
and \U$31948 ( \40466 , \14631 , \37607_nG9b8a );
and \U$31949 ( \40467 , \14628 , \37974_nG9b87 );
or \U$31950 ( \40468 , \40466 , \40467 );
xor \U$31951 ( \40469 , \14627 , \40468 );
buf \U$31952 ( \40470 , \40469 );
buf \U$31954 ( \40471 , \40470 );
xor \U$31955 ( \40472 , \40465 , \40471 );
and \U$31956 ( \40473 , \10421 , \39591_nG9b78 );
and \U$31957 ( \40474 , \10418 , \39963_nG9b75 );
or \U$31958 ( \40475 , \40473 , \40474 );
xor \U$31959 ( \40476 , \10417 , \40475 );
buf \U$31960 ( \40477 , \40476 );
buf \U$31962 ( \40478 , \40477 );
xor \U$31963 ( \40479 , \40472 , \40478 );
buf \U$31964 ( \40480 , \40479 );
xor \U$31965 ( \40481 , \40460 , \40480 );
buf \U$31966 ( \40482 , \40481 );
xor \U$31967 ( \40483 , \40353 , \40482 );
buf \U$31968 ( \40484 , \40483 );
xor \U$31969 ( \40485 , \40303 , \40484 );
and \U$31970 ( \40486 , \40213 , \40218 );
and \U$31971 ( \40487 , \40213 , \40281 );
and \U$31972 ( \40488 , \40218 , \40281 );
or \U$31973 ( \40489 , \40486 , \40487 , \40488 );
buf \U$31974 ( \40490 , \40489 );
and \U$31975 ( \40491 , \40102 , \40107 );
and \U$31976 ( \40492 , \40102 , \40211 );
and \U$31977 ( \40493 , \40107 , \40211 );
or \U$31978 ( \40494 , \40491 , \40492 , \40493 );
buf \U$31979 ( \40495 , \40494 );
and \U$31980 ( \40496 , \40087 , \40093 );
and \U$31981 ( \40497 , \40087 , \40100 );
and \U$31982 ( \40498 , \40093 , \40100 );
or \U$31983 ( \40499 , \40496 , \40497 , \40498 );
buf \U$31984 ( \40500 , \40499 );
and \U$31985 ( \40501 , \40125 , \40131 );
and \U$31986 ( \40502 , \40125 , \40209 );
and \U$31987 ( \40503 , \40131 , \40209 );
or \U$31988 ( \40504 , \40501 , \40502 , \40503 );
buf \U$31989 ( \40505 , \40504 );
xor \U$31990 ( \40506 , \40500 , \40505 );
and \U$31991 ( \40507 , \23201 , \33181_nG9bae );
and \U$31992 ( \40508 , \23198 , \33613_nG9bab );
or \U$31993 ( \40509 , \40507 , \40508 );
xor \U$31994 ( \40510 , \23197 , \40509 );
buf \U$31995 ( \40511 , \40510 );
buf \U$31997 ( \40512 , \40511 );
and \U$31998 ( \40513 , \20155 , \34643_nG9ba2 );
and \U$31999 ( \40514 , \20152 , \35094_nG9b9f );
or \U$32000 ( \40515 , \40513 , \40514 );
xor \U$32001 ( \40516 , \20151 , \40515 );
buf \U$32002 ( \40517 , \40516 );
buf \U$32004 ( \40518 , \40517 );
xor \U$32005 ( \40519 , \40512 , \40518 );
and \U$32006 ( \40520 , \18702 , \35570_nG9b9c );
and \U$32007 ( \40521 , \18699 , \35801_nG9b99 );
or \U$32008 ( \40522 , \40520 , \40521 );
xor \U$32009 ( \40523 , \18698 , \40522 );
buf \U$32010 ( \40524 , \40523 );
buf \U$32012 ( \40525 , \40524 );
xor \U$32013 ( \40526 , \40519 , \40525 );
buf \U$32014 ( \40527 , \40526 );
xor \U$32015 ( \40528 , \40506 , \40527 );
buf \U$32016 ( \40529 , \40528 );
xor \U$32017 ( \40530 , \40495 , \40529 );
and \U$32018 ( \40531 , \40258 , \40264 );
and \U$32019 ( \40532 , \40258 , \40271 );
and \U$32020 ( \40533 , \40264 , \40271 );
or \U$32021 ( \40534 , \40531 , \40532 , \40533 );
buf \U$32022 ( \40535 , \40534 );
and \U$32023 ( \40536 , \40032 , \40038 );
and \U$32024 ( \40537 , \40032 , \40045 );
and \U$32025 ( \40538 , \40038 , \40045 );
or \U$32026 ( \40539 , \40536 , \40537 , \40538 );
buf \U$32027 ( \40540 , \40539 );
xor \U$32028 ( \40541 , \40535 , \40540 );
and \U$32030 ( \40542 , \32916 , \24226_nG9bcf );
or \U$32031 ( \40543 , 1'b0 , \40542 );
xor \U$32032 ( \40544 , 1'b0 , \40543 );
buf \U$32033 ( \40545 , \40544 );
buf \U$32035 ( \40546 , \40545 );
and \U$32036 ( \40547 , \29853 , \26887_nG9bc6 );
and \U$32037 ( \40548 , \29850 , \27416_nG9bc3 );
or \U$32038 ( \40549 , \40547 , \40548 );
xor \U$32039 ( \40550 , \29849 , \40549 );
buf \U$32040 ( \40551 , \40550 );
buf \U$32042 ( \40552 , \40551 );
xor \U$32043 ( \40553 , \40546 , \40552 );
buf \U$32044 ( \40554 , \40553 );
and \U$32045 ( \40555 , \28118 , \28602_nG9bc0 );
and \U$32046 ( \40556 , \28115 , \29179_nG9bbd );
or \U$32047 ( \40557 , \40555 , \40556 );
xor \U$32048 ( \40558 , \28114 , \40557 );
buf \U$32049 ( \40559 , \40558 );
buf \U$32051 ( \40560 , \40559 );
xor \U$32052 ( \40561 , \40554 , \40560 );
and \U$32053 ( \40562 , \24792 , \32179_nG9bb4 );
and \U$32054 ( \40563 , \24789 , \32888_nG9bb1 );
or \U$32055 ( \40564 , \40562 , \40563 );
xor \U$32056 ( \40565 , \24788 , \40564 );
buf \U$32057 ( \40566 , \40565 );
buf \U$32059 ( \40567 , \40566 );
xor \U$32060 ( \40568 , \40561 , \40567 );
buf \U$32061 ( \40569 , \40568 );
xor \U$32062 ( \40570 , \40541 , \40569 );
buf \U$32063 ( \40571 , \40570 );
xor \U$32064 ( \40572 , \40530 , \40571 );
buf \U$32065 ( \40573 , \40572 );
xor \U$32066 ( \40574 , \40490 , \40573 );
and \U$32067 ( \40575 , \40010 , \40015 );
and \U$32068 ( \40576 , \40010 , \40049 );
and \U$32069 ( \40577 , \40015 , \40049 );
or \U$32070 ( \40578 , \40575 , \40576 , \40577 );
buf \U$32071 ( \40579 , \40578 );
xor \U$32072 ( \40580 , \40574 , \40579 );
buf \U$32073 ( \40581 , \40580 );
xor \U$32074 ( \40582 , \40485 , \40581 );
and \U$32075 ( \40583 , \40298 , \40582 );
and \U$32077 ( \40584 , \40292 , \40297 );
or \U$32079 ( \40585 , 1'b0 , \40584 , 1'b0 );
xor \U$32080 ( \40586 , \40583 , \40585 );
and \U$32082 ( \40587 , \40285 , \40291 );
and \U$32083 ( \40588 , \40287 , \40291 );
or \U$32084 ( \40589 , 1'b0 , \40587 , \40588 );
xor \U$32085 ( \40590 , \40586 , \40589 );
xor \U$32092 ( \40591 , \40590 , 1'b0 );
and \U$32093 ( \40592 , \40303 , \40484 );
and \U$32094 ( \40593 , \40303 , \40581 );
and \U$32095 ( \40594 , \40484 , \40581 );
or \U$32096 ( \40595 , \40592 , \40593 , \40594 );
xor \U$32097 ( \40596 , \40591 , \40595 );
and \U$32098 ( \40597 , \40347 , \40352 );
and \U$32099 ( \40598 , \40347 , \40482 );
and \U$32100 ( \40599 , \40352 , \40482 );
or \U$32101 ( \40600 , \40597 , \40598 , \40599 );
buf \U$32102 ( \40601 , \40600 );
and \U$32103 ( \40602 , \40373 , \40459 );
and \U$32104 ( \40603 , \40373 , \40480 );
and \U$32105 ( \40604 , \40459 , \40480 );
or \U$32106 ( \40605 , \40602 , \40603 , \40604 );
buf \U$32107 ( \40606 , \40605 );
and \U$32108 ( \40607 , \17297 , \36589_nG9b93 );
and \U$32109 ( \40608 , \17294 , \36986_nG9b90 );
or \U$32110 ( \40609 , \40607 , \40608 );
xor \U$32111 ( \40610 , \17293 , \40609 );
buf \U$32112 ( \40611 , \40610 );
buf \U$32114 ( \40612 , \40611 );
and \U$32115 ( \40613 , \15940 , \37250_nG9b8d );
and \U$32116 ( \40614 , \15937 , \37607_nG9b8a );
or \U$32117 ( \40615 , \40613 , \40614 );
xor \U$32118 ( \40616 , \15936 , \40615 );
buf \U$32119 ( \40617 , \40616 );
buf \U$32121 ( \40618 , \40617 );
xor \U$32122 ( \40619 , \40612 , \40618 );
and \U$32123 ( \40620 , \12157 , \39334_nG9b7b );
and \U$32124 ( \40621 , \12154 , \39591_nG9b78 );
or \U$32125 ( \40622 , \40620 , \40621 );
xor \U$32126 ( \40623 , \12153 , \40622 );
buf \U$32127 ( \40624 , \40623 );
buf \U$32129 ( \40625 , \40624 );
xor \U$32130 ( \40626 , \40619 , \40625 );
buf \U$32131 ( \40627 , \40626 );
and \U$32132 ( \40628 , \23201 , \33613_nG9bab );
and \U$32133 ( \40629 , \23198 , \34041_nG9ba8 );
or \U$32134 ( \40630 , \40628 , \40629 );
xor \U$32135 ( \40631 , \23197 , \40630 );
buf \U$32136 ( \40632 , \40631 );
buf \U$32138 ( \40633 , \40632 );
and \U$32139 ( \40634 , \20155 , \35094_nG9b9f );
and \U$32140 ( \40635 , \20152 , \35570_nG9b9c );
or \U$32141 ( \40636 , \40634 , \40635 );
xor \U$32142 ( \40637 , \20151 , \40636 );
buf \U$32143 ( \40638 , \40637 );
buf \U$32145 ( \40639 , \40638 );
xor \U$32146 ( \40640 , \40633 , \40639 );
and \U$32147 ( \40641 , \18702 , \35801_nG9b99 );
and \U$32148 ( \40642 , \18699 , \36172_nG9b96 );
or \U$32149 ( \40643 , \40641 , \40642 );
xor \U$32150 ( \40644 , \18698 , \40643 );
buf \U$32151 ( \40645 , \40644 );
buf \U$32153 ( \40646 , \40645 );
xor \U$32154 ( \40647 , \40640 , \40646 );
buf \U$32155 ( \40648 , \40647 );
xor \U$32156 ( \40649 , \40627 , \40648 );
and \U$32157 ( \40650 , \40358 , \40364 );
and \U$32158 ( \40651 , \40358 , \40371 );
and \U$32159 ( \40652 , \40364 , \40371 );
or \U$32160 ( \40653 , \40650 , \40651 , \40652 );
buf \U$32161 ( \40654 , \40653 );
xor \U$32162 ( \40655 , \40649 , \40654 );
buf \U$32163 ( \40656 , \40655 );
xor \U$32164 ( \40657 , \40606 , \40656 );
and \U$32165 ( \40658 , \40500 , \40505 );
and \U$32166 ( \40659 , \40500 , \40527 );
and \U$32167 ( \40660 , \40505 , \40527 );
or \U$32168 ( \40661 , \40658 , \40659 , \40660 );
buf \U$32169 ( \40662 , \40661 );
xor \U$32170 ( \40663 , \40657 , \40662 );
buf \U$32171 ( \40664 , \40663 );
xor \U$32172 ( \40665 , \40601 , \40664 );
and \U$32173 ( \40666 , \40379 , \40385 );
and \U$32174 ( \40667 , \40379 , \40457 );
and \U$32175 ( \40668 , \40385 , \40457 );
or \U$32176 ( \40669 , \40666 , \40667 , \40668 );
buf \U$32177 ( \40670 , \40669 );
and \U$32178 ( \40671 , \40465 , \40471 );
and \U$32179 ( \40672 , \40465 , \40478 );
and \U$32180 ( \40673 , \40471 , \40478 );
or \U$32181 ( \40674 , \40671 , \40672 , \40673 );
buf \U$32182 ( \40675 , \40674 );
xor \U$32183 ( \40676 , \40670 , \40675 );
and \U$32185 ( \40677 , \32916 , \25298_nG9bcc );
or \U$32186 ( \40678 , 1'b0 , \40677 );
xor \U$32187 ( \40679 , 1'b0 , \40678 );
buf \U$32188 ( \40680 , \40679 );
buf \U$32190 ( \40681 , \40680 );
and \U$32191 ( \40682 , \29853 , \27416_nG9bc3 );
and \U$32192 ( \40683 , \29850 , \28602_nG9bc0 );
or \U$32193 ( \40684 , \40682 , \40683 );
xor \U$32194 ( \40685 , \29849 , \40684 );
buf \U$32195 ( \40686 , \40685 );
buf \U$32197 ( \40687 , \40686 );
xor \U$32198 ( \40688 , \40681 , \40687 );
buf \U$32199 ( \40689 , \40688 );
and \U$32200 ( \40690 , \40546 , \40552 );
buf \U$32201 ( \40691 , \40690 );
xor \U$32202 ( \40692 , \40689 , \40691 );
and \U$32203 ( \40693 , \24792 , \32888_nG9bb1 );
and \U$32204 ( \40694 , \24789 , \33181_nG9bae );
or \U$32205 ( \40695 , \40693 , \40694 );
xor \U$32206 ( \40696 , \24788 , \40695 );
buf \U$32207 ( \40697 , \40696 );
buf \U$32209 ( \40698 , \40697 );
xor \U$32210 ( \40699 , \40692 , \40698 );
buf \U$32211 ( \40700 , \40699 );
xor \U$32212 ( \40701 , \40676 , \40700 );
buf \U$32213 ( \40702 , \40701 );
and \U$32214 ( \40703 , \40535 , \40540 );
and \U$32215 ( \40704 , \40535 , \40569 );
and \U$32216 ( \40705 , \40540 , \40569 );
or \U$32217 ( \40706 , \40703 , \40704 , \40705 );
buf \U$32218 ( \40707 , \40706 );
xor \U$32219 ( \40708 , \40702 , \40707 );
and \U$32220 ( \40709 , \40512 , \40518 );
and \U$32221 ( \40710 , \40512 , \40525 );
and \U$32222 ( \40711 , \40518 , \40525 );
or \U$32223 ( \40712 , \40709 , \40710 , \40711 );
buf \U$32224 ( \40713 , \40712 );
and \U$32225 ( \40714 , \40554 , \40560 );
and \U$32226 ( \40715 , \40554 , \40567 );
and \U$32227 ( \40716 , \40560 , \40567 );
or \U$32228 ( \40717 , \40714 , \40715 , \40716 );
buf \U$32229 ( \40718 , \40717 );
xor \U$32230 ( \40719 , \40713 , \40718 );
and \U$32231 ( \40720 , \31636 , \25860_nG9bc9 );
and \U$32232 ( \40721 , \31633 , \26887_nG9bc6 );
or \U$32233 ( \40722 , \40720 , \40721 );
xor \U$32234 ( \40723 , \31632 , \40722 );
buf \U$32235 ( \40724 , \40723 );
buf \U$32237 ( \40725 , \40724 );
and \U$32238 ( \40726 , \28118 , \29179_nG9bbd );
and \U$32239 ( \40727 , \28115 , \30366_nG9bba );
or \U$32240 ( \40728 , \40726 , \40727 );
xor \U$32241 ( \40729 , \28114 , \40728 );
buf \U$32242 ( \40730 , \40729 );
buf \U$32244 ( \40731 , \40730 );
xor \U$32245 ( \40732 , \40725 , \40731 );
and \U$32246 ( \40733 , \26431 , \30940_nG9bb7 );
and \U$32247 ( \40734 , \26428 , \32179_nG9bb4 );
or \U$32248 ( \40735 , \40733 , \40734 );
xor \U$32249 ( \40736 , \26427 , \40735 );
buf \U$32250 ( \40737 , \40736 );
buf \U$32252 ( \40738 , \40737 );
xor \U$32253 ( \40739 , \40732 , \40738 );
buf \U$32254 ( \40740 , \40739 );
xor \U$32255 ( \40741 , \40719 , \40740 );
buf \U$32256 ( \40742 , \40741 );
xor \U$32257 ( \40743 , \40708 , \40742 );
buf \U$32258 ( \40744 , \40743 );
xor \U$32259 ( \40745 , \40665 , \40744 );
buf \U$32260 ( \40746 , \40745 );
and \U$32261 ( \40747 , \40490 , \40573 );
and \U$32262 ( \40748 , \40490 , \40579 );
and \U$32263 ( \40749 , \40573 , \40579 );
or \U$32264 ( \40750 , \40747 , \40748 , \40749 );
buf \U$32265 ( \40751 , \40750 );
xor \U$32266 ( \40752 , \40746 , \40751 );
and \U$32267 ( \40753 , \40495 , \40529 );
and \U$32268 ( \40754 , \40495 , \40571 );
and \U$32269 ( \40755 , \40529 , \40571 );
or \U$32270 ( \40756 , \40753 , \40754 , \40755 );
buf \U$32271 ( \40757 , \40756 );
and \U$32272 ( \40758 , \40308 , \40339 );
and \U$32273 ( \40759 , \40308 , \40345 );
and \U$32274 ( \40760 , \40339 , \40345 );
or \U$32275 ( \40761 , \40758 , \40759 , \40760 );
buf \U$32276 ( \40762 , \40761 );
xor \U$32277 ( \40763 , \40757 , \40762 );
and \U$32278 ( \40764 , \40325 , \40330 );
and \U$32279 ( \40765 , \40325 , \40337 );
and \U$32280 ( \40766 , \40330 , \40337 );
or \U$32281 ( \40767 , \40764 , \40765 , \40766 );
buf \U$32282 ( \40768 , \40767 );
and \U$32283 ( \40769 , \21658 , \34294_nG9ba5 );
and \U$32284 ( \40770 , \21655 , \34643_nG9ba2 );
or \U$32285 ( \40771 , \40769 , \40770 );
xor \U$32286 ( \40772 , \21654 , \40771 );
buf \U$32287 ( \40773 , \40772 );
buf \U$32289 ( \40774 , \40773 );
and \U$32290 ( \40775 , \13370 , \38663_nG9b81 );
and \U$32291 ( \40776 , \13367 , \38968_nG9b7e );
or \U$32292 ( \40777 , \40775 , \40776 );
xor \U$32293 ( \40778 , \13366 , \40777 );
buf \U$32294 ( \40779 , \40778 );
buf \U$32296 ( \40780 , \40779 );
xor \U$32297 ( \40781 , \40774 , \40780 );
and \U$32298 ( \40782 , \10707 , \40452_nG9b6f );
and \U$32299 ( \40783 , \40427 , \40431 );
and \U$32300 ( \40784 , \40431 , \40440 );
and \U$32301 ( \40785 , \40427 , \40440 );
or \U$32302 ( \40786 , \40783 , \40784 , \40785 );
and \U$32303 ( \40787 , \40396 , \40400 );
and \U$32304 ( \40788 , \40400 , \40405 );
and \U$32305 ( \40789 , \40396 , \40405 );
or \U$32306 ( \40790 , \40787 , \40788 , \40789 );
and \U$32307 ( \40791 , \40411 , \40415 );
and \U$32308 ( \40792 , \40415 , \40420 );
and \U$32309 ( \40793 , \40411 , \40420 );
or \U$32310 ( \40794 , \40791 , \40792 , \40793 );
xor \U$32311 ( \40795 , \40790 , \40794 );
and \U$32312 ( \40796 , \32794 , \25826 );
not \U$32313 ( \40797 , \40796 );
xnor \U$32314 ( \40798 , \40797 , \25773 );
and \U$32315 ( \40799 , \27313 , \30823 );
and \U$32316 ( \40800 , \28534 , \30246 );
nor \U$32317 ( \40801 , \40799 , \40800 );
xnor \U$32318 ( \40802 , \40801 , \30813 );
xor \U$32319 ( \40803 , \40798 , \40802 );
and \U$32320 ( \40804 , \25815 , \32854 );
and \U$32321 ( \40805 , \26829 , \32067 );
nor \U$32322 ( \40806 , \40804 , \40805 );
xnor \U$32323 ( \40807 , \40806 , \32805 );
xor \U$32324 ( \40808 , \40803 , \40807 );
xor \U$32325 ( \40809 , \40795 , \40808 );
xor \U$32326 ( \40810 , \40786 , \40809 );
and \U$32327 ( \40811 , \40436 , \40437 );
and \U$32328 ( \40812 , \40437 , \40439 );
and \U$32329 ( \40813 , \40436 , \40439 );
or \U$32330 ( \40814 , \40811 , \40812 , \40813 );
and \U$32331 ( \40815 , \40395 , \40406 );
and \U$32332 ( \40816 , \40406 , \40421 );
and \U$32333 ( \40817 , \40395 , \40421 );
or \U$32334 ( \40818 , \40815 , \40816 , \40817 );
xor \U$32335 ( \40819 , \40814 , \40818 );
and \U$32336 ( \40820 , \30802 , \27397 );
and \U$32337 ( \40821 , \32054 , \26807 );
nor \U$32338 ( \40822 , \40820 , \40821 );
xnor \U$32339 ( \40823 , \40822 , \27295 );
not \U$32340 ( \40824 , \40823 );
and \U$32341 ( \40825 , \29084 , \29070 );
and \U$32342 ( \40826 , \30268 , \28526 );
nor \U$32343 ( \40827 , \40825 , \40826 );
xnor \U$32344 ( \40828 , \40827 , \29076 );
xor \U$32345 ( \40829 , \40824 , \40828 );
and \U$32346 ( \40830 , \25272 , \32802 );
xor \U$32347 ( \40831 , \40829 , \40830 );
xor \U$32348 ( \40832 , \40819 , \40831 );
xor \U$32349 ( \40833 , \40810 , \40832 );
and \U$32350 ( \40834 , \40391 , \40422 );
and \U$32351 ( \40835 , \40422 , \40441 );
and \U$32352 ( \40836 , \40391 , \40441 );
or \U$32353 ( \40837 , \40834 , \40835 , \40836 );
xor \U$32354 ( \40838 , \40833 , \40837 );
and \U$32355 ( \40839 , \40442 , \40446 );
and \U$32356 ( \40840 , \40447 , \40450 );
or \U$32357 ( \40841 , \40839 , \40840 );
xor \U$32358 ( \40842 , \40838 , \40841 );
buf g9b6c ( \40843_nG9b6c , \40842 );
and \U$32359 ( \40844 , \10704 , \40843_nG9b6c );
or \U$32360 ( \40845 , \40782 , \40844 );
xor \U$32361 ( \40846 , \10703 , \40845 );
buf \U$32362 ( \40847 , \40846 );
buf \U$32364 ( \40848 , \40847 );
xor \U$32365 ( \40849 , \40781 , \40848 );
buf \U$32366 ( \40850 , \40849 );
xor \U$32367 ( \40851 , \40768 , \40850 );
and \U$32368 ( \40852 , \40310 , \40316 );
and \U$32369 ( \40853 , \40310 , \40323 );
and \U$32370 ( \40854 , \40316 , \40323 );
or \U$32371 ( \40855 , \40852 , \40853 , \40854 );
buf \U$32372 ( \40856 , \40855 );
and \U$32373 ( \40857 , \14631 , \37974_nG9b87 );
and \U$32374 ( \40858 , \14628 , \38337_nG9b84 );
or \U$32375 ( \40859 , \40857 , \40858 );
xor \U$32376 ( \40860 , \14627 , \40859 );
buf \U$32377 ( \40861 , \40860 );
buf \U$32379 ( \40862 , \40861 );
xor \U$32380 ( \40863 , \40856 , \40862 );
and \U$32381 ( \40864 , \10421 , \39963_nG9b75 );
and \U$32382 ( \40865 , \10418 , \40204_nG9b72 );
or \U$32383 ( \40866 , \40864 , \40865 );
xor \U$32384 ( \40867 , \10417 , \40866 );
buf \U$32385 ( \40868 , \40867 );
buf \U$32387 ( \40869 , \40868 );
xor \U$32388 ( \40870 , \40863 , \40869 );
buf \U$32389 ( \40871 , \40870 );
xor \U$32390 ( \40872 , \40851 , \40871 );
buf \U$32391 ( \40873 , \40872 );
xor \U$32392 ( \40874 , \40763 , \40873 );
buf \U$32393 ( \40875 , \40874 );
xor \U$32394 ( \40876 , \40752 , \40875 );
and \U$32395 ( \40877 , \40596 , \40876 );
and \U$32397 ( \40878 , \40590 , \40595 );
or \U$32399 ( \40879 , 1'b0 , \40878 , 1'b0 );
xor \U$32400 ( \40880 , \40877 , \40879 );
and \U$32402 ( \40881 , \40583 , \40589 );
and \U$32403 ( \40882 , \40585 , \40589 );
or \U$32404 ( \40883 , 1'b0 , \40881 , \40882 );
xor \U$32405 ( \40884 , \40880 , \40883 );
xor \U$32412 ( \40885 , \40884 , 1'b0 );
and \U$32413 ( \40886 , \40746 , \40751 );
and \U$32414 ( \40887 , \40746 , \40875 );
and \U$32415 ( \40888 , \40751 , \40875 );
or \U$32416 ( \40889 , \40886 , \40887 , \40888 );
xor \U$32417 ( \40890 , \40885 , \40889 );
and \U$32418 ( \40891 , \40757 , \40762 );
and \U$32419 ( \40892 , \40757 , \40873 );
and \U$32420 ( \40893 , \40762 , \40873 );
or \U$32421 ( \40894 , \40891 , \40892 , \40893 );
buf \U$32422 ( \40895 , \40894 );
and \U$32423 ( \40896 , \40768 , \40850 );
and \U$32424 ( \40897 , \40768 , \40871 );
and \U$32425 ( \40898 , \40850 , \40871 );
or \U$32426 ( \40899 , \40896 , \40897 , \40898 );
buf \U$32427 ( \40900 , \40899 );
and \U$32428 ( \40901 , \17297 , \36986_nG9b90 );
and \U$32429 ( \40902 , \17294 , \37250_nG9b8d );
or \U$32430 ( \40903 , \40901 , \40902 );
xor \U$32431 ( \40904 , \17293 , \40903 );
buf \U$32432 ( \40905 , \40904 );
buf \U$32434 ( \40906 , \40905 );
and \U$32435 ( \40907 , \15940 , \37607_nG9b8a );
and \U$32436 ( \40908 , \15937 , \37974_nG9b87 );
or \U$32437 ( \40909 , \40907 , \40908 );
xor \U$32438 ( \40910 , \15936 , \40909 );
buf \U$32439 ( \40911 , \40910 );
buf \U$32441 ( \40912 , \40911 );
xor \U$32442 ( \40913 , \40906 , \40912 );
and \U$32443 ( \40914 , \12157 , \39591_nG9b78 );
and \U$32444 ( \40915 , \12154 , \39963_nG9b75 );
or \U$32445 ( \40916 , \40914 , \40915 );
xor \U$32446 ( \40917 , \12153 , \40916 );
buf \U$32447 ( \40918 , \40917 );
buf \U$32449 ( \40919 , \40918 );
xor \U$32450 ( \40920 , \40913 , \40919 );
buf \U$32451 ( \40921 , \40920 );
and \U$32452 ( \40922 , \23201 , \34041_nG9ba8 );
and \U$32453 ( \40923 , \23198 , \34294_nG9ba5 );
or \U$32454 ( \40924 , \40922 , \40923 );
xor \U$32455 ( \40925 , \23197 , \40924 );
buf \U$32456 ( \40926 , \40925 );
buf \U$32458 ( \40927 , \40926 );
and \U$32459 ( \40928 , \21658 , \34643_nG9ba2 );
and \U$32460 ( \40929 , \21655 , \35094_nG9b9f );
or \U$32461 ( \40930 , \40928 , \40929 );
xor \U$32462 ( \40931 , \21654 , \40930 );
buf \U$32463 ( \40932 , \40931 );
buf \U$32465 ( \40933 , \40932 );
xor \U$32466 ( \40934 , \40927 , \40933 );
and \U$32467 ( \40935 , \20155 , \35570_nG9b9c );
and \U$32468 ( \40936 , \20152 , \35801_nG9b99 );
or \U$32469 ( \40937 , \40935 , \40936 );
xor \U$32470 ( \40938 , \20151 , \40937 );
buf \U$32471 ( \40939 , \40938 );
buf \U$32473 ( \40940 , \40939 );
xor \U$32474 ( \40941 , \40934 , \40940 );
buf \U$32475 ( \40942 , \40941 );
xor \U$32476 ( \40943 , \40921 , \40942 );
and \U$32477 ( \40944 , \40612 , \40618 );
and \U$32478 ( \40945 , \40612 , \40625 );
and \U$32479 ( \40946 , \40618 , \40625 );
or \U$32480 ( \40947 , \40944 , \40945 , \40946 );
buf \U$32481 ( \40948 , \40947 );
xor \U$32482 ( \40949 , \40943 , \40948 );
buf \U$32483 ( \40950 , \40949 );
xor \U$32484 ( \40951 , \40900 , \40950 );
and \U$32485 ( \40952 , \40627 , \40648 );
and \U$32486 ( \40953 , \40627 , \40654 );
and \U$32487 ( \40954 , \40648 , \40654 );
or \U$32488 ( \40955 , \40952 , \40953 , \40954 );
buf \U$32489 ( \40956 , \40955 );
xor \U$32490 ( \40957 , \40951 , \40956 );
buf \U$32491 ( \40958 , \40957 );
xor \U$32492 ( \40959 , \40895 , \40958 );
and \U$32493 ( \40960 , \40606 , \40656 );
and \U$32494 ( \40961 , \40606 , \40662 );
and \U$32495 ( \40962 , \40656 , \40662 );
or \U$32496 ( \40963 , \40960 , \40961 , \40962 );
buf \U$32497 ( \40964 , \40963 );
xor \U$32498 ( \40965 , \40959 , \40964 );
buf \U$32499 ( \40966 , \40965 );
and \U$32500 ( \40967 , \40601 , \40664 );
and \U$32501 ( \40968 , \40601 , \40744 );
and \U$32502 ( \40969 , \40664 , \40744 );
or \U$32503 ( \40970 , \40967 , \40968 , \40969 );
buf \U$32504 ( \40971 , \40970 );
xor \U$32505 ( \40972 , \40966 , \40971 );
and \U$32506 ( \40973 , \40725 , \40731 );
and \U$32507 ( \40974 , \40725 , \40738 );
and \U$32508 ( \40975 , \40731 , \40738 );
or \U$32509 ( \40976 , \40973 , \40974 , \40975 );
buf \U$32510 ( \40977 , \40976 );
and \U$32511 ( \40978 , \14631 , \38337_nG9b84 );
and \U$32512 ( \40979 , \14628 , \38663_nG9b81 );
or \U$32513 ( \40980 , \40978 , \40979 );
xor \U$32514 ( \40981 , \14627 , \40980 );
buf \U$32515 ( \40982 , \40981 );
buf \U$32517 ( \40983 , \40982 );
xor \U$32518 ( \40984 , \40977 , \40983 );
and \U$32519 ( \40985 , \10707 , \40843_nG9b6c );
and \U$32520 ( \40986 , \40790 , \40794 );
and \U$32521 ( \40987 , \40794 , \40808 );
and \U$32522 ( \40988 , \40790 , \40808 );
or \U$32523 ( \40989 , \40986 , \40987 , \40988 );
and \U$32524 ( \40990 , \40814 , \40818 );
and \U$32525 ( \40991 , \40818 , \40831 );
and \U$32526 ( \40992 , \40814 , \40831 );
or \U$32527 ( \40993 , \40990 , \40991 , \40992 );
xor \U$32528 ( \40994 , \40989 , \40993 );
and \U$32529 ( \40995 , \40824 , \40828 );
and \U$32530 ( \40996 , \40828 , \40830 );
and \U$32531 ( \40997 , \40824 , \40830 );
or \U$32532 ( \40998 , \40995 , \40996 , \40997 );
not \U$32533 ( \40999 , \25773 );
and \U$32534 ( \41000 , \32054 , \27397 );
and \U$32535 ( \41001 , \32794 , \26807 );
nor \U$32536 ( \41002 , \41000 , \41001 );
xnor \U$32537 ( \41003 , \41002 , \27295 );
xor \U$32538 ( \41004 , \40999 , \41003 );
and \U$32539 ( \41005 , \28534 , \30823 );
and \U$32540 ( \41006 , \29084 , \30246 );
nor \U$32541 ( \41007 , \41005 , \41006 );
xnor \U$32542 ( \41008 , \41007 , \30813 );
xor \U$32543 ( \41009 , \41004 , \41008 );
xor \U$32544 ( \41010 , \40998 , \41009 );
and \U$32545 ( \41011 , \40798 , \40802 );
and \U$32546 ( \41012 , \40802 , \40807 );
and \U$32547 ( \41013 , \40798 , \40807 );
or \U$32548 ( \41014 , \41011 , \41012 , \41013 );
buf \U$32549 ( \41015 , \40823 );
xor \U$32550 ( \41016 , \41014 , \41015 );
and \U$32551 ( \41017 , \30268 , \29070 );
and \U$32552 ( \41018 , \30802 , \28526 );
nor \U$32553 ( \41019 , \41017 , \41018 );
xnor \U$32554 ( \41020 , \41019 , \29076 );
and \U$32555 ( \41021 , \26829 , \32854 );
and \U$32556 ( \41022 , \27313 , \32067 );
nor \U$32557 ( \41023 , \41021 , \41022 );
xnor \U$32558 ( \41024 , \41023 , \32805 );
xor \U$32559 ( \41025 , \41020 , \41024 );
and \U$32560 ( \41026 , \25815 , \32802 );
xor \U$32561 ( \41027 , \41025 , \41026 );
xor \U$32562 ( \41028 , \41016 , \41027 );
xor \U$32563 ( \41029 , \41010 , \41028 );
xor \U$32564 ( \41030 , \40994 , \41029 );
and \U$32565 ( \41031 , \40786 , \40809 );
and \U$32566 ( \41032 , \40809 , \40832 );
and \U$32567 ( \41033 , \40786 , \40832 );
or \U$32568 ( \41034 , \41031 , \41032 , \41033 );
xor \U$32569 ( \41035 , \41030 , \41034 );
and \U$32570 ( \41036 , \40833 , \40837 );
and \U$32571 ( \41037 , \40838 , \40841 );
or \U$32572 ( \41038 , \41036 , \41037 );
xor \U$32573 ( \41039 , \41035 , \41038 );
buf g9b69 ( \41040_nG9b69 , \41039 );
and \U$32574 ( \41041 , \10704 , \41040_nG9b69 );
or \U$32575 ( \41042 , \40985 , \41041 );
xor \U$32576 ( \41043 , \10703 , \41042 );
buf \U$32577 ( \41044 , \41043 );
buf \U$32579 ( \41045 , \41044 );
xor \U$32580 ( \41046 , \40984 , \41045 );
buf \U$32581 ( \41047 , \41046 );
and \U$32582 ( \41048 , \40713 , \40718 );
and \U$32583 ( \41049 , \40713 , \40740 );
and \U$32584 ( \41050 , \40718 , \40740 );
or \U$32585 ( \41051 , \41048 , \41049 , \41050 );
buf \U$32586 ( \41052 , \41051 );
xor \U$32587 ( \41053 , \41047 , \41052 );
and \U$32588 ( \41054 , \18702 , \36172_nG9b96 );
and \U$32589 ( \41055 , \18699 , \36589_nG9b93 );
or \U$32590 ( \41056 , \41054 , \41055 );
xor \U$32591 ( \41057 , \18698 , \41056 );
buf \U$32592 ( \41058 , \41057 );
buf \U$32594 ( \41059 , \41058 );
and \U$32595 ( \41060 , \13370 , \38968_nG9b7e );
and \U$32596 ( \41061 , \13367 , \39334_nG9b7b );
or \U$32597 ( \41062 , \41060 , \41061 );
xor \U$32598 ( \41063 , \13366 , \41062 );
buf \U$32599 ( \41064 , \41063 );
buf \U$32601 ( \41065 , \41064 );
xor \U$32602 ( \41066 , \41059 , \41065 );
and \U$32603 ( \41067 , \10421 , \40204_nG9b72 );
and \U$32604 ( \41068 , \10418 , \40452_nG9b6f );
or \U$32605 ( \41069 , \41067 , \41068 );
xor \U$32606 ( \41070 , \10417 , \41069 );
buf \U$32607 ( \41071 , \41070 );
buf \U$32609 ( \41072 , \41071 );
xor \U$32610 ( \41073 , \41066 , \41072 );
buf \U$32611 ( \41074 , \41073 );
xor \U$32612 ( \41075 , \41053 , \41074 );
buf \U$32613 ( \41076 , \41075 );
and \U$32614 ( \41077 , \40702 , \40707 );
and \U$32615 ( \41078 , \40702 , \40742 );
and \U$32616 ( \41079 , \40707 , \40742 );
or \U$32617 ( \41080 , \41077 , \41078 , \41079 );
buf \U$32618 ( \41081 , \41080 );
xor \U$32619 ( \41082 , \41076 , \41081 );
and \U$32620 ( \41083 , \40774 , \40780 );
and \U$32621 ( \41084 , \40774 , \40848 );
and \U$32622 ( \41085 , \40780 , \40848 );
or \U$32623 ( \41086 , \41083 , \41084 , \41085 );
buf \U$32624 ( \41087 , \41086 );
and \U$32625 ( \41088 , \40856 , \40862 );
and \U$32626 ( \41089 , \40856 , \40869 );
and \U$32627 ( \41090 , \40862 , \40869 );
or \U$32628 ( \41091 , \41088 , \41089 , \41090 );
buf \U$32629 ( \41092 , \41091 );
xor \U$32630 ( \41093 , \41087 , \41092 );
and \U$32632 ( \41094 , \32916 , \25860_nG9bc9 );
or \U$32633 ( \41095 , 1'b0 , \41094 );
xor \U$32634 ( \41096 , 1'b0 , \41095 );
buf \U$32635 ( \41097 , \41096 );
buf \U$32637 ( \41098 , \41097 );
and \U$32638 ( \41099 , \31636 , \26887_nG9bc6 );
and \U$32639 ( \41100 , \31633 , \27416_nG9bc3 );
or \U$32640 ( \41101 , \41099 , \41100 );
xor \U$32641 ( \41102 , \31632 , \41101 );
buf \U$32642 ( \41103 , \41102 );
buf \U$32644 ( \41104 , \41103 );
xor \U$32645 ( \41105 , \41098 , \41104 );
buf \U$32646 ( \41106 , \41105 );
and \U$32647 ( \41107 , \26431 , \32179_nG9bb4 );
and \U$32648 ( \41108 , \26428 , \32888_nG9bb1 );
or \U$32649 ( \41109 , \41107 , \41108 );
xor \U$32650 ( \41110 , \26427 , \41109 );
buf \U$32651 ( \41111 , \41110 );
buf \U$32653 ( \41112 , \41111 );
xor \U$32654 ( \41113 , \41106 , \41112 );
and \U$32655 ( \41114 , \24792 , \33181_nG9bae );
and \U$32656 ( \41115 , \24789 , \33613_nG9bab );
or \U$32657 ( \41116 , \41114 , \41115 );
xor \U$32658 ( \41117 , \24788 , \41116 );
buf \U$32659 ( \41118 , \41117 );
buf \U$32661 ( \41119 , \41118 );
xor \U$32662 ( \41120 , \41113 , \41119 );
buf \U$32663 ( \41121 , \41120 );
xor \U$32664 ( \41122 , \41093 , \41121 );
buf \U$32665 ( \41123 , \41122 );
and \U$32666 ( \41124 , \40670 , \40675 );
and \U$32667 ( \41125 , \40670 , \40700 );
and \U$32668 ( \41126 , \40675 , \40700 );
or \U$32669 ( \41127 , \41124 , \41125 , \41126 );
buf \U$32670 ( \41128 , \41127 );
xor \U$32671 ( \41129 , \41123 , \41128 );
and \U$32672 ( \41130 , \40633 , \40639 );
and \U$32673 ( \41131 , \40633 , \40646 );
and \U$32674 ( \41132 , \40639 , \40646 );
or \U$32675 ( \41133 , \41130 , \41131 , \41132 );
buf \U$32676 ( \41134 , \41133 );
and \U$32677 ( \41135 , \40689 , \40691 );
and \U$32678 ( \41136 , \40689 , \40698 );
and \U$32679 ( \41137 , \40691 , \40698 );
or \U$32680 ( \41138 , \41135 , \41136 , \41137 );
buf \U$32681 ( \41139 , \41138 );
xor \U$32682 ( \41140 , \41134 , \41139 );
and \U$32683 ( \41141 , \40681 , \40687 );
buf \U$32684 ( \41142 , \41141 );
and \U$32685 ( \41143 , \29853 , \28602_nG9bc0 );
and \U$32686 ( \41144 , \29850 , \29179_nG9bbd );
or \U$32687 ( \41145 , \41143 , \41144 );
xor \U$32688 ( \41146 , \29849 , \41145 );
buf \U$32689 ( \41147 , \41146 );
buf \U$32691 ( \41148 , \41147 );
xor \U$32692 ( \41149 , \41142 , \41148 );
and \U$32693 ( \41150 , \28118 , \30366_nG9bba );
and \U$32694 ( \41151 , \28115 , \30940_nG9bb7 );
or \U$32695 ( \41152 , \41150 , \41151 );
xor \U$32696 ( \41153 , \28114 , \41152 );
buf \U$32697 ( \41154 , \41153 );
buf \U$32699 ( \41155 , \41154 );
xor \U$32700 ( \41156 , \41149 , \41155 );
buf \U$32701 ( \41157 , \41156 );
xor \U$32702 ( \41158 , \41140 , \41157 );
buf \U$32703 ( \41159 , \41158 );
xor \U$32704 ( \41160 , \41129 , \41159 );
buf \U$32705 ( \41161 , \41160 );
xor \U$32706 ( \41162 , \41082 , \41161 );
buf \U$32707 ( \41163 , \41162 );
xor \U$32708 ( \41164 , \40972 , \41163 );
and \U$32709 ( \41165 , \40890 , \41164 );
and \U$32711 ( \41166 , \40884 , \40889 );
or \U$32713 ( \41167 , 1'b0 , \41166 , 1'b0 );
xor \U$32714 ( \41168 , \41165 , \41167 );
and \U$32716 ( \41169 , \40877 , \40883 );
and \U$32717 ( \41170 , \40879 , \40883 );
or \U$32718 ( \41171 , 1'b0 , \41169 , \41170 );
xor \U$32719 ( \41172 , \41168 , \41171 );
xor \U$32726 ( \41173 , \41172 , 1'b0 );
and \U$32727 ( \41174 , \40966 , \40971 );
and \U$32728 ( \41175 , \40966 , \41163 );
and \U$32729 ( \41176 , \40971 , \41163 );
or \U$32730 ( \41177 , \41174 , \41175 , \41176 );
xor \U$32731 ( \41178 , \41173 , \41177 );
and \U$32732 ( \41179 , \41076 , \41081 );
and \U$32733 ( \41180 , \41076 , \41161 );
and \U$32734 ( \41181 , \41081 , \41161 );
or \U$32735 ( \41182 , \41179 , \41180 , \41181 );
buf \U$32736 ( \41183 , \41182 );
and \U$32737 ( \41184 , \41047 , \41052 );
and \U$32738 ( \41185 , \41047 , \41074 );
and \U$32739 ( \41186 , \41052 , \41074 );
or \U$32740 ( \41187 , \41184 , \41185 , \41186 );
buf \U$32741 ( \41188 , \41187 );
and \U$32742 ( \41189 , \18702 , \36589_nG9b93 );
and \U$32743 ( \41190 , \18699 , \36986_nG9b90 );
or \U$32744 ( \41191 , \41189 , \41190 );
xor \U$32745 ( \41192 , \18698 , \41191 );
buf \U$32746 ( \41193 , \41192 );
buf \U$32748 ( \41194 , \41193 );
and \U$32749 ( \41195 , \13370 , \39334_nG9b7b );
and \U$32750 ( \41196 , \13367 , \39591_nG9b78 );
or \U$32751 ( \41197 , \41195 , \41196 );
xor \U$32752 ( \41198 , \13366 , \41197 );
buf \U$32753 ( \41199 , \41198 );
buf \U$32755 ( \41200 , \41199 );
xor \U$32756 ( \41201 , \41194 , \41200 );
and \U$32757 ( \41202 , \10421 , \40452_nG9b6f );
and \U$32758 ( \41203 , \10418 , \40843_nG9b6c );
or \U$32759 ( \41204 , \41202 , \41203 );
xor \U$32760 ( \41205 , \10417 , \41204 );
buf \U$32761 ( \41206 , \41205 );
buf \U$32763 ( \41207 , \41206 );
xor \U$32764 ( \41208 , \41201 , \41207 );
buf \U$32765 ( \41209 , \41208 );
and \U$32766 ( \41210 , \40906 , \40912 );
and \U$32767 ( \41211 , \40906 , \40919 );
and \U$32768 ( \41212 , \40912 , \40919 );
or \U$32769 ( \41213 , \41210 , \41211 , \41212 );
buf \U$32770 ( \41214 , \41213 );
xor \U$32771 ( \41215 , \41209 , \41214 );
and \U$32772 ( \41216 , \23201 , \34294_nG9ba5 );
and \U$32773 ( \41217 , \23198 , \34643_nG9ba2 );
or \U$32774 ( \41218 , \41216 , \41217 );
xor \U$32775 ( \41219 , \23197 , \41218 );
buf \U$32776 ( \41220 , \41219 );
buf \U$32778 ( \41221 , \41220 );
and \U$32779 ( \41222 , \21658 , \35094_nG9b9f );
and \U$32780 ( \41223 , \21655 , \35570_nG9b9c );
or \U$32781 ( \41224 , \41222 , \41223 );
xor \U$32782 ( \41225 , \21654 , \41224 );
buf \U$32783 ( \41226 , \41225 );
buf \U$32785 ( \41227 , \41226 );
xor \U$32786 ( \41228 , \41221 , \41227 );
and \U$32787 ( \41229 , \20155 , \35801_nG9b99 );
and \U$32788 ( \41230 , \20152 , \36172_nG9b96 );
or \U$32789 ( \41231 , \41229 , \41230 );
xor \U$32790 ( \41232 , \20151 , \41231 );
buf \U$32791 ( \41233 , \41232 );
buf \U$32793 ( \41234 , \41233 );
xor \U$32794 ( \41235 , \41228 , \41234 );
buf \U$32795 ( \41236 , \41235 );
xor \U$32796 ( \41237 , \41215 , \41236 );
buf \U$32797 ( \41238 , \41237 );
xor \U$32798 ( \41239 , \41188 , \41238 );
and \U$32799 ( \41240 , \40921 , \40942 );
and \U$32800 ( \41241 , \40921 , \40948 );
and \U$32801 ( \41242 , \40942 , \40948 );
or \U$32802 ( \41243 , \41240 , \41241 , \41242 );
buf \U$32803 ( \41244 , \41243 );
xor \U$32804 ( \41245 , \41239 , \41244 );
buf \U$32805 ( \41246 , \41245 );
xor \U$32806 ( \41247 , \41183 , \41246 );
and \U$32807 ( \41248 , \40900 , \40950 );
and \U$32808 ( \41249 , \40900 , \40956 );
and \U$32809 ( \41250 , \40950 , \40956 );
or \U$32810 ( \41251 , \41248 , \41249 , \41250 );
buf \U$32811 ( \41252 , \41251 );
xor \U$32812 ( \41253 , \41247 , \41252 );
buf \U$32813 ( \41254 , \41253 );
and \U$32814 ( \41255 , \40895 , \40958 );
and \U$32815 ( \41256 , \40895 , \40964 );
and \U$32816 ( \41257 , \40958 , \40964 );
or \U$32817 ( \41258 , \41255 , \41256 , \41257 );
buf \U$32818 ( \41259 , \41258 );
xor \U$32819 ( \41260 , \41254 , \41259 );
and \U$32820 ( \41261 , \41123 , \41128 );
and \U$32821 ( \41262 , \41123 , \41159 );
and \U$32822 ( \41263 , \41128 , \41159 );
or \U$32823 ( \41264 , \41261 , \41262 , \41263 );
buf \U$32824 ( \41265 , \41264 );
and \U$32825 ( \41266 , \41098 , \41104 );
buf \U$32826 ( \41267 , \41266 );
and \U$32827 ( \41268 , \29853 , \29179_nG9bbd );
and \U$32828 ( \41269 , \29850 , \30366_nG9bba );
or \U$32829 ( \41270 , \41268 , \41269 );
xor \U$32830 ( \41271 , \29849 , \41270 );
buf \U$32831 ( \41272 , \41271 );
buf \U$32833 ( \41273 , \41272 );
xor \U$32834 ( \41274 , \41267 , \41273 );
and \U$32835 ( \41275 , \28118 , \30940_nG9bb7 );
and \U$32836 ( \41276 , \28115 , \32179_nG9bb4 );
or \U$32837 ( \41277 , \41275 , \41276 );
xor \U$32838 ( \41278 , \28114 , \41277 );
buf \U$32839 ( \41279 , \41278 );
buf \U$32841 ( \41280 , \41279 );
xor \U$32842 ( \41281 , \41274 , \41280 );
buf \U$32843 ( \41282 , \41281 );
and \U$32844 ( \41283 , \40927 , \40933 );
and \U$32845 ( \41284 , \40927 , \40940 );
and \U$32846 ( \41285 , \40933 , \40940 );
or \U$32847 ( \41286 , \41283 , \41284 , \41285 );
buf \U$32848 ( \41287 , \41286 );
xor \U$32849 ( \41288 , \41282 , \41287 );
and \U$32850 ( \41289 , \41106 , \41112 );
and \U$32851 ( \41290 , \41106 , \41119 );
and \U$32852 ( \41291 , \41112 , \41119 );
or \U$32853 ( \41292 , \41289 , \41290 , \41291 );
buf \U$32854 ( \41293 , \41292 );
xor \U$32855 ( \41294 , \41288 , \41293 );
buf \U$32856 ( \41295 , \41294 );
and \U$32857 ( \41296 , \41142 , \41148 );
and \U$32858 ( \41297 , \41142 , \41155 );
and \U$32859 ( \41298 , \41148 , \41155 );
or \U$32860 ( \41299 , \41296 , \41297 , \41298 );
buf \U$32861 ( \41300 , \41299 );
and \U$32862 ( \41301 , \17297 , \37250_nG9b8d );
and \U$32863 ( \41302 , \17294 , \37607_nG9b8a );
or \U$32864 ( \41303 , \41301 , \41302 );
xor \U$32865 ( \41304 , \17293 , \41303 );
buf \U$32866 ( \41305 , \41304 );
buf \U$32868 ( \41306 , \41305 );
xor \U$32869 ( \41307 , \41300 , \41306 );
and \U$32870 ( \41308 , \12157 , \39963_nG9b75 );
and \U$32871 ( \41309 , \12154 , \40204_nG9b72 );
or \U$32872 ( \41310 , \41308 , \41309 );
xor \U$32873 ( \41311 , \12153 , \41310 );
buf \U$32874 ( \41312 , \41311 );
buf \U$32876 ( \41313 , \41312 );
xor \U$32877 ( \41314 , \41307 , \41313 );
buf \U$32878 ( \41315 , \41314 );
xor \U$32879 ( \41316 , \41295 , \41315 );
and \U$32880 ( \41317 , \15940 , \37974_nG9b87 );
and \U$32881 ( \41318 , \15937 , \38337_nG9b84 );
or \U$32882 ( \41319 , \41317 , \41318 );
xor \U$32883 ( \41320 , \15936 , \41319 );
buf \U$32884 ( \41321 , \41320 );
buf \U$32886 ( \41322 , \41321 );
and \U$32887 ( \41323 , \14631 , \38663_nG9b81 );
and \U$32888 ( \41324 , \14628 , \38968_nG9b7e );
or \U$32889 ( \41325 , \41323 , \41324 );
xor \U$32890 ( \41326 , \14627 , \41325 );
buf \U$32891 ( \41327 , \41326 );
buf \U$32893 ( \41328 , \41327 );
xor \U$32894 ( \41329 , \41322 , \41328 );
and \U$32895 ( \41330 , \10707 , \41040_nG9b69 );
and \U$32896 ( \41331 , \41014 , \41015 );
and \U$32897 ( \41332 , \41015 , \41027 );
and \U$32898 ( \41333 , \41014 , \41027 );
or \U$32899 ( \41334 , \41331 , \41332 , \41333 );
and \U$32900 ( \41335 , \40998 , \41009 );
and \U$32901 ( \41336 , \41009 , \41028 );
and \U$32902 ( \41337 , \40998 , \41028 );
or \U$32903 ( \41338 , \41335 , \41336 , \41337 );
xor \U$32904 ( \41339 , \41334 , \41338 );
and \U$32905 ( \41340 , \40999 , \41003 );
and \U$32906 ( \41341 , \41003 , \41008 );
and \U$32907 ( \41342 , \40999 , \41008 );
or \U$32908 ( \41343 , \41340 , \41341 , \41342 );
and \U$32909 ( \41344 , \32794 , \27397 );
not \U$32910 ( \41345 , \41344 );
xnor \U$32911 ( \41346 , \41345 , \27295 );
and \U$32912 ( \41347 , \27313 , \32854 );
and \U$32913 ( \41348 , \28534 , \32067 );
nor \U$32914 ( \41349 , \41347 , \41348 );
xnor \U$32915 ( \41350 , \41349 , \32805 );
xor \U$32916 ( \41351 , \41346 , \41350 );
and \U$32917 ( \41352 , \26829 , \32802 );
xor \U$32918 ( \41353 , \41351 , \41352 );
xor \U$32919 ( \41354 , \41343 , \41353 );
and \U$32920 ( \41355 , \41020 , \41024 );
and \U$32921 ( \41356 , \41024 , \41026 );
and \U$32922 ( \41357 , \41020 , \41026 );
or \U$32923 ( \41358 , \41355 , \41356 , \41357 );
and \U$32924 ( \41359 , \30802 , \29070 );
and \U$32925 ( \41360 , \32054 , \28526 );
nor \U$32926 ( \41361 , \41359 , \41360 );
xnor \U$32927 ( \41362 , \41361 , \29076 );
not \U$32928 ( \41363 , \41362 );
xor \U$32929 ( \41364 , \41358 , \41363 );
and \U$32930 ( \41365 , \29084 , \30823 );
and \U$32931 ( \41366 , \30268 , \30246 );
nor \U$32932 ( \41367 , \41365 , \41366 );
xnor \U$32933 ( \41368 , \41367 , \30813 );
xor \U$32934 ( \41369 , \41364 , \41368 );
xor \U$32935 ( \41370 , \41354 , \41369 );
xor \U$32936 ( \41371 , \41339 , \41370 );
and \U$32937 ( \41372 , \40989 , \40993 );
and \U$32938 ( \41373 , \40993 , \41029 );
and \U$32939 ( \41374 , \40989 , \41029 );
or \U$32940 ( \41375 , \41372 , \41373 , \41374 );
xor \U$32941 ( \41376 , \41371 , \41375 );
and \U$32942 ( \41377 , \41030 , \41034 );
and \U$32943 ( \41378 , \41035 , \41038 );
or \U$32944 ( \41379 , \41377 , \41378 );
xor \U$32945 ( \41380 , \41376 , \41379 );
buf g9b66 ( \41381_nG9b66 , \41380 );
and \U$32946 ( \41382 , \10704 , \41381_nG9b66 );
or \U$32947 ( \41383 , \41330 , \41382 );
xor \U$32948 ( \41384 , \10703 , \41383 );
buf \U$32949 ( \41385 , \41384 );
buf \U$32951 ( \41386 , \41385 );
xor \U$32952 ( \41387 , \41329 , \41386 );
buf \U$32953 ( \41388 , \41387 );
xor \U$32954 ( \41389 , \41316 , \41388 );
buf \U$32955 ( \41390 , \41389 );
xor \U$32956 ( \41391 , \41265 , \41390 );
and \U$32957 ( \41392 , \41087 , \41092 );
and \U$32958 ( \41393 , \41087 , \41121 );
and \U$32959 ( \41394 , \41092 , \41121 );
or \U$32960 ( \41395 , \41392 , \41393 , \41394 );
buf \U$32961 ( \41396 , \41395 );
and \U$32962 ( \41397 , \41134 , \41139 );
and \U$32963 ( \41398 , \41134 , \41157 );
and \U$32964 ( \41399 , \41139 , \41157 );
or \U$32965 ( \41400 , \41397 , \41398 , \41399 );
buf \U$32966 ( \41401 , \41400 );
xor \U$32967 ( \41402 , \41396 , \41401 );
and \U$32968 ( \41403 , \40977 , \40983 );
and \U$32969 ( \41404 , \40977 , \41045 );
and \U$32970 ( \41405 , \40983 , \41045 );
or \U$32971 ( \41406 , \41403 , \41404 , \41405 );
buf \U$32972 ( \41407 , \41406 );
and \U$32973 ( \41408 , \41059 , \41065 );
and \U$32974 ( \41409 , \41059 , \41072 );
and \U$32975 ( \41410 , \41065 , \41072 );
or \U$32976 ( \41411 , \41408 , \41409 , \41410 );
buf \U$32977 ( \41412 , \41411 );
xor \U$32978 ( \41413 , \41407 , \41412 );
and \U$32980 ( \41414 , \32916 , \26887_nG9bc6 );
or \U$32981 ( \41415 , 1'b0 , \41414 );
xor \U$32982 ( \41416 , 1'b0 , \41415 );
buf \U$32983 ( \41417 , \41416 );
buf \U$32985 ( \41418 , \41417 );
and \U$32986 ( \41419 , \31636 , \27416_nG9bc3 );
and \U$32987 ( \41420 , \31633 , \28602_nG9bc0 );
or \U$32988 ( \41421 , \41419 , \41420 );
xor \U$32989 ( \41422 , \31632 , \41421 );
buf \U$32990 ( \41423 , \41422 );
buf \U$32992 ( \41424 , \41423 );
xor \U$32993 ( \41425 , \41418 , \41424 );
buf \U$32994 ( \41426 , \41425 );
and \U$32995 ( \41427 , \26431 , \32888_nG9bb1 );
and \U$32996 ( \41428 , \26428 , \33181_nG9bae );
or \U$32997 ( \41429 , \41427 , \41428 );
xor \U$32998 ( \41430 , \26427 , \41429 );
buf \U$32999 ( \41431 , \41430 );
buf \U$33001 ( \41432 , \41431 );
xor \U$33002 ( \41433 , \41426 , \41432 );
and \U$33003 ( \41434 , \24792 , \33613_nG9bab );
and \U$33004 ( \41435 , \24789 , \34041_nG9ba8 );
or \U$33005 ( \41436 , \41434 , \41435 );
xor \U$33006 ( \41437 , \24788 , \41436 );
buf \U$33007 ( \41438 , \41437 );
buf \U$33009 ( \41439 , \41438 );
xor \U$33010 ( \41440 , \41433 , \41439 );
buf \U$33011 ( \41441 , \41440 );
xor \U$33012 ( \41442 , \41413 , \41441 );
buf \U$33013 ( \41443 , \41442 );
xor \U$33014 ( \41444 , \41402 , \41443 );
buf \U$33015 ( \41445 , \41444 );
xor \U$33016 ( \41446 , \41391 , \41445 );
buf \U$33017 ( \41447 , \41446 );
xor \U$33018 ( \41448 , \41260 , \41447 );
and \U$33019 ( \41449 , \41178 , \41448 );
and \U$33021 ( \41450 , \41172 , \41177 );
or \U$33023 ( \41451 , 1'b0 , \41450 , 1'b0 );
xor \U$33024 ( \41452 , \41449 , \41451 );
and \U$33026 ( \41453 , \41165 , \41171 );
and \U$33027 ( \41454 , \41167 , \41171 );
or \U$33028 ( \41455 , 1'b0 , \41453 , \41454 );
xor \U$33029 ( \41456 , \41452 , \41455 );
xor \U$33036 ( \41457 , \41456 , 1'b0 );
and \U$33037 ( \41458 , \41254 , \41259 );
and \U$33038 ( \41459 , \41254 , \41447 );
and \U$33039 ( \41460 , \41259 , \41447 );
or \U$33040 ( \41461 , \41458 , \41459 , \41460 );
xor \U$33041 ( \41462 , \41457 , \41461 );
and \U$33042 ( \41463 , \41265 , \41390 );
and \U$33043 ( \41464 , \41265 , \41445 );
and \U$33044 ( \41465 , \41390 , \41445 );
or \U$33045 ( \41466 , \41463 , \41464 , \41465 );
buf \U$33046 ( \41467 , \41466 );
and \U$33047 ( \41468 , \41188 , \41238 );
and \U$33048 ( \41469 , \41188 , \41244 );
and \U$33049 ( \41470 , \41238 , \41244 );
or \U$33050 ( \41471 , \41468 , \41469 , \41470 );
buf \U$33051 ( \41472 , \41471 );
xor \U$33052 ( \41473 , \41467 , \41472 );
and \U$33053 ( \41474 , \41295 , \41315 );
and \U$33054 ( \41475 , \41295 , \41388 );
and \U$33055 ( \41476 , \41315 , \41388 );
or \U$33056 ( \41477 , \41474 , \41475 , \41476 );
buf \U$33057 ( \41478 , \41477 );
and \U$33058 ( \41479 , \15940 , \38337_nG9b84 );
and \U$33059 ( \41480 , \15937 , \38663_nG9b81 );
or \U$33060 ( \41481 , \41479 , \41480 );
xor \U$33061 ( \41482 , \15936 , \41481 );
buf \U$33062 ( \41483 , \41482 );
buf \U$33064 ( \41484 , \41483 );
and \U$33065 ( \41485 , \14631 , \38968_nG9b7e );
and \U$33066 ( \41486 , \14628 , \39334_nG9b7b );
or \U$33067 ( \41487 , \41485 , \41486 );
xor \U$33068 ( \41488 , \14627 , \41487 );
buf \U$33069 ( \41489 , \41488 );
buf \U$33071 ( \41490 , \41489 );
xor \U$33072 ( \41491 , \41484 , \41490 );
and \U$33073 ( \41492 , \10421 , \40843_nG9b6c );
and \U$33074 ( \41493 , \10418 , \41040_nG9b69 );
or \U$33075 ( \41494 , \41492 , \41493 );
xor \U$33076 ( \41495 , \10417 , \41494 );
buf \U$33077 ( \41496 , \41495 );
buf \U$33079 ( \41497 , \41496 );
xor \U$33080 ( \41498 , \41491 , \41497 );
buf \U$33081 ( \41499 , \41498 );
and \U$33082 ( \41500 , \41282 , \41287 );
and \U$33083 ( \41501 , \41282 , \41293 );
and \U$33084 ( \41502 , \41287 , \41293 );
or \U$33085 ( \41503 , \41500 , \41501 , \41502 );
buf \U$33086 ( \41504 , \41503 );
xor \U$33087 ( \41505 , \41499 , \41504 );
and \U$33088 ( \41506 , \41300 , \41306 );
and \U$33089 ( \41507 , \41300 , \41313 );
and \U$33090 ( \41508 , \41306 , \41313 );
or \U$33091 ( \41509 , \41506 , \41507 , \41508 );
buf \U$33092 ( \41510 , \41509 );
xor \U$33093 ( \41511 , \41505 , \41510 );
buf \U$33094 ( \41512 , \41511 );
xor \U$33095 ( \41513 , \41478 , \41512 );
and \U$33096 ( \41514 , \41209 , \41214 );
and \U$33097 ( \41515 , \41209 , \41236 );
and \U$33098 ( \41516 , \41214 , \41236 );
or \U$33099 ( \41517 , \41514 , \41515 , \41516 );
buf \U$33100 ( \41518 , \41517 );
xor \U$33101 ( \41519 , \41513 , \41518 );
buf \U$33102 ( \41520 , \41519 );
xor \U$33103 ( \41521 , \41473 , \41520 );
buf \U$33104 ( \41522 , \41521 );
and \U$33105 ( \41523 , \41183 , \41246 );
and \U$33106 ( \41524 , \41183 , \41252 );
and \U$33107 ( \41525 , \41246 , \41252 );
or \U$33108 ( \41526 , \41523 , \41524 , \41525 );
buf \U$33109 ( \41527 , \41526 );
xor \U$33110 ( \41528 , \41522 , \41527 );
and \U$33111 ( \41529 , \24792 , \34041_nG9ba8 );
and \U$33112 ( \41530 , \24789 , \34294_nG9ba5 );
or \U$33113 ( \41531 , \41529 , \41530 );
xor \U$33114 ( \41532 , \24788 , \41531 );
buf \U$33115 ( \41533 , \41532 );
buf \U$33117 ( \41534 , \41533 );
and \U$33118 ( \41535 , \21658 , \35570_nG9b9c );
and \U$33119 ( \41536 , \21655 , \35801_nG9b99 );
or \U$33120 ( \41537 , \41535 , \41536 );
xor \U$33121 ( \41538 , \21654 , \41537 );
buf \U$33122 ( \41539 , \41538 );
buf \U$33124 ( \41540 , \41539 );
xor \U$33125 ( \41541 , \41534 , \41540 );
and \U$33126 ( \41542 , \18702 , \36986_nG9b90 );
and \U$33127 ( \41543 , \18699 , \37250_nG9b8d );
or \U$33128 ( \41544 , \41542 , \41543 );
xor \U$33129 ( \41545 , \18698 , \41544 );
buf \U$33130 ( \41546 , \41545 );
buf \U$33132 ( \41547 , \41546 );
xor \U$33133 ( \41548 , \41541 , \41547 );
buf \U$33134 ( \41549 , \41548 );
and \U$33135 ( \41550 , \41194 , \41200 );
and \U$33136 ( \41551 , \41194 , \41207 );
and \U$33137 ( \41552 , \41200 , \41207 );
or \U$33138 ( \41553 , \41550 , \41551 , \41552 );
buf \U$33139 ( \41554 , \41553 );
xor \U$33140 ( \41555 , \41549 , \41554 );
and \U$33141 ( \41556 , \41322 , \41328 );
and \U$33142 ( \41557 , \41322 , \41386 );
and \U$33143 ( \41558 , \41328 , \41386 );
or \U$33144 ( \41559 , \41556 , \41557 , \41558 );
buf \U$33145 ( \41560 , \41559 );
xor \U$33146 ( \41561 , \41555 , \41560 );
buf \U$33147 ( \41562 , \41561 );
and \U$33148 ( \41563 , \41407 , \41412 );
and \U$33149 ( \41564 , \41407 , \41441 );
and \U$33150 ( \41565 , \41412 , \41441 );
or \U$33151 ( \41566 , \41563 , \41564 , \41565 );
buf \U$33152 ( \41567 , \41566 );
xor \U$33153 ( \41568 , \41562 , \41567 );
and \U$33154 ( \41569 , \41418 , \41424 );
buf \U$33155 ( \41570 , \41569 );
and \U$33156 ( \41571 , \31636 , \28602_nG9bc0 );
and \U$33157 ( \41572 , \31633 , \29179_nG9bbd );
or \U$33158 ( \41573 , \41571 , \41572 );
xor \U$33159 ( \41574 , \31632 , \41573 );
buf \U$33160 ( \41575 , \41574 );
buf \U$33162 ( \41576 , \41575 );
xor \U$33163 ( \41577 , \41570 , \41576 );
and \U$33164 ( \41578 , \26431 , \33181_nG9bae );
and \U$33165 ( \41579 , \26428 , \33613_nG9bab );
or \U$33166 ( \41580 , \41578 , \41579 );
xor \U$33167 ( \41581 , \26427 , \41580 );
buf \U$33168 ( \41582 , \41581 );
buf \U$33170 ( \41583 , \41582 );
xor \U$33171 ( \41584 , \41577 , \41583 );
buf \U$33172 ( \41585 , \41584 );
and \U$33173 ( \41586 , \41426 , \41432 );
and \U$33174 ( \41587 , \41426 , \41439 );
and \U$33175 ( \41588 , \41432 , \41439 );
or \U$33176 ( \41589 , \41586 , \41587 , \41588 );
buf \U$33177 ( \41590 , \41589 );
xor \U$33178 ( \41591 , \41585 , \41590 );
and \U$33179 ( \41592 , \41221 , \41227 );
and \U$33180 ( \41593 , \41221 , \41234 );
and \U$33181 ( \41594 , \41227 , \41234 );
or \U$33182 ( \41595 , \41592 , \41593 , \41594 );
buf \U$33183 ( \41596 , \41595 );
xor \U$33184 ( \41597 , \41591 , \41596 );
buf \U$33185 ( \41598 , \41597 );
xor \U$33186 ( \41599 , \41568 , \41598 );
buf \U$33187 ( \41600 , \41599 );
and \U$33188 ( \41601 , \41396 , \41401 );
and \U$33189 ( \41602 , \41396 , \41443 );
and \U$33190 ( \41603 , \41401 , \41443 );
or \U$33191 ( \41604 , \41601 , \41602 , \41603 );
buf \U$33192 ( \41605 , \41604 );
xor \U$33193 ( \41606 , \41600 , \41605 );
and \U$33194 ( \41607 , \41267 , \41273 );
and \U$33195 ( \41608 , \41267 , \41280 );
and \U$33196 ( \41609 , \41273 , \41280 );
or \U$33197 ( \41610 , \41607 , \41608 , \41609 );
buf \U$33198 ( \41611 , \41610 );
and \U$33199 ( \41612 , \17297 , \37607_nG9b8a );
and \U$33200 ( \41613 , \17294 , \37974_nG9b87 );
or \U$33201 ( \41614 , \41612 , \41613 );
xor \U$33202 ( \41615 , \17293 , \41614 );
buf \U$33203 ( \41616 , \41615 );
buf \U$33205 ( \41617 , \41616 );
xor \U$33206 ( \41618 , \41611 , \41617 );
and \U$33207 ( \41619 , \12157 , \40204_nG9b72 );
and \U$33208 ( \41620 , \12154 , \40452_nG9b6f );
or \U$33209 ( \41621 , \41619 , \41620 );
xor \U$33210 ( \41622 , \12153 , \41621 );
buf \U$33211 ( \41623 , \41622 );
buf \U$33213 ( \41624 , \41623 );
xor \U$33214 ( \41625 , \41618 , \41624 );
buf \U$33215 ( \41626 , \41625 );
and \U$33216 ( \41627 , \20155 , \36172_nG9b96 );
and \U$33217 ( \41628 , \20152 , \36589_nG9b93 );
or \U$33218 ( \41629 , \41627 , \41628 );
xor \U$33219 ( \41630 , \20151 , \41629 );
buf \U$33220 ( \41631 , \41630 );
buf \U$33222 ( \41632 , \41631 );
and \U$33223 ( \41633 , \13370 , \39591_nG9b78 );
and \U$33224 ( \41634 , \13367 , \39963_nG9b75 );
or \U$33225 ( \41635 , \41633 , \41634 );
xor \U$33226 ( \41636 , \13366 , \41635 );
buf \U$33227 ( \41637 , \41636 );
buf \U$33229 ( \41638 , \41637 );
xor \U$33230 ( \41639 , \41632 , \41638 );
and \U$33231 ( \41640 , \10707 , \41381_nG9b66 );
and \U$33232 ( \41641 , \41334 , \41338 );
and \U$33233 ( \41642 , \41338 , \41370 );
and \U$33234 ( \41643 , \41334 , \41370 );
or \U$33235 ( \41644 , \41641 , \41642 , \41643 );
and \U$33236 ( \41645 , \41358 , \41363 );
and \U$33237 ( \41646 , \41363 , \41368 );
and \U$33238 ( \41647 , \41358 , \41368 );
or \U$33239 ( \41648 , \41645 , \41646 , \41647 );
and \U$33240 ( \41649 , \41343 , \41353 );
and \U$33241 ( \41650 , \41353 , \41369 );
and \U$33242 ( \41651 , \41343 , \41369 );
or \U$33243 ( \41652 , \41649 , \41650 , \41651 );
xor \U$33244 ( \41653 , \41648 , \41652 );
and \U$33245 ( \41654 , \41346 , \41350 );
and \U$33246 ( \41655 , \41350 , \41352 );
and \U$33247 ( \41656 , \41346 , \41352 );
or \U$33248 ( \41657 , \41654 , \41655 , \41656 );
not \U$33249 ( \41658 , \27295 );
and \U$33250 ( \41659 , \32054 , \29070 );
and \U$33251 ( \41660 , \32794 , \28526 );
nor \U$33252 ( \41661 , \41659 , \41660 );
xnor \U$33253 ( \41662 , \41661 , \29076 );
xor \U$33254 ( \41663 , \41658 , \41662 );
and \U$33255 ( \41664 , \28534 , \32854 );
and \U$33256 ( \41665 , \29084 , \32067 );
nor \U$33257 ( \41666 , \41664 , \41665 );
xnor \U$33258 ( \41667 , \41666 , \32805 );
xor \U$33259 ( \41668 , \41663 , \41667 );
xor \U$33260 ( \41669 , \41657 , \41668 );
buf \U$33261 ( \41670 , \41362 );
and \U$33262 ( \41671 , \30268 , \30823 );
and \U$33263 ( \41672 , \30802 , \30246 );
nor \U$33264 ( \41673 , \41671 , \41672 );
xnor \U$33265 ( \41674 , \41673 , \30813 );
xor \U$33266 ( \41675 , \41670 , \41674 );
and \U$33267 ( \41676 , \27313 , \32802 );
xor \U$33268 ( \41677 , \41675 , \41676 );
xor \U$33269 ( \41678 , \41669 , \41677 );
xor \U$33270 ( \41679 , \41653 , \41678 );
xor \U$33271 ( \41680 , \41644 , \41679 );
and \U$33272 ( \41681 , \41371 , \41375 );
and \U$33273 ( \41682 , \41376 , \41379 );
or \U$33274 ( \41683 , \41681 , \41682 );
xor \U$33275 ( \41684 , \41680 , \41683 );
buf g9b63 ( \41685_nG9b63 , \41684 );
and \U$33276 ( \41686 , \10704 , \41685_nG9b63 );
or \U$33277 ( \41687 , \41640 , \41686 );
xor \U$33278 ( \41688 , \10703 , \41687 );
buf \U$33279 ( \41689 , \41688 );
buf \U$33281 ( \41690 , \41689 );
xor \U$33282 ( \41691 , \41639 , \41690 );
buf \U$33283 ( \41692 , \41691 );
xor \U$33284 ( \41693 , \41626 , \41692 );
and \U$33286 ( \41694 , \32916 , \27416_nG9bc3 );
or \U$33287 ( \41695 , 1'b0 , \41694 );
xor \U$33288 ( \41696 , 1'b0 , \41695 );
buf \U$33289 ( \41697 , \41696 );
buf \U$33291 ( \41698 , \41697 );
and \U$33292 ( \41699 , \29853 , \30366_nG9bba );
and \U$33293 ( \41700 , \29850 , \30940_nG9bb7 );
or \U$33294 ( \41701 , \41699 , \41700 );
xor \U$33295 ( \41702 , \29849 , \41701 );
buf \U$33296 ( \41703 , \41702 );
buf \U$33298 ( \41704 , \41703 );
xor \U$33299 ( \41705 , \41698 , \41704 );
buf \U$33300 ( \41706 , \41705 );
and \U$33301 ( \41707 , \28118 , \32179_nG9bb4 );
and \U$33302 ( \41708 , \28115 , \32888_nG9bb1 );
or \U$33303 ( \41709 , \41707 , \41708 );
xor \U$33304 ( \41710 , \28114 , \41709 );
buf \U$33305 ( \41711 , \41710 );
buf \U$33307 ( \41712 , \41711 );
xor \U$33308 ( \41713 , \41706 , \41712 );
and \U$33309 ( \41714 , \23201 , \34643_nG9ba2 );
and \U$33310 ( \41715 , \23198 , \35094_nG9b9f );
or \U$33311 ( \41716 , \41714 , \41715 );
xor \U$33312 ( \41717 , \23197 , \41716 );
buf \U$33313 ( \41718 , \41717 );
buf \U$33315 ( \41719 , \41718 );
xor \U$33316 ( \41720 , \41713 , \41719 );
buf \U$33317 ( \41721 , \41720 );
xor \U$33318 ( \41722 , \41693 , \41721 );
buf \U$33319 ( \41723 , \41722 );
xor \U$33320 ( \41724 , \41606 , \41723 );
buf \U$33321 ( \41725 , \41724 );
xor \U$33322 ( \41726 , \41528 , \41725 );
and \U$33323 ( \41727 , \41462 , \41726 );
and \U$33325 ( \41728 , \41456 , \41461 );
or \U$33327 ( \41729 , 1'b0 , \41728 , 1'b0 );
xor \U$33328 ( \41730 , \41727 , \41729 );
and \U$33330 ( \41731 , \41449 , \41455 );
and \U$33331 ( \41732 , \41451 , \41455 );
or \U$33332 ( \41733 , 1'b0 , \41731 , \41732 );
xor \U$33333 ( \41734 , \41730 , \41733 );
xor \U$33340 ( \41735 , \41734 , 1'b0 );
and \U$33341 ( \41736 , \41522 , \41527 );
and \U$33342 ( \41737 , \41522 , \41725 );
and \U$33343 ( \41738 , \41527 , \41725 );
or \U$33344 ( \41739 , \41736 , \41737 , \41738 );
xor \U$33345 ( \41740 , \41735 , \41739 );
and \U$33346 ( \41741 , \41467 , \41472 );
and \U$33347 ( \41742 , \41467 , \41520 );
and \U$33348 ( \41743 , \41472 , \41520 );
or \U$33349 ( \41744 , \41741 , \41742 , \41743 );
buf \U$33350 ( \41745 , \41744 );
and \U$33351 ( \41746 , \41600 , \41605 );
and \U$33352 ( \41747 , \41600 , \41723 );
and \U$33353 ( \41748 , \41605 , \41723 );
or \U$33354 ( \41749 , \41746 , \41747 , \41748 );
buf \U$33355 ( \41750 , \41749 );
and \U$33356 ( \41751 , \41585 , \41590 );
and \U$33357 ( \41752 , \41585 , \41596 );
and \U$33358 ( \41753 , \41590 , \41596 );
or \U$33359 ( \41754 , \41751 , \41752 , \41753 );
buf \U$33360 ( \41755 , \41754 );
and \U$33361 ( \41756 , \15940 , \38663_nG9b81 );
and \U$33362 ( \41757 , \15937 , \38968_nG9b7e );
or \U$33363 ( \41758 , \41756 , \41757 );
xor \U$33364 ( \41759 , \15936 , \41758 );
buf \U$33365 ( \41760 , \41759 );
buf \U$33367 ( \41761 , \41760 );
and \U$33368 ( \41762 , \14631 , \39334_nG9b7b );
and \U$33369 ( \41763 , \14628 , \39591_nG9b78 );
or \U$33370 ( \41764 , \41762 , \41763 );
xor \U$33371 ( \41765 , \14627 , \41764 );
buf \U$33372 ( \41766 , \41765 );
buf \U$33374 ( \41767 , \41766 );
xor \U$33375 ( \41768 , \41761 , \41767 );
and \U$33376 ( \41769 , \10421 , \41040_nG9b69 );
and \U$33377 ( \41770 , \10418 , \41381_nG9b66 );
or \U$33378 ( \41771 , \41769 , \41770 );
xor \U$33379 ( \41772 , \10417 , \41771 );
buf \U$33380 ( \41773 , \41772 );
buf \U$33382 ( \41774 , \41773 );
xor \U$33383 ( \41775 , \41768 , \41774 );
buf \U$33384 ( \41776 , \41775 );
xor \U$33385 ( \41777 , \41755 , \41776 );
and \U$33386 ( \41778 , \41611 , \41617 );
and \U$33387 ( \41779 , \41611 , \41624 );
and \U$33388 ( \41780 , \41617 , \41624 );
or \U$33389 ( \41781 , \41778 , \41779 , \41780 );
buf \U$33390 ( \41782 , \41781 );
xor \U$33391 ( \41783 , \41777 , \41782 );
buf \U$33392 ( \41784 , \41783 );
and \U$33393 ( \41785 , \41499 , \41504 );
and \U$33394 ( \41786 , \41499 , \41510 );
and \U$33395 ( \41787 , \41504 , \41510 );
or \U$33396 ( \41788 , \41785 , \41786 , \41787 );
buf \U$33397 ( \41789 , \41788 );
xor \U$33398 ( \41790 , \41784 , \41789 );
and \U$33399 ( \41791 , \41626 , \41692 );
and \U$33400 ( \41792 , \41626 , \41721 );
and \U$33401 ( \41793 , \41692 , \41721 );
or \U$33402 ( \41794 , \41791 , \41792 , \41793 );
buf \U$33403 ( \41795 , \41794 );
xor \U$33404 ( \41796 , \41790 , \41795 );
buf \U$33405 ( \41797 , \41796 );
xor \U$33406 ( \41798 , \41750 , \41797 );
and \U$33407 ( \41799 , \41478 , \41512 );
and \U$33408 ( \41800 , \41478 , \41518 );
and \U$33409 ( \41801 , \41512 , \41518 );
or \U$33410 ( \41802 , \41799 , \41800 , \41801 );
buf \U$33411 ( \41803 , \41802 );
xor \U$33412 ( \41804 , \41798 , \41803 );
buf \U$33413 ( \41805 , \41804 );
xor \U$33414 ( \41806 , \41745 , \41805 );
and \U$33415 ( \41807 , \41562 , \41567 );
and \U$33416 ( \41808 , \41562 , \41598 );
and \U$33417 ( \41809 , \41567 , \41598 );
or \U$33418 ( \41810 , \41807 , \41808 , \41809 );
buf \U$33419 ( \41811 , \41810 );
and \U$33420 ( \41812 , \41549 , \41554 );
and \U$33421 ( \41813 , \41549 , \41560 );
and \U$33422 ( \41814 , \41554 , \41560 );
or \U$33423 ( \41815 , \41812 , \41813 , \41814 );
buf \U$33424 ( \41816 , \41815 );
and \U$33425 ( \41817 , \41534 , \41540 );
and \U$33426 ( \41818 , \41534 , \41547 );
and \U$33427 ( \41819 , \41540 , \41547 );
or \U$33428 ( \41820 , \41817 , \41818 , \41819 );
buf \U$33429 ( \41821 , \41820 );
and \U$33430 ( \41822 , \41706 , \41712 );
and \U$33431 ( \41823 , \41706 , \41719 );
and \U$33432 ( \41824 , \41712 , \41719 );
or \U$33433 ( \41825 , \41822 , \41823 , \41824 );
buf \U$33434 ( \41826 , \41825 );
xor \U$33435 ( \41827 , \41821 , \41826 );
and \U$33436 ( \41828 , \31636 , \29179_nG9bbd );
and \U$33437 ( \41829 , \31633 , \30366_nG9bba );
or \U$33438 ( \41830 , \41828 , \41829 );
xor \U$33439 ( \41831 , \31632 , \41830 );
buf \U$33440 ( \41832 , \41831 );
buf \U$33442 ( \41833 , \41832 );
and \U$33443 ( \41834 , \28118 , \32888_nG9bb1 );
and \U$33444 ( \41835 , \28115 , \33181_nG9bae );
or \U$33445 ( \41836 , \41834 , \41835 );
xor \U$33446 ( \41837 , \28114 , \41836 );
buf \U$33447 ( \41838 , \41837 );
buf \U$33449 ( \41839 , \41838 );
xor \U$33450 ( \41840 , \41833 , \41839 );
and \U$33451 ( \41841 , \26431 , \33613_nG9bab );
and \U$33452 ( \41842 , \26428 , \34041_nG9ba8 );
or \U$33453 ( \41843 , \41841 , \41842 );
xor \U$33454 ( \41844 , \26427 , \41843 );
buf \U$33455 ( \41845 , \41844 );
buf \U$33457 ( \41846 , \41845 );
xor \U$33458 ( \41847 , \41840 , \41846 );
buf \U$33459 ( \41848 , \41847 );
xor \U$33460 ( \41849 , \41827 , \41848 );
buf \U$33461 ( \41850 , \41849 );
xor \U$33462 ( \41851 , \41816 , \41850 );
and \U$33463 ( \41852 , \41632 , \41638 );
and \U$33464 ( \41853 , \41632 , \41690 );
and \U$33465 ( \41854 , \41638 , \41690 );
or \U$33466 ( \41855 , \41852 , \41853 , \41854 );
buf \U$33467 ( \41856 , \41855 );
and \U$33468 ( \41857 , \41484 , \41490 );
and \U$33469 ( \41858 , \41484 , \41497 );
and \U$33470 ( \41859 , \41490 , \41497 );
or \U$33471 ( \41860 , \41857 , \41858 , \41859 );
buf \U$33472 ( \41861 , \41860 );
xor \U$33473 ( \41862 , \41856 , \41861 );
and \U$33474 ( \41863 , \24792 , \34294_nG9ba5 );
and \U$33475 ( \41864 , \24789 , \34643_nG9ba2 );
or \U$33476 ( \41865 , \41863 , \41864 );
xor \U$33477 ( \41866 , \24788 , \41865 );
buf \U$33478 ( \41867 , \41866 );
buf \U$33480 ( \41868 , \41867 );
and \U$33481 ( \41869 , \21658 , \35801_nG9b99 );
and \U$33482 ( \41870 , \21655 , \36172_nG9b96 );
or \U$33483 ( \41871 , \41869 , \41870 );
xor \U$33484 ( \41872 , \21654 , \41871 );
buf \U$33485 ( \41873 , \41872 );
buf \U$33487 ( \41874 , \41873 );
xor \U$33488 ( \41875 , \41868 , \41874 );
and \U$33489 ( \41876 , \18702 , \37250_nG9b8d );
and \U$33490 ( \41877 , \18699 , \37607_nG9b8a );
or \U$33491 ( \41878 , \41876 , \41877 );
xor \U$33492 ( \41879 , \18698 , \41878 );
buf \U$33493 ( \41880 , \41879 );
buf \U$33495 ( \41881 , \41880 );
xor \U$33496 ( \41882 , \41875 , \41881 );
buf \U$33497 ( \41883 , \41882 );
xor \U$33498 ( \41884 , \41862 , \41883 );
buf \U$33499 ( \41885 , \41884 );
xor \U$33500 ( \41886 , \41851 , \41885 );
buf \U$33501 ( \41887 , \41886 );
xor \U$33502 ( \41888 , \41811 , \41887 );
and \U$33503 ( \41889 , \41570 , \41576 );
and \U$33504 ( \41890 , \41570 , \41583 );
and \U$33505 ( \41891 , \41576 , \41583 );
or \U$33506 ( \41892 , \41889 , \41890 , \41891 );
buf \U$33507 ( \41893 , \41892 );
and \U$33508 ( \41894 , \17297 , \37974_nG9b87 );
and \U$33509 ( \41895 , \17294 , \38337_nG9b84 );
or \U$33510 ( \41896 , \41894 , \41895 );
xor \U$33511 ( \41897 , \17293 , \41896 );
buf \U$33512 ( \41898 , \41897 );
buf \U$33514 ( \41899 , \41898 );
xor \U$33515 ( \41900 , \41893 , \41899 );
and \U$33516 ( \41901 , \12157 , \40452_nG9b6f );
and \U$33517 ( \41902 , \12154 , \40843_nG9b6c );
or \U$33518 ( \41903 , \41901 , \41902 );
xor \U$33519 ( \41904 , \12153 , \41903 );
buf \U$33520 ( \41905 , \41904 );
buf \U$33522 ( \41906 , \41905 );
xor \U$33523 ( \41907 , \41900 , \41906 );
buf \U$33524 ( \41908 , \41907 );
and \U$33525 ( \41909 , \20155 , \36589_nG9b93 );
and \U$33526 ( \41910 , \20152 , \36986_nG9b90 );
or \U$33527 ( \41911 , \41909 , \41910 );
xor \U$33528 ( \41912 , \20151 , \41911 );
buf \U$33529 ( \41913 , \41912 );
buf \U$33531 ( \41914 , \41913 );
and \U$33532 ( \41915 , \13370 , \39963_nG9b75 );
and \U$33533 ( \41916 , \13367 , \40204_nG9b72 );
or \U$33534 ( \41917 , \41915 , \41916 );
xor \U$33535 ( \41918 , \13366 , \41917 );
buf \U$33536 ( \41919 , \41918 );
buf \U$33538 ( \41920 , \41919 );
xor \U$33539 ( \41921 , \41914 , \41920 );
and \U$33540 ( \41922 , \10707 , \41685_nG9b63 );
and \U$33541 ( \41923 , \41670 , \41674 );
and \U$33542 ( \41924 , \41674 , \41676 );
and \U$33543 ( \41925 , \41670 , \41676 );
or \U$33544 ( \41926 , \41923 , \41924 , \41925 );
and \U$33545 ( \41927 , \41657 , \41668 );
and \U$33546 ( \41928 , \41668 , \41677 );
and \U$33547 ( \41929 , \41657 , \41677 );
or \U$33548 ( \41930 , \41927 , \41928 , \41929 );
xor \U$33549 ( \41931 , \41926 , \41930 );
and \U$33550 ( \41932 , \41658 , \41662 );
and \U$33551 ( \41933 , \41662 , \41667 );
and \U$33552 ( \41934 , \41658 , \41667 );
or \U$33553 ( \41935 , \41932 , \41933 , \41934 );
and \U$33554 ( \41936 , \32794 , \29070 );
not \U$33555 ( \41937 , \41936 );
xnor \U$33556 ( \41938 , \41937 , \29076 );
not \U$33557 ( \41939 , \41938 );
xor \U$33558 ( \41940 , \41935 , \41939 );
and \U$33559 ( \41941 , \30802 , \30823 );
and \U$33560 ( \41942 , \32054 , \30246 );
nor \U$33561 ( \41943 , \41941 , \41942 );
xnor \U$33562 ( \41944 , \41943 , \30813 );
and \U$33563 ( \41945 , \29084 , \32854 );
and \U$33564 ( \41946 , \30268 , \32067 );
nor \U$33565 ( \41947 , \41945 , \41946 );
xnor \U$33566 ( \41948 , \41947 , \32805 );
xor \U$33567 ( \41949 , \41944 , \41948 );
and \U$33568 ( \41950 , \28534 , \32802 );
xor \U$33569 ( \41951 , \41949 , \41950 );
xor \U$33570 ( \41952 , \41940 , \41951 );
xor \U$33571 ( \41953 , \41931 , \41952 );
and \U$33572 ( \41954 , \41648 , \41652 );
and \U$33573 ( \41955 , \41652 , \41678 );
and \U$33574 ( \41956 , \41648 , \41678 );
or \U$33575 ( \41957 , \41954 , \41955 , \41956 );
xor \U$33576 ( \41958 , \41953 , \41957 );
and \U$33577 ( \41959 , \41644 , \41679 );
and \U$33578 ( \41960 , \41680 , \41683 );
or \U$33579 ( \41961 , \41959 , \41960 );
xor \U$33580 ( \41962 , \41958 , \41961 );
buf g9b60 ( \41963_nG9b60 , \41962 );
and \U$33581 ( \41964 , \10704 , \41963_nG9b60 );
or \U$33582 ( \41965 , \41922 , \41964 );
xor \U$33583 ( \41966 , \10703 , \41965 );
buf \U$33584 ( \41967 , \41966 );
buf \U$33586 ( \41968 , \41967 );
xor \U$33587 ( \41969 , \41921 , \41968 );
buf \U$33588 ( \41970 , \41969 );
xor \U$33589 ( \41971 , \41908 , \41970 );
and \U$33591 ( \41972 , \32916 , \28602_nG9bc0 );
or \U$33592 ( \41973 , 1'b0 , \41972 );
xor \U$33593 ( \41974 , 1'b0 , \41973 );
buf \U$33594 ( \41975 , \41974 );
buf \U$33596 ( \41976 , \41975 );
and \U$33597 ( \41977 , \29853 , \30940_nG9bb7 );
and \U$33598 ( \41978 , \29850 , \32179_nG9bb4 );
or \U$33599 ( \41979 , \41977 , \41978 );
xor \U$33600 ( \41980 , \29849 , \41979 );
buf \U$33601 ( \41981 , \41980 );
buf \U$33603 ( \41982 , \41981 );
xor \U$33604 ( \41983 , \41976 , \41982 );
buf \U$33605 ( \41984 , \41983 );
and \U$33606 ( \41985 , \41698 , \41704 );
buf \U$33607 ( \41986 , \41985 );
xor \U$33608 ( \41987 , \41984 , \41986 );
and \U$33609 ( \41988 , \23201 , \35094_nG9b9f );
and \U$33610 ( \41989 , \23198 , \35570_nG9b9c );
or \U$33611 ( \41990 , \41988 , \41989 );
xor \U$33612 ( \41991 , \23197 , \41990 );
buf \U$33613 ( \41992 , \41991 );
buf \U$33615 ( \41993 , \41992 );
xor \U$33616 ( \41994 , \41987 , \41993 );
buf \U$33617 ( \41995 , \41994 );
xor \U$33618 ( \41996 , \41971 , \41995 );
buf \U$33619 ( \41997 , \41996 );
xor \U$33620 ( \41998 , \41888 , \41997 );
buf \U$33621 ( \41999 , \41998 );
xor \U$33622 ( \42000 , \41806 , \41999 );
and \U$33623 ( \42001 , \41740 , \42000 );
and \U$33625 ( \42002 , \41734 , \41739 );
or \U$33627 ( \42003 , 1'b0 , \42002 , 1'b0 );
xor \U$33628 ( \42004 , \42001 , \42003 );
and \U$33630 ( \42005 , \41727 , \41733 );
and \U$33631 ( \42006 , \41729 , \41733 );
or \U$33632 ( \42007 , 1'b0 , \42005 , \42006 );
xor \U$33633 ( \42008 , \42004 , \42007 );
xor \U$33640 ( \42009 , \42008 , 1'b0 );
and \U$33641 ( \42010 , \41745 , \41805 );
and \U$33642 ( \42011 , \41745 , \41999 );
and \U$33643 ( \42012 , \41805 , \41999 );
or \U$33644 ( \42013 , \42010 , \42011 , \42012 );
xor \U$33645 ( \42014 , \42009 , \42013 );
and \U$33646 ( \42015 , \41811 , \41887 );
and \U$33647 ( \42016 , \41811 , \41997 );
and \U$33648 ( \42017 , \41887 , \41997 );
or \U$33649 ( \42018 , \42015 , \42016 , \42017 );
buf \U$33650 ( \42019 , \42018 );
and \U$33651 ( \42020 , \41833 , \41839 );
and \U$33652 ( \42021 , \41833 , \41846 );
and \U$33653 ( \42022 , \41839 , \41846 );
or \U$33654 ( \42023 , \42020 , \42021 , \42022 );
buf \U$33655 ( \42024 , \42023 );
and \U$33656 ( \42025 , \17297 , \38337_nG9b84 );
and \U$33657 ( \42026 , \17294 , \38663_nG9b81 );
or \U$33658 ( \42027 , \42025 , \42026 );
xor \U$33659 ( \42028 , \17293 , \42027 );
buf \U$33660 ( \42029 , \42028 );
buf \U$33662 ( \42030 , \42029 );
xor \U$33663 ( \42031 , \42024 , \42030 );
and \U$33664 ( \42032 , \12157 , \40843_nG9b6c );
and \U$33665 ( \42033 , \12154 , \41040_nG9b69 );
or \U$33666 ( \42034 , \42032 , \42033 );
xor \U$33667 ( \42035 , \12153 , \42034 );
buf \U$33668 ( \42036 , \42035 );
buf \U$33670 ( \42037 , \42036 );
xor \U$33671 ( \42038 , \42031 , \42037 );
buf \U$33672 ( \42039 , \42038 );
and \U$33673 ( \42040 , \41893 , \41899 );
and \U$33674 ( \42041 , \41893 , \41906 );
and \U$33675 ( \42042 , \41899 , \41906 );
or \U$33676 ( \42043 , \42040 , \42041 , \42042 );
buf \U$33677 ( \42044 , \42043 );
xor \U$33678 ( \42045 , \42039 , \42044 );
and \U$33679 ( \42046 , \20155 , \36986_nG9b90 );
and \U$33680 ( \42047 , \20152 , \37250_nG9b8d );
or \U$33681 ( \42048 , \42046 , \42047 );
xor \U$33682 ( \42049 , \20151 , \42048 );
buf \U$33683 ( \42050 , \42049 );
buf \U$33685 ( \42051 , \42050 );
and \U$33686 ( \42052 , \13370 , \40204_nG9b72 );
and \U$33687 ( \42053 , \13367 , \40452_nG9b6f );
or \U$33688 ( \42054 , \42052 , \42053 );
xor \U$33689 ( \42055 , \13366 , \42054 );
buf \U$33690 ( \42056 , \42055 );
buf \U$33692 ( \42057 , \42056 );
xor \U$33693 ( \42058 , \42051 , \42057 );
and \U$33694 ( \42059 , \10421 , \41381_nG9b66 );
and \U$33695 ( \42060 , \10418 , \41685_nG9b63 );
or \U$33696 ( \42061 , \42059 , \42060 );
xor \U$33697 ( \42062 , \10417 , \42061 );
buf \U$33698 ( \42063 , \42062 );
buf \U$33700 ( \42064 , \42063 );
xor \U$33701 ( \42065 , \42058 , \42064 );
buf \U$33702 ( \42066 , \42065 );
xor \U$33703 ( \42067 , \42045 , \42066 );
buf \U$33704 ( \42068 , \42067 );
and \U$33705 ( \42069 , \41755 , \41776 );
and \U$33706 ( \42070 , \41755 , \41782 );
and \U$33707 ( \42071 , \41776 , \41782 );
or \U$33708 ( \42072 , \42069 , \42070 , \42071 );
buf \U$33709 ( \42073 , \42072 );
xor \U$33710 ( \42074 , \42068 , \42073 );
and \U$33711 ( \42075 , \41908 , \41970 );
and \U$33712 ( \42076 , \41908 , \41995 );
and \U$33713 ( \42077 , \41970 , \41995 );
or \U$33714 ( \42078 , \42075 , \42076 , \42077 );
buf \U$33715 ( \42079 , \42078 );
xor \U$33716 ( \42080 , \42074 , \42079 );
buf \U$33717 ( \42081 , \42080 );
xor \U$33718 ( \42082 , \42019 , \42081 );
and \U$33719 ( \42083 , \41784 , \41789 );
and \U$33720 ( \42084 , \41784 , \41795 );
and \U$33721 ( \42085 , \41789 , \41795 );
or \U$33722 ( \42086 , \42083 , \42084 , \42085 );
buf \U$33723 ( \42087 , \42086 );
xor \U$33724 ( \42088 , \42082 , \42087 );
buf \U$33725 ( \42089 , \42088 );
and \U$33726 ( \42090 , \41750 , \41797 );
and \U$33727 ( \42091 , \41750 , \41803 );
and \U$33728 ( \42092 , \41797 , \41803 );
or \U$33729 ( \42093 , \42090 , \42091 , \42092 );
buf \U$33730 ( \42094 , \42093 );
xor \U$33731 ( \42095 , \42089 , \42094 );
and \U$33732 ( \42096 , \41816 , \41850 );
and \U$33733 ( \42097 , \41816 , \41885 );
and \U$33734 ( \42098 , \41850 , \41885 );
or \U$33735 ( \42099 , \42096 , \42097 , \42098 );
buf \U$33736 ( \42100 , \42099 );
and \U$33737 ( \42101 , \41868 , \41874 );
and \U$33738 ( \42102 , \41868 , \41881 );
and \U$33739 ( \42103 , \41874 , \41881 );
or \U$33740 ( \42104 , \42101 , \42102 , \42103 );
buf \U$33741 ( \42105 , \42104 );
and \U$33742 ( \42106 , \41984 , \41986 );
and \U$33743 ( \42107 , \41984 , \41993 );
and \U$33744 ( \42108 , \41986 , \41993 );
or \U$33745 ( \42109 , \42106 , \42107 , \42108 );
buf \U$33746 ( \42110 , \42109 );
xor \U$33747 ( \42111 , \42105 , \42110 );
and \U$33748 ( \42112 , \41976 , \41982 );
buf \U$33749 ( \42113 , \42112 );
and \U$33750 ( \42114 , \29853 , \32179_nG9bb4 );
and \U$33751 ( \42115 , \29850 , \32888_nG9bb1 );
or \U$33752 ( \42116 , \42114 , \42115 );
xor \U$33753 ( \42117 , \29849 , \42116 );
buf \U$33754 ( \42118 , \42117 );
buf \U$33756 ( \42119 , \42118 );
xor \U$33757 ( \42120 , \42113 , \42119 );
and \U$33758 ( \42121 , \28118 , \33181_nG9bae );
and \U$33759 ( \42122 , \28115 , \33613_nG9bab );
or \U$33760 ( \42123 , \42121 , \42122 );
xor \U$33761 ( \42124 , \28114 , \42123 );
buf \U$33762 ( \42125 , \42124 );
buf \U$33764 ( \42126 , \42125 );
xor \U$33765 ( \42127 , \42120 , \42126 );
buf \U$33766 ( \42128 , \42127 );
xor \U$33767 ( \42129 , \42111 , \42128 );
buf \U$33768 ( \42130 , \42129 );
and \U$33769 ( \42131 , \21658 , \36172_nG9b96 );
and \U$33770 ( \42132 , \21655 , \36589_nG9b93 );
or \U$33771 ( \42133 , \42131 , \42132 );
xor \U$33772 ( \42134 , \21654 , \42133 );
buf \U$33773 ( \42135 , \42134 );
buf \U$33775 ( \42136 , \42135 );
and \U$33776 ( \42137 , \15940 , \38968_nG9b7e );
and \U$33777 ( \42138 , \15937 , \39334_nG9b7b );
or \U$33778 ( \42139 , \42137 , \42138 );
xor \U$33779 ( \42140 , \15936 , \42139 );
buf \U$33780 ( \42141 , \42140 );
buf \U$33782 ( \42142 , \42141 );
xor \U$33783 ( \42143 , \42136 , \42142 );
and \U$33784 ( \42144 , \14631 , \39591_nG9b78 );
and \U$33785 ( \42145 , \14628 , \39963_nG9b75 );
or \U$33786 ( \42146 , \42144 , \42145 );
xor \U$33787 ( \42147 , \14627 , \42146 );
buf \U$33788 ( \42148 , \42147 );
buf \U$33790 ( \42149 , \42148 );
xor \U$33791 ( \42150 , \42143 , \42149 );
buf \U$33792 ( \42151 , \42150 );
xor \U$33793 ( \42152 , \42130 , \42151 );
and \U$33794 ( \42153 , \24792 , \34643_nG9ba2 );
and \U$33795 ( \42154 , \24789 , \35094_nG9b9f );
or \U$33796 ( \42155 , \42153 , \42154 );
xor \U$33797 ( \42156 , \24788 , \42155 );
buf \U$33798 ( \42157 , \42156 );
buf \U$33800 ( \42158 , \42157 );
and \U$33801 ( \42159 , \18702 , \37607_nG9b8a );
and \U$33802 ( \42160 , \18699 , \37974_nG9b87 );
or \U$33803 ( \42161 , \42159 , \42160 );
xor \U$33804 ( \42162 , \18698 , \42161 );
buf \U$33805 ( \42163 , \42162 );
buf \U$33807 ( \42164 , \42163 );
xor \U$33808 ( \42165 , \42158 , \42164 );
and \U$33809 ( \42166 , \10707 , \41963_nG9b60 );
and \U$33810 ( \42167 , \41935 , \41939 );
and \U$33811 ( \42168 , \41939 , \41951 );
and \U$33812 ( \42169 , \41935 , \41951 );
or \U$33813 ( \42170 , \42167 , \42168 , \42169 );
not \U$33814 ( \42171 , \29076 );
and \U$33815 ( \42172 , \32054 , \30823 );
and \U$33816 ( \42173 , \32794 , \30246 );
nor \U$33817 ( \42174 , \42172 , \42173 );
xnor \U$33818 ( \42175 , \42174 , \30813 );
xor \U$33819 ( \42176 , \42171 , \42175 );
and \U$33820 ( \42177 , \29084 , \32802 );
xor \U$33821 ( \42178 , \42176 , \42177 );
xor \U$33822 ( \42179 , \42170 , \42178 );
and \U$33823 ( \42180 , \41944 , \41948 );
and \U$33824 ( \42181 , \41948 , \41950 );
and \U$33825 ( \42182 , \41944 , \41950 );
or \U$33826 ( \42183 , \42180 , \42181 , \42182 );
buf \U$33827 ( \42184 , \41938 );
xor \U$33828 ( \42185 , \42183 , \42184 );
and \U$33829 ( \42186 , \30268 , \32854 );
and \U$33830 ( \42187 , \30802 , \32067 );
nor \U$33831 ( \42188 , \42186 , \42187 );
xnor \U$33832 ( \42189 , \42188 , \32805 );
xor \U$33833 ( \42190 , \42185 , \42189 );
xor \U$33834 ( \42191 , \42179 , \42190 );
and \U$33835 ( \42192 , \41926 , \41930 );
and \U$33836 ( \42193 , \41930 , \41952 );
and \U$33837 ( \42194 , \41926 , \41952 );
or \U$33838 ( \42195 , \42192 , \42193 , \42194 );
xor \U$33839 ( \42196 , \42191 , \42195 );
and \U$33840 ( \42197 , \41953 , \41957 );
and \U$33841 ( \42198 , \41958 , \41961 );
or \U$33842 ( \42199 , \42197 , \42198 );
xor \U$33843 ( \42200 , \42196 , \42199 );
buf g9b5d ( \42201_nG9b5d , \42200 );
and \U$33844 ( \42202 , \10704 , \42201_nG9b5d );
or \U$33845 ( \42203 , \42166 , \42202 );
xor \U$33846 ( \42204 , \10703 , \42203 );
buf \U$33847 ( \42205 , \42204 );
buf \U$33849 ( \42206 , \42205 );
xor \U$33850 ( \42207 , \42165 , \42206 );
buf \U$33851 ( \42208 , \42207 );
xor \U$33852 ( \42209 , \42152 , \42208 );
buf \U$33853 ( \42210 , \42209 );
xor \U$33854 ( \42211 , \42100 , \42210 );
and \U$33855 ( \42212 , \41856 , \41861 );
and \U$33856 ( \42213 , \41856 , \41883 );
and \U$33857 ( \42214 , \41861 , \41883 );
or \U$33858 ( \42215 , \42212 , \42213 , \42214 );
buf \U$33859 ( \42216 , \42215 );
and \U$33861 ( \42217 , \32916 , \29179_nG9bbd );
or \U$33862 ( \42218 , 1'b0 , \42217 );
xor \U$33863 ( \42219 , 1'b0 , \42218 );
buf \U$33864 ( \42220 , \42219 );
buf \U$33866 ( \42221 , \42220 );
and \U$33867 ( \42222 , \31636 , \30366_nG9bba );
and \U$33868 ( \42223 , \31633 , \30940_nG9bb7 );
or \U$33869 ( \42224 , \42222 , \42223 );
xor \U$33870 ( \42225 , \31632 , \42224 );
buf \U$33871 ( \42226 , \42225 );
buf \U$33873 ( \42227 , \42226 );
xor \U$33874 ( \42228 , \42221 , \42227 );
buf \U$33875 ( \42229 , \42228 );
and \U$33876 ( \42230 , \26431 , \34041_nG9ba8 );
and \U$33877 ( \42231 , \26428 , \34294_nG9ba5 );
or \U$33878 ( \42232 , \42230 , \42231 );
xor \U$33879 ( \42233 , \26427 , \42232 );
buf \U$33880 ( \42234 , \42233 );
buf \U$33882 ( \42235 , \42234 );
xor \U$33883 ( \42236 , \42229 , \42235 );
and \U$33884 ( \42237 , \23201 , \35570_nG9b9c );
and \U$33885 ( \42238 , \23198 , \35801_nG9b99 );
or \U$33886 ( \42239 , \42237 , \42238 );
xor \U$33887 ( \42240 , \23197 , \42239 );
buf \U$33888 ( \42241 , \42240 );
buf \U$33890 ( \42242 , \42241 );
xor \U$33891 ( \42243 , \42236 , \42242 );
buf \U$33892 ( \42244 , \42243 );
and \U$33893 ( \42245 , \41914 , \41920 );
and \U$33894 ( \42246 , \41914 , \41968 );
and \U$33895 ( \42247 , \41920 , \41968 );
or \U$33896 ( \42248 , \42245 , \42246 , \42247 );
buf \U$33897 ( \42249 , \42248 );
xor \U$33898 ( \42250 , \42244 , \42249 );
and \U$33899 ( \42251 , \41761 , \41767 );
and \U$33900 ( \42252 , \41761 , \41774 );
and \U$33901 ( \42253 , \41767 , \41774 );
or \U$33902 ( \42254 , \42251 , \42252 , \42253 );
buf \U$33903 ( \42255 , \42254 );
xor \U$33904 ( \42256 , \42250 , \42255 );
buf \U$33905 ( \42257 , \42256 );
xor \U$33906 ( \42258 , \42216 , \42257 );
and \U$33907 ( \42259 , \41821 , \41826 );
and \U$33908 ( \42260 , \41821 , \41848 );
and \U$33909 ( \42261 , \41826 , \41848 );
or \U$33910 ( \42262 , \42259 , \42260 , \42261 );
buf \U$33911 ( \42263 , \42262 );
xor \U$33912 ( \42264 , \42258 , \42263 );
buf \U$33913 ( \42265 , \42264 );
xor \U$33914 ( \42266 , \42211 , \42265 );
buf \U$33915 ( \42267 , \42266 );
xor \U$33916 ( \42268 , \42095 , \42267 );
and \U$33917 ( \42269 , \42014 , \42268 );
and \U$33919 ( \42270 , \42008 , \42013 );
or \U$33921 ( \42271 , 1'b0 , \42270 , 1'b0 );
xor \U$33922 ( \42272 , \42269 , \42271 );
and \U$33924 ( \42273 , \42001 , \42007 );
and \U$33925 ( \42274 , \42003 , \42007 );
or \U$33926 ( \42275 , 1'b0 , \42273 , \42274 );
xor \U$33927 ( \42276 , \42272 , \42275 );
xor \U$33934 ( \42277 , \42276 , 1'b0 );
and \U$33935 ( \42278 , \42089 , \42094 );
and \U$33936 ( \42279 , \42089 , \42267 );
and \U$33937 ( \42280 , \42094 , \42267 );
or \U$33938 ( \42281 , \42278 , \42279 , \42280 );
xor \U$33939 ( \42282 , \42277 , \42281 );
and \U$33940 ( \42283 , \42100 , \42210 );
and \U$33941 ( \42284 , \42100 , \42265 );
and \U$33942 ( \42285 , \42210 , \42265 );
or \U$33943 ( \42286 , \42283 , \42284 , \42285 );
buf \U$33944 ( \42287 , \42286 );
and \U$33945 ( \42288 , \42221 , \42227 );
buf \U$33946 ( \42289 , \42288 );
and \U$33947 ( \42290 , \29853 , \32888_nG9bb1 );
and \U$33948 ( \42291 , \29850 , \33181_nG9bae );
or \U$33949 ( \42292 , \42290 , \42291 );
xor \U$33950 ( \42293 , \29849 , \42292 );
buf \U$33951 ( \42294 , \42293 );
buf \U$33953 ( \42295 , \42294 );
xor \U$33954 ( \42296 , \42289 , \42295 );
and \U$33955 ( \42297 , \28118 , \33613_nG9bab );
and \U$33956 ( \42298 , \28115 , \34041_nG9ba8 );
or \U$33957 ( \42299 , \42297 , \42298 );
xor \U$33958 ( \42300 , \28114 , \42299 );
buf \U$33959 ( \42301 , \42300 );
buf \U$33961 ( \42302 , \42301 );
xor \U$33962 ( \42303 , \42296 , \42302 );
buf \U$33963 ( \42304 , \42303 );
and \U$33964 ( \42305 , \42229 , \42235 );
and \U$33965 ( \42306 , \42229 , \42242 );
and \U$33966 ( \42307 , \42235 , \42242 );
or \U$33967 ( \42308 , \42305 , \42306 , \42307 );
buf \U$33968 ( \42309 , \42308 );
xor \U$33969 ( \42310 , \42304 , \42309 );
and \U$33970 ( \42311 , \42158 , \42164 );
and \U$33971 ( \42312 , \42158 , \42206 );
and \U$33972 ( \42313 , \42164 , \42206 );
or \U$33973 ( \42314 , \42311 , \42312 , \42313 );
buf \U$33974 ( \42315 , \42314 );
xor \U$33975 ( \42316 , \42310 , \42315 );
buf \U$33976 ( \42317 , \42316 );
and \U$33977 ( \42318 , \42113 , \42119 );
and \U$33978 ( \42319 , \42113 , \42126 );
and \U$33979 ( \42320 , \42119 , \42126 );
or \U$33980 ( \42321 , \42318 , \42319 , \42320 );
buf \U$33981 ( \42322 , \42321 );
and \U$33982 ( \42323 , \17297 , \38663_nG9b81 );
and \U$33983 ( \42324 , \17294 , \38968_nG9b7e );
or \U$33984 ( \42325 , \42323 , \42324 );
xor \U$33985 ( \42326 , \17293 , \42325 );
buf \U$33986 ( \42327 , \42326 );
buf \U$33988 ( \42328 , \42327 );
xor \U$33989 ( \42329 , \42322 , \42328 );
and \U$33990 ( \42330 , \12157 , \41040_nG9b69 );
and \U$33991 ( \42331 , \12154 , \41381_nG9b66 );
or \U$33992 ( \42332 , \42330 , \42331 );
xor \U$33993 ( \42333 , \12153 , \42332 );
buf \U$33994 ( \42334 , \42333 );
buf \U$33996 ( \42335 , \42334 );
xor \U$33997 ( \42336 , \42329 , \42335 );
buf \U$33998 ( \42337 , \42336 );
xor \U$33999 ( \42338 , \42317 , \42337 );
and \U$34000 ( \42339 , \21658 , \36589_nG9b93 );
and \U$34001 ( \42340 , \21655 , \36986_nG9b90 );
or \U$34002 ( \42341 , \42339 , \42340 );
xor \U$34003 ( \42342 , \21654 , \42341 );
buf \U$34004 ( \42343 , \42342 );
buf \U$34006 ( \42344 , \42343 );
and \U$34007 ( \42345 , \15940 , \39334_nG9b7b );
and \U$34008 ( \42346 , \15937 , \39591_nG9b78 );
or \U$34009 ( \42347 , \42345 , \42346 );
xor \U$34010 ( \42348 , \15936 , \42347 );
buf \U$34011 ( \42349 , \42348 );
buf \U$34013 ( \42350 , \42349 );
xor \U$34014 ( \42351 , \42344 , \42350 );
and \U$34015 ( \42352 , \14631 , \39963_nG9b75 );
and \U$34016 ( \42353 , \14628 , \40204_nG9b72 );
or \U$34017 ( \42354 , \42352 , \42353 );
xor \U$34018 ( \42355 , \14627 , \42354 );
buf \U$34019 ( \42356 , \42355 );
buf \U$34021 ( \42357 , \42356 );
xor \U$34022 ( \42358 , \42351 , \42357 );
buf \U$34023 ( \42359 , \42358 );
xor \U$34024 ( \42360 , \42338 , \42359 );
buf \U$34025 ( \42361 , \42360 );
and \U$34026 ( \42362 , \42024 , \42030 );
and \U$34027 ( \42363 , \42024 , \42037 );
and \U$34028 ( \42364 , \42030 , \42037 );
or \U$34029 ( \42365 , \42362 , \42363 , \42364 );
buf \U$34030 ( \42366 , \42365 );
and \U$34031 ( \42367 , \20155 , \37250_nG9b8d );
and \U$34032 ( \42368 , \20152 , \37607_nG9b8a );
or \U$34033 ( \42369 , \42367 , \42368 );
xor \U$34034 ( \42370 , \20151 , \42369 );
buf \U$34035 ( \42371 , \42370 );
buf \U$34037 ( \42372 , \42371 );
and \U$34038 ( \42373 , \13370 , \40452_nG9b6f );
and \U$34039 ( \42374 , \13367 , \40843_nG9b6c );
or \U$34040 ( \42375 , \42373 , \42374 );
xor \U$34041 ( \42376 , \13366 , \42375 );
buf \U$34042 ( \42377 , \42376 );
buf \U$34044 ( \42378 , \42377 );
xor \U$34045 ( \42379 , \42372 , \42378 );
and \U$34046 ( \42380 , \10421 , \41685_nG9b63 );
and \U$34047 ( \42381 , \10418 , \41963_nG9b60 );
or \U$34048 ( \42382 , \42380 , \42381 );
xor \U$34049 ( \42383 , \10417 , \42382 );
buf \U$34050 ( \42384 , \42383 );
buf \U$34052 ( \42385 , \42384 );
xor \U$34053 ( \42386 , \42379 , \42385 );
buf \U$34054 ( \42387 , \42386 );
xor \U$34055 ( \42388 , \42366 , \42387 );
and \U$34056 ( \42389 , \24792 , \35094_nG9b9f );
and \U$34057 ( \42390 , \24789 , \35570_nG9b9c );
or \U$34058 ( \42391 , \42389 , \42390 );
xor \U$34059 ( \42392 , \24788 , \42391 );
buf \U$34060 ( \42393 , \42392 );
buf \U$34062 ( \42394 , \42393 );
and \U$34063 ( \42395 , \18702 , \37974_nG9b87 );
and \U$34064 ( \42396 , \18699 , \38337_nG9b84 );
or \U$34065 ( \42397 , \42395 , \42396 );
xor \U$34066 ( \42398 , \18698 , \42397 );
buf \U$34067 ( \42399 , \42398 );
buf \U$34069 ( \42400 , \42399 );
xor \U$34070 ( \42401 , \42394 , \42400 );
and \U$34071 ( \42402 , \10707 , \42201_nG9b5d );
and \U$34072 ( \42403 , \42171 , \42175 );
and \U$34073 ( \42404 , \42175 , \42177 );
and \U$34074 ( \42405 , \42171 , \42177 );
or \U$34075 ( \42406 , \42403 , \42404 , \42405 );
and \U$34076 ( \42407 , \42183 , \42184 );
and \U$34077 ( \42408 , \42184 , \42189 );
and \U$34078 ( \42409 , \42183 , \42189 );
or \U$34079 ( \42410 , \42407 , \42408 , \42409 );
xor \U$34080 ( \42411 , \42406 , \42410 );
and \U$34081 ( \42412 , \32794 , \30823 );
not \U$34082 ( \42413 , \42412 );
xnor \U$34083 ( \42414 , \42413 , \30813 );
not \U$34084 ( \42415 , \42414 );
and \U$34085 ( \42416 , \30802 , \32854 );
and \U$34086 ( \42417 , \32054 , \32067 );
nor \U$34087 ( \42418 , \42416 , \42417 );
xnor \U$34088 ( \42419 , \42418 , \32805 );
xor \U$34089 ( \42420 , \42415 , \42419 );
and \U$34090 ( \42421 , \30268 , \32802 );
xor \U$34091 ( \42422 , \42420 , \42421 );
xor \U$34092 ( \42423 , \42411 , \42422 );
and \U$34093 ( \42424 , \42170 , \42178 );
and \U$34094 ( \42425 , \42178 , \42190 );
and \U$34095 ( \42426 , \42170 , \42190 );
or \U$34096 ( \42427 , \42424 , \42425 , \42426 );
xor \U$34097 ( \42428 , \42423 , \42427 );
and \U$34098 ( \42429 , \42191 , \42195 );
and \U$34099 ( \42430 , \42196 , \42199 );
or \U$34100 ( \42431 , \42429 , \42430 );
xor \U$34101 ( \42432 , \42428 , \42431 );
buf g9b5a ( \42433_nG9b5a , \42432 );
and \U$34102 ( \42434 , \10704 , \42433_nG9b5a );
or \U$34103 ( \42435 , \42402 , \42434 );
xor \U$34104 ( \42436 , \10703 , \42435 );
buf \U$34105 ( \42437 , \42436 );
buf \U$34107 ( \42438 , \42437 );
xor \U$34108 ( \42439 , \42401 , \42438 );
buf \U$34109 ( \42440 , \42439 );
xor \U$34110 ( \42441 , \42388 , \42440 );
buf \U$34111 ( \42442 , \42441 );
xor \U$34112 ( \42443 , \42361 , \42442 );
and \U$34113 ( \42444 , \42039 , \42044 );
and \U$34114 ( \42445 , \42039 , \42066 );
and \U$34115 ( \42446 , \42044 , \42066 );
or \U$34116 ( \42447 , \42444 , \42445 , \42446 );
buf \U$34117 ( \42448 , \42447 );
xor \U$34118 ( \42449 , \42443 , \42448 );
buf \U$34119 ( \42450 , \42449 );
xor \U$34120 ( \42451 , \42287 , \42450 );
and \U$34121 ( \42452 , \42068 , \42073 );
and \U$34122 ( \42453 , \42068 , \42079 );
and \U$34123 ( \42454 , \42073 , \42079 );
or \U$34124 ( \42455 , \42452 , \42453 , \42454 );
buf \U$34125 ( \42456 , \42455 );
xor \U$34126 ( \42457 , \42451 , \42456 );
buf \U$34127 ( \42458 , \42457 );
and \U$34128 ( \42459 , \42019 , \42081 );
and \U$34129 ( \42460 , \42019 , \42087 );
and \U$34130 ( \42461 , \42081 , \42087 );
or \U$34131 ( \42462 , \42459 , \42460 , \42461 );
buf \U$34132 ( \42463 , \42462 );
xor \U$34133 ( \42464 , \42458 , \42463 );
and \U$34134 ( \42465 , \42216 , \42257 );
and \U$34135 ( \42466 , \42216 , \42263 );
and \U$34136 ( \42467 , \42257 , \42263 );
or \U$34137 ( \42468 , \42465 , \42466 , \42467 );
buf \U$34138 ( \42469 , \42468 );
and \U$34140 ( \42470 , \32916 , \30366_nG9bba );
or \U$34141 ( \42471 , 1'b0 , \42470 );
xor \U$34142 ( \42472 , 1'b0 , \42471 );
buf \U$34143 ( \42473 , \42472 );
buf \U$34145 ( \42474 , \42473 );
and \U$34146 ( \42475 , \31636 , \30940_nG9bb7 );
and \U$34147 ( \42476 , \31633 , \32179_nG9bb4 );
or \U$34148 ( \42477 , \42475 , \42476 );
xor \U$34149 ( \42478 , \31632 , \42477 );
buf \U$34150 ( \42479 , \42478 );
buf \U$34152 ( \42480 , \42479 );
xor \U$34153 ( \42481 , \42474 , \42480 );
buf \U$34154 ( \42482 , \42481 );
and \U$34155 ( \42483 , \26431 , \34294_nG9ba5 );
and \U$34156 ( \42484 , \26428 , \34643_nG9ba2 );
or \U$34157 ( \42485 , \42483 , \42484 );
xor \U$34158 ( \42486 , \26427 , \42485 );
buf \U$34159 ( \42487 , \42486 );
buf \U$34161 ( \42488 , \42487 );
xor \U$34162 ( \42489 , \42482 , \42488 );
and \U$34163 ( \42490 , \23201 , \35801_nG9b99 );
and \U$34164 ( \42491 , \23198 , \36172_nG9b96 );
or \U$34165 ( \42492 , \42490 , \42491 );
xor \U$34166 ( \42493 , \23197 , \42492 );
buf \U$34167 ( \42494 , \42493 );
buf \U$34169 ( \42495 , \42494 );
xor \U$34170 ( \42496 , \42489 , \42495 );
buf \U$34171 ( \42497 , \42496 );
and \U$34172 ( \42498 , \42051 , \42057 );
and \U$34173 ( \42499 , \42051 , \42064 );
and \U$34174 ( \42500 , \42057 , \42064 );
or \U$34175 ( \42501 , \42498 , \42499 , \42500 );
buf \U$34176 ( \42502 , \42501 );
xor \U$34177 ( \42503 , \42497 , \42502 );
and \U$34178 ( \42504 , \42136 , \42142 );
and \U$34179 ( \42505 , \42136 , \42149 );
and \U$34180 ( \42506 , \42142 , \42149 );
or \U$34181 ( \42507 , \42504 , \42505 , \42506 );
buf \U$34182 ( \42508 , \42507 );
xor \U$34183 ( \42509 , \42503 , \42508 );
buf \U$34184 ( \42510 , \42509 );
and \U$34185 ( \42511 , \42244 , \42249 );
and \U$34186 ( \42512 , \42244 , \42255 );
and \U$34187 ( \42513 , \42249 , \42255 );
or \U$34188 ( \42514 , \42511 , \42512 , \42513 );
buf \U$34189 ( \42515 , \42514 );
xor \U$34190 ( \42516 , \42510 , \42515 );
and \U$34191 ( \42517 , \42105 , \42110 );
and \U$34192 ( \42518 , \42105 , \42128 );
and \U$34193 ( \42519 , \42110 , \42128 );
or \U$34194 ( \42520 , \42517 , \42518 , \42519 );
buf \U$34195 ( \42521 , \42520 );
xor \U$34196 ( \42522 , \42516 , \42521 );
buf \U$34197 ( \42523 , \42522 );
xor \U$34198 ( \42524 , \42469 , \42523 );
and \U$34199 ( \42525 , \42130 , \42151 );
and \U$34200 ( \42526 , \42130 , \42208 );
and \U$34201 ( \42527 , \42151 , \42208 );
or \U$34202 ( \42528 , \42525 , \42526 , \42527 );
buf \U$34203 ( \42529 , \42528 );
xor \U$34204 ( \42530 , \42524 , \42529 );
buf \U$34205 ( \42531 , \42530 );
xor \U$34206 ( \42532 , \42464 , \42531 );
and \U$34207 ( \42533 , \42282 , \42532 );
and \U$34209 ( \42534 , \42276 , \42281 );
or \U$34211 ( \42535 , 1'b0 , \42534 , 1'b0 );
xor \U$34212 ( \42536 , \42533 , \42535 );
and \U$34214 ( \42537 , \42269 , \42275 );
and \U$34215 ( \42538 , \42271 , \42275 );
or \U$34216 ( \42539 , 1'b0 , \42537 , \42538 );
xor \U$34217 ( \42540 , \42536 , \42539 );
xor \U$34224 ( \42541 , \42540 , 1'b0 );
and \U$34225 ( \42542 , \42458 , \42463 );
and \U$34226 ( \42543 , \42458 , \42531 );
and \U$34227 ( \42544 , \42463 , \42531 );
or \U$34228 ( \42545 , \42542 , \42543 , \42544 );
xor \U$34229 ( \42546 , \42541 , \42545 );
and \U$34230 ( \42547 , \42469 , \42523 );
and \U$34231 ( \42548 , \42469 , \42529 );
and \U$34232 ( \42549 , \42523 , \42529 );
or \U$34233 ( \42550 , \42547 , \42548 , \42549 );
buf \U$34234 ( \42551 , \42550 );
and \U$34235 ( \42552 , \42361 , \42442 );
and \U$34236 ( \42553 , \42361 , \42448 );
and \U$34237 ( \42554 , \42442 , \42448 );
or \U$34238 ( \42555 , \42552 , \42553 , \42554 );
buf \U$34239 ( \42556 , \42555 );
xor \U$34240 ( \42557 , \42551 , \42556 );
and \U$34241 ( \42558 , \42317 , \42337 );
and \U$34242 ( \42559 , \42317 , \42359 );
and \U$34243 ( \42560 , \42337 , \42359 );
or \U$34244 ( \42561 , \42558 , \42559 , \42560 );
buf \U$34245 ( \42562 , \42561 );
and \U$34247 ( \42563 , \32916 , \30940_nG9bb7 );
or \U$34248 ( \42564 , 1'b0 , \42563 );
xor \U$34249 ( \42565 , 1'b0 , \42564 );
buf \U$34250 ( \42566 , \42565 );
buf \U$34252 ( \42567 , \42566 );
and \U$34253 ( \42568 , \29853 , \33181_nG9bae );
and \U$34254 ( \42569 , \29850 , \33613_nG9bab );
or \U$34255 ( \42570 , \42568 , \42569 );
xor \U$34256 ( \42571 , \29849 , \42570 );
buf \U$34257 ( \42572 , \42571 );
buf \U$34259 ( \42573 , \42572 );
xor \U$34260 ( \42574 , \42567 , \42573 );
buf \U$34261 ( \42575 , \42574 );
and \U$34262 ( \42576 , \20155 , \37607_nG9b8a );
and \U$34263 ( \42577 , \20152 , \37974_nG9b87 );
or \U$34264 ( \42578 , \42576 , \42577 );
xor \U$34265 ( \42579 , \20151 , \42578 );
buf \U$34266 ( \42580 , \42579 );
buf \U$34268 ( \42581 , \42580 );
xor \U$34269 ( \42582 , \42575 , \42581 );
and \U$34270 ( \42583 , \18702 , \38337_nG9b84 );
and \U$34271 ( \42584 , \18699 , \38663_nG9b81 );
or \U$34272 ( \42585 , \42583 , \42584 );
xor \U$34273 ( \42586 , \18698 , \42585 );
buf \U$34274 ( \42587 , \42586 );
buf \U$34276 ( \42588 , \42587 );
xor \U$34277 ( \42589 , \42582 , \42588 );
buf \U$34278 ( \42590 , \42589 );
and \U$34279 ( \42591 , \23201 , \36172_nG9b96 );
and \U$34280 ( \42592 , \23198 , \36589_nG9b93 );
or \U$34281 ( \42593 , \42591 , \42592 );
xor \U$34282 ( \42594 , \23197 , \42593 );
buf \U$34283 ( \42595 , \42594 );
buf \U$34285 ( \42596 , \42595 );
and \U$34286 ( \42597 , \21658 , \36986_nG9b90 );
and \U$34287 ( \42598 , \21655 , \37250_nG9b8d );
or \U$34288 ( \42599 , \42597 , \42598 );
xor \U$34289 ( \42600 , \21654 , \42599 );
buf \U$34290 ( \42601 , \42600 );
buf \U$34292 ( \42602 , \42601 );
xor \U$34293 ( \42603 , \42596 , \42602 );
and \U$34294 ( \42604 , \14631 , \40204_nG9b72 );
and \U$34295 ( \42605 , \14628 , \40452_nG9b6f );
or \U$34296 ( \42606 , \42604 , \42605 );
xor \U$34297 ( \42607 , \14627 , \42606 );
buf \U$34298 ( \42608 , \42607 );
buf \U$34300 ( \42609 , \42608 );
xor \U$34301 ( \42610 , \42603 , \42609 );
buf \U$34302 ( \42611 , \42610 );
xor \U$34303 ( \42612 , \42590 , \42611 );
and \U$34304 ( \42613 , \15940 , \39591_nG9b78 );
and \U$34305 ( \42614 , \15937 , \39963_nG9b75 );
or \U$34306 ( \42615 , \42613 , \42614 );
xor \U$34307 ( \42616 , \15936 , \42615 );
buf \U$34308 ( \42617 , \42616 );
buf \U$34310 ( \42618 , \42617 );
and \U$34311 ( \42619 , \12157 , \41381_nG9b66 );
and \U$34312 ( \42620 , \12154 , \41685_nG9b63 );
or \U$34313 ( \42621 , \42619 , \42620 );
xor \U$34314 ( \42622 , \12153 , \42621 );
buf \U$34315 ( \42623 , \42622 );
buf \U$34317 ( \42624 , \42623 );
xor \U$34318 ( \42625 , \42618 , \42624 );
and \U$34319 ( \42626 , \10421 , \41963_nG9b60 );
and \U$34320 ( \42627 , \10418 , \42201_nG9b5d );
or \U$34321 ( \42628 , \42626 , \42627 );
xor \U$34322 ( \42629 , \10417 , \42628 );
buf \U$34323 ( \42630 , \42629 );
buf \U$34325 ( \42631 , \42630 );
xor \U$34326 ( \42632 , \42625 , \42631 );
buf \U$34327 ( \42633 , \42632 );
xor \U$34328 ( \42634 , \42612 , \42633 );
buf \U$34329 ( \42635 , \42634 );
xor \U$34330 ( \42636 , \42562 , \42635 );
and \U$34331 ( \42637 , \42366 , \42387 );
and \U$34332 ( \42638 , \42366 , \42440 );
and \U$34333 ( \42639 , \42387 , \42440 );
or \U$34334 ( \42640 , \42637 , \42638 , \42639 );
buf \U$34335 ( \42641 , \42640 );
xor \U$34336 ( \42642 , \42636 , \42641 );
buf \U$34337 ( \42643 , \42642 );
xor \U$34338 ( \42644 , \42557 , \42643 );
buf \U$34339 ( \42645 , \42644 );
and \U$34340 ( \42646 , \42287 , \42450 );
and \U$34341 ( \42647 , \42287 , \42456 );
and \U$34342 ( \42648 , \42450 , \42456 );
or \U$34343 ( \42649 , \42646 , \42647 , \42648 );
buf \U$34344 ( \42650 , \42649 );
xor \U$34345 ( \42651 , \42645 , \42650 );
and \U$34346 ( \42652 , \42344 , \42350 );
and \U$34347 ( \42653 , \42344 , \42357 );
and \U$34348 ( \42654 , \42350 , \42357 );
or \U$34349 ( \42655 , \42652 , \42653 , \42654 );
buf \U$34350 ( \42656 , \42655 );
and \U$34351 ( \42657 , \28118 , \34041_nG9ba8 );
and \U$34352 ( \42658 , \28115 , \34294_nG9ba5 );
or \U$34353 ( \42659 , \42657 , \42658 );
xor \U$34354 ( \42660 , \28114 , \42659 );
buf \U$34355 ( \42661 , \42660 );
buf \U$34357 ( \42662 , \42661 );
and \U$34358 ( \42663 , \26431 , \34643_nG9ba2 );
and \U$34359 ( \42664 , \26428 , \35094_nG9b9f );
or \U$34360 ( \42665 , \42663 , \42664 );
xor \U$34361 ( \42666 , \26427 , \42665 );
buf \U$34362 ( \42667 , \42666 );
buf \U$34364 ( \42668 , \42667 );
xor \U$34365 ( \42669 , \42662 , \42668 );
and \U$34366 ( \42670 , \13370 , \40843_nG9b6c );
and \U$34367 ( \42671 , \13367 , \41040_nG9b69 );
or \U$34368 ( \42672 , \42670 , \42671 );
xor \U$34369 ( \42673 , \13366 , \42672 );
buf \U$34370 ( \42674 , \42673 );
buf \U$34372 ( \42675 , \42674 );
xor \U$34373 ( \42676 , \42669 , \42675 );
buf \U$34374 ( \42677 , \42676 );
xor \U$34375 ( \42678 , \42656 , \42677 );
and \U$34376 ( \42679 , \42474 , \42480 );
buf \U$34377 ( \42680 , \42679 );
and \U$34378 ( \42681 , \31636 , \32179_nG9bb4 );
and \U$34379 ( \42682 , \31633 , \32888_nG9bb1 );
or \U$34380 ( \42683 , \42681 , \42682 );
xor \U$34381 ( \42684 , \31632 , \42683 );
buf \U$34382 ( \42685 , \42684 );
buf \U$34384 ( \42686 , \42685 );
xor \U$34385 ( \42687 , \42680 , \42686 );
and \U$34386 ( \42688 , \24792 , \35570_nG9b9c );
and \U$34387 ( \42689 , \24789 , \35801_nG9b99 );
or \U$34388 ( \42690 , \42688 , \42689 );
xor \U$34389 ( \42691 , \24788 , \42690 );
buf \U$34390 ( \42692 , \42691 );
buf \U$34392 ( \42693 , \42692 );
xor \U$34393 ( \42694 , \42687 , \42693 );
buf \U$34394 ( \42695 , \42694 );
xor \U$34395 ( \42696 , \42678 , \42695 );
buf \U$34396 ( \42697 , \42696 );
and \U$34397 ( \42698 , \42394 , \42400 );
and \U$34398 ( \42699 , \42394 , \42438 );
and \U$34399 ( \42700 , \42400 , \42438 );
or \U$34400 ( \42701 , \42698 , \42699 , \42700 );
buf \U$34401 ( \42702 , \42701 );
and \U$34402 ( \42703 , \42372 , \42378 );
and \U$34403 ( \42704 , \42372 , \42385 );
and \U$34404 ( \42705 , \42378 , \42385 );
or \U$34405 ( \42706 , \42703 , \42704 , \42705 );
buf \U$34406 ( \42707 , \42706 );
xor \U$34407 ( \42708 , \42702 , \42707 );
and \U$34408 ( \42709 , \42482 , \42488 );
and \U$34409 ( \42710 , \42482 , \42495 );
and \U$34410 ( \42711 , \42488 , \42495 );
or \U$34411 ( \42712 , \42709 , \42710 , \42711 );
buf \U$34412 ( \42713 , \42712 );
xor \U$34413 ( \42714 , \42708 , \42713 );
buf \U$34414 ( \42715 , \42714 );
xor \U$34415 ( \42716 , \42697 , \42715 );
and \U$34416 ( \42717 , \42497 , \42502 );
and \U$34417 ( \42718 , \42497 , \42508 );
and \U$34418 ( \42719 , \42502 , \42508 );
or \U$34419 ( \42720 , \42717 , \42718 , \42719 );
buf \U$34420 ( \42721 , \42720 );
xor \U$34421 ( \42722 , \42716 , \42721 );
buf \U$34422 ( \42723 , \42722 );
and \U$34423 ( \42724 , \42304 , \42309 );
and \U$34424 ( \42725 , \42304 , \42315 );
and \U$34425 ( \42726 , \42309 , \42315 );
or \U$34426 ( \42727 , \42724 , \42725 , \42726 );
buf \U$34427 ( \42728 , \42727 );
and \U$34428 ( \42729 , \42289 , \42295 );
and \U$34429 ( \42730 , \42289 , \42302 );
and \U$34430 ( \42731 , \42295 , \42302 );
or \U$34431 ( \42732 , \42729 , \42730 , \42731 );
buf \U$34432 ( \42733 , \42732 );
and \U$34433 ( \42734 , \17297 , \38968_nG9b7e );
and \U$34434 ( \42735 , \17294 , \39334_nG9b7b );
or \U$34435 ( \42736 , \42734 , \42735 );
xor \U$34436 ( \42737 , \17293 , \42736 );
buf \U$34437 ( \42738 , \42737 );
buf \U$34439 ( \42739 , \42738 );
xor \U$34440 ( \42740 , \42733 , \42739 );
and \U$34441 ( \42741 , \10707 , \42433_nG9b5a );
and \U$34442 ( \42742 , \42415 , \42419 );
and \U$34443 ( \42743 , \42419 , \42421 );
and \U$34444 ( \42744 , \42415 , \42421 );
or \U$34445 ( \42745 , \42742 , \42743 , \42744 );
buf \U$34446 ( \42746 , \42414 );
xor \U$34447 ( \42747 , \42745 , \42746 );
not \U$34448 ( \42748 , \30813 );
and \U$34449 ( \42749 , \32054 , \32854 );
and \U$34450 ( \42750 , \32794 , \32067 );
nor \U$34451 ( \42751 , \42749 , \42750 );
xnor \U$34452 ( \42752 , \42751 , \32805 );
xor \U$34453 ( \42753 , \42748 , \42752 );
and \U$34454 ( \42754 , \30802 , \32802 );
xor \U$34455 ( \42755 , \42753 , \42754 );
xor \U$34456 ( \42756 , \42747 , \42755 );
and \U$34457 ( \42757 , \42406 , \42410 );
and \U$34458 ( \42758 , \42410 , \42422 );
and \U$34459 ( \42759 , \42406 , \42422 );
or \U$34460 ( \42760 , \42757 , \42758 , \42759 );
xor \U$34461 ( \42761 , \42756 , \42760 );
and \U$34462 ( \42762 , \42423 , \42427 );
and \U$34463 ( \42763 , \42428 , \42431 );
or \U$34464 ( \42764 , \42762 , \42763 );
xor \U$34465 ( \42765 , \42761 , \42764 );
buf g9b57 ( \42766_nG9b57 , \42765 );
and \U$34466 ( \42767 , \10704 , \42766_nG9b57 );
or \U$34467 ( \42768 , \42741 , \42767 );
xor \U$34468 ( \42769 , \10703 , \42768 );
buf \U$34469 ( \42770 , \42769 );
buf \U$34471 ( \42771 , \42770 );
xor \U$34472 ( \42772 , \42740 , \42771 );
buf \U$34473 ( \42773 , \42772 );
xor \U$34474 ( \42774 , \42728 , \42773 );
and \U$34475 ( \42775 , \42322 , \42328 );
and \U$34476 ( \42776 , \42322 , \42335 );
and \U$34477 ( \42777 , \42328 , \42335 );
or \U$34478 ( \42778 , \42775 , \42776 , \42777 );
buf \U$34479 ( \42779 , \42778 );
xor \U$34480 ( \42780 , \42774 , \42779 );
buf \U$34481 ( \42781 , \42780 );
xor \U$34482 ( \42782 , \42723 , \42781 );
and \U$34483 ( \42783 , \42510 , \42515 );
and \U$34484 ( \42784 , \42510 , \42521 );
and \U$34485 ( \42785 , \42515 , \42521 );
or \U$34486 ( \42786 , \42783 , \42784 , \42785 );
buf \U$34487 ( \42787 , \42786 );
xor \U$34488 ( \42788 , \42782 , \42787 );
buf \U$34489 ( \42789 , \42788 );
xor \U$34490 ( \42790 , \42651 , \42789 );
and \U$34491 ( \42791 , \42546 , \42790 );
and \U$34493 ( \42792 , \42540 , \42545 );
or \U$34495 ( \42793 , 1'b0 , \42792 , 1'b0 );
xor \U$34496 ( \42794 , \42791 , \42793 );
and \U$34498 ( \42795 , \42533 , \42539 );
and \U$34499 ( \42796 , \42535 , \42539 );
or \U$34500 ( \42797 , 1'b0 , \42795 , \42796 );
xor \U$34501 ( \42798 , \42794 , \42797 );
xor \U$34508 ( \42799 , \42798 , 1'b0 );
and \U$34509 ( \42800 , \42645 , \42650 );
and \U$34510 ( \42801 , \42645 , \42789 );
and \U$34511 ( \42802 , \42650 , \42789 );
or \U$34512 ( \42803 , \42800 , \42801 , \42802 );
xor \U$34513 ( \42804 , \42799 , \42803 );
and \U$34514 ( \42805 , \42551 , \42556 );
and \U$34515 ( \42806 , \42551 , \42643 );
and \U$34516 ( \42807 , \42556 , \42643 );
or \U$34517 ( \42808 , \42805 , \42806 , \42807 );
buf \U$34518 ( \42809 , \42808 );
and \U$34519 ( \42810 , \42562 , \42635 );
and \U$34520 ( \42811 , \42562 , \42641 );
and \U$34521 ( \42812 , \42635 , \42641 );
or \U$34522 ( \42813 , \42810 , \42811 , \42812 );
buf \U$34523 ( \42814 , \42813 );
and \U$34524 ( \42815 , \42680 , \42686 );
and \U$34525 ( \42816 , \42680 , \42693 );
and \U$34526 ( \42817 , \42686 , \42693 );
or \U$34527 ( \42818 , \42815 , \42816 , \42817 );
buf \U$34528 ( \42819 , \42818 );
and \U$34529 ( \42820 , \17297 , \39334_nG9b7b );
and \U$34530 ( \42821 , \17294 , \39591_nG9b78 );
or \U$34531 ( \42822 , \42820 , \42821 );
xor \U$34532 ( \42823 , \17293 , \42822 );
buf \U$34533 ( \42824 , \42823 );
buf \U$34535 ( \42825 , \42824 );
xor \U$34536 ( \42826 , \42819 , \42825 );
and \U$34537 ( \42827 , \10707 , \42766_nG9b57 );
and \U$34538 ( \42828 , \42748 , \42752 );
and \U$34539 ( \42829 , \42752 , \42754 );
and \U$34540 ( \42830 , \42748 , \42754 );
or \U$34541 ( \42831 , \42828 , \42829 , \42830 );
and \U$34542 ( \42832 , \32794 , \32854 );
not \U$34543 ( \42833 , \42832 );
xnor \U$34544 ( \42834 , \42833 , \32805 );
xor \U$34545 ( \42835 , \42831 , \42834 );
and \U$34546 ( \42836 , \32054 , \32802 );
not \U$34547 ( \42837 , \42836 );
xor \U$34548 ( \42838 , \42835 , \42837 );
and \U$34549 ( \42839 , \42745 , \42746 );
and \U$34550 ( \42840 , \42746 , \42755 );
and \U$34551 ( \42841 , \42745 , \42755 );
or \U$34552 ( \42842 , \42839 , \42840 , \42841 );
xor \U$34553 ( \42843 , \42838 , \42842 );
and \U$34554 ( \42844 , \42756 , \42760 );
and \U$34555 ( \42845 , \42761 , \42764 );
or \U$34556 ( \42846 , \42844 , \42845 );
xor \U$34557 ( \42847 , \42843 , \42846 );
buf g9b54 ( \42848_nG9b54 , \42847 );
and \U$34558 ( \42849 , \10704 , \42848_nG9b54 );
or \U$34559 ( \42850 , \42827 , \42849 );
xor \U$34560 ( \42851 , \10703 , \42850 );
buf \U$34561 ( \42852 , \42851 );
buf \U$34563 ( \42853 , \42852 );
xor \U$34564 ( \42854 , \42826 , \42853 );
buf \U$34565 ( \42855 , \42854 );
and \U$34566 ( \42856 , \42733 , \42739 );
and \U$34567 ( \42857 , \42733 , \42771 );
and \U$34568 ( \42858 , \42739 , \42771 );
or \U$34569 ( \42859 , \42856 , \42857 , \42858 );
buf \U$34570 ( \42860 , \42859 );
xor \U$34571 ( \42861 , \42855 , \42860 );
and \U$34572 ( \42862 , \42702 , \42707 );
and \U$34573 ( \42863 , \42702 , \42713 );
and \U$34574 ( \42864 , \42707 , \42713 );
or \U$34575 ( \42865 , \42862 , \42863 , \42864 );
buf \U$34576 ( \42866 , \42865 );
xor \U$34577 ( \42867 , \42861 , \42866 );
buf \U$34578 ( \42868 , \42867 );
and \U$34579 ( \42869 , \28118 , \34294_nG9ba5 );
and \U$34580 ( \42870 , \28115 , \34643_nG9ba2 );
or \U$34581 ( \42871 , \42869 , \42870 );
xor \U$34582 ( \42872 , \28114 , \42871 );
buf \U$34583 ( \42873 , \42872 );
buf \U$34585 ( \42874 , \42873 );
and \U$34586 ( \42875 , \18702 , \38663_nG9b81 );
and \U$34587 ( \42876 , \18699 , \38968_nG9b7e );
or \U$34588 ( \42877 , \42875 , \42876 );
xor \U$34589 ( \42878 , \18698 , \42877 );
buf \U$34590 ( \42879 , \42878 );
buf \U$34592 ( \42880 , \42879 );
xor \U$34593 ( \42881 , \42874 , \42880 );
and \U$34594 ( \42882 , \13370 , \41040_nG9b69 );
and \U$34595 ( \42883 , \13367 , \41381_nG9b66 );
or \U$34596 ( \42884 , \42882 , \42883 );
xor \U$34597 ( \42885 , \13366 , \42884 );
buf \U$34598 ( \42886 , \42885 );
buf \U$34600 ( \42887 , \42886 );
xor \U$34601 ( \42888 , \42881 , \42887 );
buf \U$34602 ( \42889 , \42888 );
and \U$34603 ( \42890 , \42567 , \42573 );
buf \U$34604 ( \42891 , \42890 );
and \U$34606 ( \42892 , \32916 , \32179_nG9bb4 );
or \U$34607 ( \42893 , 1'b0 , \42892 );
xor \U$34608 ( \42894 , 1'b0 , \42893 );
buf \U$34609 ( \42895 , \42894 );
buf \U$34611 ( \42896 , \42895 );
and \U$34612 ( \42897 , \29853 , \33613_nG9bab );
and \U$34613 ( \42898 , \29850 , \34041_nG9ba8 );
or \U$34614 ( \42899 , \42897 , \42898 );
xor \U$34615 ( \42900 , \29849 , \42899 );
buf \U$34616 ( \42901 , \42900 );
buf \U$34618 ( \42902 , \42901 );
xor \U$34619 ( \42903 , \42896 , \42902 );
buf \U$34620 ( \42904 , \42903 );
xor \U$34621 ( \42905 , \42891 , \42904 );
and \U$34622 ( \42906 , \20155 , \37974_nG9b87 );
and \U$34623 ( \42907 , \20152 , \38337_nG9b84 );
or \U$34624 ( \42908 , \42906 , \42907 );
xor \U$34625 ( \42909 , \20151 , \42908 );
buf \U$34626 ( \42910 , \42909 );
buf \U$34628 ( \42911 , \42910 );
xor \U$34629 ( \42912 , \42905 , \42911 );
buf \U$34630 ( \42913 , \42912 );
xor \U$34631 ( \42914 , \42889 , \42913 );
and \U$34632 ( \42915 , \23201 , \36589_nG9b93 );
and \U$34633 ( \42916 , \23198 , \36986_nG9b90 );
or \U$34634 ( \42917 , \42915 , \42916 );
xor \U$34635 ( \42918 , \23197 , \42917 );
buf \U$34636 ( \42919 , \42918 );
buf \U$34638 ( \42920 , \42919 );
and \U$34639 ( \42921 , \21658 , \37250_nG9b8d );
and \U$34640 ( \42922 , \21655 , \37607_nG9b8a );
or \U$34641 ( \42923 , \42921 , \42922 );
xor \U$34642 ( \42924 , \21654 , \42923 );
buf \U$34643 ( \42925 , \42924 );
buf \U$34645 ( \42926 , \42925 );
xor \U$34646 ( \42927 , \42920 , \42926 );
and \U$34647 ( \42928 , \14631 , \40452_nG9b6f );
and \U$34648 ( \42929 , \14628 , \40843_nG9b6c );
or \U$34649 ( \42930 , \42928 , \42929 );
xor \U$34650 ( \42931 , \14627 , \42930 );
buf \U$34651 ( \42932 , \42931 );
buf \U$34653 ( \42933 , \42932 );
xor \U$34654 ( \42934 , \42927 , \42933 );
buf \U$34655 ( \42935 , \42934 );
xor \U$34656 ( \42936 , \42914 , \42935 );
buf \U$34657 ( \42937 , \42936 );
xor \U$34658 ( \42938 , \42868 , \42937 );
and \U$34659 ( \42939 , \42590 , \42611 );
and \U$34660 ( \42940 , \42590 , \42633 );
and \U$34661 ( \42941 , \42611 , \42633 );
or \U$34662 ( \42942 , \42939 , \42940 , \42941 );
buf \U$34663 ( \42943 , \42942 );
xor \U$34664 ( \42944 , \42938 , \42943 );
buf \U$34665 ( \42945 , \42944 );
xor \U$34666 ( \42946 , \42814 , \42945 );
and \U$34667 ( \42947 , \42723 , \42781 );
and \U$34668 ( \42948 , \42723 , \42787 );
and \U$34669 ( \42949 , \42781 , \42787 );
or \U$34670 ( \42950 , \42947 , \42948 , \42949 );
buf \U$34671 ( \42951 , \42950 );
xor \U$34672 ( \42952 , \42946 , \42951 );
buf \U$34673 ( \42953 , \42952 );
xor \U$34674 ( \42954 , \42809 , \42953 );
and \U$34675 ( \42955 , \42575 , \42581 );
and \U$34676 ( \42956 , \42575 , \42588 );
and \U$34677 ( \42957 , \42581 , \42588 );
or \U$34678 ( \42958 , \42955 , \42956 , \42957 );
buf \U$34679 ( \42959 , \42958 );
and \U$34680 ( \42960 , \42596 , \42602 );
and \U$34681 ( \42961 , \42596 , \42609 );
and \U$34682 ( \42962 , \42602 , \42609 );
or \U$34683 ( \42963 , \42960 , \42961 , \42962 );
buf \U$34684 ( \42964 , \42963 );
xor \U$34685 ( \42965 , \42959 , \42964 );
and \U$34686 ( \42966 , \42662 , \42668 );
and \U$34687 ( \42967 , \42662 , \42675 );
and \U$34688 ( \42968 , \42668 , \42675 );
or \U$34689 ( \42969 , \42966 , \42967 , \42968 );
buf \U$34690 ( \42970 , \42969 );
xor \U$34691 ( \42971 , \42965 , \42970 );
buf \U$34692 ( \42972 , \42971 );
and \U$34693 ( \42973 , \42656 , \42677 );
and \U$34694 ( \42974 , \42656 , \42695 );
and \U$34695 ( \42975 , \42677 , \42695 );
or \U$34696 ( \42976 , \42973 , \42974 , \42975 );
buf \U$34697 ( \42977 , \42976 );
xor \U$34698 ( \42978 , \42972 , \42977 );
and \U$34699 ( \42979 , \15940 , \39963_nG9b75 );
and \U$34700 ( \42980 , \15937 , \40204_nG9b72 );
or \U$34701 ( \42981 , \42979 , \42980 );
xor \U$34702 ( \42982 , \15936 , \42981 );
buf \U$34703 ( \42983 , \42982 );
buf \U$34705 ( \42984 , \42983 );
and \U$34706 ( \42985 , \12157 , \41685_nG9b63 );
and \U$34707 ( \42986 , \12154 , \41963_nG9b60 );
or \U$34708 ( \42987 , \42985 , \42986 );
xor \U$34709 ( \42988 , \12153 , \42987 );
buf \U$34710 ( \42989 , \42988 );
buf \U$34712 ( \42990 , \42989 );
xor \U$34713 ( \42991 , \42984 , \42990 );
and \U$34714 ( \42992 , \10421 , \42201_nG9b5d );
and \U$34715 ( \42993 , \10418 , \42433_nG9b5a );
or \U$34716 ( \42994 , \42992 , \42993 );
xor \U$34717 ( \42995 , \10417 , \42994 );
buf \U$34718 ( \42996 , \42995 );
buf \U$34720 ( \42997 , \42996 );
xor \U$34721 ( \42998 , \42991 , \42997 );
buf \U$34722 ( \42999 , \42998 );
and \U$34723 ( \43000 , \31636 , \32888_nG9bb1 );
and \U$34724 ( \43001 , \31633 , \33181_nG9bae );
or \U$34725 ( \43002 , \43000 , \43001 );
xor \U$34726 ( \43003 , \31632 , \43002 );
buf \U$34727 ( \43004 , \43003 );
buf \U$34729 ( \43005 , \43004 );
and \U$34730 ( \43006 , \26431 , \35094_nG9b9f );
and \U$34731 ( \43007 , \26428 , \35570_nG9b9c );
or \U$34732 ( \43008 , \43006 , \43007 );
xor \U$34733 ( \43009 , \26427 , \43008 );
buf \U$34734 ( \43010 , \43009 );
buf \U$34736 ( \43011 , \43010 );
xor \U$34737 ( \43012 , \43005 , \43011 );
and \U$34738 ( \43013 , \24792 , \35801_nG9b99 );
and \U$34739 ( \43014 , \24789 , \36172_nG9b96 );
or \U$34740 ( \43015 , \43013 , \43014 );
xor \U$34741 ( \43016 , \24788 , \43015 );
buf \U$34742 ( \43017 , \43016 );
buf \U$34744 ( \43018 , \43017 );
xor \U$34745 ( \43019 , \43012 , \43018 );
buf \U$34746 ( \43020 , \43019 );
xor \U$34747 ( \43021 , \42999 , \43020 );
and \U$34748 ( \43022 , \42618 , \42624 );
and \U$34749 ( \43023 , \42618 , \42631 );
and \U$34750 ( \43024 , \42624 , \42631 );
or \U$34751 ( \43025 , \43022 , \43023 , \43024 );
buf \U$34752 ( \43026 , \43025 );
xor \U$34753 ( \43027 , \43021 , \43026 );
buf \U$34754 ( \43028 , \43027 );
xor \U$34755 ( \43029 , \42978 , \43028 );
buf \U$34756 ( \43030 , \43029 );
and \U$34757 ( \43031 , \42697 , \42715 );
and \U$34758 ( \43032 , \42697 , \42721 );
and \U$34759 ( \43033 , \42715 , \42721 );
or \U$34760 ( \43034 , \43031 , \43032 , \43033 );
buf \U$34761 ( \43035 , \43034 );
xor \U$34762 ( \43036 , \43030 , \43035 );
and \U$34763 ( \43037 , \42728 , \42773 );
and \U$34764 ( \43038 , \42728 , \42779 );
and \U$34765 ( \43039 , \42773 , \42779 );
or \U$34766 ( \43040 , \43037 , \43038 , \43039 );
buf \U$34767 ( \43041 , \43040 );
xor \U$34768 ( \43042 , \43036 , \43041 );
buf \U$34769 ( \43043 , \43042 );
xor \U$34770 ( \43044 , \42954 , \43043 );
and \U$34771 ( \43045 , \42804 , \43044 );
and \U$34773 ( \43046 , \42798 , \42803 );
or \U$34775 ( \43047 , 1'b0 , \43046 , 1'b0 );
xor \U$34776 ( \43048 , \43045 , \43047 );
and \U$34778 ( \43049 , \42791 , \42797 );
and \U$34779 ( \43050 , \42793 , \42797 );
or \U$34780 ( \43051 , 1'b0 , \43049 , \43050 );
xor \U$34781 ( \43052 , \43048 , \43051 );
xor \U$34788 ( \43053 , \43052 , 1'b0 );
and \U$34789 ( \43054 , \42809 , \42953 );
and \U$34790 ( \43055 , \42809 , \43043 );
and \U$34791 ( \43056 , \42953 , \43043 );
or \U$34792 ( \43057 , \43054 , \43055 , \43056 );
xor \U$34793 ( \43058 , \43053 , \43057 );
and \U$34794 ( \43059 , \42999 , \43020 );
and \U$34795 ( \43060 , \42999 , \43026 );
and \U$34796 ( \43061 , \43020 , \43026 );
or \U$34797 ( \43062 , \43059 , \43060 , \43061 );
buf \U$34798 ( \43063 , \43062 );
and \U$34799 ( \43064 , \42891 , \42904 );
and \U$34800 ( \43065 , \42891 , \42911 );
and \U$34801 ( \43066 , \42904 , \42911 );
or \U$34802 ( \43067 , \43064 , \43065 , \43066 );
buf \U$34803 ( \43068 , \43067 );
and \U$34804 ( \43069 , \42874 , \42880 );
and \U$34805 ( \43070 , \42874 , \42887 );
and \U$34806 ( \43071 , \42880 , \42887 );
or \U$34807 ( \43072 , \43069 , \43070 , \43071 );
buf \U$34808 ( \43073 , \43072 );
xor \U$34809 ( \43074 , \43068 , \43073 );
and \U$34810 ( \43075 , \29853 , \34041_nG9ba8 );
and \U$34811 ( \43076 , \29850 , \34294_nG9ba5 );
or \U$34812 ( \43077 , \43075 , \43076 );
xor \U$34813 ( \43078 , \29849 , \43077 );
buf \U$34814 ( \43079 , \43078 );
buf \U$34816 ( \43080 , \43079 );
and \U$34817 ( \43081 , \28118 , \34643_nG9ba2 );
and \U$34818 ( \43082 , \28115 , \35094_nG9b9f );
or \U$34819 ( \43083 , \43081 , \43082 );
xor \U$34820 ( \43084 , \28114 , \43083 );
buf \U$34821 ( \43085 , \43084 );
buf \U$34823 ( \43086 , \43085 );
xor \U$34824 ( \43087 , \43080 , \43086 );
and \U$34825 ( \43088 , \26431 , \35570_nG9b9c );
and \U$34826 ( \43089 , \26428 , \35801_nG9b99 );
or \U$34827 ( \43090 , \43088 , \43089 );
xor \U$34828 ( \43091 , \26427 , \43090 );
buf \U$34829 ( \43092 , \43091 );
buf \U$34831 ( \43093 , \43092 );
xor \U$34832 ( \43094 , \43087 , \43093 );
buf \U$34833 ( \43095 , \43094 );
xor \U$34834 ( \43096 , \43074 , \43095 );
buf \U$34835 ( \43097 , \43096 );
xor \U$34836 ( \43098 , \43063 , \43097 );
and \U$34837 ( \43099 , \24792 , \36172_nG9b96 );
and \U$34838 ( \43100 , \24789 , \36589_nG9b93 );
or \U$34839 ( \43101 , \43099 , \43100 );
xor \U$34840 ( \43102 , \24788 , \43101 );
buf \U$34841 ( \43103 , \43102 );
buf \U$34843 ( \43104 , \43103 );
and \U$34844 ( \43105 , \17297 , \39591_nG9b78 );
and \U$34845 ( \43106 , \17294 , \39963_nG9b75 );
or \U$34846 ( \43107 , \43105 , \43106 );
xor \U$34847 ( \43108 , \17293 , \43107 );
buf \U$34848 ( \43109 , \43108 );
buf \U$34850 ( \43110 , \43109 );
xor \U$34851 ( \43111 , \43104 , \43110 );
and \U$34852 ( \43112 , \15940 , \40204_nG9b72 );
and \U$34853 ( \43113 , \15937 , \40452_nG9b6f );
or \U$34854 ( \43114 , \43112 , \43113 );
xor \U$34855 ( \43115 , \15936 , \43114 );
buf \U$34856 ( \43116 , \43115 );
buf \U$34858 ( \43117 , \43116 );
xor \U$34859 ( \43118 , \43111 , \43117 );
buf \U$34860 ( \43119 , \43118 );
and \U$34861 ( \43120 , \42984 , \42990 );
and \U$34862 ( \43121 , \42984 , \42997 );
and \U$34863 ( \43122 , \42990 , \42997 );
or \U$34864 ( \43123 , \43120 , \43121 , \43122 );
buf \U$34865 ( \43124 , \43123 );
xor \U$34866 ( \43125 , \43119 , \43124 );
and \U$34867 ( \43126 , \42920 , \42926 );
and \U$34868 ( \43127 , \42920 , \42933 );
and \U$34869 ( \43128 , \42926 , \42933 );
or \U$34870 ( \43129 , \43126 , \43127 , \43128 );
buf \U$34871 ( \43130 , \43129 );
xor \U$34872 ( \43131 , \43125 , \43130 );
buf \U$34873 ( \43132 , \43131 );
xor \U$34874 ( \43133 , \43098 , \43132 );
buf \U$34875 ( \43134 , \43133 );
and \U$34876 ( \43135 , \42972 , \42977 );
and \U$34877 ( \43136 , \42972 , \43028 );
and \U$34878 ( \43137 , \42977 , \43028 );
or \U$34879 ( \43138 , \43135 , \43136 , \43137 );
buf \U$34880 ( \43139 , \43138 );
xor \U$34881 ( \43140 , \43134 , \43139 );
and \U$34882 ( \43141 , \42855 , \42860 );
and \U$34883 ( \43142 , \42855 , \42866 );
and \U$34884 ( \43143 , \42860 , \42866 );
or \U$34885 ( \43144 , \43141 , \43142 , \43143 );
buf \U$34886 ( \43145 , \43144 );
xor \U$34887 ( \43146 , \43140 , \43145 );
buf \U$34888 ( \43147 , \43146 );
and \U$34889 ( \43148 , \42868 , \42937 );
and \U$34890 ( \43149 , \42868 , \42943 );
and \U$34891 ( \43150 , \42937 , \42943 );
or \U$34892 ( \43151 , \43148 , \43149 , \43150 );
buf \U$34893 ( \43152 , \43151 );
xor \U$34894 ( \43153 , \43147 , \43152 );
and \U$34895 ( \43154 , \42959 , \42964 );
and \U$34896 ( \43155 , \42959 , \42970 );
and \U$34897 ( \43156 , \42964 , \42970 );
or \U$34898 ( \43157 , \43154 , \43155 , \43156 );
buf \U$34899 ( \43158 , \43157 );
and \U$34900 ( \43159 , \43005 , \43011 );
and \U$34901 ( \43160 , \43005 , \43018 );
and \U$34902 ( \43161 , \43011 , \43018 );
or \U$34903 ( \43162 , \43159 , \43160 , \43161 );
buf \U$34904 ( \43163 , \43162 );
and \U$34905 ( \43164 , \10707 , \42848_nG9b54 );
and \U$34906 ( \43165 , \42831 , \42834 );
and \U$34907 ( \43166 , \42834 , \42837 );
and \U$34908 ( \43167 , \42831 , \42837 );
or \U$34909 ( \43168 , \43165 , \43166 , \43167 );
buf \U$34910 ( \43169 , \42836 );
not \U$34911 ( \43170 , \32805 );
xor \U$34912 ( \43171 , \43169 , \43170 );
and \U$34913 ( \43172 , \32794 , \32802 );
xor \U$34914 ( \43173 , \43171 , \43172 );
xor \U$34915 ( \43174 , \43168 , \43173 );
and \U$34916 ( \43175 , \42838 , \42842 );
and \U$34917 ( \43176 , \42843 , \42846 );
or \U$34918 ( \43177 , \43175 , \43176 );
xor \U$34919 ( \43178 , \43174 , \43177 );
buf g9b51 ( \43179_nG9b51 , \43178 );
and \U$34920 ( \43180 , \10704 , \43179_nG9b51 );
or \U$34921 ( \43181 , \43164 , \43180 );
xor \U$34922 ( \43182 , \10703 , \43181 );
buf \U$34923 ( \43183 , \43182 );
buf \U$34925 ( \43184 , \43183 );
xor \U$34926 ( \43185 , \43163 , \43184 );
and \U$34927 ( \43186 , \10421 , \42433_nG9b5a );
and \U$34928 ( \43187 , \10418 , \42766_nG9b57 );
or \U$34929 ( \43188 , \43186 , \43187 );
xor \U$34930 ( \43189 , \10417 , \43188 );
buf \U$34931 ( \43190 , \43189 );
buf \U$34933 ( \43191 , \43190 );
xor \U$34934 ( \43192 , \43185 , \43191 );
buf \U$34935 ( \43193 , \43192 );
xor \U$34936 ( \43194 , \43158 , \43193 );
and \U$34937 ( \43195 , \42819 , \42825 );
and \U$34938 ( \43196 , \42819 , \42853 );
and \U$34939 ( \43197 , \42825 , \42853 );
or \U$34940 ( \43198 , \43195 , \43196 , \43197 );
buf \U$34941 ( \43199 , \43198 );
xor \U$34942 ( \43200 , \43194 , \43199 );
buf \U$34943 ( \43201 , \43200 );
and \U$34944 ( \43202 , \42889 , \42913 );
and \U$34945 ( \43203 , \42889 , \42935 );
and \U$34946 ( \43204 , \42913 , \42935 );
or \U$34947 ( \43205 , \43202 , \43203 , \43204 );
buf \U$34948 ( \43206 , \43205 );
xor \U$34949 ( \43207 , \43201 , \43206 );
and \U$34951 ( \43208 , \32916 , \32888_nG9bb1 );
or \U$34952 ( \43209 , 1'b0 , \43208 );
xor \U$34953 ( \43210 , 1'b0 , \43209 );
buf \U$34954 ( \43211 , \43210 );
buf \U$34956 ( \43212 , \43211 );
and \U$34957 ( \43213 , \31636 , \33181_nG9bae );
and \U$34958 ( \43214 , \31633 , \33613_nG9bab );
or \U$34959 ( \43215 , \43213 , \43214 );
xor \U$34960 ( \43216 , \31632 , \43215 );
buf \U$34961 ( \43217 , \43216 );
buf \U$34963 ( \43218 , \43217 );
xor \U$34964 ( \43219 , \43212 , \43218 );
buf \U$34965 ( \43220 , \43219 );
and \U$34966 ( \43221 , \18702 , \38968_nG9b7e );
and \U$34967 ( \43222 , \18699 , \39334_nG9b7b );
or \U$34968 ( \43223 , \43221 , \43222 );
xor \U$34969 ( \43224 , \18698 , \43223 );
buf \U$34970 ( \43225 , \43224 );
buf \U$34972 ( \43226 , \43225 );
xor \U$34973 ( \43227 , \43220 , \43226 );
and \U$34974 ( \43228 , \13370 , \41381_nG9b66 );
and \U$34975 ( \43229 , \13367 , \41685_nG9b63 );
or \U$34976 ( \43230 , \43228 , \43229 );
xor \U$34977 ( \43231 , \13366 , \43230 );
buf \U$34978 ( \43232 , \43231 );
buf \U$34980 ( \43233 , \43232 );
xor \U$34981 ( \43234 , \43227 , \43233 );
buf \U$34982 ( \43235 , \43234 );
and \U$34983 ( \43236 , \23201 , \36986_nG9b90 );
and \U$34984 ( \43237 , \23198 , \37250_nG9b8d );
or \U$34985 ( \43238 , \43236 , \43237 );
xor \U$34986 ( \43239 , \23197 , \43238 );
buf \U$34987 ( \43240 , \43239 );
buf \U$34989 ( \43241 , \43240 );
and \U$34990 ( \43242 , \21658 , \37607_nG9b8a );
and \U$34991 ( \43243 , \21655 , \37974_nG9b87 );
or \U$34992 ( \43244 , \43242 , \43243 );
xor \U$34993 ( \43245 , \21654 , \43244 );
buf \U$34994 ( \43246 , \43245 );
buf \U$34996 ( \43247 , \43246 );
xor \U$34997 ( \43248 , \43241 , \43247 );
and \U$34998 ( \43249 , \12157 , \41963_nG9b60 );
and \U$34999 ( \43250 , \12154 , \42201_nG9b5d );
or \U$35000 ( \43251 , \43249 , \43250 );
xor \U$35001 ( \43252 , \12153 , \43251 );
buf \U$35002 ( \43253 , \43252 );
buf \U$35004 ( \43254 , \43253 );
xor \U$35005 ( \43255 , \43248 , \43254 );
buf \U$35006 ( \43256 , \43255 );
xor \U$35007 ( \43257 , \43235 , \43256 );
and \U$35008 ( \43258 , \42896 , \42902 );
buf \U$35009 ( \43259 , \43258 );
and \U$35010 ( \43260 , \20155 , \38337_nG9b84 );
and \U$35011 ( \43261 , \20152 , \38663_nG9b81 );
or \U$35012 ( \43262 , \43260 , \43261 );
xor \U$35013 ( \43263 , \20151 , \43262 );
buf \U$35014 ( \43264 , \43263 );
buf \U$35016 ( \43265 , \43264 );
xor \U$35017 ( \43266 , \43259 , \43265 );
and \U$35018 ( \43267 , \14631 , \40843_nG9b6c );
and \U$35019 ( \43268 , \14628 , \41040_nG9b69 );
or \U$35020 ( \43269 , \43267 , \43268 );
xor \U$35021 ( \43270 , \14627 , \43269 );
buf \U$35022 ( \43271 , \43270 );
buf \U$35024 ( \43272 , \43271 );
xor \U$35025 ( \43273 , \43266 , \43272 );
buf \U$35026 ( \43274 , \43273 );
xor \U$35027 ( \43275 , \43257 , \43274 );
buf \U$35028 ( \43276 , \43275 );
xor \U$35029 ( \43277 , \43207 , \43276 );
buf \U$35030 ( \43278 , \43277 );
xor \U$35031 ( \43279 , \43153 , \43278 );
buf \U$35032 ( \43280 , \43279 );
and \U$35033 ( \43281 , \42814 , \42945 );
and \U$35034 ( \43282 , \42814 , \42951 );
and \U$35035 ( \43283 , \42945 , \42951 );
or \U$35036 ( \43284 , \43281 , \43282 , \43283 );
buf \U$35037 ( \43285 , \43284 );
xor \U$35038 ( \43286 , \43280 , \43285 );
and \U$35039 ( \43287 , \43030 , \43035 );
and \U$35040 ( \43288 , \43030 , \43041 );
and \U$35041 ( \43289 , \43035 , \43041 );
or \U$35042 ( \43290 , \43287 , \43288 , \43289 );
buf \U$35043 ( \43291 , \43290 );
xor \U$35044 ( \43292 , \43286 , \43291 );
and \U$35045 ( \43293 , \43058 , \43292 );
and \U$35047 ( \43294 , \43052 , \43057 );
or \U$35049 ( \43295 , 1'b0 , \43294 , 1'b0 );
xor \U$35050 ( \43296 , \43293 , \43295 );
and \U$35052 ( \43297 , \43045 , \43051 );
and \U$35053 ( \43298 , \43047 , \43051 );
or \U$35054 ( \43299 , 1'b0 , \43297 , \43298 );
xor \U$35055 ( \43300 , \43296 , \43299 );
xor \U$35062 ( \43301 , \43300 , 1'b0 );
and \U$35063 ( \43302 , \43280 , \43285 );
and \U$35064 ( \43303 , \43280 , \43291 );
and \U$35065 ( \43304 , \43285 , \43291 );
or \U$35066 ( \43305 , \43302 , \43303 , \43304 );
xor \U$35067 ( \43306 , \43301 , \43305 );
and \U$35068 ( \43307 , \43147 , \43152 );
and \U$35069 ( \43308 , \43147 , \43278 );
and \U$35070 ( \43309 , \43152 , \43278 );
or \U$35071 ( \43310 , \43307 , \43308 , \43309 );
buf \U$35072 ( \43311 , \43310 );
and \U$35073 ( \43312 , \43134 , \43139 );
and \U$35074 ( \43313 , \43134 , \43145 );
and \U$35075 ( \43314 , \43139 , \43145 );
or \U$35076 ( \43315 , \43312 , \43313 , \43314 );
buf \U$35077 ( \43316 , \43315 );
xor \U$35078 ( \43317 , \43311 , \43316 );
and \U$35079 ( \43318 , \43201 , \43206 );
and \U$35080 ( \43319 , \43201 , \43276 );
and \U$35081 ( \43320 , \43206 , \43276 );
or \U$35082 ( \43321 , \43318 , \43319 , \43320 );
buf \U$35083 ( \43322 , \43321 );
and \U$35085 ( \43323 , \32916 , \33181_nG9bae );
or \U$35086 ( \43324 , 1'b0 , \43323 );
xor \U$35087 ( \43325 , 1'b0 , \43324 );
buf \U$35088 ( \43326 , \43325 );
buf \U$35090 ( \43327 , \43326 );
and \U$35091 ( \43328 , \31636 , \33613_nG9bab );
and \U$35092 ( \43329 , \31633 , \34041_nG9ba8 );
or \U$35093 ( \43330 , \43328 , \43329 );
xor \U$35094 ( \43331 , \31632 , \43330 );
buf \U$35095 ( \43332 , \43331 );
buf \U$35097 ( \43333 , \43332 );
xor \U$35098 ( \43334 , \43327 , \43333 );
buf \U$35099 ( \43335 , \43334 );
and \U$35100 ( \43336 , \18702 , \39334_nG9b7b );
and \U$35101 ( \43337 , \18699 , \39591_nG9b78 );
or \U$35102 ( \43338 , \43336 , \43337 );
xor \U$35103 ( \43339 , \18698 , \43338 );
buf \U$35104 ( \43340 , \43339 );
buf \U$35106 ( \43341 , \43340 );
xor \U$35107 ( \43342 , \43335 , \43341 );
and \U$35108 ( \43343 , \13370 , \41685_nG9b63 );
and \U$35109 ( \43344 , \13367 , \41963_nG9b60 );
or \U$35110 ( \43345 , \43343 , \43344 );
xor \U$35111 ( \43346 , \13366 , \43345 );
buf \U$35112 ( \43347 , \43346 );
buf \U$35114 ( \43348 , \43347 );
xor \U$35115 ( \43349 , \43342 , \43348 );
buf \U$35116 ( \43350 , \43349 );
and \U$35117 ( \43351 , \23201 , \37250_nG9b8d );
and \U$35118 ( \43352 , \23198 , \37607_nG9b8a );
or \U$35119 ( \43353 , \43351 , \43352 );
xor \U$35120 ( \43354 , \23197 , \43353 );
buf \U$35121 ( \43355 , \43354 );
buf \U$35123 ( \43356 , \43355 );
and \U$35124 ( \43357 , \21658 , \37974_nG9b87 );
and \U$35125 ( \43358 , \21655 , \38337_nG9b84 );
or \U$35126 ( \43359 , \43357 , \43358 );
xor \U$35127 ( \43360 , \21654 , \43359 );
buf \U$35128 ( \43361 , \43360 );
buf \U$35130 ( \43362 , \43361 );
xor \U$35131 ( \43363 , \43356 , \43362 );
and \U$35132 ( \43364 , \12157 , \42201_nG9b5d );
and \U$35133 ( \43365 , \12154 , \42433_nG9b5a );
or \U$35134 ( \43366 , \43364 , \43365 );
xor \U$35135 ( \43367 , \12153 , \43366 );
buf \U$35136 ( \43368 , \43367 );
buf \U$35138 ( \43369 , \43368 );
xor \U$35139 ( \43370 , \43363 , \43369 );
buf \U$35140 ( \43371 , \43370 );
xor \U$35141 ( \43372 , \43350 , \43371 );
and \U$35142 ( \43373 , \43212 , \43218 );
buf \U$35143 ( \43374 , \43373 );
and \U$35144 ( \43375 , \20155 , \38663_nG9b81 );
and \U$35145 ( \43376 , \20152 , \38968_nG9b7e );
or \U$35146 ( \43377 , \43375 , \43376 );
xor \U$35147 ( \43378 , \20151 , \43377 );
buf \U$35148 ( \43379 , \43378 );
buf \U$35150 ( \43380 , \43379 );
xor \U$35151 ( \43381 , \43374 , \43380 );
and \U$35152 ( \43382 , \14631 , \41040_nG9b69 );
and \U$35153 ( \43383 , \14628 , \41381_nG9b66 );
or \U$35154 ( \43384 , \43382 , \43383 );
xor \U$35155 ( \43385 , \14627 , \43384 );
buf \U$35156 ( \43386 , \43385 );
buf \U$35158 ( \43387 , \43386 );
xor \U$35159 ( \43388 , \43381 , \43387 );
buf \U$35160 ( \43389 , \43388 );
xor \U$35161 ( \43390 , \43372 , \43389 );
buf \U$35162 ( \43391 , \43390 );
and \U$35163 ( \43392 , \43068 , \43073 );
and \U$35164 ( \43393 , \43068 , \43095 );
and \U$35165 ( \43394 , \43073 , \43095 );
or \U$35166 ( \43395 , \43392 , \43393 , \43394 );
buf \U$35167 ( \43396 , \43395 );
and \U$35168 ( \43397 , \43080 , \43086 );
and \U$35169 ( \43398 , \43080 , \43093 );
and \U$35170 ( \43399 , \43086 , \43093 );
or \U$35171 ( \43400 , \43397 , \43398 , \43399 );
buf \U$35172 ( \43401 , \43400 );
and \U$35173 ( \43402 , \10707 , \43179_nG9b51 );
or \U$35176 ( \43403 , \43402 , 1'b0 );
xor \U$35177 ( \43404 , \10703 , \43403 );
buf \U$35178 ( \43405 , \43404 );
buf \U$35180 ( \43406 , \43405 );
xor \U$35181 ( \43407 , \43401 , \43406 );
and \U$35182 ( \43408 , \10421 , \42766_nG9b57 );
and \U$35183 ( \43409 , \10418 , \42848_nG9b54 );
or \U$35184 ( \43410 , \43408 , \43409 );
xor \U$35185 ( \43411 , \10417 , \43410 );
buf \U$35186 ( \43412 , \43411 );
buf \U$35188 ( \43413 , \43412 );
xor \U$35189 ( \43414 , \43407 , \43413 );
buf \U$35190 ( \43415 , \43414 );
xor \U$35191 ( \43416 , \43396 , \43415 );
and \U$35192 ( \43417 , \43163 , \43184 );
and \U$35193 ( \43418 , \43163 , \43191 );
and \U$35194 ( \43419 , \43184 , \43191 );
or \U$35195 ( \43420 , \43417 , \43418 , \43419 );
buf \U$35196 ( \43421 , \43420 );
xor \U$35197 ( \43422 , \43416 , \43421 );
buf \U$35198 ( \43423 , \43422 );
xor \U$35199 ( \43424 , \43391 , \43423 );
and \U$35200 ( \43425 , \43235 , \43256 );
and \U$35201 ( \43426 , \43235 , \43274 );
and \U$35202 ( \43427 , \43256 , \43274 );
or \U$35203 ( \43428 , \43425 , \43426 , \43427 );
buf \U$35204 ( \43429 , \43428 );
xor \U$35205 ( \43430 , \43424 , \43429 );
buf \U$35206 ( \43431 , \43430 );
xor \U$35207 ( \43432 , \43322 , \43431 );
and \U$35208 ( \43433 , \43158 , \43193 );
and \U$35209 ( \43434 , \43158 , \43199 );
and \U$35210 ( \43435 , \43193 , \43199 );
or \U$35211 ( \43436 , \43433 , \43434 , \43435 );
buf \U$35212 ( \43437 , \43436 );
and \U$35213 ( \43438 , \43063 , \43097 );
and \U$35214 ( \43439 , \43063 , \43132 );
and \U$35215 ( \43440 , \43097 , \43132 );
or \U$35216 ( \43441 , \43438 , \43439 , \43440 );
buf \U$35217 ( \43442 , \43441 );
xor \U$35218 ( \43443 , \43437 , \43442 );
and \U$35219 ( \43444 , \43119 , \43124 );
and \U$35220 ( \43445 , \43119 , \43130 );
and \U$35221 ( \43446 , \43124 , \43130 );
or \U$35222 ( \43447 , \43444 , \43445 , \43446 );
buf \U$35223 ( \43448 , \43447 );
and \U$35224 ( \43449 , \43259 , \43265 );
and \U$35225 ( \43450 , \43259 , \43272 );
and \U$35226 ( \43451 , \43265 , \43272 );
or \U$35227 ( \43452 , \43449 , \43450 , \43451 );
buf \U$35228 ( \43453 , \43452 );
and \U$35229 ( \43454 , \29853 , \34294_nG9ba5 );
and \U$35230 ( \43455 , \29850 , \34643_nG9ba2 );
or \U$35231 ( \43456 , \43454 , \43455 );
xor \U$35232 ( \43457 , \29849 , \43456 );
buf \U$35233 ( \43458 , \43457 );
buf \U$35235 ( \43459 , \43458 );
and \U$35236 ( \43460 , \28118 , \35094_nG9b9f );
and \U$35237 ( \43461 , \28115 , \35570_nG9b9c );
or \U$35238 ( \43462 , \43460 , \43461 );
xor \U$35239 ( \43463 , \28114 , \43462 );
buf \U$35240 ( \43464 , \43463 );
buf \U$35242 ( \43465 , \43464 );
xor \U$35243 ( \43466 , \43459 , \43465 );
and \U$35244 ( \43467 , \26431 , \35801_nG9b99 );
and \U$35245 ( \43468 , \26428 , \36172_nG9b96 );
or \U$35246 ( \43469 , \43467 , \43468 );
xor \U$35247 ( \43470 , \26427 , \43469 );
buf \U$35248 ( \43471 , \43470 );
buf \U$35250 ( \43472 , \43471 );
xor \U$35251 ( \43473 , \43466 , \43472 );
buf \U$35252 ( \43474 , \43473 );
xor \U$35253 ( \43475 , \43453 , \43474 );
and \U$35254 ( \43476 , \43220 , \43226 );
and \U$35255 ( \43477 , \43220 , \43233 );
and \U$35256 ( \43478 , \43226 , \43233 );
or \U$35257 ( \43479 , \43476 , \43477 , \43478 );
buf \U$35258 ( \43480 , \43479 );
xor \U$35259 ( \43481 , \43475 , \43480 );
buf \U$35260 ( \43482 , \43481 );
xor \U$35261 ( \43483 , \43448 , \43482 );
and \U$35262 ( \43484 , \43104 , \43110 );
and \U$35263 ( \43485 , \43104 , \43117 );
and \U$35264 ( \43486 , \43110 , \43117 );
or \U$35265 ( \43487 , \43484 , \43485 , \43486 );
buf \U$35266 ( \43488 , \43487 );
and \U$35267 ( \43489 , \24792 , \36589_nG9b93 );
and \U$35268 ( \43490 , \24789 , \36986_nG9b90 );
or \U$35269 ( \43491 , \43489 , \43490 );
xor \U$35270 ( \43492 , \24788 , \43491 );
buf \U$35271 ( \43493 , \43492 );
buf \U$35273 ( \43494 , \43493 );
and \U$35274 ( \43495 , \17297 , \39963_nG9b75 );
and \U$35275 ( \43496 , \17294 , \40204_nG9b72 );
or \U$35276 ( \43497 , \43495 , \43496 );
xor \U$35277 ( \43498 , \17293 , \43497 );
buf \U$35278 ( \43499 , \43498 );
buf \U$35280 ( \43500 , \43499 );
xor \U$35281 ( \43501 , \43494 , \43500 );
and \U$35282 ( \43502 , \15940 , \40452_nG9b6f );
and \U$35283 ( \43503 , \15937 , \40843_nG9b6c );
or \U$35284 ( \43504 , \43502 , \43503 );
xor \U$35285 ( \43505 , \15936 , \43504 );
buf \U$35286 ( \43506 , \43505 );
buf \U$35288 ( \43507 , \43506 );
xor \U$35289 ( \43508 , \43501 , \43507 );
buf \U$35290 ( \43509 , \43508 );
xor \U$35291 ( \43510 , \43488 , \43509 );
and \U$35292 ( \43511 , \43241 , \43247 );
and \U$35293 ( \43512 , \43241 , \43254 );
and \U$35294 ( \43513 , \43247 , \43254 );
or \U$35295 ( \43514 , \43511 , \43512 , \43513 );
buf \U$35296 ( \43515 , \43514 );
xor \U$35297 ( \43516 , \43510 , \43515 );
buf \U$35298 ( \43517 , \43516 );
xor \U$35299 ( \43518 , \43483 , \43517 );
buf \U$35300 ( \43519 , \43518 );
xor \U$35301 ( \43520 , \43443 , \43519 );
buf \U$35302 ( \43521 , \43520 );
xor \U$35303 ( \43522 , \43432 , \43521 );
buf \U$35304 ( \43523 , \43522 );
xor \U$35305 ( \43524 , \43317 , \43523 );
and \U$35306 ( \43525 , \43306 , \43524 );
and \U$35308 ( \43526 , \43300 , \43305 );
or \U$35310 ( \43527 , 1'b0 , \43526 , 1'b0 );
xor \U$35311 ( \43528 , \43525 , \43527 );
and \U$35313 ( \43529 , \43293 , \43299 );
and \U$35314 ( \43530 , \43295 , \43299 );
or \U$35315 ( \43531 , 1'b0 , \43529 , \43530 );
xor \U$35316 ( \43532 , \43528 , \43531 );
xor \U$35323 ( \43533 , \43532 , 1'b0 );
and \U$35324 ( \43534 , \43311 , \43316 );
and \U$35325 ( \43535 , \43311 , \43523 );
and \U$35326 ( \43536 , \43316 , \43523 );
or \U$35327 ( \43537 , \43534 , \43535 , \43536 );
xor \U$35328 ( \43538 , \43533 , \43537 );
and \U$35329 ( \43539 , \43322 , \43431 );
and \U$35330 ( \43540 , \43322 , \43521 );
and \U$35331 ( \43541 , \43431 , \43521 );
or \U$35332 ( \43542 , \43539 , \43540 , \43541 );
buf \U$35333 ( \43543 , \43542 );
and \U$35334 ( \43544 , \43437 , \43442 );
and \U$35335 ( \43545 , \43437 , \43519 );
and \U$35336 ( \43546 , \43442 , \43519 );
or \U$35337 ( \43547 , \43544 , \43545 , \43546 );
buf \U$35338 ( \43548 , \43547 );
and \U$35339 ( \43549 , \43350 , \43371 );
and \U$35340 ( \43550 , \43350 , \43389 );
and \U$35341 ( \43551 , \43371 , \43389 );
or \U$35342 ( \43552 , \43549 , \43550 , \43551 );
buf \U$35343 ( \43553 , \43552 );
and \U$35344 ( \43554 , \43453 , \43474 );
and \U$35345 ( \43555 , \43453 , \43480 );
and \U$35346 ( \43556 , \43474 , \43480 );
or \U$35347 ( \43557 , \43554 , \43555 , \43556 );
buf \U$35348 ( \43558 , \43557 );
and \U$35349 ( \43559 , \43459 , \43465 );
and \U$35350 ( \43560 , \43459 , \43472 );
and \U$35351 ( \43561 , \43465 , \43472 );
or \U$35352 ( \43562 , \43559 , \43560 , \43561 );
buf \U$35353 ( \43563 , \43562 );
xor \U$35358 ( \43564 , \10703 , 1'b0 );
not \U$35359 ( \43565 , \43564 );
buf \U$35360 ( \43566 , \43565 );
buf \U$35362 ( \43567 , \43566 );
xor \U$35363 ( \43568 , 1'b1 , \43567 );
and \U$35365 ( \43569 , \32916 , \33613_nG9bab );
or \U$35366 ( \43570 , 1'b0 , \43569 );
xor \U$35367 ( \43571 , 1'b0 , \43570 );
buf \U$35368 ( \43572 , \43571 );
buf \U$35370 ( \43573 , \43572 );
xor \U$35371 ( \43574 , \43568 , \43573 );
buf \U$35372 ( \43575 , \43574 );
xor \U$35373 ( \43576 , \43563 , \43575 );
and \U$35374 ( \43577 , \12157 , \42433_nG9b5a );
and \U$35375 ( \43578 , \12154 , \42766_nG9b57 );
or \U$35376 ( \43579 , \43577 , \43578 );
xor \U$35377 ( \43580 , \12153 , \43579 );
buf \U$35378 ( \43581 , \43580 );
buf \U$35380 ( \43582 , \43581 );
xor \U$35381 ( \43583 , \43576 , \43582 );
buf \U$35382 ( \43584 , \43583 );
xor \U$35383 ( \43585 , \43558 , \43584 );
and \U$35384 ( \43586 , \43401 , \43406 );
and \U$35385 ( \43587 , \43401 , \43413 );
and \U$35386 ( \43588 , \43406 , \43413 );
or \U$35387 ( \43589 , \43586 , \43587 , \43588 );
buf \U$35388 ( \43590 , \43589 );
xor \U$35389 ( \43591 , \43585 , \43590 );
buf \U$35390 ( \43592 , \43591 );
xor \U$35391 ( \43593 , \43553 , \43592 );
and \U$35392 ( \43594 , \43327 , \43333 );
buf \U$35393 ( \43595 , \43594 );
and \U$35394 ( \43596 , \20155 , \38968_nG9b7e );
and \U$35395 ( \43597 , \20152 , \39334_nG9b7b );
or \U$35396 ( \43598 , \43596 , \43597 );
xor \U$35397 ( \43599 , \20151 , \43598 );
buf \U$35398 ( \43600 , \43599 );
buf \U$35400 ( \43601 , \43600 );
xor \U$35401 ( \43602 , \43595 , \43601 );
and \U$35402 ( \43603 , \14631 , \41381_nG9b66 );
and \U$35403 ( \43604 , \14628 , \41685_nG9b63 );
or \U$35404 ( \43605 , \43603 , \43604 );
xor \U$35405 ( \43606 , \14627 , \43605 );
buf \U$35406 ( \43607 , \43606 );
buf \U$35408 ( \43608 , \43607 );
xor \U$35409 ( \43609 , \43602 , \43608 );
buf \U$35410 ( \43610 , \43609 );
and \U$35411 ( \43611 , \10421 , \42848_nG9b54 );
and \U$35412 ( \43612 , \10418 , \43179_nG9b51 );
or \U$35413 ( \43613 , \43611 , \43612 );
xor \U$35414 ( \43614 , \10417 , \43613 );
buf \U$35415 ( \43615 , \43614 );
buf \U$35417 ( \43616 , \43615 );
and \U$35418 ( \43617 , \18702 , \39591_nG9b78 );
and \U$35419 ( \43618 , \18699 , \39963_nG9b75 );
or \U$35420 ( \43619 , \43617 , \43618 );
xor \U$35421 ( \43620 , \18698 , \43619 );
buf \U$35422 ( \43621 , \43620 );
buf \U$35424 ( \43622 , \43621 );
xor \U$35425 ( \43623 , \43616 , \43622 );
and \U$35426 ( \43624 , \13370 , \41963_nG9b60 );
and \U$35427 ( \43625 , \13367 , \42201_nG9b5d );
or \U$35428 ( \43626 , \43624 , \43625 );
xor \U$35429 ( \43627 , \13366 , \43626 );
buf \U$35430 ( \43628 , \43627 );
buf \U$35432 ( \43629 , \43628 );
xor \U$35433 ( \43630 , \43623 , \43629 );
buf \U$35434 ( \43631 , \43630 );
xor \U$35435 ( \43632 , \43610 , \43631 );
and \U$35436 ( \43633 , \24792 , \36986_nG9b90 );
and \U$35437 ( \43634 , \24789 , \37250_nG9b8d );
or \U$35438 ( \43635 , \43633 , \43634 );
xor \U$35439 ( \43636 , \24788 , \43635 );
buf \U$35440 ( \43637 , \43636 );
buf \U$35442 ( \43638 , \43637 );
and \U$35443 ( \43639 , \23201 , \37607_nG9b8a );
and \U$35444 ( \43640 , \23198 , \37974_nG9b87 );
or \U$35445 ( \43641 , \43639 , \43640 );
xor \U$35446 ( \43642 , \23197 , \43641 );
buf \U$35447 ( \43643 , \43642 );
buf \U$35449 ( \43644 , \43643 );
xor \U$35450 ( \43645 , \43638 , \43644 );
and \U$35451 ( \43646 , \21658 , \38337_nG9b84 );
and \U$35452 ( \43647 , \21655 , \38663_nG9b81 );
or \U$35453 ( \43648 , \43646 , \43647 );
xor \U$35454 ( \43649 , \21654 , \43648 );
buf \U$35455 ( \43650 , \43649 );
buf \U$35457 ( \43651 , \43650 );
xor \U$35458 ( \43652 , \43645 , \43651 );
buf \U$35459 ( \43653 , \43652 );
xor \U$35460 ( \43654 , \43632 , \43653 );
buf \U$35461 ( \43655 , \43654 );
xor \U$35462 ( \43656 , \43593 , \43655 );
buf \U$35463 ( \43657 , \43656 );
xor \U$35464 ( \43658 , \43548 , \43657 );
and \U$35465 ( \43659 , \43391 , \43423 );
and \U$35466 ( \43660 , \43391 , \43429 );
and \U$35467 ( \43661 , \43423 , \43429 );
or \U$35468 ( \43662 , \43659 , \43660 , \43661 );
buf \U$35469 ( \43663 , \43662 );
xor \U$35470 ( \43664 , \43658 , \43663 );
buf \U$35471 ( \43665 , \43664 );
xor \U$35472 ( \43666 , \43543 , \43665 );
and \U$35473 ( \43667 , \43448 , \43482 );
and \U$35474 ( \43668 , \43448 , \43517 );
and \U$35475 ( \43669 , \43482 , \43517 );
or \U$35476 ( \43670 , \43667 , \43668 , \43669 );
buf \U$35477 ( \43671 , \43670 );
and \U$35478 ( \43672 , \43396 , \43415 );
and \U$35479 ( \43673 , \43396 , \43421 );
and \U$35480 ( \43674 , \43415 , \43421 );
or \U$35481 ( \43675 , \43672 , \43673 , \43674 );
buf \U$35482 ( \43676 , \43675 );
xor \U$35483 ( \43677 , \43671 , \43676 );
and \U$35484 ( \43678 , \43488 , \43509 );
and \U$35485 ( \43679 , \43488 , \43515 );
and \U$35486 ( \43680 , \43509 , \43515 );
or \U$35487 ( \43681 , \43678 , \43679 , \43680 );
buf \U$35488 ( \43682 , \43681 );
and \U$35489 ( \43683 , \26431 , \36172_nG9b96 );
and \U$35490 ( \43684 , \26428 , \36589_nG9b93 );
or \U$35491 ( \43685 , \43683 , \43684 );
xor \U$35492 ( \43686 , \26427 , \43685 );
buf \U$35493 ( \43687 , \43686 );
buf \U$35495 ( \43688 , \43687 );
and \U$35496 ( \43689 , \17297 , \40204_nG9b72 );
and \U$35497 ( \43690 , \17294 , \40452_nG9b6f );
or \U$35498 ( \43691 , \43689 , \43690 );
xor \U$35499 ( \43692 , \17293 , \43691 );
buf \U$35500 ( \43693 , \43692 );
buf \U$35502 ( \43694 , \43693 );
xor \U$35503 ( \43695 , \43688 , \43694 );
and \U$35504 ( \43696 , \15940 , \40843_nG9b6c );
and \U$35505 ( \43697 , \15937 , \41040_nG9b69 );
or \U$35506 ( \43698 , \43696 , \43697 );
xor \U$35507 ( \43699 , \15936 , \43698 );
buf \U$35508 ( \43700 , \43699 );
buf \U$35510 ( \43701 , \43700 );
xor \U$35511 ( \43702 , \43695 , \43701 );
buf \U$35512 ( \43703 , \43702 );
and \U$35513 ( \43704 , \43494 , \43500 );
and \U$35514 ( \43705 , \43494 , \43507 );
and \U$35515 ( \43706 , \43500 , \43507 );
or \U$35516 ( \43707 , \43704 , \43705 , \43706 );
buf \U$35517 ( \43708 , \43707 );
xor \U$35518 ( \43709 , \43703 , \43708 );
and \U$35519 ( \43710 , \43356 , \43362 );
and \U$35520 ( \43711 , \43356 , \43369 );
and \U$35521 ( \43712 , \43362 , \43369 );
or \U$35522 ( \43713 , \43710 , \43711 , \43712 );
buf \U$35523 ( \43714 , \43713 );
xor \U$35524 ( \43715 , \43709 , \43714 );
buf \U$35525 ( \43716 , \43715 );
xor \U$35526 ( \43717 , \43682 , \43716 );
and \U$35527 ( \43718 , \43335 , \43341 );
and \U$35528 ( \43719 , \43335 , \43348 );
and \U$35529 ( \43720 , \43341 , \43348 );
or \U$35530 ( \43721 , \43718 , \43719 , \43720 );
buf \U$35531 ( \43722 , \43721 );
and \U$35532 ( \43723 , \31636 , \34041_nG9ba8 );
and \U$35533 ( \43724 , \31633 , \34294_nG9ba5 );
or \U$35534 ( \43725 , \43723 , \43724 );
xor \U$35535 ( \43726 , \31632 , \43725 );
buf \U$35536 ( \43727 , \43726 );
buf \U$35538 ( \43728 , \43727 );
and \U$35539 ( \43729 , \29853 , \34643_nG9ba2 );
and \U$35540 ( \43730 , \29850 , \35094_nG9b9f );
or \U$35541 ( \43731 , \43729 , \43730 );
xor \U$35542 ( \43732 , \29849 , \43731 );
buf \U$35543 ( \43733 , \43732 );
buf \U$35545 ( \43734 , \43733 );
xor \U$35546 ( \43735 , \43728 , \43734 );
and \U$35547 ( \43736 , \28118 , \35570_nG9b9c );
and \U$35548 ( \43737 , \28115 , \35801_nG9b99 );
or \U$35549 ( \43738 , \43736 , \43737 );
xor \U$35550 ( \43739 , \28114 , \43738 );
buf \U$35551 ( \43740 , \43739 );
buf \U$35553 ( \43741 , \43740 );
xor \U$35554 ( \43742 , \43735 , \43741 );
buf \U$35555 ( \43743 , \43742 );
xor \U$35556 ( \43744 , \43722 , \43743 );
and \U$35557 ( \43745 , \43374 , \43380 );
and \U$35558 ( \43746 , \43374 , \43387 );
and \U$35559 ( \43747 , \43380 , \43387 );
or \U$35560 ( \43748 , \43745 , \43746 , \43747 );
buf \U$35561 ( \43749 , \43748 );
xor \U$35562 ( \43750 , \43744 , \43749 );
buf \U$35563 ( \43751 , \43750 );
xor \U$35564 ( \43752 , \43717 , \43751 );
buf \U$35565 ( \43753 , \43752 );
xor \U$35566 ( \43754 , \43677 , \43753 );
buf \U$35567 ( \43755 , \43754 );
xor \U$35568 ( \43756 , \43666 , \43755 );
and \U$35569 ( \43757 , \43538 , \43756 );
and \U$35571 ( \43758 , \43532 , \43537 );
or \U$35573 ( \43759 , 1'b0 , \43758 , 1'b0 );
xor \U$35574 ( \43760 , \43757 , \43759 );
and \U$35576 ( \43761 , \43525 , \43531 );
and \U$35577 ( \43762 , \43527 , \43531 );
or \U$35578 ( \43763 , 1'b0 , \43761 , \43762 );
xor \U$35579 ( \43764 , \43760 , \43763 );
xor \U$35586 ( \43765 , \43764 , 1'b0 );
and \U$35587 ( \43766 , \43543 , \43665 );
and \U$35588 ( \43767 , \43543 , \43755 );
and \U$35589 ( \43768 , \43665 , \43755 );
or \U$35590 ( \43769 , \43766 , \43767 , \43768 );
xor \U$35591 ( \43770 , \43765 , \43769 );
and \U$35592 ( \43771 , \43671 , \43676 );
and \U$35593 ( \43772 , \43671 , \43753 );
and \U$35594 ( \43773 , \43676 , \43753 );
or \U$35595 ( \43774 , \43771 , \43772 , \43773 );
buf \U$35596 ( \43775 , \43774 );
and \U$35597 ( \43776 , \43553 , \43592 );
and \U$35598 ( \43777 , \43553 , \43655 );
and \U$35599 ( \43778 , \43592 , \43655 );
or \U$35600 ( \43779 , \43776 , \43777 , \43778 );
buf \U$35601 ( \43780 , \43779 );
xor \U$35602 ( \43781 , \43775 , \43780 );
and \U$35603 ( \43782 , \43703 , \43708 );
and \U$35604 ( \43783 , \43703 , \43714 );
and \U$35605 ( \43784 , \43708 , \43714 );
or \U$35606 ( \43785 , \43782 , \43783 , \43784 );
buf \U$35607 ( \43786 , \43785 );
and \U$35608 ( \43787 , \43722 , \43743 );
and \U$35609 ( \43788 , \43722 , \43749 );
and \U$35610 ( \43789 , \43743 , \43749 );
or \U$35611 ( \43790 , \43787 , \43788 , \43789 );
buf \U$35612 ( \43791 , \43790 );
and \U$35613 ( \43792 , \43728 , \43734 );
and \U$35614 ( \43793 , \43728 , \43741 );
and \U$35615 ( \43794 , \43734 , \43741 );
or \U$35616 ( \43795 , \43792 , \43793 , \43794 );
buf \U$35617 ( \43796 , \43795 );
and \U$35618 ( \43797 , 1'b1 , \43567 );
and \U$35619 ( \43798 , 1'b1 , \43573 );
and \U$35620 ( \43799 , \43567 , \43573 );
or \U$35621 ( \43800 , \43797 , \43798 , \43799 );
buf \U$35622 ( \43801 , \43800 );
xor \U$35623 ( \43802 , \43796 , \43801 );
and \U$35624 ( \43803 , \12157 , \42766_nG9b57 );
and \U$35625 ( \43804 , \12154 , \42848_nG9b54 );
or \U$35626 ( \43805 , \43803 , \43804 );
xor \U$35627 ( \43806 , \12153 , \43805 );
buf \U$35628 ( \43807 , \43806 );
buf \U$35630 ( \43808 , \43807 );
xor \U$35631 ( \43809 , \43802 , \43808 );
buf \U$35632 ( \43810 , \43809 );
xor \U$35633 ( \43811 , \43791 , \43810 );
and \U$35634 ( \43812 , \43563 , \43575 );
and \U$35635 ( \43813 , \43563 , \43582 );
and \U$35636 ( \43814 , \43575 , \43582 );
or \U$35637 ( \43815 , \43812 , \43813 , \43814 );
buf \U$35638 ( \43816 , \43815 );
xor \U$35639 ( \43817 , \43811 , \43816 );
buf \U$35640 ( \43818 , \43817 );
xor \U$35641 ( \43819 , \43786 , \43818 );
and \U$35642 ( \43820 , \23201 , \37974_nG9b87 );
and \U$35643 ( \43821 , \23198 , \38337_nG9b84 );
or \U$35644 ( \43822 , \43820 , \43821 );
xor \U$35645 ( \43823 , \23197 , \43822 );
buf \U$35646 ( \43824 , \43823 );
buf \U$35648 ( \43825 , \43824 );
and \U$35649 ( \43826 , \21658 , \38663_nG9b81 );
and \U$35650 ( \43827 , \21655 , \38968_nG9b7e );
or \U$35651 ( \43828 , \43826 , \43827 );
xor \U$35652 ( \43829 , \21654 , \43828 );
buf \U$35653 ( \43830 , \43829 );
buf \U$35655 ( \43831 , \43830 );
xor \U$35656 ( \43832 , \43825 , \43831 );
and \U$35657 ( \43833 , \15940 , \41040_nG9b69 );
and \U$35658 ( \43834 , \15937 , \41381_nG9b66 );
or \U$35659 ( \43835 , \43833 , \43834 );
xor \U$35660 ( \43836 , \15936 , \43835 );
buf \U$35661 ( \43837 , \43836 );
buf \U$35663 ( \43838 , \43837 );
xor \U$35664 ( \43839 , \43832 , \43838 );
buf \U$35665 ( \43840 , \43839 );
and \U$35666 ( \43841 , \26431 , \36589_nG9b93 );
and \U$35667 ( \43842 , \26428 , \36986_nG9b90 );
or \U$35668 ( \43843 , \43841 , \43842 );
xor \U$35669 ( \43844 , \26427 , \43843 );
buf \U$35670 ( \43845 , \43844 );
buf \U$35672 ( \43846 , \43845 );
and \U$35673 ( \43847 , \24792 , \37250_nG9b8d );
and \U$35674 ( \43848 , \24789 , \37607_nG9b8a );
or \U$35675 ( \43849 , \43847 , \43848 );
xor \U$35676 ( \43850 , \24788 , \43849 );
buf \U$35677 ( \43851 , \43850 );
buf \U$35679 ( \43852 , \43851 );
xor \U$35680 ( \43853 , \43846 , \43852 );
and \U$35681 ( \43854 , \13370 , \42201_nG9b5d );
and \U$35682 ( \43855 , \13367 , \42433_nG9b5a );
or \U$35683 ( \43856 , \43854 , \43855 );
xor \U$35684 ( \43857 , \13366 , \43856 );
buf \U$35685 ( \43858 , \43857 );
buf \U$35687 ( \43859 , \43858 );
xor \U$35688 ( \43860 , \43853 , \43859 );
buf \U$35689 ( \43861 , \43860 );
xor \U$35690 ( \43862 , \43840 , \43861 );
and \U$35692 ( \43863 , \32916 , \34041_nG9ba8 );
or \U$35693 ( \43864 , 1'b0 , \43863 );
xor \U$35694 ( \43865 , 1'b0 , \43864 );
buf \U$35695 ( \43866 , \43865 );
buf \U$35696 ( \43867 , \43866 );
not \U$35697 ( \43868 , \43867 );
and \U$35698 ( \43869 , \20155 , \39334_nG9b7b );
and \U$35699 ( \43870 , \20152 , \39591_nG9b78 );
or \U$35700 ( \43871 , \43869 , \43870 );
xor \U$35701 ( \43872 , \20151 , \43871 );
buf \U$35702 ( \43873 , \43872 );
buf \U$35704 ( \43874 , \43873 );
xor \U$35705 ( \43875 , \43868 , \43874 );
and \U$35706 ( \43876 , \14631 , \41685_nG9b63 );
and \U$35707 ( \43877 , \14628 , \41963_nG9b60 );
or \U$35708 ( \43878 , \43876 , \43877 );
xor \U$35709 ( \43879 , \14627 , \43878 );
buf \U$35710 ( \43880 , \43879 );
buf \U$35712 ( \43881 , \43880 );
xor \U$35713 ( \43882 , \43875 , \43881 );
buf \U$35714 ( \43883 , \43882 );
xor \U$35715 ( \43884 , \43862 , \43883 );
buf \U$35716 ( \43885 , \43884 );
xor \U$35717 ( \43886 , \43819 , \43885 );
buf \U$35718 ( \43887 , \43886 );
xor \U$35719 ( \43888 , \43781 , \43887 );
buf \U$35720 ( \43889 , \43888 );
and \U$35721 ( \43890 , \43548 , \43657 );
and \U$35722 ( \43891 , \43548 , \43663 );
and \U$35723 ( \43892 , \43657 , \43663 );
or \U$35724 ( \43893 , \43890 , \43891 , \43892 );
buf \U$35725 ( \43894 , \43893 );
xor \U$35726 ( \43895 , \43889 , \43894 );
and \U$35727 ( \43896 , \43610 , \43631 );
and \U$35728 ( \43897 , \43610 , \43653 );
and \U$35729 ( \43898 , \43631 , \43653 );
or \U$35730 ( \43899 , \43896 , \43897 , \43898 );
buf \U$35731 ( \43900 , \43899 );
and \U$35732 ( \43901 , \10421 , \43179_nG9b51 );
or \U$35734 ( \43902 , \43901 , 1'b0 );
xor \U$35735 ( \43903 , \10417 , \43902 );
buf \U$35736 ( \43904 , \43903 );
buf \U$35738 ( \43905 , \43904 );
and \U$35739 ( \43906 , \18702 , \39963_nG9b75 );
and \U$35740 ( \43907 , \18699 , \40204_nG9b72 );
or \U$35741 ( \43908 , \43906 , \43907 );
xor \U$35742 ( \43909 , \18698 , \43908 );
buf \U$35743 ( \43910 , \43909 );
buf \U$35745 ( \43911 , \43910 );
xor \U$35746 ( \43912 , \43905 , \43911 );
and \U$35747 ( \43913 , \17297 , \40452_nG9b6f );
and \U$35748 ( \43914 , \17294 , \40843_nG9b6c );
or \U$35749 ( \43915 , \43913 , \43914 );
xor \U$35750 ( \43916 , \17293 , \43915 );
buf \U$35751 ( \43917 , \43916 );
buf \U$35753 ( \43918 , \43917 );
xor \U$35754 ( \43919 , \43912 , \43918 );
buf \U$35755 ( \43920 , \43919 );
and \U$35756 ( \43921 , \43688 , \43694 );
and \U$35757 ( \43922 , \43688 , \43701 );
and \U$35758 ( \43923 , \43694 , \43701 );
or \U$35759 ( \43924 , \43921 , \43922 , \43923 );
buf \U$35760 ( \43925 , \43924 );
xor \U$35761 ( \43926 , \43920 , \43925 );
and \U$35762 ( \43927 , \43638 , \43644 );
and \U$35763 ( \43928 , \43638 , \43651 );
and \U$35764 ( \43929 , \43644 , \43651 );
or \U$35765 ( \43930 , \43927 , \43928 , \43929 );
buf \U$35766 ( \43931 , \43930 );
xor \U$35767 ( \43932 , \43926 , \43931 );
buf \U$35768 ( \43933 , \43932 );
xor \U$35769 ( \43934 , \43900 , \43933 );
and \U$35770 ( \43935 , \43595 , \43601 );
and \U$35771 ( \43936 , \43595 , \43608 );
and \U$35772 ( \43937 , \43601 , \43608 );
or \U$35773 ( \43938 , \43935 , \43936 , \43937 );
buf \U$35774 ( \43939 , \43938 );
and \U$35775 ( \43940 , \31636 , \34294_nG9ba5 );
and \U$35776 ( \43941 , \31633 , \34643_nG9ba2 );
or \U$35777 ( \43942 , \43940 , \43941 );
xor \U$35778 ( \43943 , \31632 , \43942 );
buf \U$35779 ( \43944 , \43943 );
buf \U$35781 ( \43945 , \43944 );
and \U$35782 ( \43946 , \29853 , \35094_nG9b9f );
and \U$35783 ( \43947 , \29850 , \35570_nG9b9c );
or \U$35784 ( \43948 , \43946 , \43947 );
xor \U$35785 ( \43949 , \29849 , \43948 );
buf \U$35786 ( \43950 , \43949 );
buf \U$35788 ( \43951 , \43950 );
xor \U$35789 ( \43952 , \43945 , \43951 );
and \U$35790 ( \43953 , \28118 , \35801_nG9b99 );
and \U$35791 ( \43954 , \28115 , \36172_nG9b96 );
or \U$35792 ( \43955 , \43953 , \43954 );
xor \U$35793 ( \43956 , \28114 , \43955 );
buf \U$35794 ( \43957 , \43956 );
buf \U$35796 ( \43958 , \43957 );
xor \U$35797 ( \43959 , \43952 , \43958 );
buf \U$35798 ( \43960 , \43959 );
xor \U$35799 ( \43961 , \43939 , \43960 );
and \U$35800 ( \43962 , \43616 , \43622 );
and \U$35801 ( \43963 , \43616 , \43629 );
and \U$35802 ( \43964 , \43622 , \43629 );
or \U$35803 ( \43965 , \43962 , \43963 , \43964 );
buf \U$35804 ( \43966 , \43965 );
xor \U$35805 ( \43967 , \43961 , \43966 );
buf \U$35806 ( \43968 , \43967 );
xor \U$35807 ( \43969 , \43934 , \43968 );
buf \U$35808 ( \43970 , \43969 );
and \U$35809 ( \43971 , \43558 , \43584 );
and \U$35810 ( \43972 , \43558 , \43590 );
and \U$35811 ( \43973 , \43584 , \43590 );
or \U$35812 ( \43974 , \43971 , \43972 , \43973 );
buf \U$35813 ( \43975 , \43974 );
xor \U$35814 ( \43976 , \43970 , \43975 );
and \U$35815 ( \43977 , \43682 , \43716 );
and \U$35816 ( \43978 , \43682 , \43751 );
and \U$35817 ( \43979 , \43716 , \43751 );
or \U$35818 ( \43980 , \43977 , \43978 , \43979 );
buf \U$35819 ( \43981 , \43980 );
xor \U$35820 ( \43982 , \43976 , \43981 );
buf \U$35821 ( \43983 , \43982 );
xor \U$35822 ( \43984 , \43895 , \43983 );
and \U$35823 ( \43985 , \43770 , \43984 );
and \U$35825 ( \43986 , \43764 , \43769 );
or \U$35827 ( \43987 , 1'b0 , \43986 , 1'b0 );
xor \U$35828 ( \43988 , \43985 , \43987 );
and \U$35830 ( \43989 , \43757 , \43763 );
and \U$35831 ( \43990 , \43759 , \43763 );
or \U$35832 ( \43991 , 1'b0 , \43989 , \43990 );
xor \U$35833 ( \43992 , \43988 , \43991 );
xor \U$35840 ( \43993 , \43992 , 1'b0 );
and \U$35841 ( \43994 , \43889 , \43894 );
and \U$35842 ( \43995 , \43889 , \43983 );
and \U$35843 ( \43996 , \43894 , \43983 );
or \U$35844 ( \43997 , \43994 , \43995 , \43996 );
xor \U$35845 ( \43998 , \43993 , \43997 );
and \U$35846 ( \43999 , \43775 , \43780 );
and \U$35847 ( \44000 , \43775 , \43887 );
and \U$35848 ( \44001 , \43780 , \43887 );
or \U$35849 ( \44002 , \43999 , \44000 , \44001 );
buf \U$35850 ( \44003 , \44002 );
and \U$35851 ( \44004 , \43939 , \43960 );
and \U$35852 ( \44005 , \43939 , \43966 );
and \U$35853 ( \44006 , \43960 , \43966 );
or \U$35854 ( \44007 , \44004 , \44005 , \44006 );
buf \U$35855 ( \44008 , \44007 );
and \U$35856 ( \44009 , \43796 , \43801 );
and \U$35857 ( \44010 , \43796 , \43808 );
and \U$35858 ( \44011 , \43801 , \43808 );
or \U$35859 ( \44012 , \44009 , \44010 , \44011 );
buf \U$35860 ( \44013 , \44012 );
xor \U$35861 ( \44014 , \44008 , \44013 );
and \U$35862 ( \44015 , \43945 , \43951 );
and \U$35863 ( \44016 , \43945 , \43958 );
and \U$35864 ( \44017 , \43951 , \43958 );
or \U$35865 ( \44018 , \44015 , \44016 , \44017 );
buf \U$35866 ( \44019 , \44018 );
and \U$35867 ( \44020 , \17297 , \40843_nG9b6c );
and \U$35868 ( \44021 , \17294 , \41040_nG9b69 );
or \U$35869 ( \44022 , \44020 , \44021 );
xor \U$35870 ( \44023 , \17293 , \44022 );
buf \U$35871 ( \44024 , \44023 );
buf \U$35873 ( \44025 , \44024 );
xor \U$35874 ( \44026 , \44019 , \44025 );
and \U$35875 ( \44027 , \13370 , \42433_nG9b5a );
and \U$35876 ( \44028 , \13367 , \42766_nG9b57 );
or \U$35877 ( \44029 , \44027 , \44028 );
xor \U$35878 ( \44030 , \13366 , \44029 );
buf \U$35879 ( \44031 , \44030 );
buf \U$35881 ( \44032 , \44031 );
xor \U$35882 ( \44033 , \44026 , \44032 );
buf \U$35883 ( \44034 , \44033 );
xor \U$35884 ( \44035 , \44014 , \44034 );
buf \U$35885 ( \44036 , \44035 );
and \U$35886 ( \44037 , \43840 , \43861 );
and \U$35887 ( \44038 , \43840 , \43883 );
and \U$35888 ( \44039 , \43861 , \43883 );
or \U$35889 ( \44040 , \44037 , \44038 , \44039 );
buf \U$35890 ( \44041 , \44040 );
and \U$35891 ( \44042 , \28118 , \36172_nG9b96 );
and \U$35892 ( \44043 , \28115 , \36589_nG9b93 );
or \U$35893 ( \44044 , \44042 , \44043 );
xor \U$35894 ( \44045 , \28114 , \44044 );
buf \U$35895 ( \44046 , \44045 );
buf \U$35897 ( \44047 , \44046 );
and \U$35898 ( \44048 , \26431 , \36986_nG9b90 );
and \U$35899 ( \44049 , \26428 , \37250_nG9b8d );
or \U$35900 ( \44050 , \44048 , \44049 );
xor \U$35901 ( \44051 , \26427 , \44050 );
buf \U$35902 ( \44052 , \44051 );
buf \U$35904 ( \44053 , \44052 );
xor \U$35905 ( \44054 , \44047 , \44053 );
and \U$35906 ( \44055 , \18702 , \40204_nG9b72 );
and \U$35907 ( \44056 , \18699 , \40452_nG9b6f );
or \U$35908 ( \44057 , \44055 , \44056 );
xor \U$35909 ( \44058 , \18698 , \44057 );
buf \U$35910 ( \44059 , \44058 );
buf \U$35912 ( \44060 , \44059 );
xor \U$35913 ( \44061 , \44054 , \44060 );
buf \U$35914 ( \44062 , \44061 );
and \U$35915 ( \44063 , \43905 , \43911 );
and \U$35916 ( \44064 , \43905 , \43918 );
and \U$35917 ( \44065 , \43911 , \43918 );
or \U$35918 ( \44066 , \44063 , \44064 , \44065 );
buf \U$35919 ( \44067 , \44066 );
xor \U$35920 ( \44068 , \44062 , \44067 );
and \U$35921 ( \44069 , \43846 , \43852 );
and \U$35922 ( \44070 , \43846 , \43859 );
and \U$35923 ( \44071 , \43852 , \43859 );
or \U$35924 ( \44072 , \44069 , \44070 , \44071 );
buf \U$35925 ( \44073 , \44072 );
xor \U$35926 ( \44074 , \44068 , \44073 );
buf \U$35927 ( \44075 , \44074 );
xor \U$35928 ( \44076 , \44041 , \44075 );
and \U$35929 ( \44077 , \43920 , \43925 );
and \U$35930 ( \44078 , \43920 , \43931 );
and \U$35931 ( \44079 , \43925 , \43931 );
or \U$35932 ( \44080 , \44077 , \44078 , \44079 );
buf \U$35933 ( \44081 , \44080 );
xor \U$35934 ( \44082 , \44076 , \44081 );
buf \U$35935 ( \44083 , \44082 );
xor \U$35936 ( \44084 , \44036 , \44083 );
and \U$35937 ( \44085 , \43900 , \43933 );
and \U$35938 ( \44086 , \43900 , \43968 );
and \U$35939 ( \44087 , \43933 , \43968 );
or \U$35940 ( \44088 , \44085 , \44086 , \44087 );
buf \U$35941 ( \44089 , \44088 );
xor \U$35942 ( \44090 , \44084 , \44089 );
buf \U$35943 ( \44091 , \44090 );
xor \U$35944 ( \44092 , \44003 , \44091 );
and \U$35945 ( \44093 , \43970 , \43975 );
and \U$35946 ( \44094 , \43970 , \43981 );
and \U$35947 ( \44095 , \43975 , \43981 );
or \U$35948 ( \44096 , \44093 , \44094 , \44095 );
buf \U$35949 ( \44097 , \44096 );
and \U$35950 ( \44098 , \43791 , \43810 );
and \U$35951 ( \44099 , \43791 , \43816 );
and \U$35952 ( \44100 , \43810 , \43816 );
or \U$35953 ( \44101 , \44098 , \44099 , \44100 );
buf \U$35954 ( \44102 , \44101 );
buf \U$35955 ( \44103 , \43867 );
and \U$35956 ( \44104 , \21658 , \38968_nG9b7e );
and \U$35957 ( \44105 , \21655 , \39334_nG9b7b );
or \U$35958 ( \44106 , \44104 , \44105 );
xor \U$35959 ( \44107 , \21654 , \44106 );
buf \U$35960 ( \44108 , \44107 );
buf \U$35962 ( \44109 , \44108 );
xor \U$35963 ( \44110 , \44103 , \44109 );
and \U$35964 ( \44111 , \20155 , \39591_nG9b78 );
and \U$35965 ( \44112 , \20152 , \39963_nG9b75 );
or \U$35966 ( \44113 , \44111 , \44112 );
xor \U$35967 ( \44114 , \20151 , \44113 );
buf \U$35968 ( \44115 , \44114 );
buf \U$35970 ( \44116 , \44115 );
xor \U$35971 ( \44117 , \44110 , \44116 );
buf \U$35972 ( \44118 , \44117 );
and \U$35973 ( \44119 , \12157 , \42848_nG9b54 );
and \U$35974 ( \44120 , \12154 , \43179_nG9b51 );
or \U$35975 ( \44121 , \44119 , \44120 );
xor \U$35976 ( \44122 , \12153 , \44121 );
buf \U$35977 ( \44123 , \44122 );
buf \U$35979 ( \44124 , \44123 );
and \U$35980 ( \44125 , \31636 , \34643_nG9ba2 );
and \U$35981 ( \44126 , \31633 , \35094_nG9b9f );
or \U$35982 ( \44127 , \44125 , \44126 );
xor \U$35983 ( \44128 , \31632 , \44127 );
buf \U$35984 ( \44129 , \44128 );
buf \U$35986 ( \44130 , \44129 );
xor \U$35987 ( \44131 , \44124 , \44130 );
and \U$35988 ( \44132 , \14631 , \41963_nG9b60 );
and \U$35989 ( \44133 , \14628 , \42201_nG9b5d );
or \U$35990 ( \44134 , \44132 , \44133 );
xor \U$35991 ( \44135 , \14627 , \44134 );
buf \U$35992 ( \44136 , \44135 );
buf \U$35994 ( \44137 , \44136 );
xor \U$35995 ( \44138 , \44131 , \44137 );
buf \U$35996 ( \44139 , \44138 );
xor \U$35997 ( \44140 , \44118 , \44139 );
and \U$35998 ( \44141 , \24792 , \37607_nG9b8a );
and \U$35999 ( \44142 , \24789 , \37974_nG9b87 );
or \U$36000 ( \44143 , \44141 , \44142 );
xor \U$36001 ( \44144 , \24788 , \44143 );
buf \U$36002 ( \44145 , \44144 );
buf \U$36004 ( \44146 , \44145 );
and \U$36005 ( \44147 , \23201 , \38337_nG9b84 );
and \U$36006 ( \44148 , \23198 , \38663_nG9b81 );
or \U$36007 ( \44149 , \44147 , \44148 );
xor \U$36008 ( \44150 , \23197 , \44149 );
buf \U$36009 ( \44151 , \44150 );
buf \U$36011 ( \44152 , \44151 );
xor \U$36012 ( \44153 , \44146 , \44152 );
and \U$36013 ( \44154 , \15940 , \41381_nG9b66 );
and \U$36014 ( \44155 , \15937 , \41685_nG9b63 );
or \U$36015 ( \44156 , \44154 , \44155 );
xor \U$36016 ( \44157 , \15936 , \44156 );
buf \U$36017 ( \44158 , \44157 );
buf \U$36019 ( \44159 , \44158 );
xor \U$36020 ( \44160 , \44153 , \44159 );
buf \U$36021 ( \44161 , \44160 );
xor \U$36022 ( \44162 , \44140 , \44161 );
buf \U$36023 ( \44163 , \44162 );
xor \U$36024 ( \44164 , \44102 , \44163 );
and \U$36025 ( \44165 , \43825 , \43831 );
and \U$36026 ( \44166 , \43825 , \43838 );
and \U$36027 ( \44167 , \43831 , \43838 );
or \U$36028 ( \44168 , \44165 , \44166 , \44167 );
buf \U$36029 ( \44169 , \44168 );
and \U$36030 ( \44170 , \43868 , \43874 );
and \U$36031 ( \44171 , \43868 , \43881 );
and \U$36032 ( \44172 , \43874 , \43881 );
or \U$36033 ( \44173 , \44170 , \44171 , \44172 );
buf \U$36034 ( \44174 , \44173 );
xor \U$36035 ( \44175 , \44169 , \44174 );
xor \U$36039 ( \44176 , \10417 , 1'b0 );
not \U$36040 ( \44177 , \44176 );
buf \U$36041 ( \44178 , \44177 );
buf \U$36043 ( \44179 , \44178 );
and \U$36045 ( \44180 , \32916 , \34294_nG9ba5 );
or \U$36046 ( \44181 , 1'b0 , \44180 );
xor \U$36047 ( \44182 , 1'b0 , \44181 );
buf \U$36048 ( \44183 , \44182 );
buf \U$36050 ( \44184 , \44183 );
xor \U$36051 ( \44185 , \44179 , \44184 );
and \U$36052 ( \44186 , \29853 , \35570_nG9b9c );
and \U$36053 ( \44187 , \29850 , \35801_nG9b99 );
or \U$36054 ( \44188 , \44186 , \44187 );
xor \U$36055 ( \44189 , \29849 , \44188 );
buf \U$36056 ( \44190 , \44189 );
buf \U$36058 ( \44191 , \44190 );
xor \U$36059 ( \44192 , \44185 , \44191 );
buf \U$36060 ( \44193 , \44192 );
xor \U$36061 ( \44194 , \44175 , \44193 );
buf \U$36062 ( \44195 , \44194 );
xor \U$36063 ( \44196 , \44164 , \44195 );
buf \U$36064 ( \44197 , \44196 );
xor \U$36065 ( \44198 , \44097 , \44197 );
and \U$36066 ( \44199 , \43786 , \43818 );
and \U$36067 ( \44200 , \43786 , \43885 );
and \U$36068 ( \44201 , \43818 , \43885 );
or \U$36069 ( \44202 , \44199 , \44200 , \44201 );
buf \U$36070 ( \44203 , \44202 );
xor \U$36071 ( \44204 , \44198 , \44203 );
buf \U$36072 ( \44205 , \44204 );
xor \U$36073 ( \44206 , \44092 , \44205 );
and \U$36074 ( \44207 , \43998 , \44206 );
and \U$36076 ( \44208 , \43992 , \43997 );
or \U$36078 ( \44209 , 1'b0 , \44208 , 1'b0 );
xor \U$36079 ( \44210 , \44207 , \44209 );
and \U$36081 ( \44211 , \43985 , \43991 );
and \U$36082 ( \44212 , \43987 , \43991 );
or \U$36083 ( \44213 , 1'b0 , \44211 , \44212 );
xor \U$36084 ( \44214 , \44210 , \44213 );
xor \U$36091 ( \44215 , \44214 , 1'b0 );
and \U$36092 ( \44216 , \44003 , \44091 );
and \U$36093 ( \44217 , \44003 , \44205 );
and \U$36094 ( \44218 , \44091 , \44205 );
or \U$36095 ( \44219 , \44216 , \44217 , \44218 );
xor \U$36096 ( \44220 , \44215 , \44219 );
and \U$36097 ( \44221 , \44097 , \44197 );
and \U$36098 ( \44222 , \44097 , \44203 );
and \U$36099 ( \44223 , \44197 , \44203 );
or \U$36100 ( \44224 , \44221 , \44222 , \44223 );
buf \U$36101 ( \44225 , \44224 );
and \U$36102 ( \44226 , \44041 , \44075 );
and \U$36103 ( \44227 , \44041 , \44081 );
and \U$36104 ( \44228 , \44075 , \44081 );
or \U$36105 ( \44229 , \44226 , \44227 , \44228 );
buf \U$36106 ( \44230 , \44229 );
and \U$36107 ( \44231 , \44118 , \44139 );
and \U$36108 ( \44232 , \44118 , \44161 );
and \U$36109 ( \44233 , \44139 , \44161 );
or \U$36110 ( \44234 , \44231 , \44232 , \44233 );
buf \U$36111 ( \44235 , \44234 );
and \U$36113 ( \44236 , \32916 , \34643_nG9ba2 );
or \U$36114 ( \44237 , 1'b0 , \44236 );
xor \U$36115 ( \44238 , 1'b0 , \44237 );
buf \U$36116 ( \44239 , \44238 );
buf \U$36118 ( \44240 , \44239 );
and \U$36119 ( \44241 , \31636 , \35094_nG9b9f );
and \U$36120 ( \44242 , \31633 , \35570_nG9b9c );
or \U$36121 ( \44243 , \44241 , \44242 );
xor \U$36122 ( \44244 , \31632 , \44243 );
buf \U$36123 ( \44245 , \44244 );
buf \U$36125 ( \44246 , \44245 );
xor \U$36126 ( \44247 , \44240 , \44246 );
and \U$36127 ( \44248 , \15940 , \41685_nG9b63 );
and \U$36128 ( \44249 , \15937 , \41963_nG9b60 );
or \U$36129 ( \44250 , \44248 , \44249 );
xor \U$36130 ( \44251 , \15936 , \44250 );
buf \U$36131 ( \44252 , \44251 );
buf \U$36133 ( \44253 , \44252 );
xor \U$36134 ( \44254 , \44247 , \44253 );
buf \U$36135 ( \44255 , \44254 );
and \U$36136 ( \44256 , \44146 , \44152 );
and \U$36137 ( \44257 , \44146 , \44159 );
and \U$36138 ( \44258 , \44152 , \44159 );
or \U$36139 ( \44259 , \44256 , \44257 , \44258 );
buf \U$36140 ( \44260 , \44259 );
xor \U$36141 ( \44261 , \44255 , \44260 );
and \U$36142 ( \44262 , \44047 , \44053 );
and \U$36143 ( \44263 , \44047 , \44060 );
and \U$36144 ( \44264 , \44053 , \44060 );
or \U$36145 ( \44265 , \44262 , \44263 , \44264 );
buf \U$36146 ( \44266 , \44265 );
xor \U$36147 ( \44267 , \44261 , \44266 );
buf \U$36148 ( \44268 , \44267 );
xor \U$36149 ( \44269 , \44235 , \44268 );
and \U$36150 ( \44270 , \44124 , \44130 );
and \U$36151 ( \44271 , \44124 , \44137 );
and \U$36152 ( \44272 , \44130 , \44137 );
or \U$36153 ( \44273 , \44270 , \44271 , \44272 );
buf \U$36154 ( \44274 , \44273 );
and \U$36155 ( \44275 , \44179 , \44184 );
and \U$36156 ( \44276 , \44179 , \44191 );
and \U$36157 ( \44277 , \44184 , \44191 );
or \U$36158 ( \44278 , \44275 , \44276 , \44277 );
buf \U$36159 ( \44279 , \44278 );
xor \U$36160 ( \44280 , \44274 , \44279 );
and \U$36161 ( \44281 , \44103 , \44109 );
and \U$36162 ( \44282 , \44103 , \44116 );
and \U$36163 ( \44283 , \44109 , \44116 );
or \U$36164 ( \44284 , \44281 , \44282 , \44283 );
buf \U$36165 ( \44285 , \44284 );
xor \U$36166 ( \44286 , \44280 , \44285 );
buf \U$36167 ( \44287 , \44286 );
xor \U$36168 ( \44288 , \44269 , \44287 );
buf \U$36169 ( \44289 , \44288 );
xor \U$36170 ( \44290 , \44230 , \44289 );
and \U$36171 ( \44291 , \12157 , \43179_nG9b51 );
or \U$36173 ( \44292 , \44291 , 1'b0 );
xor \U$36174 ( \44293 , \12153 , \44292 );
buf \U$36175 ( \44294 , \44293 );
buf \U$36177 ( \44295 , \44294 );
and \U$36178 ( \44296 , \29853 , \35801_nG9b99 );
and \U$36179 ( \44297 , \29850 , \36172_nG9b96 );
or \U$36180 ( \44298 , \44296 , \44297 );
xor \U$36181 ( \44299 , \29849 , \44298 );
buf \U$36182 ( \44300 , \44299 );
buf \U$36183 ( \44301 , \44300 );
not \U$36184 ( \44302 , \44301 );
xor \U$36185 ( \44303 , \44295 , \44302 );
and \U$36186 ( \44304 , \13370 , \42766_nG9b57 );
and \U$36187 ( \44305 , \13367 , \42848_nG9b54 );
or \U$36188 ( \44306 , \44304 , \44305 );
xor \U$36189 ( \44307 , \13366 , \44306 );
buf \U$36190 ( \44308 , \44307 );
buf \U$36192 ( \44309 , \44308 );
xor \U$36193 ( \44310 , \44303 , \44309 );
buf \U$36194 ( \44311 , \44310 );
and \U$36195 ( \44312 , \44019 , \44025 );
and \U$36196 ( \44313 , \44019 , \44032 );
and \U$36197 ( \44314 , \44025 , \44032 );
or \U$36198 ( \44315 , \44312 , \44313 , \44314 );
buf \U$36199 ( \44316 , \44315 );
xor \U$36200 ( \44317 , \44311 , \44316 );
and \U$36201 ( \44318 , \44169 , \44174 );
and \U$36202 ( \44319 , \44169 , \44193 );
and \U$36203 ( \44320 , \44174 , \44193 );
or \U$36204 ( \44321 , \44318 , \44319 , \44320 );
buf \U$36205 ( \44322 , \44321 );
xor \U$36206 ( \44323 , \44317 , \44322 );
buf \U$36207 ( \44324 , \44323 );
xor \U$36208 ( \44325 , \44290 , \44324 );
buf \U$36209 ( \44326 , \44325 );
and \U$36210 ( \44327 , \44102 , \44163 );
and \U$36211 ( \44328 , \44102 , \44195 );
and \U$36212 ( \44329 , \44163 , \44195 );
or \U$36213 ( \44330 , \44327 , \44328 , \44329 );
buf \U$36214 ( \44331 , \44330 );
xor \U$36215 ( \44332 , \44326 , \44331 );
and \U$36216 ( \44333 , \44008 , \44013 );
and \U$36217 ( \44334 , \44008 , \44034 );
and \U$36218 ( \44335 , \44013 , \44034 );
or \U$36219 ( \44336 , \44333 , \44334 , \44335 );
buf \U$36220 ( \44337 , \44336 );
and \U$36221 ( \44338 , \28118 , \36589_nG9b93 );
and \U$36222 ( \44339 , \28115 , \36986_nG9b90 );
or \U$36223 ( \44340 , \44338 , \44339 );
xor \U$36224 ( \44341 , \28114 , \44340 );
buf \U$36225 ( \44342 , \44341 );
buf \U$36227 ( \44343 , \44342 );
and \U$36228 ( \44344 , \20155 , \39963_nG9b75 );
and \U$36229 ( \44345 , \20152 , \40204_nG9b72 );
or \U$36230 ( \44346 , \44344 , \44345 );
xor \U$36231 ( \44347 , \20151 , \44346 );
buf \U$36232 ( \44348 , \44347 );
buf \U$36234 ( \44349 , \44348 );
xor \U$36235 ( \44350 , \44343 , \44349 );
and \U$36236 ( \44351 , \18702 , \40452_nG9b6f );
and \U$36237 ( \44352 , \18699 , \40843_nG9b6c );
or \U$36238 ( \44353 , \44351 , \44352 );
xor \U$36239 ( \44354 , \18698 , \44353 );
buf \U$36240 ( \44355 , \44354 );
buf \U$36242 ( \44356 , \44355 );
xor \U$36243 ( \44357 , \44350 , \44356 );
buf \U$36244 ( \44358 , \44357 );
and \U$36245 ( \44359 , \23201 , \38663_nG9b81 );
and \U$36246 ( \44360 , \23198 , \38968_nG9b7e );
or \U$36247 ( \44361 , \44359 , \44360 );
xor \U$36248 ( \44362 , \23197 , \44361 );
buf \U$36249 ( \44363 , \44362 );
buf \U$36251 ( \44364 , \44363 );
and \U$36252 ( \44365 , \21658 , \39334_nG9b7b );
and \U$36253 ( \44366 , \21655 , \39591_nG9b78 );
or \U$36254 ( \44367 , \44365 , \44366 );
xor \U$36255 ( \44368 , \21654 , \44367 );
buf \U$36256 ( \44369 , \44368 );
buf \U$36258 ( \44370 , \44369 );
xor \U$36259 ( \44371 , \44364 , \44370 );
and \U$36260 ( \44372 , \17297 , \41040_nG9b69 );
and \U$36261 ( \44373 , \17294 , \41381_nG9b66 );
or \U$36262 ( \44374 , \44372 , \44373 );
xor \U$36263 ( \44375 , \17293 , \44374 );
buf \U$36264 ( \44376 , \44375 );
buf \U$36266 ( \44377 , \44376 );
xor \U$36267 ( \44378 , \44371 , \44377 );
buf \U$36268 ( \44379 , \44378 );
xor \U$36269 ( \44380 , \44358 , \44379 );
and \U$36270 ( \44381 , \26431 , \37250_nG9b8d );
and \U$36271 ( \44382 , \26428 , \37607_nG9b8a );
or \U$36272 ( \44383 , \44381 , \44382 );
xor \U$36273 ( \44384 , \26427 , \44383 );
buf \U$36274 ( \44385 , \44384 );
buf \U$36276 ( \44386 , \44385 );
and \U$36277 ( \44387 , \24792 , \37974_nG9b87 );
and \U$36278 ( \44388 , \24789 , \38337_nG9b84 );
or \U$36279 ( \44389 , \44387 , \44388 );
xor \U$36280 ( \44390 , \24788 , \44389 );
buf \U$36281 ( \44391 , \44390 );
buf \U$36283 ( \44392 , \44391 );
xor \U$36284 ( \44393 , \44386 , \44392 );
and \U$36285 ( \44394 , \14631 , \42201_nG9b5d );
and \U$36286 ( \44395 , \14628 , \42433_nG9b5a );
or \U$36287 ( \44396 , \44394 , \44395 );
xor \U$36288 ( \44397 , \14627 , \44396 );
buf \U$36289 ( \44398 , \44397 );
buf \U$36291 ( \44399 , \44398 );
xor \U$36292 ( \44400 , \44393 , \44399 );
buf \U$36293 ( \44401 , \44400 );
xor \U$36294 ( \44402 , \44380 , \44401 );
buf \U$36295 ( \44403 , \44402 );
xor \U$36296 ( \44404 , \44337 , \44403 );
and \U$36297 ( \44405 , \44062 , \44067 );
and \U$36298 ( \44406 , \44062 , \44073 );
and \U$36299 ( \44407 , \44067 , \44073 );
or \U$36300 ( \44408 , \44405 , \44406 , \44407 );
buf \U$36301 ( \44409 , \44408 );
xor \U$36302 ( \44410 , \44404 , \44409 );
buf \U$36303 ( \44411 , \44410 );
xor \U$36304 ( \44412 , \44332 , \44411 );
buf \U$36305 ( \44413 , \44412 );
xor \U$36306 ( \44414 , \44225 , \44413 );
and \U$36307 ( \44415 , \44036 , \44083 );
and \U$36308 ( \44416 , \44036 , \44089 );
and \U$36309 ( \44417 , \44083 , \44089 );
or \U$36310 ( \44418 , \44415 , \44416 , \44417 );
buf \U$36311 ( \44419 , \44418 );
xor \U$36312 ( \44420 , \44414 , \44419 );
and \U$36313 ( \44421 , \44220 , \44420 );
and \U$36315 ( \44422 , \44214 , \44219 );
or \U$36317 ( \44423 , 1'b0 , \44422 , 1'b0 );
xor \U$36318 ( \44424 , \44421 , \44423 );
and \U$36320 ( \44425 , \44207 , \44213 );
and \U$36321 ( \44426 , \44209 , \44213 );
or \U$36322 ( \44427 , 1'b0 , \44425 , \44426 );
xor \U$36323 ( \44428 , \44424 , \44427 );
xor \U$36330 ( \44429 , \44428 , 1'b0 );
and \U$36331 ( \44430 , \44225 , \44413 );
and \U$36332 ( \44431 , \44225 , \44419 );
and \U$36333 ( \44432 , \44413 , \44419 );
or \U$36334 ( \44433 , \44430 , \44431 , \44432 );
xor \U$36335 ( \44434 , \44429 , \44433 );
and \U$36336 ( \44435 , \44326 , \44331 );
and \U$36337 ( \44436 , \44326 , \44411 );
and \U$36338 ( \44437 , \44331 , \44411 );
or \U$36339 ( \44438 , \44435 , \44436 , \44437 );
buf \U$36340 ( \44439 , \44438 );
and \U$36341 ( \44440 , \44311 , \44316 );
and \U$36342 ( \44441 , \44311 , \44322 );
and \U$36343 ( \44442 , \44316 , \44322 );
or \U$36344 ( \44443 , \44440 , \44441 , \44442 );
buf \U$36345 ( \44444 , \44443 );
and \U$36346 ( \44445 , \44240 , \44246 );
and \U$36347 ( \44446 , \44240 , \44253 );
and \U$36348 ( \44447 , \44246 , \44253 );
or \U$36349 ( \44448 , \44445 , \44446 , \44447 );
buf \U$36350 ( \44449 , \44448 );
and \U$36351 ( \44450 , \44364 , \44370 );
and \U$36352 ( \44451 , \44364 , \44377 );
and \U$36353 ( \44452 , \44370 , \44377 );
or \U$36354 ( \44453 , \44450 , \44451 , \44452 );
buf \U$36355 ( \44454 , \44453 );
xor \U$36356 ( \44455 , \44449 , \44454 );
and \U$36357 ( \44456 , \14631 , \42433_nG9b5a );
and \U$36358 ( \44457 , \14628 , \42766_nG9b57 );
or \U$36359 ( \44458 , \44456 , \44457 );
xor \U$36360 ( \44459 , \14627 , \44458 );
buf \U$36361 ( \44460 , \44459 );
buf \U$36363 ( \44461 , \44460 );
xor \U$36364 ( \44462 , \44455 , \44461 );
buf \U$36365 ( \44463 , \44462 );
xor \U$36366 ( \44464 , \44444 , \44463 );
and \U$36367 ( \44465 , \29853 , \36172_nG9b96 );
and \U$36368 ( \44466 , \29850 , \36589_nG9b93 );
or \U$36369 ( \44467 , \44465 , \44466 );
xor \U$36370 ( \44468 , \29849 , \44467 );
buf \U$36371 ( \44469 , \44468 );
buf \U$36373 ( \44470 , \44469 );
and \U$36374 ( \44471 , \28118 , \36986_nG9b90 );
and \U$36375 ( \44472 , \28115 , \37250_nG9b8d );
or \U$36376 ( \44473 , \44471 , \44472 );
xor \U$36377 ( \44474 , \28114 , \44473 );
buf \U$36378 ( \44475 , \44474 );
buf \U$36380 ( \44476 , \44475 );
xor \U$36381 ( \44477 , \44470 , \44476 );
and \U$36382 ( \44478 , \26431 , \37607_nG9b8a );
and \U$36383 ( \44479 , \26428 , \37974_nG9b87 );
or \U$36384 ( \44480 , \44478 , \44479 );
xor \U$36385 ( \44481 , \26427 , \44480 );
buf \U$36386 ( \44482 , \44481 );
buf \U$36388 ( \44483 , \44482 );
xor \U$36389 ( \44484 , \44477 , \44483 );
buf \U$36390 ( \44485 , \44484 );
buf \U$36391 ( \44486 , \44301 );
and \U$36392 ( \44487 , \20155 , \40204_nG9b72 );
and \U$36393 ( \44488 , \20152 , \40452_nG9b6f );
or \U$36394 ( \44489 , \44487 , \44488 );
xor \U$36395 ( \44490 , \20151 , \44489 );
buf \U$36396 ( \44491 , \44490 );
buf \U$36398 ( \44492 , \44491 );
xor \U$36399 ( \44493 , \44486 , \44492 );
and \U$36400 ( \44494 , \18702 , \40843_nG9b6c );
and \U$36401 ( \44495 , \18699 , \41040_nG9b69 );
or \U$36402 ( \44496 , \44494 , \44495 );
xor \U$36403 ( \44497 , \18698 , \44496 );
buf \U$36404 ( \44498 , \44497 );
buf \U$36406 ( \44499 , \44498 );
xor \U$36407 ( \44500 , \44493 , \44499 );
buf \U$36408 ( \44501 , \44500 );
xor \U$36409 ( \44502 , \44485 , \44501 );
and \U$36410 ( \44503 , \44295 , \44302 );
and \U$36411 ( \44504 , \44295 , \44309 );
and \U$36412 ( \44505 , \44302 , \44309 );
or \U$36413 ( \44506 , \44503 , \44504 , \44505 );
buf \U$36414 ( \44507 , \44506 );
xor \U$36415 ( \44508 , \44502 , \44507 );
buf \U$36416 ( \44509 , \44508 );
xor \U$36417 ( \44510 , \44464 , \44509 );
buf \U$36418 ( \44511 , \44510 );
and \U$36419 ( \44512 , \44337 , \44403 );
and \U$36420 ( \44513 , \44337 , \44409 );
and \U$36421 ( \44514 , \44403 , \44409 );
or \U$36422 ( \44515 , \44512 , \44513 , \44514 );
buf \U$36423 ( \44516 , \44515 );
xor \U$36424 ( \44517 , \44511 , \44516 );
and \U$36425 ( \44518 , \44230 , \44289 );
and \U$36426 ( \44519 , \44230 , \44324 );
and \U$36427 ( \44520 , \44289 , \44324 );
or \U$36428 ( \44521 , \44518 , \44519 , \44520 );
buf \U$36429 ( \44522 , \44521 );
xor \U$36430 ( \44523 , \44517 , \44522 );
buf \U$36431 ( \44524 , \44523 );
xor \U$36432 ( \44525 , \44439 , \44524 );
and \U$36433 ( \44526 , \44235 , \44268 );
and \U$36434 ( \44527 , \44235 , \44287 );
and \U$36435 ( \44528 , \44268 , \44287 );
or \U$36436 ( \44529 , \44526 , \44527 , \44528 );
buf \U$36437 ( \44530 , \44529 );
and \U$36438 ( \44531 , \44358 , \44379 );
and \U$36439 ( \44532 , \44358 , \44401 );
and \U$36440 ( \44533 , \44379 , \44401 );
or \U$36441 ( \44534 , \44531 , \44532 , \44533 );
buf \U$36442 ( \44535 , \44534 );
and \U$36443 ( \44536 , \44343 , \44349 );
and \U$36444 ( \44537 , \44343 , \44356 );
and \U$36445 ( \44538 , \44349 , \44356 );
or \U$36446 ( \44539 , \44536 , \44537 , \44538 );
buf \U$36447 ( \44540 , \44539 );
and \U$36448 ( \44541 , \44386 , \44392 );
and \U$36449 ( \44542 , \44386 , \44399 );
and \U$36450 ( \44543 , \44392 , \44399 );
or \U$36451 ( \44544 , \44541 , \44542 , \44543 );
buf \U$36452 ( \44545 , \44544 );
xor \U$36453 ( \44546 , \44540 , \44545 );
xor \U$36457 ( \44547 , \12153 , 1'b0 );
not \U$36458 ( \44548 , \44547 );
buf \U$36459 ( \44549 , \44548 );
buf \U$36461 ( \44550 , \44549 );
and \U$36463 ( \44551 , \32916 , \35094_nG9b9f );
or \U$36464 ( \44552 , 1'b0 , \44551 );
xor \U$36465 ( \44553 , 1'b0 , \44552 );
buf \U$36466 ( \44554 , \44553 );
buf \U$36468 ( \44555 , \44554 );
xor \U$36469 ( \44556 , \44550 , \44555 );
and \U$36470 ( \44557 , \31636 , \35570_nG9b9c );
and \U$36471 ( \44558 , \31633 , \35801_nG9b99 );
or \U$36472 ( \44559 , \44557 , \44558 );
xor \U$36473 ( \44560 , \31632 , \44559 );
buf \U$36474 ( \44561 , \44560 );
buf \U$36476 ( \44562 , \44561 );
xor \U$36477 ( \44563 , \44556 , \44562 );
buf \U$36478 ( \44564 , \44563 );
xor \U$36479 ( \44565 , \44546 , \44564 );
buf \U$36480 ( \44566 , \44565 );
xor \U$36481 ( \44567 , \44535 , \44566 );
and \U$36482 ( \44568 , \44255 , \44260 );
and \U$36483 ( \44569 , \44255 , \44266 );
and \U$36484 ( \44570 , \44260 , \44266 );
or \U$36485 ( \44571 , \44568 , \44569 , \44570 );
buf \U$36486 ( \44572 , \44571 );
xor \U$36487 ( \44573 , \44567 , \44572 );
buf \U$36488 ( \44574 , \44573 );
xor \U$36489 ( \44575 , \44530 , \44574 );
and \U$36490 ( \44576 , \44274 , \44279 );
and \U$36491 ( \44577 , \44274 , \44285 );
and \U$36492 ( \44578 , \44279 , \44285 );
or \U$36493 ( \44579 , \44576 , \44577 , \44578 );
buf \U$36494 ( \44580 , \44579 );
and \U$36495 ( \44581 , \24792 , \38337_nG9b84 );
and \U$36496 ( \44582 , \24789 , \38663_nG9b81 );
or \U$36497 ( \44583 , \44581 , \44582 );
xor \U$36498 ( \44584 , \24788 , \44583 );
buf \U$36499 ( \44585 , \44584 );
buf \U$36501 ( \44586 , \44585 );
and \U$36502 ( \44587 , \23201 , \38968_nG9b7e );
and \U$36503 ( \44588 , \23198 , \39334_nG9b7b );
or \U$36504 ( \44589 , \44587 , \44588 );
xor \U$36505 ( \44590 , \23197 , \44589 );
buf \U$36506 ( \44591 , \44590 );
buf \U$36508 ( \44592 , \44591 );
xor \U$36509 ( \44593 , \44586 , \44592 );
and \U$36510 ( \44594 , \17297 , \41381_nG9b66 );
and \U$36511 ( \44595 , \17294 , \41685_nG9b63 );
or \U$36512 ( \44596 , \44594 , \44595 );
xor \U$36513 ( \44597 , \17293 , \44596 );
buf \U$36514 ( \44598 , \44597 );
buf \U$36516 ( \44599 , \44598 );
xor \U$36517 ( \44600 , \44593 , \44599 );
buf \U$36518 ( \44601 , \44600 );
xor \U$36519 ( \44602 , \44580 , \44601 );
and \U$36520 ( \44603 , \13370 , \42848_nG9b54 );
and \U$36521 ( \44604 , \13367 , \43179_nG9b51 );
or \U$36522 ( \44605 , \44603 , \44604 );
xor \U$36523 ( \44606 , \13366 , \44605 );
buf \U$36524 ( \44607 , \44606 );
buf \U$36526 ( \44608 , \44607 );
and \U$36527 ( \44609 , \21658 , \39591_nG9b78 );
and \U$36528 ( \44610 , \21655 , \39963_nG9b75 );
or \U$36529 ( \44611 , \44609 , \44610 );
xor \U$36530 ( \44612 , \21654 , \44611 );
buf \U$36531 ( \44613 , \44612 );
buf \U$36533 ( \44614 , \44613 );
xor \U$36534 ( \44615 , \44608 , \44614 );
and \U$36535 ( \44616 , \15940 , \41963_nG9b60 );
and \U$36536 ( \44617 , \15937 , \42201_nG9b5d );
or \U$36537 ( \44618 , \44616 , \44617 );
xor \U$36538 ( \44619 , \15936 , \44618 );
buf \U$36539 ( \44620 , \44619 );
buf \U$36541 ( \44621 , \44620 );
xor \U$36542 ( \44622 , \44615 , \44621 );
buf \U$36543 ( \44623 , \44622 );
xor \U$36544 ( \44624 , \44602 , \44623 );
buf \U$36545 ( \44625 , \44624 );
xor \U$36546 ( \44626 , \44575 , \44625 );
buf \U$36547 ( \44627 , \44626 );
xor \U$36548 ( \44628 , \44525 , \44627 );
and \U$36549 ( \44629 , \44434 , \44628 );
and \U$36551 ( \44630 , \44428 , \44433 );
or \U$36553 ( \44631 , 1'b0 , \44630 , 1'b0 );
xor \U$36554 ( \44632 , \44629 , \44631 );
and \U$36556 ( \44633 , \44421 , \44427 );
and \U$36557 ( \44634 , \44423 , \44427 );
or \U$36558 ( \44635 , 1'b0 , \44633 , \44634 );
xor \U$36559 ( \44636 , \44632 , \44635 );
xor \U$36566 ( \44637 , \44636 , 1'b0 );
and \U$36567 ( \44638 , \44439 , \44524 );
and \U$36568 ( \44639 , \44439 , \44627 );
and \U$36569 ( \44640 , \44524 , \44627 );
or \U$36570 ( \44641 , \44638 , \44639 , \44640 );
xor \U$36571 ( \44642 , \44637 , \44641 );
and \U$36572 ( \44643 , \44511 , \44516 );
and \U$36573 ( \44644 , \44511 , \44522 );
and \U$36574 ( \44645 , \44516 , \44522 );
or \U$36575 ( \44646 , \44643 , \44644 , \44645 );
buf \U$36576 ( \44647 , \44646 );
and \U$36577 ( \44648 , \44530 , \44574 );
and \U$36578 ( \44649 , \44530 , \44625 );
and \U$36579 ( \44650 , \44574 , \44625 );
or \U$36580 ( \44651 , \44648 , \44649 , \44650 );
buf \U$36581 ( \44652 , \44651 );
and \U$36582 ( \44653 , \44444 , \44463 );
and \U$36583 ( \44654 , \44444 , \44509 );
and \U$36584 ( \44655 , \44463 , \44509 );
or \U$36585 ( \44656 , \44653 , \44654 , \44655 );
buf \U$36586 ( \44657 , \44656 );
xor \U$36587 ( \44658 , \44652 , \44657 );
and \U$36588 ( \44659 , \44550 , \44555 );
and \U$36589 ( \44660 , \44550 , \44562 );
and \U$36590 ( \44661 , \44555 , \44562 );
or \U$36591 ( \44662 , \44659 , \44660 , \44661 );
buf \U$36592 ( \44663 , \44662 );
and \U$36593 ( \44664 , \31636 , \35801_nG9b99 );
and \U$36594 ( \44665 , \31633 , \36172_nG9b96 );
or \U$36595 ( \44666 , \44664 , \44665 );
xor \U$36596 ( \44667 , \31632 , \44666 );
buf \U$36597 ( \44668 , \44667 );
buf \U$36598 ( \44669 , \44668 );
not \U$36599 ( \44670 , \44669 );
xor \U$36600 ( \44671 , \44663 , \44670 );
and \U$36601 ( \44672 , \14631 , \42766_nG9b57 );
and \U$36602 ( \44673 , \14628 , \42848_nG9b54 );
or \U$36603 ( \44674 , \44672 , \44673 );
xor \U$36604 ( \44675 , \14627 , \44674 );
buf \U$36605 ( \44676 , \44675 );
buf \U$36607 ( \44677 , \44676 );
xor \U$36608 ( \44678 , \44671 , \44677 );
buf \U$36609 ( \44679 , \44678 );
and \U$36610 ( \44680 , \26431 , \37974_nG9b87 );
and \U$36611 ( \44681 , \26428 , \38337_nG9b84 );
or \U$36612 ( \44682 , \44680 , \44681 );
xor \U$36613 ( \44683 , \26427 , \44682 );
buf \U$36614 ( \44684 , \44683 );
buf \U$36616 ( \44685 , \44684 );
and \U$36617 ( \44686 , \24792 , \38663_nG9b81 );
and \U$36618 ( \44687 , \24789 , \38968_nG9b7e );
or \U$36619 ( \44688 , \44686 , \44687 );
xor \U$36620 ( \44689 , \24788 , \44688 );
buf \U$36621 ( \44690 , \44689 );
buf \U$36623 ( \44691 , \44690 );
xor \U$36624 ( \44692 , \44685 , \44691 );
and \U$36625 ( \44693 , \18702 , \41040_nG9b69 );
and \U$36626 ( \44694 , \18699 , \41381_nG9b66 );
or \U$36627 ( \44695 , \44693 , \44694 );
xor \U$36628 ( \44696 , \18698 , \44695 );
buf \U$36629 ( \44697 , \44696 );
buf \U$36631 ( \44698 , \44697 );
xor \U$36632 ( \44699 , \44692 , \44698 );
buf \U$36633 ( \44700 , \44699 );
xor \U$36634 ( \44701 , \44679 , \44700 );
and \U$36635 ( \44702 , \29853 , \36589_nG9b93 );
and \U$36636 ( \44703 , \29850 , \36986_nG9b90 );
or \U$36637 ( \44704 , \44702 , \44703 );
xor \U$36638 ( \44705 , \29849 , \44704 );
buf \U$36639 ( \44706 , \44705 );
buf \U$36641 ( \44707 , \44706 );
and \U$36642 ( \44708 , \28118 , \37250_nG9b8d );
and \U$36643 ( \44709 , \28115 , \37607_nG9b8a );
or \U$36644 ( \44710 , \44708 , \44709 );
xor \U$36645 ( \44711 , \28114 , \44710 );
buf \U$36646 ( \44712 , \44711 );
buf \U$36648 ( \44713 , \44712 );
xor \U$36649 ( \44714 , \44707 , \44713 );
and \U$36650 ( \44715 , \15940 , \42201_nG9b5d );
and \U$36651 ( \44716 , \15937 , \42433_nG9b5a );
or \U$36652 ( \44717 , \44715 , \44716 );
xor \U$36653 ( \44718 , \15936 , \44717 );
buf \U$36654 ( \44719 , \44718 );
buf \U$36656 ( \44720 , \44719 );
xor \U$36657 ( \44721 , \44714 , \44720 );
buf \U$36658 ( \44722 , \44721 );
xor \U$36659 ( \44723 , \44701 , \44722 );
buf \U$36660 ( \44724 , \44723 );
and \U$36661 ( \44725 , \13370 , \43179_nG9b51 );
or \U$36663 ( \44726 , \44725 , 1'b0 );
xor \U$36664 ( \44727 , \13366 , \44726 );
buf \U$36665 ( \44728 , \44727 );
buf \U$36667 ( \44729 , \44728 );
and \U$36668 ( \44730 , \21658 , \39963_nG9b75 );
and \U$36669 ( \44731 , \21655 , \40204_nG9b72 );
or \U$36670 ( \44732 , \44730 , \44731 );
xor \U$36671 ( \44733 , \21654 , \44732 );
buf \U$36672 ( \44734 , \44733 );
buf \U$36674 ( \44735 , \44734 );
xor \U$36675 ( \44736 , \44729 , \44735 );
and \U$36676 ( \44737 , \20155 , \40452_nG9b6f );
and \U$36677 ( \44738 , \20152 , \40843_nG9b6c );
or \U$36678 ( \44739 , \44737 , \44738 );
xor \U$36679 ( \44740 , \20151 , \44739 );
buf \U$36680 ( \44741 , \44740 );
buf \U$36682 ( \44742 , \44741 );
xor \U$36683 ( \44743 , \44736 , \44742 );
buf \U$36684 ( \44744 , \44743 );
and \U$36685 ( \44745 , \44486 , \44492 );
and \U$36686 ( \44746 , \44486 , \44499 );
and \U$36687 ( \44747 , \44492 , \44499 );
or \U$36688 ( \44748 , \44745 , \44746 , \44747 );
buf \U$36689 ( \44749 , \44748 );
xor \U$36690 ( \44750 , \44744 , \44749 );
and \U$36692 ( \44751 , \32916 , \35570_nG9b9c );
or \U$36693 ( \44752 , 1'b0 , \44751 );
xor \U$36694 ( \44753 , 1'b0 , \44752 );
buf \U$36695 ( \44754 , \44753 );
buf \U$36697 ( \44755 , \44754 );
and \U$36698 ( \44756 , \23201 , \39334_nG9b7b );
and \U$36699 ( \44757 , \23198 , \39591_nG9b78 );
or \U$36700 ( \44758 , \44756 , \44757 );
xor \U$36701 ( \44759 , \23197 , \44758 );
buf \U$36702 ( \44760 , \44759 );
buf \U$36704 ( \44761 , \44760 );
xor \U$36705 ( \44762 , \44755 , \44761 );
and \U$36706 ( \44763 , \17297 , \41685_nG9b63 );
and \U$36707 ( \44764 , \17294 , \41963_nG9b60 );
or \U$36708 ( \44765 , \44763 , \44764 );
xor \U$36709 ( \44766 , \17293 , \44765 );
buf \U$36710 ( \44767 , \44766 );
buf \U$36712 ( \44768 , \44767 );
xor \U$36713 ( \44769 , \44762 , \44768 );
buf \U$36714 ( \44770 , \44769 );
xor \U$36715 ( \44771 , \44750 , \44770 );
buf \U$36716 ( \44772 , \44771 );
xor \U$36717 ( \44773 , \44724 , \44772 );
and \U$36718 ( \44774 , \44485 , \44501 );
and \U$36719 ( \44775 , \44485 , \44507 );
and \U$36720 ( \44776 , \44501 , \44507 );
or \U$36721 ( \44777 , \44774 , \44775 , \44776 );
buf \U$36722 ( \44778 , \44777 );
xor \U$36723 ( \44779 , \44773 , \44778 );
buf \U$36724 ( \44780 , \44779 );
xor \U$36725 ( \44781 , \44658 , \44780 );
buf \U$36726 ( \44782 , \44781 );
xor \U$36727 ( \44783 , \44647 , \44782 );
and \U$36728 ( \44784 , \44535 , \44566 );
and \U$36729 ( \44785 , \44535 , \44572 );
and \U$36730 ( \44786 , \44566 , \44572 );
or \U$36731 ( \44787 , \44784 , \44785 , \44786 );
buf \U$36732 ( \44788 , \44787 );
and \U$36733 ( \44789 , \44580 , \44601 );
and \U$36734 ( \44790 , \44580 , \44623 );
and \U$36735 ( \44791 , \44601 , \44623 );
or \U$36736 ( \44792 , \44789 , \44790 , \44791 );
buf \U$36737 ( \44793 , \44792 );
xor \U$36738 ( \44794 , \44788 , \44793 );
and \U$36739 ( \44795 , \44540 , \44545 );
and \U$36740 ( \44796 , \44540 , \44564 );
and \U$36741 ( \44797 , \44545 , \44564 );
or \U$36742 ( \44798 , \44795 , \44796 , \44797 );
buf \U$36743 ( \44799 , \44798 );
and \U$36744 ( \44800 , \44449 , \44454 );
and \U$36745 ( \44801 , \44449 , \44461 );
and \U$36746 ( \44802 , \44454 , \44461 );
or \U$36747 ( \44803 , \44800 , \44801 , \44802 );
buf \U$36748 ( \44804 , \44803 );
xor \U$36749 ( \44805 , \44799 , \44804 );
and \U$36750 ( \44806 , \44608 , \44614 );
and \U$36751 ( \44807 , \44608 , \44621 );
and \U$36752 ( \44808 , \44614 , \44621 );
or \U$36753 ( \44809 , \44806 , \44807 , \44808 );
buf \U$36754 ( \44810 , \44809 );
and \U$36755 ( \44811 , \44470 , \44476 );
and \U$36756 ( \44812 , \44470 , \44483 );
and \U$36757 ( \44813 , \44476 , \44483 );
or \U$36758 ( \44814 , \44811 , \44812 , \44813 );
buf \U$36759 ( \44815 , \44814 );
xor \U$36760 ( \44816 , \44810 , \44815 );
and \U$36761 ( \44817 , \44586 , \44592 );
and \U$36762 ( \44818 , \44586 , \44599 );
and \U$36763 ( \44819 , \44592 , \44599 );
or \U$36764 ( \44820 , \44817 , \44818 , \44819 );
buf \U$36765 ( \44821 , \44820 );
xor \U$36766 ( \44822 , \44816 , \44821 );
buf \U$36767 ( \44823 , \44822 );
xor \U$36768 ( \44824 , \44805 , \44823 );
buf \U$36769 ( \44825 , \44824 );
xor \U$36770 ( \44826 , \44794 , \44825 );
buf \U$36771 ( \44827 , \44826 );
xor \U$36772 ( \44828 , \44783 , \44827 );
and \U$36773 ( \44829 , \44642 , \44828 );
and \U$36775 ( \44830 , \44636 , \44641 );
or \U$36777 ( \44831 , 1'b0 , \44830 , 1'b0 );
xor \U$36778 ( \44832 , \44829 , \44831 );
and \U$36780 ( \44833 , \44629 , \44635 );
and \U$36781 ( \44834 , \44631 , \44635 );
or \U$36782 ( \44835 , 1'b0 , \44833 , \44834 );
xor \U$36783 ( \44836 , \44832 , \44835 );
xor \U$36790 ( \44837 , \44836 , 1'b0 );
and \U$36791 ( \44838 , \44652 , \44657 );
and \U$36792 ( \44839 , \44652 , \44780 );
and \U$36793 ( \44840 , \44657 , \44780 );
or \U$36794 ( \44841 , \44838 , \44839 , \44840 );
buf \U$36795 ( \44842 , \44841 );
and \U$36796 ( \44843 , \44810 , \44815 );
and \U$36797 ( \44844 , \44810 , \44821 );
and \U$36798 ( \44845 , \44815 , \44821 );
or \U$36799 ( \44846 , \44843 , \44844 , \44845 );
buf \U$36800 ( \44847 , \44846 );
and \U$36801 ( \44848 , \24792 , \38968_nG9b7e );
and \U$36802 ( \44849 , \24789 , \39334_nG9b7b );
or \U$36803 ( \44850 , \44848 , \44849 );
xor \U$36804 ( \44851 , \24788 , \44850 );
buf \U$36805 ( \44852 , \44851 );
buf \U$36807 ( \44853 , \44852 );
and \U$36808 ( \44854 , \23201 , \39591_nG9b78 );
and \U$36809 ( \44855 , \23198 , \39963_nG9b75 );
or \U$36810 ( \44856 , \44854 , \44855 );
xor \U$36811 ( \44857 , \23197 , \44856 );
buf \U$36812 ( \44858 , \44857 );
buf \U$36814 ( \44859 , \44858 );
xor \U$36815 ( \44860 , \44853 , \44859 );
and \U$36816 ( \44861 , \17297 , \41963_nG9b60 );
and \U$36817 ( \44862 , \17294 , \42201_nG9b5d );
or \U$36818 ( \44863 , \44861 , \44862 );
xor \U$36819 ( \44864 , \17293 , \44863 );
buf \U$36820 ( \44865 , \44864 );
buf \U$36822 ( \44866 , \44865 );
xor \U$36823 ( \44867 , \44860 , \44866 );
buf \U$36824 ( \44868 , \44867 );
and \U$36825 ( \44869 , \44729 , \44735 );
and \U$36826 ( \44870 , \44729 , \44742 );
and \U$36827 ( \44871 , \44735 , \44742 );
or \U$36828 ( \44872 , \44869 , \44870 , \44871 );
buf \U$36829 ( \44873 , \44872 );
xor \U$36830 ( \44874 , \44868 , \44873 );
and \U$36831 ( \44875 , \14631 , \42848_nG9b54 );
and \U$36832 ( \44876 , \14628 , \43179_nG9b51 );
or \U$36833 ( \44877 , \44875 , \44876 );
xor \U$36834 ( \44878 , \14627 , \44877 );
buf \U$36835 ( \44879 , \44878 );
buf \U$36837 ( \44880 , \44879 );
xor \U$36841 ( \44881 , \13366 , 1'b0 );
not \U$36842 ( \44882 , \44881 );
buf \U$36843 ( \44883 , \44882 );
buf \U$36845 ( \44884 , \44883 );
xor \U$36846 ( \44885 , \44880 , \44884 );
and \U$36848 ( \44886 , \32916 , \35801_nG9b99 );
or \U$36849 ( \44887 , 1'b0 , \44886 );
xor \U$36850 ( \44888 , 1'b0 , \44887 );
buf \U$36851 ( \44889 , \44888 );
buf \U$36853 ( \44890 , \44889 );
xor \U$36854 ( \44891 , \44885 , \44890 );
buf \U$36855 ( \44892 , \44891 );
xor \U$36856 ( \44893 , \44874 , \44892 );
buf \U$36857 ( \44894 , \44893 );
xor \U$36858 ( \44895 , \44847 , \44894 );
and \U$36859 ( \44896 , \44663 , \44670 );
and \U$36860 ( \44897 , \44663 , \44677 );
and \U$36861 ( \44898 , \44670 , \44677 );
or \U$36862 ( \44899 , \44896 , \44897 , \44898 );
buf \U$36863 ( \44900 , \44899 );
xor \U$36864 ( \44901 , \44895 , \44900 );
buf \U$36865 ( \44902 , \44901 );
and \U$36866 ( \44903 , \44799 , \44804 );
and \U$36867 ( \44904 , \44799 , \44823 );
and \U$36868 ( \44905 , \44804 , \44823 );
or \U$36869 ( \44906 , \44903 , \44904 , \44905 );
buf \U$36870 ( \44907 , \44906 );
xor \U$36871 ( \44908 , \44902 , \44907 );
and \U$36872 ( \44909 , \28118 , \37607_nG9b8a );
and \U$36873 ( \44910 , \28115 , \37974_nG9b87 );
or \U$36874 ( \44911 , \44909 , \44910 );
xor \U$36875 ( \44912 , \28114 , \44911 );
buf \U$36876 ( \44913 , \44912 );
buf \U$36878 ( \44914 , \44913 );
and \U$36879 ( \44915 , \26431 , \38337_nG9b84 );
and \U$36880 ( \44916 , \26428 , \38663_nG9b81 );
or \U$36881 ( \44917 , \44915 , \44916 );
xor \U$36882 ( \44918 , \26427 , \44917 );
buf \U$36883 ( \44919 , \44918 );
buf \U$36885 ( \44920 , \44919 );
xor \U$36886 ( \44921 , \44914 , \44920 );
and \U$36887 ( \44922 , \18702 , \41381_nG9b66 );
and \U$36888 ( \44923 , \18699 , \41685_nG9b63 );
or \U$36889 ( \44924 , \44922 , \44923 );
xor \U$36890 ( \44925 , \18698 , \44924 );
buf \U$36891 ( \44926 , \44925 );
buf \U$36893 ( \44927 , \44926 );
xor \U$36894 ( \44928 , \44921 , \44927 );
buf \U$36895 ( \44929 , \44928 );
buf \U$36896 ( \44930 , \44669 );
and \U$36897 ( \44931 , \21658 , \40204_nG9b72 );
and \U$36898 ( \44932 , \21655 , \40452_nG9b6f );
or \U$36899 ( \44933 , \44931 , \44932 );
xor \U$36900 ( \44934 , \21654 , \44933 );
buf \U$36901 ( \44935 , \44934 );
buf \U$36903 ( \44936 , \44935 );
xor \U$36904 ( \44937 , \44930 , \44936 );
and \U$36905 ( \44938 , \15940 , \42433_nG9b5a );
and \U$36906 ( \44939 , \15937 , \42766_nG9b57 );
or \U$36907 ( \44940 , \44938 , \44939 );
xor \U$36908 ( \44941 , \15936 , \44940 );
buf \U$36909 ( \44942 , \44941 );
buf \U$36911 ( \44943 , \44942 );
xor \U$36912 ( \44944 , \44937 , \44943 );
buf \U$36913 ( \44945 , \44944 );
xor \U$36914 ( \44946 , \44929 , \44945 );
and \U$36915 ( \44947 , \31636 , \36172_nG9b96 );
and \U$36916 ( \44948 , \31633 , \36589_nG9b93 );
or \U$36917 ( \44949 , \44947 , \44948 );
xor \U$36918 ( \44950 , \31632 , \44949 );
buf \U$36919 ( \44951 , \44950 );
buf \U$36921 ( \44952 , \44951 );
and \U$36922 ( \44953 , \29853 , \36986_nG9b90 );
and \U$36923 ( \44954 , \29850 , \37250_nG9b8d );
or \U$36924 ( \44955 , \44953 , \44954 );
xor \U$36925 ( \44956 , \29849 , \44955 );
buf \U$36926 ( \44957 , \44956 );
buf \U$36928 ( \44958 , \44957 );
xor \U$36929 ( \44959 , \44952 , \44958 );
and \U$36930 ( \44960 , \20155 , \40843_nG9b6c );
and \U$36931 ( \44961 , \20152 , \41040_nG9b69 );
or \U$36932 ( \44962 , \44960 , \44961 );
xor \U$36933 ( \44963 , \20151 , \44962 );
buf \U$36934 ( \44964 , \44963 );
buf \U$36936 ( \44965 , \44964 );
xor \U$36937 ( \44966 , \44959 , \44965 );
buf \U$36938 ( \44967 , \44966 );
xor \U$36939 ( \44968 , \44946 , \44967 );
buf \U$36940 ( \44969 , \44968 );
xor \U$36941 ( \44970 , \44908 , \44969 );
buf \U$36942 ( \44971 , \44970 );
xor \U$36943 ( \44972 , \44842 , \44971 );
and \U$36944 ( \44973 , \44788 , \44793 );
and \U$36945 ( \44974 , \44788 , \44825 );
and \U$36946 ( \44975 , \44793 , \44825 );
or \U$36947 ( \44976 , \44973 , \44974 , \44975 );
buf \U$36948 ( \44977 , \44976 );
and \U$36949 ( \44978 , \44724 , \44772 );
and \U$36950 ( \44979 , \44724 , \44778 );
and \U$36951 ( \44980 , \44772 , \44778 );
or \U$36952 ( \44981 , \44978 , \44979 , \44980 );
buf \U$36953 ( \44982 , \44981 );
xor \U$36954 ( \44983 , \44977 , \44982 );
and \U$36955 ( \44984 , \44744 , \44749 );
and \U$36956 ( \44985 , \44744 , \44770 );
and \U$36957 ( \44986 , \44749 , \44770 );
or \U$36958 ( \44987 , \44984 , \44985 , \44986 );
buf \U$36959 ( \44988 , \44987 );
and \U$36960 ( \44989 , \44685 , \44691 );
and \U$36961 ( \44990 , \44685 , \44698 );
and \U$36962 ( \44991 , \44691 , \44698 );
or \U$36963 ( \44992 , \44989 , \44990 , \44991 );
buf \U$36964 ( \44993 , \44992 );
and \U$36965 ( \44994 , \44755 , \44761 );
and \U$36966 ( \44995 , \44755 , \44768 );
and \U$36967 ( \44996 , \44761 , \44768 );
or \U$36968 ( \44997 , \44994 , \44995 , \44996 );
buf \U$36969 ( \44998 , \44997 );
xor \U$36970 ( \44999 , \44993 , \44998 );
and \U$36971 ( \45000 , \44707 , \44713 );
and \U$36972 ( \45001 , \44707 , \44720 );
and \U$36973 ( \45002 , \44713 , \44720 );
or \U$36974 ( \45003 , \45000 , \45001 , \45002 );
buf \U$36975 ( \45004 , \45003 );
xor \U$36976 ( \45005 , \44999 , \45004 );
buf \U$36977 ( \45006 , \45005 );
xor \U$36978 ( \45007 , \44988 , \45006 );
and \U$36979 ( \45008 , \44679 , \44700 );
and \U$36980 ( \45009 , \44679 , \44722 );
and \U$36981 ( \45010 , \44700 , \44722 );
or \U$36982 ( \45011 , \45008 , \45009 , \45010 );
buf \U$36983 ( \45012 , \45011 );
xor \U$36984 ( \45013 , \45007 , \45012 );
buf \U$36985 ( \45014 , \45013 );
xor \U$36986 ( \45015 , \44983 , \45014 );
buf \U$36987 ( \45016 , \45015 );
xor \U$36988 ( \45017 , \44972 , \45016 );
xor \U$36989 ( \45018 , \44837 , \45017 );
and \U$36990 ( \45019 , \44647 , \44782 );
and \U$36991 ( \45020 , \44647 , \44827 );
and \U$36992 ( \45021 , \44782 , \44827 );
or \U$36993 ( \45022 , \45019 , \45020 , \45021 );
and \U$36994 ( \45023 , \45018 , \45022 );
and \U$36996 ( \45024 , \44836 , \45017 );
or \U$36998 ( \45025 , 1'b0 , \45024 , 1'b0 );
xor \U$36999 ( \45026 , \45023 , \45025 );
and \U$37001 ( \45027 , \44829 , \44835 );
and \U$37002 ( \45028 , \44831 , \44835 );
or \U$37003 ( \45029 , 1'b0 , \45027 , \45028 );
xor \U$37004 ( \45030 , \45026 , \45029 );
xor \U$37011 ( \45031 , \45030 , 1'b0 );
and \U$37012 ( \45032 , \44842 , \44971 );
and \U$37013 ( \45033 , \44842 , \45016 );
and \U$37014 ( \45034 , \44971 , \45016 );
or \U$37015 ( \45035 , \45032 , \45033 , \45034 );
xor \U$37016 ( \45036 , \45031 , \45035 );
and \U$37017 ( \45037 , \44977 , \44982 );
and \U$37018 ( \45038 , \44977 , \45014 );
and \U$37019 ( \45039 , \44982 , \45014 );
or \U$37020 ( \45040 , \45037 , \45038 , \45039 );
buf \U$37021 ( \45041 , \45040 );
and \U$37022 ( \45042 , \44902 , \44907 );
and \U$37023 ( \45043 , \44902 , \44969 );
and \U$37024 ( \45044 , \44907 , \44969 );
or \U$37025 ( \45045 , \45042 , \45043 , \45044 );
buf \U$37026 ( \45046 , \45045 );
and \U$37027 ( \45047 , \31636 , \36589_nG9b93 );
and \U$37028 ( \45048 , \31633 , \36986_nG9b90 );
or \U$37029 ( \45049 , \45047 , \45048 );
xor \U$37030 ( \45050 , \31632 , \45049 );
buf \U$37031 ( \45051 , \45050 );
buf \U$37033 ( \45052 , \45051 );
and \U$37034 ( \45053 , \21658 , \40452_nG9b6f );
and \U$37035 ( \45054 , \21655 , \40843_nG9b6c );
or \U$37036 ( \45055 , \45053 , \45054 );
xor \U$37037 ( \45056 , \21654 , \45055 );
buf \U$37038 ( \45057 , \45056 );
buf \U$37040 ( \45058 , \45057 );
xor \U$37041 ( \45059 , \45052 , \45058 );
and \U$37042 ( \45060 , \17297 , \42201_nG9b5d );
and \U$37043 ( \45061 , \17294 , \42433_nG9b5a );
or \U$37044 ( \45062 , \45060 , \45061 );
xor \U$37045 ( \45063 , \17293 , \45062 );
buf \U$37046 ( \45064 , \45063 );
buf \U$37048 ( \45065 , \45064 );
xor \U$37049 ( \45066 , \45059 , \45065 );
buf \U$37050 ( \45067 , \45066 );
and \U$37051 ( \45068 , \29853 , \37250_nG9b8d );
and \U$37052 ( \45069 , \29850 , \37607_nG9b8a );
or \U$37053 ( \45070 , \45068 , \45069 );
xor \U$37054 ( \45071 , \29849 , \45070 );
buf \U$37055 ( \45072 , \45071 );
buf \U$37057 ( \45073 , \45072 );
and \U$37058 ( \45074 , \28118 , \37974_nG9b87 );
and \U$37059 ( \45075 , \28115 , \38337_nG9b84 );
or \U$37060 ( \45076 , \45074 , \45075 );
xor \U$37061 ( \45077 , \28114 , \45076 );
buf \U$37062 ( \45078 , \45077 );
buf \U$37064 ( \45079 , \45078 );
xor \U$37065 ( \45080 , \45073 , \45079 );
and \U$37066 ( \45081 , \20155 , \41040_nG9b69 );
and \U$37067 ( \45082 , \20152 , \41381_nG9b66 );
or \U$37068 ( \45083 , \45081 , \45082 );
xor \U$37069 ( \45084 , \20151 , \45083 );
buf \U$37070 ( \45085 , \45084 );
buf \U$37072 ( \45086 , \45085 );
xor \U$37073 ( \45087 , \45080 , \45086 );
buf \U$37074 ( \45088 , \45087 );
xor \U$37075 ( \45089 , \45067 , \45088 );
and \U$37076 ( \45090 , \14631 , \43179_nG9b51 );
or \U$37078 ( \45091 , \45090 , 1'b0 );
xor \U$37079 ( \45092 , \14627 , \45091 );
buf \U$37080 ( \45093 , \45092 );
buf \U$37082 ( \45094 , \45093 );
and \U$37084 ( \45095 , \32916 , \36172_nG9b96 );
or \U$37085 ( \45096 , 1'b0 , \45095 );
xor \U$37086 ( \45097 , 1'b0 , \45096 );
buf \U$37087 ( \45098 , \45097 );
buf \U$37088 ( \45099 , \45098 );
not \U$37089 ( \45100 , \45099 );
xor \U$37090 ( \45101 , \45094 , \45100 );
and \U$37091 ( \45102 , \23201 , \39963_nG9b75 );
and \U$37092 ( \45103 , \23198 , \40204_nG9b72 );
or \U$37093 ( \45104 , \45102 , \45103 );
xor \U$37094 ( \45105 , \23197 , \45104 );
buf \U$37095 ( \45106 , \45105 );
buf \U$37097 ( \45107 , \45106 );
xor \U$37098 ( \45108 , \45101 , \45107 );
buf \U$37099 ( \45109 , \45108 );
xor \U$37100 ( \45110 , \45089 , \45109 );
buf \U$37101 ( \45111 , \45110 );
and \U$37102 ( \45112 , \44868 , \44873 );
and \U$37103 ( \45113 , \44868 , \44892 );
and \U$37104 ( \45114 , \44873 , \44892 );
or \U$37105 ( \45115 , \45112 , \45113 , \45114 );
buf \U$37106 ( \45116 , \45115 );
xor \U$37107 ( \45117 , \45111 , \45116 );
and \U$37108 ( \45118 , \44930 , \44936 );
and \U$37109 ( \45119 , \44930 , \44943 );
and \U$37110 ( \45120 , \44936 , \44943 );
or \U$37111 ( \45121 , \45118 , \45119 , \45120 );
buf \U$37112 ( \45122 , \45121 );
and \U$37113 ( \45123 , \44880 , \44884 );
and \U$37114 ( \45124 , \44880 , \44890 );
and \U$37115 ( \45125 , \44884 , \44890 );
or \U$37116 ( \45126 , \45123 , \45124 , \45125 );
buf \U$37117 ( \45127 , \45126 );
xor \U$37118 ( \45128 , \45122 , \45127 );
and \U$37119 ( \45129 , \44952 , \44958 );
and \U$37120 ( \45130 , \44952 , \44965 );
and \U$37121 ( \45131 , \44958 , \44965 );
or \U$37122 ( \45132 , \45129 , \45130 , \45131 );
buf \U$37123 ( \45133 , \45132 );
xor \U$37124 ( \45134 , \45128 , \45133 );
buf \U$37125 ( \45135 , \45134 );
xor \U$37126 ( \45136 , \45117 , \45135 );
buf \U$37127 ( \45137 , \45136 );
xor \U$37128 ( \45138 , \45046 , \45137 );
and \U$37129 ( \45139 , \44988 , \45006 );
and \U$37130 ( \45140 , \44988 , \45012 );
and \U$37131 ( \45141 , \45006 , \45012 );
or \U$37132 ( \45142 , \45139 , \45140 , \45141 );
buf \U$37133 ( \45143 , \45142 );
xor \U$37134 ( \45144 , \45138 , \45143 );
buf \U$37135 ( \45145 , \45144 );
xor \U$37136 ( \45146 , \45041 , \45145 );
and \U$37137 ( \45147 , \44847 , \44894 );
and \U$37138 ( \45148 , \44847 , \44900 );
and \U$37139 ( \45149 , \44894 , \44900 );
or \U$37140 ( \45150 , \45147 , \45148 , \45149 );
buf \U$37141 ( \45151 , \45150 );
and \U$37142 ( \45152 , \44853 , \44859 );
and \U$37143 ( \45153 , \44853 , \44866 );
and \U$37144 ( \45154 , \44859 , \44866 );
or \U$37145 ( \45155 , \45152 , \45153 , \45154 );
buf \U$37146 ( \45156 , \45155 );
and \U$37147 ( \45157 , \44914 , \44920 );
and \U$37148 ( \45158 , \44914 , \44927 );
and \U$37149 ( \45159 , \44920 , \44927 );
or \U$37150 ( \45160 , \45157 , \45158 , \45159 );
buf \U$37151 ( \45161 , \45160 );
xor \U$37152 ( \45162 , \45156 , \45161 );
and \U$37153 ( \45163 , \15940 , \42766_nG9b57 );
and \U$37154 ( \45164 , \15937 , \42848_nG9b54 );
or \U$37155 ( \45165 , \45163 , \45164 );
xor \U$37156 ( \45166 , \15936 , \45165 );
buf \U$37157 ( \45167 , \45166 );
buf \U$37159 ( \45168 , \45167 );
xor \U$37160 ( \45169 , \45162 , \45168 );
buf \U$37161 ( \45170 , \45169 );
and \U$37162 ( \45171 , \44993 , \44998 );
and \U$37163 ( \45172 , \44993 , \45004 );
and \U$37164 ( \45173 , \44998 , \45004 );
or \U$37165 ( \45174 , \45171 , \45172 , \45173 );
buf \U$37166 ( \45175 , \45174 );
xor \U$37167 ( \45176 , \45170 , \45175 );
and \U$37168 ( \45177 , \26431 , \38663_nG9b81 );
and \U$37169 ( \45178 , \26428 , \38968_nG9b7e );
or \U$37170 ( \45179 , \45177 , \45178 );
xor \U$37171 ( \45180 , \26427 , \45179 );
buf \U$37172 ( \45181 , \45180 );
buf \U$37174 ( \45182 , \45181 );
and \U$37175 ( \45183 , \24792 , \39334_nG9b7b );
and \U$37176 ( \45184 , \24789 , \39591_nG9b78 );
or \U$37177 ( \45185 , \45183 , \45184 );
xor \U$37178 ( \45186 , \24788 , \45185 );
buf \U$37179 ( \45187 , \45186 );
buf \U$37181 ( \45188 , \45187 );
xor \U$37182 ( \45189 , \45182 , \45188 );
and \U$37183 ( \45190 , \18702 , \41685_nG9b63 );
and \U$37184 ( \45191 , \18699 , \41963_nG9b60 );
or \U$37185 ( \45192 , \45190 , \45191 );
xor \U$37186 ( \45193 , \18698 , \45192 );
buf \U$37187 ( \45194 , \45193 );
buf \U$37189 ( \45195 , \45194 );
xor \U$37190 ( \45196 , \45189 , \45195 );
buf \U$37191 ( \45197 , \45196 );
xor \U$37192 ( \45198 , \45176 , \45197 );
buf \U$37193 ( \45199 , \45198 );
xor \U$37194 ( \45200 , \45151 , \45199 );
and \U$37195 ( \45201 , \44929 , \44945 );
and \U$37196 ( \45202 , \44929 , \44967 );
and \U$37197 ( \45203 , \44945 , \44967 );
or \U$37198 ( \45204 , \45201 , \45202 , \45203 );
buf \U$37199 ( \45205 , \45204 );
xor \U$37200 ( \45206 , \45200 , \45205 );
buf \U$37201 ( \45207 , \45206 );
xor \U$37202 ( \45208 , \45146 , \45207 );
and \U$37203 ( \45209 , \45036 , \45208 );
and \U$37205 ( \45210 , \45030 , \45035 );
or \U$37207 ( \45211 , 1'b0 , \45210 , 1'b0 );
xor \U$37208 ( \45212 , \45209 , \45211 );
and \U$37210 ( \45213 , \45023 , \45029 );
and \U$37211 ( \45214 , \45025 , \45029 );
or \U$37212 ( \45215 , 1'b0 , \45213 , \45214 );
xor \U$37213 ( \45216 , \45212 , \45215 );
xor \U$37220 ( \45217 , \45216 , 1'b0 );
and \U$37221 ( \45218 , \45041 , \45145 );
and \U$37222 ( \45219 , \45041 , \45207 );
and \U$37223 ( \45220 , \45145 , \45207 );
or \U$37224 ( \45221 , \45218 , \45219 , \45220 );
xor \U$37225 ( \45222 , \45217 , \45221 );
and \U$37226 ( \45223 , \45067 , \45088 );
and \U$37227 ( \45224 , \45067 , \45109 );
and \U$37228 ( \45225 , \45088 , \45109 );
or \U$37229 ( \45226 , \45223 , \45224 , \45225 );
buf \U$37230 ( \45227 , \45226 );
and \U$37231 ( \45228 , \45052 , \45058 );
and \U$37232 ( \45229 , \45052 , \45065 );
and \U$37233 ( \45230 , \45058 , \45065 );
or \U$37234 ( \45231 , \45228 , \45229 , \45230 );
buf \U$37235 ( \45232 , \45231 );
and \U$37236 ( \45233 , \45094 , \45100 );
and \U$37237 ( \45234 , \45094 , \45107 );
and \U$37238 ( \45235 , \45100 , \45107 );
or \U$37239 ( \45236 , \45233 , \45234 , \45235 );
buf \U$37240 ( \45237 , \45236 );
xor \U$37241 ( \45238 , \45232 , \45237 );
and \U$37242 ( \45239 , \45182 , \45188 );
and \U$37243 ( \45240 , \45182 , \45195 );
and \U$37244 ( \45241 , \45188 , \45195 );
or \U$37245 ( \45242 , \45239 , \45240 , \45241 );
buf \U$37246 ( \45243 , \45242 );
xor \U$37247 ( \45244 , \45238 , \45243 );
buf \U$37248 ( \45245 , \45244 );
xor \U$37249 ( \45246 , \45227 , \45245 );
and \U$37250 ( \45247 , \45122 , \45127 );
and \U$37251 ( \45248 , \45122 , \45133 );
and \U$37252 ( \45249 , \45127 , \45133 );
or \U$37253 ( \45250 , \45247 , \45248 , \45249 );
buf \U$37254 ( \45251 , \45250 );
xor \U$37255 ( \45252 , \45246 , \45251 );
buf \U$37256 ( \45253 , \45252 );
and \U$37257 ( \45254 , \45111 , \45116 );
and \U$37258 ( \45255 , \45111 , \45135 );
and \U$37259 ( \45256 , \45116 , \45135 );
or \U$37260 ( \45257 , \45254 , \45255 , \45256 );
buf \U$37261 ( \45258 , \45257 );
xor \U$37262 ( \45259 , \45253 , \45258 );
and \U$37263 ( \45260 , \45151 , \45199 );
and \U$37264 ( \45261 , \45151 , \45205 );
and \U$37265 ( \45262 , \45199 , \45205 );
or \U$37266 ( \45263 , \45260 , \45261 , \45262 );
buf \U$37267 ( \45264 , \45263 );
xor \U$37268 ( \45265 , \45259 , \45264 );
buf \U$37269 ( \45266 , \45265 );
and \U$37270 ( \45267 , \45046 , \45137 );
and \U$37271 ( \45268 , \45046 , \45143 );
and \U$37272 ( \45269 , \45137 , \45143 );
or \U$37273 ( \45270 , \45267 , \45268 , \45269 );
buf \U$37274 ( \45271 , \45270 );
xor \U$37275 ( \45272 , \45266 , \45271 );
and \U$37276 ( \45273 , \45073 , \45079 );
and \U$37277 ( \45274 , \45073 , \45086 );
and \U$37278 ( \45275 , \45079 , \45086 );
or \U$37279 ( \45276 , \45273 , \45274 , \45275 );
buf \U$37280 ( \45277 , \45276 );
buf \U$37281 ( \45278 , \45099 );
xor \U$37282 ( \45279 , \45277 , \45278 );
and \U$37283 ( \45280 , \17297 , \42433_nG9b5a );
and \U$37284 ( \45281 , \17294 , \42766_nG9b57 );
or \U$37285 ( \45282 , \45280 , \45281 );
xor \U$37286 ( \45283 , \17293 , \45282 );
buf \U$37287 ( \45284 , \45283 );
buf \U$37289 ( \45285 , \45284 );
xor \U$37290 ( \45286 , \45279 , \45285 );
buf \U$37291 ( \45287 , \45286 );
and \U$37292 ( \45288 , \45156 , \45161 );
and \U$37293 ( \45289 , \45156 , \45168 );
and \U$37294 ( \45290 , \45161 , \45168 );
or \U$37295 ( \45291 , \45288 , \45289 , \45290 );
buf \U$37296 ( \45292 , \45291 );
xor \U$37297 ( \45293 , \45287 , \45292 );
and \U$37299 ( \45294 , \32916 , \36589_nG9b93 );
or \U$37300 ( \45295 , 1'b0 , \45294 );
xor \U$37301 ( \45296 , 1'b0 , \45295 );
buf \U$37302 ( \45297 , \45296 );
buf \U$37304 ( \45298 , \45297 );
and \U$37305 ( \45299 , \31636 , \36986_nG9b90 );
and \U$37306 ( \45300 , \31633 , \37250_nG9b8d );
or \U$37307 ( \45301 , \45299 , \45300 );
xor \U$37308 ( \45302 , \31632 , \45301 );
buf \U$37309 ( \45303 , \45302 );
buf \U$37311 ( \45304 , \45303 );
xor \U$37312 ( \45305 , \45298 , \45304 );
and \U$37313 ( \45306 , \23201 , \40204_nG9b72 );
and \U$37314 ( \45307 , \23198 , \40452_nG9b6f );
or \U$37315 ( \45308 , \45306 , \45307 );
xor \U$37316 ( \45309 , \23197 , \45308 );
buf \U$37317 ( \45310 , \45309 );
buf \U$37319 ( \45311 , \45310 );
xor \U$37320 ( \45312 , \45305 , \45311 );
buf \U$37321 ( \45313 , \45312 );
xor \U$37322 ( \45314 , \45293 , \45313 );
buf \U$37323 ( \45315 , \45314 );
and \U$37324 ( \45316 , \45170 , \45175 );
and \U$37325 ( \45317 , \45170 , \45197 );
and \U$37326 ( \45318 , \45175 , \45197 );
or \U$37327 ( \45319 , \45316 , \45317 , \45318 );
buf \U$37328 ( \45320 , \45319 );
xor \U$37329 ( \45321 , \45315 , \45320 );
and \U$37330 ( \45322 , \26431 , \38968_nG9b7e );
and \U$37331 ( \45323 , \26428 , \39334_nG9b7b );
or \U$37332 ( \45324 , \45322 , \45323 );
xor \U$37333 ( \45325 , \26427 , \45324 );
buf \U$37334 ( \45326 , \45325 );
buf \U$37336 ( \45327 , \45326 );
and \U$37337 ( \45328 , \24792 , \39591_nG9b78 );
and \U$37338 ( \45329 , \24789 , \39963_nG9b75 );
or \U$37339 ( \45330 , \45328 , \45329 );
xor \U$37340 ( \45331 , \24788 , \45330 );
buf \U$37341 ( \45332 , \45331 );
buf \U$37343 ( \45333 , \45332 );
xor \U$37344 ( \45334 , \45327 , \45333 );
and \U$37345 ( \45335 , \20155 , \41381_nG9b66 );
and \U$37346 ( \45336 , \20152 , \41685_nG9b63 );
or \U$37347 ( \45337 , \45335 , \45336 );
xor \U$37348 ( \45338 , \20151 , \45337 );
buf \U$37349 ( \45339 , \45338 );
buf \U$37351 ( \45340 , \45339 );
xor \U$37352 ( \45341 , \45334 , \45340 );
buf \U$37353 ( \45342 , \45341 );
and \U$37354 ( \45343 , \15940 , \42848_nG9b54 );
and \U$37355 ( \45344 , \15937 , \43179_nG9b51 );
or \U$37356 ( \45345 , \45343 , \45344 );
xor \U$37357 ( \45346 , \15936 , \45345 );
buf \U$37358 ( \45347 , \45346 );
buf \U$37360 ( \45348 , \45347 );
xor \U$37364 ( \45349 , \14627 , 1'b0 );
not \U$37365 ( \45350 , \45349 );
buf \U$37366 ( \45351 , \45350 );
buf \U$37368 ( \45352 , \45351 );
xor \U$37369 ( \45353 , \45348 , \45352 );
and \U$37370 ( \45354 , \18702 , \41963_nG9b60 );
and \U$37371 ( \45355 , \18699 , \42201_nG9b5d );
or \U$37372 ( \45356 , \45354 , \45355 );
xor \U$37373 ( \45357 , \18698 , \45356 );
buf \U$37374 ( \45358 , \45357 );
buf \U$37376 ( \45359 , \45358 );
xor \U$37377 ( \45360 , \45353 , \45359 );
buf \U$37378 ( \45361 , \45360 );
xor \U$37379 ( \45362 , \45342 , \45361 );
and \U$37380 ( \45363 , \29853 , \37607_nG9b8a );
and \U$37381 ( \45364 , \29850 , \37974_nG9b87 );
or \U$37382 ( \45365 , \45363 , \45364 );
xor \U$37383 ( \45366 , \29849 , \45365 );
buf \U$37384 ( \45367 , \45366 );
buf \U$37386 ( \45368 , \45367 );
and \U$37387 ( \45369 , \28118 , \38337_nG9b84 );
and \U$37388 ( \45370 , \28115 , \38663_nG9b81 );
or \U$37389 ( \45371 , \45369 , \45370 );
xor \U$37390 ( \45372 , \28114 , \45371 );
buf \U$37391 ( \45373 , \45372 );
buf \U$37393 ( \45374 , \45373 );
xor \U$37394 ( \45375 , \45368 , \45374 );
and \U$37395 ( \45376 , \21658 , \40843_nG9b6c );
and \U$37396 ( \45377 , \21655 , \41040_nG9b69 );
or \U$37397 ( \45378 , \45376 , \45377 );
xor \U$37398 ( \45379 , \21654 , \45378 );
buf \U$37399 ( \45380 , \45379 );
buf \U$37401 ( \45381 , \45380 );
xor \U$37402 ( \45382 , \45375 , \45381 );
buf \U$37403 ( \45383 , \45382 );
xor \U$37404 ( \45384 , \45362 , \45383 );
buf \U$37405 ( \45385 , \45384 );
xor \U$37406 ( \45386 , \45321 , \45385 );
buf \U$37407 ( \45387 , \45386 );
xor \U$37408 ( \45388 , \45272 , \45387 );
and \U$37409 ( \45389 , \45222 , \45388 );
and \U$37411 ( \45390 , \45216 , \45221 );
or \U$37413 ( \45391 , 1'b0 , \45390 , 1'b0 );
xor \U$37414 ( \45392 , \45389 , \45391 );
and \U$37416 ( \45393 , \45209 , \45215 );
and \U$37417 ( \45394 , \45211 , \45215 );
or \U$37418 ( \45395 , 1'b0 , \45393 , \45394 );
xor \U$37419 ( \45396 , \45392 , \45395 );
xor \U$37426 ( \45397 , \45396 , 1'b0 );
and \U$37427 ( \45398 , \45266 , \45271 );
and \U$37428 ( \45399 , \45266 , \45387 );
and \U$37429 ( \45400 , \45271 , \45387 );
or \U$37430 ( \45401 , \45398 , \45399 , \45400 );
xor \U$37431 ( \45402 , \45397 , \45401 );
and \U$37432 ( \45403 , \45277 , \45278 );
and \U$37433 ( \45404 , \45277 , \45285 );
and \U$37434 ( \45405 , \45278 , \45285 );
or \U$37435 ( \45406 , \45403 , \45404 , \45405 );
buf \U$37436 ( \45407 , \45406 );
and \U$37437 ( \45408 , \24792 , \39963_nG9b75 );
and \U$37438 ( \45409 , \24789 , \40204_nG9b72 );
or \U$37439 ( \45410 , \45408 , \45409 );
xor \U$37440 ( \45411 , \24788 , \45410 );
buf \U$37441 ( \45412 , \45411 );
buf \U$37443 ( \45413 , \45412 );
and \U$37444 ( \45414 , \20155 , \41685_nG9b63 );
and \U$37445 ( \45415 , \20152 , \41963_nG9b60 );
or \U$37446 ( \45416 , \45414 , \45415 );
xor \U$37447 ( \45417 , \20151 , \45416 );
buf \U$37448 ( \45418 , \45417 );
buf \U$37449 ( \45419 , \45418 );
not \U$37450 ( \45420 , \45419 );
xor \U$37451 ( \45421 , \45413 , \45420 );
and \U$37452 ( \45422 , \17297 , \42766_nG9b57 );
and \U$37453 ( \45423 , \17294 , \42848_nG9b54 );
or \U$37454 ( \45424 , \45422 , \45423 );
xor \U$37455 ( \45425 , \17293 , \45424 );
buf \U$37456 ( \45426 , \45425 );
buf \U$37458 ( \45427 , \45426 );
xor \U$37459 ( \45428 , \45421 , \45427 );
buf \U$37460 ( \45429 , \45428 );
xor \U$37461 ( \45430 , \45407 , \45429 );
and \U$37462 ( \45431 , \28118 , \38663_nG9b81 );
and \U$37463 ( \45432 , \28115 , \38968_nG9b7e );
or \U$37464 ( \45433 , \45431 , \45432 );
xor \U$37465 ( \45434 , \28114 , \45433 );
buf \U$37466 ( \45435 , \45434 );
buf \U$37468 ( \45436 , \45435 );
and \U$37469 ( \45437 , \26431 , \39334_nG9b7b );
and \U$37470 ( \45438 , \26428 , \39591_nG9b78 );
or \U$37471 ( \45439 , \45437 , \45438 );
xor \U$37472 ( \45440 , \26427 , \45439 );
buf \U$37473 ( \45441 , \45440 );
buf \U$37475 ( \45442 , \45441 );
xor \U$37476 ( \45443 , \45436 , \45442 );
and \U$37477 ( \45444 , \21658 , \41040_nG9b69 );
and \U$37478 ( \45445 , \21655 , \41381_nG9b66 );
or \U$37479 ( \45446 , \45444 , \45445 );
xor \U$37480 ( \45447 , \21654 , \45446 );
buf \U$37481 ( \45448 , \45447 );
buf \U$37483 ( \45449 , \45448 );
xor \U$37484 ( \45450 , \45443 , \45449 );
buf \U$37485 ( \45451 , \45450 );
xor \U$37486 ( \45452 , \45430 , \45451 );
buf \U$37487 ( \45453 , \45452 );
and \U$37488 ( \45454 , \45287 , \45292 );
and \U$37489 ( \45455 , \45287 , \45313 );
and \U$37490 ( \45456 , \45292 , \45313 );
or \U$37491 ( \45457 , \45454 , \45455 , \45456 );
buf \U$37492 ( \45458 , \45457 );
xor \U$37493 ( \45459 , \45453 , \45458 );
and \U$37494 ( \45460 , \15940 , \43179_nG9b51 );
or \U$37496 ( \45461 , \45460 , 1'b0 );
xor \U$37497 ( \45462 , \15936 , \45461 );
buf \U$37498 ( \45463 , \45462 );
buf \U$37500 ( \45464 , \45463 );
and \U$37501 ( \45465 , \31636 , \37250_nG9b8d );
and \U$37502 ( \45466 , \31633 , \37607_nG9b8a );
or \U$37503 ( \45467 , \45465 , \45466 );
xor \U$37504 ( \45468 , \31632 , \45467 );
buf \U$37505 ( \45469 , \45468 );
buf \U$37507 ( \45470 , \45469 );
xor \U$37508 ( \45471 , \45464 , \45470 );
and \U$37509 ( \45472 , \29853 , \37974_nG9b87 );
and \U$37510 ( \45473 , \29850 , \38337_nG9b84 );
or \U$37511 ( \45474 , \45472 , \45473 );
xor \U$37512 ( \45475 , \29849 , \45474 );
buf \U$37513 ( \45476 , \45475 );
buf \U$37515 ( \45477 , \45476 );
xor \U$37516 ( \45478 , \45471 , \45477 );
buf \U$37517 ( \45479 , \45478 );
and \U$37519 ( \45480 , \32916 , \36986_nG9b90 );
or \U$37520 ( \45481 , 1'b0 , \45480 );
xor \U$37521 ( \45482 , 1'b0 , \45481 );
buf \U$37522 ( \45483 , \45482 );
buf \U$37524 ( \45484 , \45483 );
and \U$37525 ( \45485 , \23201 , \40452_nG9b6f );
and \U$37526 ( \45486 , \23198 , \40843_nG9b6c );
or \U$37527 ( \45487 , \45485 , \45486 );
xor \U$37528 ( \45488 , \23197 , \45487 );
buf \U$37529 ( \45489 , \45488 );
buf \U$37531 ( \45490 , \45489 );
xor \U$37532 ( \45491 , \45484 , \45490 );
and \U$37533 ( \45492 , \18702 , \42201_nG9b5d );
and \U$37534 ( \45493 , \18699 , \42433_nG9b5a );
or \U$37535 ( \45494 , \45492 , \45493 );
xor \U$37536 ( \45495 , \18698 , \45494 );
buf \U$37537 ( \45496 , \45495 );
buf \U$37539 ( \45497 , \45496 );
xor \U$37540 ( \45498 , \45491 , \45497 );
buf \U$37541 ( \45499 , \45498 );
xor \U$37542 ( \45500 , \45479 , \45499 );
and \U$37543 ( \45501 , \45327 , \45333 );
and \U$37544 ( \45502 , \45327 , \45340 );
and \U$37545 ( \45503 , \45333 , \45340 );
or \U$37546 ( \45504 , \45501 , \45502 , \45503 );
buf \U$37547 ( \45505 , \45504 );
xor \U$37548 ( \45506 , \45500 , \45505 );
buf \U$37549 ( \45507 , \45506 );
xor \U$37550 ( \45508 , \45459 , \45507 );
buf \U$37551 ( \45509 , \45508 );
and \U$37552 ( \45510 , \45342 , \45361 );
and \U$37553 ( \45511 , \45342 , \45383 );
and \U$37554 ( \45512 , \45361 , \45383 );
or \U$37555 ( \45513 , \45510 , \45511 , \45512 );
buf \U$37556 ( \45514 , \45513 );
and \U$37557 ( \45515 , \45348 , \45352 );
and \U$37558 ( \45516 , \45348 , \45359 );
and \U$37559 ( \45517 , \45352 , \45359 );
or \U$37560 ( \45518 , \45515 , \45516 , \45517 );
buf \U$37561 ( \45519 , \45518 );
and \U$37562 ( \45520 , \45368 , \45374 );
and \U$37563 ( \45521 , \45368 , \45381 );
and \U$37564 ( \45522 , \45374 , \45381 );
or \U$37565 ( \45523 , \45520 , \45521 , \45522 );
buf \U$37566 ( \45524 , \45523 );
xor \U$37567 ( \45525 , \45519 , \45524 );
and \U$37568 ( \45526 , \45298 , \45304 );
and \U$37569 ( \45527 , \45298 , \45311 );
and \U$37570 ( \45528 , \45304 , \45311 );
or \U$37571 ( \45529 , \45526 , \45527 , \45528 );
buf \U$37572 ( \45530 , \45529 );
xor \U$37573 ( \45531 , \45525 , \45530 );
buf \U$37574 ( \45532 , \45531 );
xor \U$37575 ( \45533 , \45514 , \45532 );
and \U$37576 ( \45534 , \45232 , \45237 );
and \U$37577 ( \45535 , \45232 , \45243 );
and \U$37578 ( \45536 , \45237 , \45243 );
or \U$37579 ( \45537 , \45534 , \45535 , \45536 );
buf \U$37580 ( \45538 , \45537 );
xor \U$37581 ( \45539 , \45533 , \45538 );
buf \U$37582 ( \45540 , \45539 );
xor \U$37583 ( \45541 , \45509 , \45540 );
and \U$37584 ( \45542 , \45227 , \45245 );
and \U$37585 ( \45543 , \45227 , \45251 );
and \U$37586 ( \45544 , \45245 , \45251 );
or \U$37587 ( \45545 , \45542 , \45543 , \45544 );
buf \U$37588 ( \45546 , \45545 );
xor \U$37589 ( \45547 , \45541 , \45546 );
buf \U$37590 ( \45548 , \45547 );
and \U$37591 ( \45549 , \45253 , \45258 );
and \U$37592 ( \45550 , \45253 , \45264 );
and \U$37593 ( \45551 , \45258 , \45264 );
or \U$37594 ( \45552 , \45549 , \45550 , \45551 );
buf \U$37595 ( \45553 , \45552 );
xor \U$37596 ( \45554 , \45548 , \45553 );
and \U$37597 ( \45555 , \45315 , \45320 );
and \U$37598 ( \45556 , \45315 , \45385 );
and \U$37599 ( \45557 , \45320 , \45385 );
or \U$37600 ( \45558 , \45555 , \45556 , \45557 );
buf \U$37601 ( \45559 , \45558 );
xor \U$37602 ( \45560 , \45554 , \45559 );
and \U$37603 ( \45561 , \45402 , \45560 );
and \U$37605 ( \45562 , \45396 , \45401 );
or \U$37607 ( \45563 , 1'b0 , \45562 , 1'b0 );
xor \U$37608 ( \45564 , \45561 , \45563 );
and \U$37610 ( \45565 , \45389 , \45395 );
and \U$37611 ( \45566 , \45391 , \45395 );
or \U$37612 ( \45567 , 1'b0 , \45565 , \45566 );
xor \U$37613 ( \45568 , \45564 , \45567 );
xor \U$37620 ( \45569 , \45568 , 1'b0 );
and \U$37621 ( \45570 , \45548 , \45553 );
and \U$37622 ( \45571 , \45548 , \45559 );
and \U$37623 ( \45572 , \45553 , \45559 );
or \U$37624 ( \45573 , \45570 , \45571 , \45572 );
xor \U$37625 ( \45574 , \45569 , \45573 );
and \U$37626 ( \45575 , \45407 , \45429 );
and \U$37627 ( \45576 , \45407 , \45451 );
and \U$37628 ( \45577 , \45429 , \45451 );
or \U$37629 ( \45578 , \45575 , \45576 , \45577 );
buf \U$37630 ( \45579 , \45578 );
and \U$37631 ( \45580 , \45413 , \45420 );
and \U$37632 ( \45581 , \45413 , \45427 );
and \U$37633 ( \45582 , \45420 , \45427 );
or \U$37634 ( \45583 , \45580 , \45581 , \45582 );
buf \U$37635 ( \45584 , \45583 );
and \U$37636 ( \45585 , \28118 , \38968_nG9b7e );
and \U$37637 ( \45586 , \28115 , \39334_nG9b7b );
or \U$37638 ( \45587 , \45585 , \45586 );
xor \U$37639 ( \45588 , \28114 , \45587 );
buf \U$37640 ( \45589 , \45588 );
buf \U$37642 ( \45590 , \45589 );
and \U$37643 ( \45591 , \26431 , \39591_nG9b78 );
and \U$37644 ( \45592 , \26428 , \39963_nG9b75 );
or \U$37645 ( \45593 , \45591 , \45592 );
xor \U$37646 ( \45594 , \26427 , \45593 );
buf \U$37647 ( \45595 , \45594 );
buf \U$37649 ( \45596 , \45595 );
xor \U$37650 ( \45597 , \45590 , \45596 );
and \U$37651 ( \45598 , \21658 , \41381_nG9b66 );
and \U$37652 ( \45599 , \21655 , \41685_nG9b63 );
or \U$37653 ( \45600 , \45598 , \45599 );
xor \U$37654 ( \45601 , \21654 , \45600 );
buf \U$37655 ( \45602 , \45601 );
buf \U$37657 ( \45603 , \45602 );
xor \U$37658 ( \45604 , \45597 , \45603 );
buf \U$37659 ( \45605 , \45604 );
xor \U$37660 ( \45606 , \45584 , \45605 );
and \U$37661 ( \45607 , \17297 , \42848_nG9b54 );
and \U$37662 ( \45608 , \17294 , \43179_nG9b51 );
or \U$37663 ( \45609 , \45607 , \45608 );
xor \U$37664 ( \45610 , \17293 , \45609 );
buf \U$37665 ( \45611 , \45610 );
buf \U$37667 ( \45612 , \45611 );
xor \U$37671 ( \45613 , \15936 , 1'b0 );
not \U$37672 ( \45614 , \45613 );
buf \U$37673 ( \45615 , \45614 );
buf \U$37675 ( \45616 , \45615 );
xor \U$37676 ( \45617 , \45612 , \45616 );
and \U$37677 ( \45618 , \20155 , \41963_nG9b60 );
and \U$37678 ( \45619 , \20152 , \42201_nG9b5d );
or \U$37679 ( \45620 , \45618 , \45619 );
xor \U$37680 ( \45621 , \20151 , \45620 );
buf \U$37681 ( \45622 , \45621 );
buf \U$37683 ( \45623 , \45622 );
xor \U$37684 ( \45624 , \45617 , \45623 );
buf \U$37685 ( \45625 , \45624 );
xor \U$37686 ( \45626 , \45606 , \45625 );
buf \U$37687 ( \45627 , \45626 );
xor \U$37688 ( \45628 , \45579 , \45627 );
and \U$37690 ( \45629 , \32916 , \37250_nG9b8d );
or \U$37691 ( \45630 , 1'b0 , \45629 );
xor \U$37692 ( \45631 , 1'b0 , \45630 );
buf \U$37693 ( \45632 , \45631 );
buf \U$37695 ( \45633 , \45632 );
and \U$37696 ( \45634 , \24792 , \40204_nG9b72 );
and \U$37697 ( \45635 , \24789 , \40452_nG9b6f );
or \U$37698 ( \45636 , \45634 , \45635 );
xor \U$37699 ( \45637 , \24788 , \45636 );
buf \U$37700 ( \45638 , \45637 );
buf \U$37702 ( \45639 , \45638 );
xor \U$37703 ( \45640 , \45633 , \45639 );
and \U$37704 ( \45641 , \18702 , \42433_nG9b5a );
and \U$37705 ( \45642 , \18699 , \42766_nG9b57 );
or \U$37706 ( \45643 , \45641 , \45642 );
xor \U$37707 ( \45644 , \18698 , \45643 );
buf \U$37708 ( \45645 , \45644 );
buf \U$37710 ( \45646 , \45645 );
xor \U$37711 ( \45647 , \45640 , \45646 );
buf \U$37712 ( \45648 , \45647 );
and \U$37713 ( \45649 , \31636 , \37607_nG9b8a );
and \U$37714 ( \45650 , \31633 , \37974_nG9b87 );
or \U$37715 ( \45651 , \45649 , \45650 );
xor \U$37716 ( \45652 , \31632 , \45651 );
buf \U$37717 ( \45653 , \45652 );
buf \U$37719 ( \45654 , \45653 );
and \U$37720 ( \45655 , \29853 , \38337_nG9b84 );
and \U$37721 ( \45656 , \29850 , \38663_nG9b81 );
or \U$37722 ( \45657 , \45655 , \45656 );
xor \U$37723 ( \45658 , \29849 , \45657 );
buf \U$37724 ( \45659 , \45658 );
buf \U$37726 ( \45660 , \45659 );
xor \U$37727 ( \45661 , \45654 , \45660 );
and \U$37728 ( \45662 , \23201 , \40843_nG9b6c );
and \U$37729 ( \45663 , \23198 , \41040_nG9b69 );
or \U$37730 ( \45664 , \45662 , \45663 );
xor \U$37731 ( \45665 , \23197 , \45664 );
buf \U$37732 ( \45666 , \45665 );
buf \U$37734 ( \45667 , \45666 );
xor \U$37735 ( \45668 , \45661 , \45667 );
buf \U$37736 ( \45669 , \45668 );
xor \U$37737 ( \45670 , \45648 , \45669 );
and \U$37738 ( \45671 , \45464 , \45470 );
and \U$37739 ( \45672 , \45464 , \45477 );
and \U$37740 ( \45673 , \45470 , \45477 );
or \U$37741 ( \45674 , \45671 , \45672 , \45673 );
buf \U$37742 ( \45675 , \45674 );
xor \U$37743 ( \45676 , \45670 , \45675 );
buf \U$37744 ( \45677 , \45676 );
xor \U$37745 ( \45678 , \45628 , \45677 );
buf \U$37746 ( \45679 , \45678 );
and \U$37747 ( \45680 , \45479 , \45499 );
and \U$37748 ( \45681 , \45479 , \45505 );
and \U$37749 ( \45682 , \45499 , \45505 );
or \U$37750 ( \45683 , \45680 , \45681 , \45682 );
buf \U$37751 ( \45684 , \45683 );
and \U$37752 ( \45685 , \45519 , \45524 );
and \U$37753 ( \45686 , \45519 , \45530 );
and \U$37754 ( \45687 , \45524 , \45530 );
or \U$37755 ( \45688 , \45685 , \45686 , \45687 );
buf \U$37756 ( \45689 , \45688 );
xor \U$37757 ( \45690 , \45684 , \45689 );
and \U$37758 ( \45691 , \45484 , \45490 );
and \U$37759 ( \45692 , \45484 , \45497 );
and \U$37760 ( \45693 , \45490 , \45497 );
or \U$37761 ( \45694 , \45691 , \45692 , \45693 );
buf \U$37762 ( \45695 , \45694 );
and \U$37763 ( \45696 , \45436 , \45442 );
and \U$37764 ( \45697 , \45436 , \45449 );
and \U$37765 ( \45698 , \45442 , \45449 );
or \U$37766 ( \45699 , \45696 , \45697 , \45698 );
buf \U$37767 ( \45700 , \45699 );
xor \U$37768 ( \45701 , \45695 , \45700 );
buf \U$37769 ( \45702 , \45419 );
xor \U$37770 ( \45703 , \45701 , \45702 );
buf \U$37771 ( \45704 , \45703 );
xor \U$37772 ( \45705 , \45690 , \45704 );
buf \U$37773 ( \45706 , \45705 );
xor \U$37774 ( \45707 , \45679 , \45706 );
and \U$37775 ( \45708 , \45514 , \45532 );
and \U$37776 ( \45709 , \45514 , \45538 );
and \U$37777 ( \45710 , \45532 , \45538 );
or \U$37778 ( \45711 , \45708 , \45709 , \45710 );
buf \U$37779 ( \45712 , \45711 );
xor \U$37780 ( \45713 , \45707 , \45712 );
buf \U$37781 ( \45714 , \45713 );
and \U$37782 ( \45715 , \45509 , \45540 );
and \U$37783 ( \45716 , \45509 , \45546 );
and \U$37784 ( \45717 , \45540 , \45546 );
or \U$37785 ( \45718 , \45715 , \45716 , \45717 );
buf \U$37786 ( \45719 , \45718 );
xor \U$37787 ( \45720 , \45714 , \45719 );
and \U$37788 ( \45721 , \45453 , \45458 );
and \U$37789 ( \45722 , \45453 , \45507 );
and \U$37790 ( \45723 , \45458 , \45507 );
or \U$37791 ( \45724 , \45721 , \45722 , \45723 );
buf \U$37792 ( \45725 , \45724 );
xor \U$37793 ( \45726 , \45720 , \45725 );
and \U$37794 ( \45727 , \45574 , \45726 );
and \U$37796 ( \45728 , \45568 , \45573 );
or \U$37798 ( \45729 , 1'b0 , \45728 , 1'b0 );
xor \U$37799 ( \45730 , \45727 , \45729 );
and \U$37801 ( \45731 , \45561 , \45567 );
and \U$37802 ( \45732 , \45563 , \45567 );
or \U$37803 ( \45733 , 1'b0 , \45731 , \45732 );
xor \U$37804 ( \45734 , \45730 , \45733 );
xor \U$37811 ( \45735 , \45734 , 1'b0 );
and \U$37812 ( \45736 , \45714 , \45719 );
and \U$37813 ( \45737 , \45714 , \45725 );
and \U$37814 ( \45738 , \45719 , \45725 );
or \U$37815 ( \45739 , \45736 , \45737 , \45738 );
xor \U$37816 ( \45740 , \45735 , \45739 );
and \U$37817 ( \45741 , \45679 , \45706 );
and \U$37818 ( \45742 , \45679 , \45712 );
and \U$37819 ( \45743 , \45706 , \45712 );
or \U$37820 ( \45744 , \45741 , \45742 , \45743 );
buf \U$37821 ( \45745 , \45744 );
and \U$37822 ( \45746 , \26431 , \39963_nG9b75 );
and \U$37823 ( \45747 , \26428 , \40204_nG9b72 );
or \U$37824 ( \45748 , \45746 , \45747 );
xor \U$37825 ( \45749 , \26427 , \45748 );
buf \U$37826 ( \45750 , \45749 );
buf \U$37828 ( \45751 , \45750 );
and \U$37829 ( \45752 , \24792 , \40452_nG9b6f );
and \U$37830 ( \45753 , \24789 , \40843_nG9b6c );
or \U$37831 ( \45754 , \45752 , \45753 );
xor \U$37832 ( \45755 , \24788 , \45754 );
buf \U$37833 ( \45756 , \45755 );
buf \U$37835 ( \45757 , \45756 );
xor \U$37836 ( \45758 , \45751 , \45757 );
and \U$37837 ( \45759 , \20155 , \42201_nG9b5d );
and \U$37838 ( \45760 , \20152 , \42433_nG9b5a );
or \U$37839 ( \45761 , \45759 , \45760 );
xor \U$37840 ( \45762 , \20151 , \45761 );
buf \U$37841 ( \45763 , \45762 );
buf \U$37843 ( \45764 , \45763 );
xor \U$37844 ( \45765 , \45758 , \45764 );
buf \U$37845 ( \45766 , \45765 );
and \U$37846 ( \45767 , \29853 , \38663_nG9b81 );
and \U$37847 ( \45768 , \29850 , \38968_nG9b7e );
or \U$37848 ( \45769 , \45767 , \45768 );
xor \U$37849 ( \45770 , \29849 , \45769 );
buf \U$37850 ( \45771 , \45770 );
buf \U$37852 ( \45772 , \45771 );
and \U$37853 ( \45773 , \28118 , \39334_nG9b7b );
and \U$37854 ( \45774 , \28115 , \39591_nG9b78 );
or \U$37855 ( \45775 , \45773 , \45774 );
xor \U$37856 ( \45776 , \28114 , \45775 );
buf \U$37857 ( \45777 , \45776 );
buf \U$37859 ( \45778 , \45777 );
xor \U$37860 ( \45779 , \45772 , \45778 );
and \U$37861 ( \45780 , \23201 , \41040_nG9b69 );
and \U$37862 ( \45781 , \23198 , \41381_nG9b66 );
or \U$37863 ( \45782 , \45780 , \45781 );
xor \U$37864 ( \45783 , \23197 , \45782 );
buf \U$37865 ( \45784 , \45783 );
buf \U$37867 ( \45785 , \45784 );
xor \U$37868 ( \45786 , \45779 , \45785 );
buf \U$37869 ( \45787 , \45786 );
xor \U$37870 ( \45788 , \45766 , \45787 );
and \U$37871 ( \45789 , \17297 , \43179_nG9b51 );
or \U$37873 ( \45790 , \45789 , 1'b0 );
xor \U$37874 ( \45791 , \17293 , \45790 );
buf \U$37875 ( \45792 , \45791 );
buf \U$37877 ( \45793 , \45792 );
and \U$37879 ( \45794 , \32916 , \37607_nG9b8a );
or \U$37880 ( \45795 , 1'b0 , \45794 );
xor \U$37881 ( \45796 , 1'b0 , \45795 );
buf \U$37882 ( \45797 , \45796 );
buf \U$37884 ( \45798 , \45797 );
xor \U$37885 ( \45799 , \45793 , \45798 );
and \U$37886 ( \45800 , \31636 , \37974_nG9b87 );
and \U$37887 ( \45801 , \31633 , \38337_nG9b84 );
or \U$37888 ( \45802 , \45800 , \45801 );
xor \U$37889 ( \45803 , \31632 , \45802 );
buf \U$37890 ( \45804 , \45803 );
buf \U$37892 ( \45805 , \45804 );
xor \U$37893 ( \45806 , \45799 , \45805 );
buf \U$37894 ( \45807 , \45806 );
xor \U$37895 ( \45808 , \45788 , \45807 );
buf \U$37896 ( \45809 , \45808 );
and \U$37897 ( \45810 , \45648 , \45669 );
and \U$37898 ( \45811 , \45648 , \45675 );
and \U$37899 ( \45812 , \45669 , \45675 );
or \U$37900 ( \45813 , \45810 , \45811 , \45812 );
buf \U$37901 ( \45814 , \45813 );
xor \U$37902 ( \45815 , \45809 , \45814 );
and \U$37903 ( \45816 , \45584 , \45605 );
and \U$37904 ( \45817 , \45584 , \45625 );
and \U$37905 ( \45818 , \45605 , \45625 );
or \U$37906 ( \45819 , \45816 , \45817 , \45818 );
buf \U$37907 ( \45820 , \45819 );
xor \U$37908 ( \45821 , \45815 , \45820 );
buf \U$37909 ( \45822 , \45821 );
and \U$37910 ( \45823 , \45633 , \45639 );
and \U$37911 ( \45824 , \45633 , \45646 );
and \U$37912 ( \45825 , \45639 , \45646 );
or \U$37913 ( \45826 , \45823 , \45824 , \45825 );
buf \U$37914 ( \45827 , \45826 );
and \U$37915 ( \45828 , \45612 , \45616 );
and \U$37916 ( \45829 , \45612 , \45623 );
and \U$37917 ( \45830 , \45616 , \45623 );
or \U$37918 ( \45831 , \45828 , \45829 , \45830 );
buf \U$37919 ( \45832 , \45831 );
xor \U$37920 ( \45833 , \45827 , \45832 );
and \U$37921 ( \45834 , \45590 , \45596 );
and \U$37922 ( \45835 , \45590 , \45603 );
and \U$37923 ( \45836 , \45596 , \45603 );
or \U$37924 ( \45837 , \45834 , \45835 , \45836 );
buf \U$37925 ( \45838 , \45837 );
xor \U$37926 ( \45839 , \45833 , \45838 );
buf \U$37927 ( \45840 , \45839 );
and \U$37928 ( \45841 , \45695 , \45700 );
and \U$37929 ( \45842 , \45695 , \45702 );
and \U$37930 ( \45843 , \45700 , \45702 );
or \U$37931 ( \45844 , \45841 , \45842 , \45843 );
buf \U$37932 ( \45845 , \45844 );
xor \U$37933 ( \45846 , \45840 , \45845 );
and \U$37934 ( \45847 , \45654 , \45660 );
and \U$37935 ( \45848 , \45654 , \45667 );
and \U$37936 ( \45849 , \45660 , \45667 );
or \U$37937 ( \45850 , \45847 , \45848 , \45849 );
buf \U$37938 ( \45851 , \45850 );
and \U$37939 ( \45852 , \21658 , \41685_nG9b63 );
and \U$37940 ( \45853 , \21655 , \41963_nG9b60 );
or \U$37941 ( \45854 , \45852 , \45853 );
xor \U$37942 ( \45855 , \21654 , \45854 );
buf \U$37943 ( \45856 , \45855 );
buf \U$37944 ( \45857 , \45856 );
not \U$37945 ( \45858 , \45857 );
xor \U$37946 ( \45859 , \45851 , \45858 );
and \U$37947 ( \45860 , \18702 , \42766_nG9b57 );
and \U$37948 ( \45861 , \18699 , \42848_nG9b54 );
or \U$37949 ( \45862 , \45860 , \45861 );
xor \U$37950 ( \45863 , \18698 , \45862 );
buf \U$37951 ( \45864 , \45863 );
buf \U$37953 ( \45865 , \45864 );
xor \U$37954 ( \45866 , \45859 , \45865 );
buf \U$37955 ( \45867 , \45866 );
xor \U$37956 ( \45868 , \45846 , \45867 );
buf \U$37957 ( \45869 , \45868 );
xor \U$37958 ( \45870 , \45822 , \45869 );
and \U$37959 ( \45871 , \45684 , \45689 );
and \U$37960 ( \45872 , \45684 , \45704 );
and \U$37961 ( \45873 , \45689 , \45704 );
or \U$37962 ( \45874 , \45871 , \45872 , \45873 );
buf \U$37963 ( \45875 , \45874 );
xor \U$37964 ( \45876 , \45870 , \45875 );
buf \U$37965 ( \45877 , \45876 );
xor \U$37966 ( \45878 , \45745 , \45877 );
and \U$37967 ( \45879 , \45579 , \45627 );
and \U$37968 ( \45880 , \45579 , \45677 );
and \U$37969 ( \45881 , \45627 , \45677 );
or \U$37970 ( \45882 , \45879 , \45880 , \45881 );
buf \U$37971 ( \45883 , \45882 );
xor \U$37972 ( \45884 , \45878 , \45883 );
and \U$37973 ( \45885 , \45740 , \45884 );
and \U$37975 ( \45886 , \45734 , \45739 );
or \U$37977 ( \45887 , 1'b0 , \45886 , 1'b0 );
xor \U$37978 ( \45888 , \45885 , \45887 );
and \U$37980 ( \45889 , \45727 , \45733 );
and \U$37981 ( \45890 , \45729 , \45733 );
or \U$37982 ( \45891 , 1'b0 , \45889 , \45890 );
xor \U$37983 ( \45892 , \45888 , \45891 );
xor \U$37990 ( \45893 , \45892 , 1'b0 );
and \U$37991 ( \45894 , \45745 , \45877 );
and \U$37992 ( \45895 , \45745 , \45883 );
and \U$37993 ( \45896 , \45877 , \45883 );
or \U$37994 ( \45897 , \45894 , \45895 , \45896 );
xor \U$37995 ( \45898 , \45893 , \45897 );
and \U$37996 ( \45899 , \45822 , \45869 );
and \U$37997 ( \45900 , \45822 , \45875 );
and \U$37998 ( \45901 , \45869 , \45875 );
or \U$37999 ( \45902 , \45899 , \45900 , \45901 );
buf \U$38000 ( \45903 , \45902 );
and \U$38001 ( \45904 , \18702 , \42848_nG9b54 );
and \U$38002 ( \45905 , \18699 , \43179_nG9b51 );
or \U$38003 ( \45906 , \45904 , \45905 );
xor \U$38004 ( \45907 , \18698 , \45906 );
buf \U$38005 ( \45908 , \45907 );
buf \U$38007 ( \45909 , \45908 );
xor \U$38011 ( \45910 , \17293 , 1'b0 );
not \U$38012 ( \45911 , \45910 );
buf \U$38013 ( \45912 , \45911 );
buf \U$38015 ( \45913 , \45912 );
xor \U$38016 ( \45914 , \45909 , \45913 );
and \U$38017 ( \45915 , \21658 , \41963_nG9b60 );
and \U$38018 ( \45916 , \21655 , \42201_nG9b5d );
or \U$38019 ( \45917 , \45915 , \45916 );
xor \U$38020 ( \45918 , \21654 , \45917 );
buf \U$38021 ( \45919 , \45918 );
buf \U$38023 ( \45920 , \45919 );
xor \U$38024 ( \45921 , \45914 , \45920 );
buf \U$38025 ( \45922 , \45921 );
and \U$38026 ( \45923 , \29853 , \38968_nG9b7e );
and \U$38027 ( \45924 , \29850 , \39334_nG9b7b );
or \U$38028 ( \45925 , \45923 , \45924 );
xor \U$38029 ( \45926 , \29849 , \45925 );
buf \U$38030 ( \45927 , \45926 );
buf \U$38032 ( \45928 , \45927 );
and \U$38033 ( \45929 , \28118 , \39591_nG9b78 );
and \U$38034 ( \45930 , \28115 , \39963_nG9b75 );
or \U$38035 ( \45931 , \45929 , \45930 );
xor \U$38036 ( \45932 , \28114 , \45931 );
buf \U$38037 ( \45933 , \45932 );
buf \U$38039 ( \45934 , \45933 );
xor \U$38040 ( \45935 , \45928 , \45934 );
and \U$38041 ( \45936 , \23201 , \41381_nG9b66 );
and \U$38042 ( \45937 , \23198 , \41685_nG9b63 );
or \U$38043 ( \45938 , \45936 , \45937 );
xor \U$38044 ( \45939 , \23197 , \45938 );
buf \U$38045 ( \45940 , \45939 );
buf \U$38047 ( \45941 , \45940 );
xor \U$38048 ( \45942 , \45935 , \45941 );
buf \U$38049 ( \45943 , \45942 );
xor \U$38050 ( \45944 , \45922 , \45943 );
and \U$38052 ( \45945 , \32916 , \37974_nG9b87 );
or \U$38053 ( \45946 , 1'b0 , \45945 );
xor \U$38054 ( \45947 , 1'b0 , \45946 );
buf \U$38055 ( \45948 , \45947 );
buf \U$38057 ( \45949 , \45948 );
and \U$38058 ( \45950 , \31636 , \38337_nG9b84 );
and \U$38059 ( \45951 , \31633 , \38663_nG9b81 );
or \U$38060 ( \45952 , \45950 , \45951 );
xor \U$38061 ( \45953 , \31632 , \45952 );
buf \U$38062 ( \45954 , \45953 );
buf \U$38064 ( \45955 , \45954 );
xor \U$38065 ( \45956 , \45949 , \45955 );
and \U$38066 ( \45957 , \24792 , \40843_nG9b6c );
and \U$38067 ( \45958 , \24789 , \41040_nG9b69 );
or \U$38068 ( \45959 , \45957 , \45958 );
xor \U$38069 ( \45960 , \24788 , \45959 );
buf \U$38070 ( \45961 , \45960 );
buf \U$38072 ( \45962 , \45961 );
xor \U$38073 ( \45963 , \45956 , \45962 );
buf \U$38074 ( \45964 , \45963 );
xor \U$38075 ( \45965 , \45944 , \45964 );
buf \U$38076 ( \45966 , \45965 );
and \U$38077 ( \45967 , \45751 , \45757 );
and \U$38078 ( \45968 , \45751 , \45764 );
and \U$38079 ( \45969 , \45757 , \45764 );
or \U$38080 ( \45970 , \45967 , \45968 , \45969 );
buf \U$38081 ( \45971 , \45970 );
and \U$38082 ( \45972 , \45793 , \45798 );
and \U$38083 ( \45973 , \45793 , \45805 );
and \U$38084 ( \45974 , \45798 , \45805 );
or \U$38085 ( \45975 , \45972 , \45973 , \45974 );
buf \U$38086 ( \45976 , \45975 );
xor \U$38087 ( \45977 , \45971 , \45976 );
and \U$38088 ( \45978 , \45772 , \45778 );
and \U$38089 ( \45979 , \45772 , \45785 );
and \U$38090 ( \45980 , \45778 , \45785 );
or \U$38091 ( \45981 , \45978 , \45979 , \45980 );
buf \U$38092 ( \45982 , \45981 );
xor \U$38093 ( \45983 , \45977 , \45982 );
buf \U$38094 ( \45984 , \45983 );
xor \U$38095 ( \45985 , \45966 , \45984 );
and \U$38096 ( \45986 , \45827 , \45832 );
and \U$38097 ( \45987 , \45827 , \45838 );
and \U$38098 ( \45988 , \45832 , \45838 );
or \U$38099 ( \45989 , \45986 , \45987 , \45988 );
buf \U$38100 ( \45990 , \45989 );
xor \U$38101 ( \45991 , \45985 , \45990 );
buf \U$38102 ( \45992 , \45991 );
and \U$38103 ( \45993 , \45840 , \45845 );
and \U$38104 ( \45994 , \45840 , \45867 );
and \U$38105 ( \45995 , \45845 , \45867 );
or \U$38106 ( \45996 , \45993 , \45994 , \45995 );
buf \U$38107 ( \45997 , \45996 );
xor \U$38108 ( \45998 , \45992 , \45997 );
and \U$38109 ( \45999 , \45766 , \45787 );
and \U$38110 ( \46000 , \45766 , \45807 );
and \U$38111 ( \46001 , \45787 , \45807 );
or \U$38112 ( \46002 , \45999 , \46000 , \46001 );
buf \U$38113 ( \46003 , \46002 );
and \U$38114 ( \46004 , \26431 , \40204_nG9b72 );
and \U$38115 ( \46005 , \26428 , \40452_nG9b6f );
or \U$38116 ( \46006 , \46004 , \46005 );
xor \U$38117 ( \46007 , \26427 , \46006 );
buf \U$38118 ( \46008 , \46007 );
buf \U$38120 ( \46009 , \46008 );
buf \U$38121 ( \46010 , \45857 );
xor \U$38122 ( \46011 , \46009 , \46010 );
and \U$38123 ( \46012 , \20155 , \42433_nG9b5a );
and \U$38124 ( \46013 , \20152 , \42766_nG9b57 );
or \U$38125 ( \46014 , \46012 , \46013 );
xor \U$38126 ( \46015 , \20151 , \46014 );
buf \U$38127 ( \46016 , \46015 );
buf \U$38129 ( \46017 , \46016 );
xor \U$38130 ( \46018 , \46011 , \46017 );
buf \U$38131 ( \46019 , \46018 );
xor \U$38132 ( \46020 , \46003 , \46019 );
and \U$38133 ( \46021 , \45851 , \45858 );
and \U$38134 ( \46022 , \45851 , \45865 );
and \U$38135 ( \46023 , \45858 , \45865 );
or \U$38136 ( \46024 , \46021 , \46022 , \46023 );
buf \U$38137 ( \46025 , \46024 );
xor \U$38138 ( \46026 , \46020 , \46025 );
buf \U$38139 ( \46027 , \46026 );
xor \U$38140 ( \46028 , \45998 , \46027 );
buf \U$38141 ( \46029 , \46028 );
xor \U$38142 ( \46030 , \45903 , \46029 );
and \U$38143 ( \46031 , \45809 , \45814 );
and \U$38144 ( \46032 , \45809 , \45820 );
and \U$38145 ( \46033 , \45814 , \45820 );
or \U$38146 ( \46034 , \46031 , \46032 , \46033 );
buf \U$38147 ( \46035 , \46034 );
xor \U$38148 ( \46036 , \46030 , \46035 );
and \U$38149 ( \46037 , \45898 , \46036 );
and \U$38151 ( \46038 , \45892 , \45897 );
or \U$38153 ( \46039 , 1'b0 , \46038 , 1'b0 );
xor \U$38154 ( \46040 , \46037 , \46039 );
and \U$38156 ( \46041 , \45885 , \45891 );
and \U$38157 ( \46042 , \45887 , \45891 );
or \U$38158 ( \46043 , 1'b0 , \46041 , \46042 );
xor \U$38159 ( \46044 , \46040 , \46043 );
xor \U$38166 ( \46045 , \46044 , 1'b0 );
and \U$38167 ( \46046 , \45992 , \45997 );
and \U$38168 ( \46047 , \45992 , \46027 );
and \U$38169 ( \46048 , \45997 , \46027 );
or \U$38170 ( \46049 , \46046 , \46047 , \46048 );
buf \U$38171 ( \46050 , \46049 );
and \U$38172 ( \46051 , \45971 , \45976 );
and \U$38173 ( \46052 , \45971 , \45982 );
and \U$38174 ( \46053 , \45976 , \45982 );
or \U$38175 ( \46054 , \46051 , \46052 , \46053 );
buf \U$38176 ( \46055 , \46054 );
and \U$38177 ( \46056 , \46009 , \46010 );
and \U$38178 ( \46057 , \46009 , \46017 );
and \U$38179 ( \46058 , \46010 , \46017 );
or \U$38180 ( \46059 , \46056 , \46057 , \46058 );
buf \U$38181 ( \46060 , \46059 );
xor \U$38182 ( \46061 , \46055 , \46060 );
and \U$38183 ( \46062 , \28118 , \39963_nG9b75 );
and \U$38184 ( \46063 , \28115 , \40204_nG9b72 );
or \U$38185 ( \46064 , \46062 , \46063 );
xor \U$38186 ( \46065 , \28114 , \46064 );
buf \U$38187 ( \46066 , \46065 );
buf \U$38189 ( \46067 , \46066 );
and \U$38190 ( \46068 , \26431 , \40452_nG9b6f );
and \U$38191 ( \46069 , \26428 , \40843_nG9b6c );
or \U$38192 ( \46070 , \46068 , \46069 );
xor \U$38193 ( \46071 , \26427 , \46070 );
buf \U$38194 ( \46072 , \46071 );
buf \U$38196 ( \46073 , \46072 );
xor \U$38197 ( \46074 , \46067 , \46073 );
and \U$38198 ( \46075 , \20155 , \42766_nG9b57 );
and \U$38199 ( \46076 , \20152 , \42848_nG9b54 );
or \U$38200 ( \46077 , \46075 , \46076 );
xor \U$38201 ( \46078 , \20151 , \46077 );
buf \U$38202 ( \46079 , \46078 );
buf \U$38204 ( \46080 , \46079 );
xor \U$38205 ( \46081 , \46074 , \46080 );
buf \U$38206 ( \46082 , \46081 );
xor \U$38207 ( \46083 , \46061 , \46082 );
buf \U$38208 ( \46084 , \46083 );
and \U$38209 ( \46085 , \46003 , \46019 );
and \U$38210 ( \46086 , \46003 , \46025 );
and \U$38211 ( \46087 , \46019 , \46025 );
or \U$38212 ( \46088 , \46085 , \46086 , \46087 );
buf \U$38213 ( \46089 , \46088 );
xor \U$38214 ( \46090 , \46084 , \46089 );
and \U$38215 ( \46091 , \45966 , \45984 );
and \U$38216 ( \46092 , \45966 , \45990 );
and \U$38217 ( \46093 , \45984 , \45990 );
or \U$38218 ( \46094 , \46091 , \46092 , \46093 );
buf \U$38219 ( \46095 , \46094 );
xor \U$38220 ( \46096 , \46090 , \46095 );
buf \U$38221 ( \46097 , \46096 );
xor \U$38222 ( \46098 , \46050 , \46097 );
and \U$38223 ( \46099 , \31636 , \38663_nG9b81 );
and \U$38224 ( \46100 , \31633 , \38968_nG9b7e );
or \U$38225 ( \46101 , \46099 , \46100 );
xor \U$38226 ( \46102 , \31632 , \46101 );
buf \U$38227 ( \46103 , \46102 );
buf \U$38229 ( \46104 , \46103 );
and \U$38230 ( \46105 , \29853 , \39334_nG9b7b );
and \U$38231 ( \46106 , \29850 , \39591_nG9b78 );
or \U$38232 ( \46107 , \46105 , \46106 );
xor \U$38233 ( \46108 , \29849 , \46107 );
buf \U$38234 ( \46109 , \46108 );
buf \U$38236 ( \46110 , \46109 );
xor \U$38237 ( \46111 , \46104 , \46110 );
and \U$38238 ( \46112 , \23201 , \41685_nG9b63 );
and \U$38239 ( \46113 , \23198 , \41963_nG9b60 );
or \U$38240 ( \46114 , \46112 , \46113 );
xor \U$38241 ( \46115 , \23197 , \46114 );
buf \U$38242 ( \46116 , \46115 );
buf \U$38244 ( \46117 , \46116 );
xor \U$38245 ( \46118 , \46111 , \46117 );
buf \U$38246 ( \46119 , \46118 );
and \U$38248 ( \46120 , \32916 , \38337_nG9b84 );
or \U$38249 ( \46121 , 1'b0 , \46120 );
xor \U$38250 ( \46122 , 1'b0 , \46121 );
buf \U$38251 ( \46123 , \46122 );
buf \U$38253 ( \46124 , \46123 );
and \U$38254 ( \46125 , \24792 , \41040_nG9b69 );
and \U$38255 ( \46126 , \24789 , \41381_nG9b66 );
or \U$38256 ( \46127 , \46125 , \46126 );
xor \U$38257 ( \46128 , \24788 , \46127 );
buf \U$38258 ( \46129 , \46128 );
buf \U$38260 ( \46130 , \46129 );
xor \U$38261 ( \46131 , \46124 , \46130 );
and \U$38262 ( \46132 , \21658 , \42201_nG9b5d );
and \U$38263 ( \46133 , \21655 , \42433_nG9b5a );
or \U$38264 ( \46134 , \46132 , \46133 );
xor \U$38265 ( \46135 , \21654 , \46134 );
buf \U$38266 ( \46136 , \46135 );
buf \U$38268 ( \46137 , \46136 );
xor \U$38269 ( \46138 , \46131 , \46137 );
buf \U$38270 ( \46139 , \46138 );
xor \U$38271 ( \46140 , \46119 , \46139 );
and \U$38272 ( \46141 , \45949 , \45955 );
and \U$38273 ( \46142 , \45949 , \45962 );
and \U$38274 ( \46143 , \45955 , \45962 );
or \U$38275 ( \46144 , \46141 , \46142 , \46143 );
buf \U$38276 ( \46145 , \46144 );
xor \U$38277 ( \46146 , \46140 , \46145 );
buf \U$38278 ( \46147 , \46146 );
and \U$38279 ( \46148 , \45922 , \45943 );
and \U$38280 ( \46149 , \45922 , \45964 );
and \U$38281 ( \46150 , \45943 , \45964 );
or \U$38282 ( \46151 , \46148 , \46149 , \46150 );
buf \U$38283 ( \46152 , \46151 );
xor \U$38284 ( \46153 , \46147 , \46152 );
and \U$38285 ( \46154 , \45909 , \45913 );
and \U$38286 ( \46155 , \45909 , \45920 );
and \U$38287 ( \46156 , \45913 , \45920 );
or \U$38288 ( \46157 , \46154 , \46155 , \46156 );
buf \U$38289 ( \46158 , \46157 );
and \U$38290 ( \46159 , \45928 , \45934 );
and \U$38291 ( \46160 , \45928 , \45941 );
and \U$38292 ( \46161 , \45934 , \45941 );
or \U$38293 ( \46162 , \46159 , \46160 , \46161 );
buf \U$38294 ( \46163 , \46162 );
xor \U$38295 ( \46164 , \46158 , \46163 );
and \U$38296 ( \46165 , \18702 , \43179_nG9b51 );
or \U$38298 ( \46166 , \46165 , 1'b0 );
xor \U$38299 ( \46167 , \18698 , \46166 );
buf \U$38300 ( \46168 , \46167 );
buf \U$38301 ( \46169 , \46168 );
not \U$38302 ( \46170 , \46169 );
xor \U$38303 ( \46171 , \46164 , \46170 );
buf \U$38304 ( \46172 , \46171 );
xor \U$38305 ( \46173 , \46153 , \46172 );
buf \U$38306 ( \46174 , \46173 );
xor \U$38307 ( \46175 , \46098 , \46174 );
xor \U$38308 ( \46176 , \46045 , \46175 );
and \U$38309 ( \46177 , \45903 , \46029 );
and \U$38310 ( \46178 , \45903 , \46035 );
and \U$38311 ( \46179 , \46029 , \46035 );
or \U$38312 ( \46180 , \46177 , \46178 , \46179 );
and \U$38313 ( \46181 , \46176 , \46180 );
and \U$38315 ( \46182 , \46044 , \46175 );
or \U$38317 ( \46183 , 1'b0 , \46182 , 1'b0 );
xor \U$38318 ( \46184 , \46181 , \46183 );
and \U$38320 ( \46185 , \46037 , \46043 );
and \U$38321 ( \46186 , \46039 , \46043 );
or \U$38322 ( \46187 , 1'b0 , \46185 , \46186 );
xor \U$38323 ( \46188 , \46184 , \46187 );
xor \U$38330 ( \46189 , \46188 , 1'b0 );
and \U$38331 ( \46190 , \46084 , \46089 );
and \U$38332 ( \46191 , \46084 , \46095 );
and \U$38333 ( \46192 , \46089 , \46095 );
or \U$38334 ( \46193 , \46190 , \46191 , \46192 );
buf \U$38335 ( \46194 , \46193 );
and \U$38336 ( \46195 , \20155 , \42848_nG9b54 );
and \U$38337 ( \46196 , \20152 , \43179_nG9b51 );
or \U$38338 ( \46197 , \46195 , \46196 );
xor \U$38339 ( \46198 , \20151 , \46197 );
buf \U$38340 ( \46199 , \46198 );
buf \U$38342 ( \46200 , \46199 );
xor \U$38346 ( \46201 , \18698 , 1'b0 );
not \U$38347 ( \46202 , \46201 );
buf \U$38348 ( \46203 , \46202 );
buf \U$38350 ( \46204 , \46203 );
xor \U$38351 ( \46205 , \46200 , \46204 );
and \U$38352 ( \46206 , \23201 , \41963_nG9b60 );
and \U$38353 ( \46207 , \23198 , \42201_nG9b5d );
or \U$38354 ( \46208 , \46206 , \46207 );
xor \U$38355 ( \46209 , \23197 , \46208 );
buf \U$38356 ( \46210 , \46209 );
buf \U$38358 ( \46211 , \46210 );
xor \U$38359 ( \46212 , \46205 , \46211 );
buf \U$38360 ( \46213 , \46212 );
and \U$38362 ( \46214 , \32916 , \38663_nG9b81 );
or \U$38363 ( \46215 , 1'b0 , \46214 );
xor \U$38364 ( \46216 , 1'b0 , \46215 );
buf \U$38365 ( \46217 , \46216 );
buf \U$38367 ( \46218 , \46217 );
and \U$38368 ( \46219 , \28118 , \40204_nG9b72 );
and \U$38369 ( \46220 , \28115 , \40452_nG9b6f );
or \U$38370 ( \46221 , \46219 , \46220 );
xor \U$38371 ( \46222 , \28114 , \46221 );
buf \U$38372 ( \46223 , \46222 );
buf \U$38374 ( \46224 , \46223 );
xor \U$38375 ( \46225 , \46218 , \46224 );
and \U$38376 ( \46226 , \26431 , \40843_nG9b6c );
and \U$38377 ( \46227 , \26428 , \41040_nG9b69 );
or \U$38378 ( \46228 , \46226 , \46227 );
xor \U$38379 ( \46229 , \26427 , \46228 );
buf \U$38380 ( \46230 , \46229 );
buf \U$38382 ( \46231 , \46230 );
xor \U$38383 ( \46232 , \46225 , \46231 );
buf \U$38384 ( \46233 , \46232 );
xor \U$38385 ( \46234 , \46213 , \46233 );
and \U$38386 ( \46235 , \46124 , \46130 );
and \U$38387 ( \46236 , \46124 , \46137 );
and \U$38388 ( \46237 , \46130 , \46137 );
or \U$38389 ( \46238 , \46235 , \46236 , \46237 );
buf \U$38390 ( \46239 , \46238 );
xor \U$38391 ( \46240 , \46234 , \46239 );
buf \U$38392 ( \46241 , \46240 );
and \U$38393 ( \46242 , \46158 , \46163 );
and \U$38394 ( \46243 , \46158 , \46170 );
and \U$38395 ( \46244 , \46163 , \46170 );
or \U$38396 ( \46245 , \46242 , \46243 , \46244 );
buf \U$38397 ( \46246 , \46245 );
xor \U$38398 ( \46247 , \46241 , \46246 );
and \U$38399 ( \46248 , \46119 , \46139 );
and \U$38400 ( \46249 , \46119 , \46145 );
and \U$38401 ( \46250 , \46139 , \46145 );
or \U$38402 ( \46251 , \46248 , \46249 , \46250 );
buf \U$38403 ( \46252 , \46251 );
xor \U$38404 ( \46253 , \46247 , \46252 );
buf \U$38405 ( \46254 , \46253 );
xor \U$38406 ( \46255 , \46194 , \46254 );
and \U$38407 ( \46256 , \46055 , \46060 );
and \U$38408 ( \46257 , \46055 , \46082 );
and \U$38409 ( \46258 , \46060 , \46082 );
or \U$38410 ( \46259 , \46256 , \46257 , \46258 );
buf \U$38411 ( \46260 , \46259 );
and \U$38412 ( \46261 , \46104 , \46110 );
and \U$38413 ( \46262 , \46104 , \46117 );
and \U$38414 ( \46263 , \46110 , \46117 );
or \U$38415 ( \46264 , \46261 , \46262 , \46263 );
buf \U$38416 ( \46265 , \46264 );
buf \U$38417 ( \46266 , \46169 );
xor \U$38418 ( \46267 , \46265 , \46266 );
and \U$38419 ( \46268 , \21658 , \42433_nG9b5a );
and \U$38420 ( \46269 , \21655 , \42766_nG9b57 );
or \U$38421 ( \46270 , \46268 , \46269 );
xor \U$38422 ( \46271 , \21654 , \46270 );
buf \U$38423 ( \46272 , \46271 );
buf \U$38425 ( \46273 , \46272 );
xor \U$38426 ( \46274 , \46267 , \46273 );
buf \U$38427 ( \46275 , \46274 );
and \U$38428 ( \46276 , \31636 , \38968_nG9b7e );
and \U$38429 ( \46277 , \31633 , \39334_nG9b7b );
or \U$38430 ( \46278 , \46276 , \46277 );
xor \U$38431 ( \46279 , \31632 , \46278 );
buf \U$38432 ( \46280 , \46279 );
buf \U$38434 ( \46281 , \46280 );
and \U$38435 ( \46282 , \29853 , \39591_nG9b78 );
and \U$38436 ( \46283 , \29850 , \39963_nG9b75 );
or \U$38437 ( \46284 , \46282 , \46283 );
xor \U$38438 ( \46285 , \29849 , \46284 );
buf \U$38439 ( \46286 , \46285 );
buf \U$38441 ( \46287 , \46286 );
xor \U$38442 ( \46288 , \46281 , \46287 );
and \U$38443 ( \46289 , \24792 , \41381_nG9b66 );
and \U$38444 ( \46290 , \24789 , \41685_nG9b63 );
or \U$38445 ( \46291 , \46289 , \46290 );
xor \U$38446 ( \46292 , \24788 , \46291 );
buf \U$38447 ( \46293 , \46292 );
buf \U$38449 ( \46294 , \46293 );
xor \U$38450 ( \46295 , \46288 , \46294 );
buf \U$38451 ( \46296 , \46295 );
xor \U$38452 ( \46297 , \46275 , \46296 );
and \U$38453 ( \46298 , \46067 , \46073 );
and \U$38454 ( \46299 , \46067 , \46080 );
and \U$38455 ( \46300 , \46073 , \46080 );
or \U$38456 ( \46301 , \46298 , \46299 , \46300 );
buf \U$38457 ( \46302 , \46301 );
xor \U$38458 ( \46303 , \46297 , \46302 );
buf \U$38459 ( \46304 , \46303 );
xor \U$38460 ( \46305 , \46260 , \46304 );
and \U$38461 ( \46306 , \46147 , \46152 );
and \U$38462 ( \46307 , \46147 , \46172 );
and \U$38463 ( \46308 , \46152 , \46172 );
or \U$38464 ( \46309 , \46306 , \46307 , \46308 );
buf \U$38465 ( \46310 , \46309 );
xor \U$38466 ( \46311 , \46305 , \46310 );
buf \U$38467 ( \46312 , \46311 );
xor \U$38468 ( \46313 , \46255 , \46312 );
xor \U$38469 ( \46314 , \46189 , \46313 );
and \U$38470 ( \46315 , \46050 , \46097 );
and \U$38471 ( \46316 , \46050 , \46174 );
and \U$38472 ( \46317 , \46097 , \46174 );
or \U$38473 ( \46318 , \46315 , \46316 , \46317 );
and \U$38474 ( \46319 , \46314 , \46318 );
and \U$38476 ( \46320 , \46188 , \46313 );
or \U$38478 ( \46321 , 1'b0 , \46320 , 1'b0 );
xor \U$38479 ( \46322 , \46319 , \46321 );
and \U$38481 ( \46323 , \46181 , \46187 );
and \U$38482 ( \46324 , \46183 , \46187 );
or \U$38483 ( \46325 , 1'b0 , \46323 , \46324 );
xor \U$38484 ( \46326 , \46322 , \46325 );
xor \U$38491 ( \46327 , \46326 , 1'b0 );
and \U$38492 ( \46328 , \46194 , \46254 );
and \U$38493 ( \46329 , \46194 , \46312 );
and \U$38494 ( \46330 , \46254 , \46312 );
or \U$38495 ( \46331 , \46328 , \46329 , \46330 );
xor \U$38496 ( \46332 , \46327 , \46331 );
and \U$38497 ( \46333 , \28118 , \40452_nG9b6f );
and \U$38498 ( \46334 , \28115 , \40843_nG9b6c );
or \U$38499 ( \46335 , \46333 , \46334 );
xor \U$38500 ( \46336 , \28114 , \46335 );
buf \U$38501 ( \46337 , \46336 );
buf \U$38503 ( \46338 , \46337 );
and \U$38504 ( \46339 , \26431 , \41040_nG9b69 );
and \U$38505 ( \46340 , \26428 , \41381_nG9b66 );
or \U$38506 ( \46341 , \46339 , \46340 );
xor \U$38507 ( \46342 , \26427 , \46341 );
buf \U$38508 ( \46343 , \46342 );
buf \U$38510 ( \46344 , \46343 );
xor \U$38511 ( \46345 , \46338 , \46344 );
and \U$38512 ( \46346 , \23201 , \42201_nG9b5d );
and \U$38513 ( \46347 , \23198 , \42433_nG9b5a );
or \U$38514 ( \46348 , \46346 , \46347 );
xor \U$38515 ( \46349 , \23197 , \46348 );
buf \U$38516 ( \46350 , \46349 );
buf \U$38518 ( \46351 , \46350 );
xor \U$38519 ( \46352 , \46345 , \46351 );
buf \U$38520 ( \46353 , \46352 );
and \U$38521 ( \46354 , \20155 , \43179_nG9b51 );
or \U$38523 ( \46355 , \46354 , 1'b0 );
xor \U$38524 ( \46356 , \20151 , \46355 );
buf \U$38525 ( \46357 , \46356 );
buf \U$38526 ( \46358 , \46357 );
not \U$38527 ( \46359 , \46358 );
and \U$38528 ( \46360 , \29853 , \39963_nG9b75 );
and \U$38529 ( \46361 , \29850 , \40204_nG9b72 );
or \U$38530 ( \46362 , \46360 , \46361 );
xor \U$38531 ( \46363 , \29849 , \46362 );
buf \U$38532 ( \46364 , \46363 );
buf \U$38534 ( \46365 , \46364 );
xor \U$38535 ( \46366 , \46359 , \46365 );
and \U$38536 ( \46367 , \21658 , \42766_nG9b57 );
and \U$38537 ( \46368 , \21655 , \42848_nG9b54 );
or \U$38538 ( \46369 , \46367 , \46368 );
xor \U$38539 ( \46370 , \21654 , \46369 );
buf \U$38540 ( \46371 , \46370 );
buf \U$38542 ( \46372 , \46371 );
xor \U$38543 ( \46373 , \46366 , \46372 );
buf \U$38544 ( \46374 , \46373 );
xor \U$38545 ( \46375 , \46353 , \46374 );
and \U$38547 ( \46376 , \32916 , \38968_nG9b7e );
or \U$38548 ( \46377 , 1'b0 , \46376 );
xor \U$38549 ( \46378 , 1'b0 , \46377 );
buf \U$38550 ( \46379 , \46378 );
buf \U$38552 ( \46380 , \46379 );
and \U$38553 ( \46381 , \31636 , \39334_nG9b7b );
and \U$38554 ( \46382 , \31633 , \39591_nG9b78 );
or \U$38555 ( \46383 , \46381 , \46382 );
xor \U$38556 ( \46384 , \31632 , \46383 );
buf \U$38557 ( \46385 , \46384 );
buf \U$38559 ( \46386 , \46385 );
xor \U$38560 ( \46387 , \46380 , \46386 );
and \U$38561 ( \46388 , \24792 , \41685_nG9b63 );
and \U$38562 ( \46389 , \24789 , \41963_nG9b60 );
or \U$38563 ( \46390 , \46388 , \46389 );
xor \U$38564 ( \46391 , \24788 , \46390 );
buf \U$38565 ( \46392 , \46391 );
buf \U$38567 ( \46393 , \46392 );
xor \U$38568 ( \46394 , \46387 , \46393 );
buf \U$38569 ( \46395 , \46394 );
xor \U$38570 ( \46396 , \46375 , \46395 );
buf \U$38571 ( \46397 , \46396 );
and \U$38572 ( \46398 , \46275 , \46296 );
and \U$38573 ( \46399 , \46275 , \46302 );
and \U$38574 ( \46400 , \46296 , \46302 );
or \U$38575 ( \46401 , \46398 , \46399 , \46400 );
buf \U$38576 ( \46402 , \46401 );
xor \U$38577 ( \46403 , \46397 , \46402 );
and \U$38578 ( \46404 , \46213 , \46233 );
and \U$38579 ( \46405 , \46213 , \46239 );
and \U$38580 ( \46406 , \46233 , \46239 );
or \U$38581 ( \46407 , \46404 , \46405 , \46406 );
buf \U$38582 ( \46408 , \46407 );
and \U$38583 ( \46409 , \46200 , \46204 );
and \U$38584 ( \46410 , \46200 , \46211 );
and \U$38585 ( \46411 , \46204 , \46211 );
or \U$38586 ( \46412 , \46409 , \46410 , \46411 );
buf \U$38587 ( \46413 , \46412 );
and \U$38588 ( \46414 , \46218 , \46224 );
and \U$38589 ( \46415 , \46218 , \46231 );
and \U$38590 ( \46416 , \46224 , \46231 );
or \U$38591 ( \46417 , \46414 , \46415 , \46416 );
buf \U$38592 ( \46418 , \46417 );
xor \U$38593 ( \46419 , \46413 , \46418 );
and \U$38594 ( \46420 , \46281 , \46287 );
and \U$38595 ( \46421 , \46281 , \46294 );
and \U$38596 ( \46422 , \46287 , \46294 );
or \U$38597 ( \46423 , \46420 , \46421 , \46422 );
buf \U$38598 ( \46424 , \46423 );
xor \U$38599 ( \46425 , \46419 , \46424 );
buf \U$38600 ( \46426 , \46425 );
xor \U$38601 ( \46427 , \46408 , \46426 );
and \U$38602 ( \46428 , \46265 , \46266 );
and \U$38603 ( \46429 , \46265 , \46273 );
and \U$38604 ( \46430 , \46266 , \46273 );
or \U$38605 ( \46431 , \46428 , \46429 , \46430 );
buf \U$38606 ( \46432 , \46431 );
xor \U$38607 ( \46433 , \46427 , \46432 );
buf \U$38608 ( \46434 , \46433 );
xor \U$38609 ( \46435 , \46403 , \46434 );
buf \U$38610 ( \46436 , \46435 );
and \U$38611 ( \46437 , \46260 , \46304 );
and \U$38612 ( \46438 , \46260 , \46310 );
and \U$38613 ( \46439 , \46304 , \46310 );
or \U$38614 ( \46440 , \46437 , \46438 , \46439 );
buf \U$38615 ( \46441 , \46440 );
xor \U$38616 ( \46442 , \46436 , \46441 );
and \U$38617 ( \46443 , \46241 , \46246 );
and \U$38618 ( \46444 , \46241 , \46252 );
and \U$38619 ( \46445 , \46246 , \46252 );
or \U$38620 ( \46446 , \46443 , \46444 , \46445 );
buf \U$38621 ( \46447 , \46446 );
xor \U$38622 ( \46448 , \46442 , \46447 );
and \U$38623 ( \46449 , \46332 , \46448 );
and \U$38625 ( \46450 , \46326 , \46331 );
or \U$38627 ( \46451 , 1'b0 , \46450 , 1'b0 );
xor \U$38628 ( \46452 , \46449 , \46451 );
and \U$38630 ( \46453 , \46319 , \46325 );
and \U$38631 ( \46454 , \46321 , \46325 );
or \U$38632 ( \46455 , 1'b0 , \46453 , \46454 );
xor \U$38633 ( \46456 , \46452 , \46455 );
xor \U$38640 ( \46457 , \46456 , 1'b0 );
and \U$38641 ( \46458 , \46436 , \46441 );
and \U$38642 ( \46459 , \46436 , \46447 );
and \U$38643 ( \46460 , \46441 , \46447 );
or \U$38644 ( \46461 , \46458 , \46459 , \46460 );
xor \U$38645 ( \46462 , \46457 , \46461 );
and \U$38646 ( \46463 , \46397 , \46402 );
and \U$38647 ( \46464 , \46397 , \46434 );
and \U$38648 ( \46465 , \46402 , \46434 );
or \U$38649 ( \46466 , \46463 , \46464 , \46465 );
buf \U$38650 ( \46467 , \46466 );
and \U$38651 ( \46468 , \29853 , \40204_nG9b72 );
and \U$38652 ( \46469 , \29850 , \40452_nG9b6f );
or \U$38653 ( \46470 , \46468 , \46469 );
xor \U$38654 ( \46471 , \29849 , \46470 );
buf \U$38655 ( \46472 , \46471 );
buf \U$38657 ( \46473 , \46472 );
and \U$38658 ( \46474 , \28118 , \40843_nG9b6c );
and \U$38659 ( \46475 , \28115 , \41040_nG9b69 );
or \U$38660 ( \46476 , \46474 , \46475 );
xor \U$38661 ( \46477 , \28114 , \46476 );
buf \U$38662 ( \46478 , \46477 );
buf \U$38664 ( \46479 , \46478 );
xor \U$38665 ( \46480 , \46473 , \46479 );
and \U$38666 ( \46481 , \23201 , \42433_nG9b5a );
and \U$38667 ( \46482 , \23198 , \42766_nG9b57 );
or \U$38668 ( \46483 , \46481 , \46482 );
xor \U$38669 ( \46484 , \23197 , \46483 );
buf \U$38670 ( \46485 , \46484 );
buf \U$38672 ( \46486 , \46485 );
xor \U$38673 ( \46487 , \46480 , \46486 );
buf \U$38674 ( \46488 , \46487 );
and \U$38676 ( \46489 , \32916 , \39334_nG9b7b );
or \U$38677 ( \46490 , 1'b0 , \46489 );
xor \U$38678 ( \46491 , 1'b0 , \46490 );
buf \U$38679 ( \46492 , \46491 );
buf \U$38681 ( \46493 , \46492 );
and \U$38682 ( \46494 , \31636 , \39591_nG9b78 );
and \U$38683 ( \46495 , \31633 , \39963_nG9b75 );
or \U$38684 ( \46496 , \46494 , \46495 );
xor \U$38685 ( \46497 , \31632 , \46496 );
buf \U$38686 ( \46498 , \46497 );
buf \U$38688 ( \46499 , \46498 );
xor \U$38689 ( \46500 , \46493 , \46499 );
and \U$38690 ( \46501 , \26431 , \41381_nG9b66 );
and \U$38691 ( \46502 , \26428 , \41685_nG9b63 );
or \U$38692 ( \46503 , \46501 , \46502 );
xor \U$38693 ( \46504 , \26427 , \46503 );
buf \U$38694 ( \46505 , \46504 );
buf \U$38696 ( \46506 , \46505 );
xor \U$38697 ( \46507 , \46500 , \46506 );
buf \U$38698 ( \46508 , \46507 );
xor \U$38699 ( \46509 , \46488 , \46508 );
and \U$38700 ( \46510 , \21658 , \42848_nG9b54 );
and \U$38701 ( \46511 , \21655 , \43179_nG9b51 );
or \U$38702 ( \46512 , \46510 , \46511 );
xor \U$38703 ( \46513 , \21654 , \46512 );
buf \U$38704 ( \46514 , \46513 );
buf \U$38706 ( \46515 , \46514 );
xor \U$38710 ( \46516 , \20151 , 1'b0 );
not \U$38711 ( \46517 , \46516 );
buf \U$38712 ( \46518 , \46517 );
buf \U$38714 ( \46519 , \46518 );
xor \U$38715 ( \46520 , \46515 , \46519 );
and \U$38716 ( \46521 , \24792 , \41963_nG9b60 );
and \U$38717 ( \46522 , \24789 , \42201_nG9b5d );
or \U$38718 ( \46523 , \46521 , \46522 );
xor \U$38719 ( \46524 , \24788 , \46523 );
buf \U$38720 ( \46525 , \46524 );
buf \U$38722 ( \46526 , \46525 );
xor \U$38723 ( \46527 , \46520 , \46526 );
buf \U$38724 ( \46528 , \46527 );
xor \U$38725 ( \46529 , \46509 , \46528 );
buf \U$38726 ( \46530 , \46529 );
and \U$38727 ( \46531 , \46353 , \46374 );
and \U$38728 ( \46532 , \46353 , \46395 );
and \U$38729 ( \46533 , \46374 , \46395 );
or \U$38730 ( \46534 , \46531 , \46532 , \46533 );
buf \U$38731 ( \46535 , \46534 );
xor \U$38732 ( \46536 , \46530 , \46535 );
and \U$38733 ( \46537 , \46408 , \46426 );
and \U$38734 ( \46538 , \46408 , \46432 );
and \U$38735 ( \46539 , \46426 , \46432 );
or \U$38736 ( \46540 , \46537 , \46538 , \46539 );
buf \U$38737 ( \46541 , \46540 );
xor \U$38738 ( \46542 , \46536 , \46541 );
buf \U$38739 ( \46543 , \46542 );
xor \U$38740 ( \46544 , \46467 , \46543 );
and \U$38741 ( \46545 , \46413 , \46418 );
and \U$38742 ( \46546 , \46413 , \46424 );
and \U$38743 ( \46547 , \46418 , \46424 );
or \U$38744 ( \46548 , \46545 , \46546 , \46547 );
buf \U$38745 ( \46549 , \46548 );
and \U$38746 ( \46550 , \46380 , \46386 );
and \U$38747 ( \46551 , \46380 , \46393 );
and \U$38748 ( \46552 , \46386 , \46393 );
or \U$38749 ( \46553 , \46550 , \46551 , \46552 );
buf \U$38750 ( \46554 , \46553 );
and \U$38751 ( \46555 , \46338 , \46344 );
and \U$38752 ( \46556 , \46338 , \46351 );
and \U$38753 ( \46557 , \46344 , \46351 );
or \U$38754 ( \46558 , \46555 , \46556 , \46557 );
buf \U$38755 ( \46559 , \46558 );
xor \U$38756 ( \46560 , \46554 , \46559 );
buf \U$38757 ( \46561 , \46358 );
xor \U$38758 ( \46562 , \46560 , \46561 );
buf \U$38759 ( \46563 , \46562 );
xor \U$38760 ( \46564 , \46549 , \46563 );
and \U$38761 ( \46565 , \46359 , \46365 );
and \U$38762 ( \46566 , \46359 , \46372 );
and \U$38763 ( \46567 , \46365 , \46372 );
or \U$38764 ( \46568 , \46565 , \46566 , \46567 );
buf \U$38765 ( \46569 , \46568 );
xor \U$38766 ( \46570 , \46564 , \46569 );
buf \U$38767 ( \46571 , \46570 );
xor \U$38768 ( \46572 , \46544 , \46571 );
and \U$38769 ( \46573 , \46462 , \46572 );
and \U$38771 ( \46574 , \46456 , \46461 );
or \U$38773 ( \46575 , 1'b0 , \46574 , 1'b0 );
xor \U$38774 ( \46576 , \46573 , \46575 );
and \U$38776 ( \46577 , \46449 , \46455 );
and \U$38777 ( \46578 , \46451 , \46455 );
or \U$38778 ( \46579 , 1'b0 , \46577 , \46578 );
xor \U$38779 ( \46580 , \46576 , \46579 );
xor \U$38786 ( \46581 , \46580 , 1'b0 );
and \U$38787 ( \46582 , \46467 , \46543 );
and \U$38788 ( \46583 , \46467 , \46571 );
and \U$38789 ( \46584 , \46543 , \46571 );
or \U$38790 ( \46585 , \46582 , \46583 , \46584 );
xor \U$38791 ( \46586 , \46581 , \46585 );
and \U$38792 ( \46587 , \46530 , \46535 );
and \U$38793 ( \46588 , \46530 , \46541 );
and \U$38794 ( \46589 , \46535 , \46541 );
or \U$38795 ( \46590 , \46587 , \46588 , \46589 );
buf \U$38796 ( \46591 , \46590 );
and \U$38797 ( \46592 , \46488 , \46508 );
and \U$38798 ( \46593 , \46488 , \46528 );
and \U$38799 ( \46594 , \46508 , \46528 );
or \U$38800 ( \46595 , \46592 , \46593 , \46594 );
buf \U$38801 ( \46596 , \46595 );
and \U$38802 ( \46597 , \46554 , \46559 );
and \U$38803 ( \46598 , \46554 , \46561 );
and \U$38804 ( \46599 , \46559 , \46561 );
or \U$38805 ( \46600 , \46597 , \46598 , \46599 );
buf \U$38806 ( \46601 , \46600 );
and \U$38807 ( \46602 , \46515 , \46519 );
and \U$38808 ( \46603 , \46515 , \46526 );
and \U$38809 ( \46604 , \46519 , \46526 );
or \U$38810 ( \46605 , \46602 , \46603 , \46604 );
buf \U$38811 ( \46606 , \46605 );
and \U$38812 ( \46607 , \21658 , \43179_nG9b51 );
or \U$38814 ( \46608 , \46607 , 1'b0 );
xor \U$38815 ( \46609 , \21654 , \46608 );
buf \U$38816 ( \46610 , \46609 );
buf \U$38817 ( \46611 , \46610 );
not \U$38818 ( \46612 , \46611 );
xor \U$38819 ( \46613 , \46606 , \46612 );
and \U$38820 ( \46614 , \23201 , \42766_nG9b57 );
and \U$38821 ( \46615 , \23198 , \42848_nG9b54 );
or \U$38822 ( \46616 , \46614 , \46615 );
xor \U$38823 ( \46617 , \23197 , \46616 );
buf \U$38824 ( \46618 , \46617 );
buf \U$38826 ( \46619 , \46618 );
xor \U$38827 ( \46620 , \46613 , \46619 );
buf \U$38828 ( \46621 , \46620 );
xor \U$38829 ( \46622 , \46601 , \46621 );
and \U$38831 ( \46623 , \32916 , \39591_nG9b78 );
or \U$38832 ( \46624 , 1'b0 , \46623 );
xor \U$38833 ( \46625 , 1'b0 , \46624 );
buf \U$38834 ( \46626 , \46625 );
buf \U$38836 ( \46627 , \46626 );
and \U$38837 ( \46628 , \28118 , \41040_nG9b69 );
and \U$38838 ( \46629 , \28115 , \41381_nG9b66 );
or \U$38839 ( \46630 , \46628 , \46629 );
xor \U$38840 ( \46631 , \28114 , \46630 );
buf \U$38841 ( \46632 , \46631 );
buf \U$38843 ( \46633 , \46632 );
xor \U$38844 ( \46634 , \46627 , \46633 );
and \U$38845 ( \46635 , \26431 , \41685_nG9b63 );
and \U$38846 ( \46636 , \26428 , \41963_nG9b60 );
or \U$38847 ( \46637 , \46635 , \46636 );
xor \U$38848 ( \46638 , \26427 , \46637 );
buf \U$38849 ( \46639 , \46638 );
buf \U$38851 ( \46640 , \46639 );
xor \U$38852 ( \46641 , \46634 , \46640 );
buf \U$38853 ( \46642 , \46641 );
xor \U$38854 ( \46643 , \46622 , \46642 );
buf \U$38855 ( \46644 , \46643 );
xor \U$38856 ( \46645 , \46596 , \46644 );
and \U$38857 ( \46646 , \46493 , \46499 );
and \U$38858 ( \46647 , \46493 , \46506 );
and \U$38859 ( \46648 , \46499 , \46506 );
or \U$38860 ( \46649 , \46646 , \46647 , \46648 );
buf \U$38861 ( \46650 , \46649 );
and \U$38862 ( \46651 , \31636 , \39963_nG9b75 );
and \U$38863 ( \46652 , \31633 , \40204_nG9b72 );
or \U$38864 ( \46653 , \46651 , \46652 );
xor \U$38865 ( \46654 , \31632 , \46653 );
buf \U$38866 ( \46655 , \46654 );
buf \U$38868 ( \46656 , \46655 );
and \U$38869 ( \46657 , \29853 , \40452_nG9b6f );
and \U$38870 ( \46658 , \29850 , \40843_nG9b6c );
or \U$38871 ( \46659 , \46657 , \46658 );
xor \U$38872 ( \46660 , \29849 , \46659 );
buf \U$38873 ( \46661 , \46660 );
buf \U$38875 ( \46662 , \46661 );
xor \U$38876 ( \46663 , \46656 , \46662 );
and \U$38877 ( \46664 , \24792 , \42201_nG9b5d );
and \U$38878 ( \46665 , \24789 , \42433_nG9b5a );
or \U$38879 ( \46666 , \46664 , \46665 );
xor \U$38880 ( \46667 , \24788 , \46666 );
buf \U$38881 ( \46668 , \46667 );
buf \U$38883 ( \46669 , \46668 );
xor \U$38884 ( \46670 , \46663 , \46669 );
buf \U$38885 ( \46671 , \46670 );
xor \U$38886 ( \46672 , \46650 , \46671 );
and \U$38887 ( \46673 , \46473 , \46479 );
and \U$38888 ( \46674 , \46473 , \46486 );
and \U$38889 ( \46675 , \46479 , \46486 );
or \U$38890 ( \46676 , \46673 , \46674 , \46675 );
buf \U$38891 ( \46677 , \46676 );
xor \U$38892 ( \46678 , \46672 , \46677 );
buf \U$38893 ( \46679 , \46678 );
xor \U$38894 ( \46680 , \46645 , \46679 );
buf \U$38895 ( \46681 , \46680 );
xor \U$38896 ( \46682 , \46591 , \46681 );
and \U$38897 ( \46683 , \46549 , \46563 );
and \U$38898 ( \46684 , \46549 , \46569 );
and \U$38899 ( \46685 , \46563 , \46569 );
or \U$38900 ( \46686 , \46683 , \46684 , \46685 );
buf \U$38901 ( \46687 , \46686 );
xor \U$38902 ( \46688 , \46682 , \46687 );
and \U$38903 ( \46689 , \46586 , \46688 );
and \U$38905 ( \46690 , \46580 , \46585 );
or \U$38907 ( \46691 , 1'b0 , \46690 , 1'b0 );
xor \U$38908 ( \46692 , \46689 , \46691 );
and \U$38910 ( \46693 , \46573 , \46579 );
and \U$38911 ( \46694 , \46575 , \46579 );
or \U$38912 ( \46695 , 1'b0 , \46693 , \46694 );
xor \U$38913 ( \46696 , \46692 , \46695 );
xor \U$38920 ( \46697 , \46696 , 1'b0 );
and \U$38921 ( \46698 , \46591 , \46681 );
and \U$38922 ( \46699 , \46591 , \46687 );
and \U$38923 ( \46700 , \46681 , \46687 );
or \U$38924 ( \46701 , \46698 , \46699 , \46700 );
xor \U$38925 ( \46702 , \46697 , \46701 );
and \U$38926 ( \46703 , \46596 , \46644 );
and \U$38927 ( \46704 , \46596 , \46679 );
and \U$38928 ( \46705 , \46644 , \46679 );
or \U$38929 ( \46706 , \46703 , \46704 , \46705 );
buf \U$38930 ( \46707 , \46706 );
and \U$38931 ( \46708 , \46601 , \46621 );
and \U$38932 ( \46709 , \46601 , \46642 );
and \U$38933 ( \46710 , \46621 , \46642 );
or \U$38934 ( \46711 , \46708 , \46709 , \46710 );
buf \U$38935 ( \46712 , \46711 );
and \U$38936 ( \46713 , \23201 , \42848_nG9b54 );
and \U$38937 ( \46714 , \23198 , \43179_nG9b51 );
or \U$38938 ( \46715 , \46713 , \46714 );
xor \U$38939 ( \46716 , \23197 , \46715 );
buf \U$38940 ( \46717 , \46716 );
buf \U$38942 ( \46718 , \46717 );
xor \U$38946 ( \46719 , \21654 , 1'b0 );
not \U$38947 ( \46720 , \46719 );
buf \U$38948 ( \46721 , \46720 );
buf \U$38950 ( \46722 , \46721 );
xor \U$38951 ( \46723 , \46718 , \46722 );
and \U$38952 ( \46724 , \26431 , \41963_nG9b60 );
and \U$38953 ( \46725 , \26428 , \42201_nG9b5d );
or \U$38954 ( \46726 , \46724 , \46725 );
xor \U$38955 ( \46727 , \26427 , \46726 );
buf \U$38956 ( \46728 , \46727 );
buf \U$38958 ( \46729 , \46728 );
xor \U$38959 ( \46730 , \46723 , \46729 );
buf \U$38960 ( \46731 , \46730 );
and \U$38961 ( \46732 , \46656 , \46662 );
and \U$38962 ( \46733 , \46656 , \46669 );
and \U$38963 ( \46734 , \46662 , \46669 );
or \U$38964 ( \46735 , \46732 , \46733 , \46734 );
buf \U$38965 ( \46736 , \46735 );
xor \U$38966 ( \46737 , \46731 , \46736 );
and \U$38967 ( \46738 , \46627 , \46633 );
and \U$38968 ( \46739 , \46627 , \46640 );
and \U$38969 ( \46740 , \46633 , \46640 );
or \U$38970 ( \46741 , \46738 , \46739 , \46740 );
buf \U$38971 ( \46742 , \46741 );
xor \U$38972 ( \46743 , \46737 , \46742 );
buf \U$38973 ( \46744 , \46743 );
xor \U$38974 ( \46745 , \46712 , \46744 );
and \U$38975 ( \46746 , \46650 , \46671 );
and \U$38976 ( \46747 , \46650 , \46677 );
and \U$38977 ( \46748 , \46671 , \46677 );
or \U$38978 ( \46749 , \46746 , \46747 , \46748 );
buf \U$38979 ( \46750 , \46749 );
xor \U$38980 ( \46751 , \46745 , \46750 );
buf \U$38981 ( \46752 , \46751 );
xor \U$38982 ( \46753 , \46707 , \46752 );
and \U$38983 ( \46754 , \46606 , \46612 );
and \U$38984 ( \46755 , \46606 , \46619 );
and \U$38985 ( \46756 , \46612 , \46619 );
or \U$38986 ( \46757 , \46754 , \46755 , \46756 );
buf \U$38987 ( \46758 , \46757 );
buf \U$38988 ( \46759 , \46611 );
and \U$38989 ( \46760 , \31636 , \40204_nG9b72 );
and \U$38990 ( \46761 , \31633 , \40452_nG9b6f );
or \U$38991 ( \46762 , \46760 , \46761 );
xor \U$38992 ( \46763 , \31632 , \46762 );
buf \U$38993 ( \46764 , \46763 );
buf \U$38995 ( \46765 , \46764 );
xor \U$38996 ( \46766 , \46759 , \46765 );
and \U$38997 ( \46767 , \24792 , \42433_nG9b5a );
and \U$38998 ( \46768 , \24789 , \42766_nG9b57 );
or \U$38999 ( \46769 , \46767 , \46768 );
xor \U$39000 ( \46770 , \24788 , \46769 );
buf \U$39001 ( \46771 , \46770 );
buf \U$39003 ( \46772 , \46771 );
xor \U$39004 ( \46773 , \46766 , \46772 );
buf \U$39005 ( \46774 , \46773 );
xor \U$39006 ( \46775 , \46758 , \46774 );
and \U$39008 ( \46776 , \32916 , \39963_nG9b75 );
or \U$39009 ( \46777 , 1'b0 , \46776 );
xor \U$39010 ( \46778 , 1'b0 , \46777 );
buf \U$39011 ( \46779 , \46778 );
buf \U$39013 ( \46780 , \46779 );
and \U$39014 ( \46781 , \29853 , \40843_nG9b6c );
and \U$39015 ( \46782 , \29850 , \41040_nG9b69 );
or \U$39016 ( \46783 , \46781 , \46782 );
xor \U$39017 ( \46784 , \29849 , \46783 );
buf \U$39018 ( \46785 , \46784 );
buf \U$39020 ( \46786 , \46785 );
xor \U$39021 ( \46787 , \46780 , \46786 );
and \U$39022 ( \46788 , \28118 , \41381_nG9b66 );
and \U$39023 ( \46789 , \28115 , \41685_nG9b63 );
or \U$39024 ( \46790 , \46788 , \46789 );
xor \U$39025 ( \46791 , \28114 , \46790 );
buf \U$39026 ( \46792 , \46791 );
buf \U$39028 ( \46793 , \46792 );
xor \U$39029 ( \46794 , \46787 , \46793 );
buf \U$39030 ( \46795 , \46794 );
xor \U$39031 ( \46796 , \46775 , \46795 );
buf \U$39032 ( \46797 , \46796 );
xor \U$39033 ( \46798 , \46753 , \46797 );
and \U$39034 ( \46799 , \46702 , \46798 );
and \U$39036 ( \46800 , \46696 , \46701 );
or \U$39038 ( \46801 , 1'b0 , \46800 , 1'b0 );
xor \U$39039 ( \46802 , \46799 , \46801 );
and \U$39041 ( \46803 , \46689 , \46695 );
and \U$39042 ( \46804 , \46691 , \46695 );
or \U$39043 ( \46805 , 1'b0 , \46803 , \46804 );
xor \U$39044 ( \46806 , \46802 , \46805 );
xor \U$39051 ( \46807 , \46806 , 1'b0 );
and \U$39052 ( \46808 , \46707 , \46752 );
and \U$39053 ( \46809 , \46707 , \46797 );
and \U$39054 ( \46810 , \46752 , \46797 );
or \U$39055 ( \46811 , \46808 , \46809 , \46810 );
xor \U$39056 ( \46812 , \46807 , \46811 );
and \U$39057 ( \46813 , \46712 , \46744 );
and \U$39058 ( \46814 , \46712 , \46750 );
and \U$39059 ( \46815 , \46744 , \46750 );
or \U$39060 ( \46816 , \46813 , \46814 , \46815 );
buf \U$39061 ( \46817 , \46816 );
and \U$39062 ( \46818 , \29853 , \41040_nG9b69 );
and \U$39063 ( \46819 , \29850 , \41381_nG9b66 );
or \U$39064 ( \46820 , \46818 , \46819 );
xor \U$39065 ( \46821 , \29849 , \46820 );
buf \U$39066 ( \46822 , \46821 );
buf \U$39068 ( \46823 , \46822 );
and \U$39069 ( \46824 , \28118 , \41685_nG9b63 );
and \U$39070 ( \46825 , \28115 , \41963_nG9b60 );
or \U$39071 ( \46826 , \46824 , \46825 );
xor \U$39072 ( \46827 , \28114 , \46826 );
buf \U$39073 ( \46828 , \46827 );
buf \U$39075 ( \46829 , \46828 );
xor \U$39076 ( \46830 , \46823 , \46829 );
and \U$39077 ( \46831 , \26431 , \42201_nG9b5d );
and \U$39078 ( \46832 , \26428 , \42433_nG9b5a );
or \U$39079 ( \46833 , \46831 , \46832 );
xor \U$39080 ( \46834 , \26427 , \46833 );
buf \U$39081 ( \46835 , \46834 );
buf \U$39083 ( \46836 , \46835 );
xor \U$39084 ( \46837 , \46830 , \46836 );
buf \U$39085 ( \46838 , \46837 );
and \U$39087 ( \46839 , \32916 , \40204_nG9b72 );
or \U$39088 ( \46840 , 1'b0 , \46839 );
xor \U$39089 ( \46841 , 1'b0 , \46840 );
buf \U$39090 ( \46842 , \46841 );
buf \U$39092 ( \46843 , \46842 );
and \U$39093 ( \46844 , \31636 , \40452_nG9b6f );
and \U$39094 ( \46845 , \31633 , \40843_nG9b6c );
or \U$39095 ( \46846 , \46844 , \46845 );
xor \U$39096 ( \46847 , \31632 , \46846 );
buf \U$39097 ( \46848 , \46847 );
buf \U$39099 ( \46849 , \46848 );
xor \U$39100 ( \46850 , \46843 , \46849 );
and \U$39101 ( \46851 , \24792 , \42766_nG9b57 );
and \U$39102 ( \46852 , \24789 , \42848_nG9b54 );
or \U$39103 ( \46853 , \46851 , \46852 );
xor \U$39104 ( \46854 , \24788 , \46853 );
buf \U$39105 ( \46855 , \46854 );
buf \U$39107 ( \46856 , \46855 );
xor \U$39108 ( \46857 , \46850 , \46856 );
buf \U$39109 ( \46858 , \46857 );
xor \U$39110 ( \46859 , \46838 , \46858 );
and \U$39111 ( \46860 , \46759 , \46765 );
and \U$39112 ( \46861 , \46759 , \46772 );
and \U$39113 ( \46862 , \46765 , \46772 );
or \U$39114 ( \46863 , \46860 , \46861 , \46862 );
buf \U$39115 ( \46864 , \46863 );
xor \U$39116 ( \46865 , \46859 , \46864 );
buf \U$39117 ( \46866 , \46865 );
and \U$39118 ( \46867 , \46731 , \46736 );
and \U$39119 ( \46868 , \46731 , \46742 );
and \U$39120 ( \46869 , \46736 , \46742 );
or \U$39121 ( \46870 , \46867 , \46868 , \46869 );
buf \U$39122 ( \46871 , \46870 );
xor \U$39123 ( \46872 , \46866 , \46871 );
and \U$39124 ( \46873 , \46718 , \46722 );
and \U$39125 ( \46874 , \46718 , \46729 );
and \U$39126 ( \46875 , \46722 , \46729 );
or \U$39127 ( \46876 , \46873 , \46874 , \46875 );
buf \U$39128 ( \46877 , \46876 );
and \U$39129 ( \46878 , \46780 , \46786 );
and \U$39130 ( \46879 , \46780 , \46793 );
and \U$39131 ( \46880 , \46786 , \46793 );
or \U$39132 ( \46881 , \46878 , \46879 , \46880 );
buf \U$39133 ( \46882 , \46881 );
xor \U$39134 ( \46883 , \46877 , \46882 );
and \U$39135 ( \46884 , \23201 , \43179_nG9b51 );
or \U$39137 ( \46885 , \46884 , 1'b0 );
xor \U$39138 ( \46886 , \23197 , \46885 );
buf \U$39139 ( \46887 , \46886 );
buf \U$39140 ( \46888 , \46887 );
not \U$39141 ( \46889 , \46888 );
xor \U$39142 ( \46890 , \46883 , \46889 );
buf \U$39143 ( \46891 , \46890 );
xor \U$39144 ( \46892 , \46872 , \46891 );
buf \U$39145 ( \46893 , \46892 );
xor \U$39146 ( \46894 , \46817 , \46893 );
and \U$39147 ( \46895 , \46758 , \46774 );
and \U$39148 ( \46896 , \46758 , \46795 );
and \U$39149 ( \46897 , \46774 , \46795 );
or \U$39150 ( \46898 , \46895 , \46896 , \46897 );
buf \U$39151 ( \46899 , \46898 );
xor \U$39152 ( \46900 , \46894 , \46899 );
and \U$39153 ( \46901 , \46812 , \46900 );
and \U$39155 ( \46902 , \46806 , \46811 );
or \U$39157 ( \46903 , 1'b0 , \46902 , 1'b0 );
xor \U$39158 ( \46904 , \46901 , \46903 );
and \U$39160 ( \46905 , \46799 , \46805 );
and \U$39161 ( \46906 , \46801 , \46805 );
or \U$39162 ( \46907 , 1'b0 , \46905 , \46906 );
xor \U$39163 ( \46908 , \46904 , \46907 );
xor \U$39170 ( \46909 , \46908 , 1'b0 );
and \U$39171 ( \46910 , \46817 , \46893 );
and \U$39172 ( \46911 , \46817 , \46899 );
and \U$39173 ( \46912 , \46893 , \46899 );
or \U$39174 ( \46913 , \46910 , \46911 , \46912 );
xor \U$39175 ( \46914 , \46909 , \46913 );
and \U$39176 ( \46915 , \46866 , \46871 );
and \U$39177 ( \46916 , \46866 , \46891 );
and \U$39178 ( \46917 , \46871 , \46891 );
or \U$39179 ( \46918 , \46915 , \46916 , \46917 );
buf \U$39180 ( \46919 , \46918 );
and \U$39181 ( \46920 , \46838 , \46858 );
and \U$39182 ( \46921 , \46838 , \46864 );
and \U$39183 ( \46922 , \46858 , \46864 );
or \U$39184 ( \46923 , \46920 , \46921 , \46922 );
buf \U$39185 ( \46924 , \46923 );
and \U$39186 ( \46925 , \46877 , \46882 );
and \U$39187 ( \46926 , \46877 , \46889 );
and \U$39188 ( \46927 , \46882 , \46889 );
or \U$39189 ( \46928 , \46925 , \46926 , \46927 );
buf \U$39190 ( \46929 , \46928 );
xor \U$39191 ( \46930 , \46924 , \46929 );
and \U$39192 ( \46931 , \46823 , \46829 );
and \U$39193 ( \46932 , \46823 , \46836 );
and \U$39194 ( \46933 , \46829 , \46836 );
or \U$39195 ( \46934 , \46931 , \46932 , \46933 );
buf \U$39196 ( \46935 , \46934 );
buf \U$39197 ( \46936 , \46888 );
xor \U$39198 ( \46937 , \46935 , \46936 );
and \U$39199 ( \46938 , \26431 , \42433_nG9b5a );
and \U$39200 ( \46939 , \26428 , \42766_nG9b57 );
or \U$39201 ( \46940 , \46938 , \46939 );
xor \U$39202 ( \46941 , \26427 , \46940 );
buf \U$39203 ( \46942 , \46941 );
buf \U$39205 ( \46943 , \46942 );
xor \U$39206 ( \46944 , \46937 , \46943 );
buf \U$39207 ( \46945 , \46944 );
xor \U$39208 ( \46946 , \46930 , \46945 );
buf \U$39209 ( \46947 , \46946 );
xor \U$39210 ( \46948 , \46919 , \46947 );
and \U$39212 ( \46949 , \32916 , \40452_nG9b6f );
or \U$39213 ( \46950 , 1'b0 , \46949 );
xor \U$39214 ( \46951 , 1'b0 , \46950 );
buf \U$39215 ( \46952 , \46951 );
buf \U$39217 ( \46953 , \46952 );
and \U$39218 ( \46954 , \31636 , \40843_nG9b6c );
and \U$39219 ( \46955 , \31633 , \41040_nG9b69 );
or \U$39220 ( \46956 , \46954 , \46955 );
xor \U$39221 ( \46957 , \31632 , \46956 );
buf \U$39222 ( \46958 , \46957 );
buf \U$39224 ( \46959 , \46958 );
xor \U$39225 ( \46960 , \46953 , \46959 );
and \U$39226 ( \46961 , \29853 , \41381_nG9b66 );
and \U$39227 ( \46962 , \29850 , \41685_nG9b63 );
or \U$39228 ( \46963 , \46961 , \46962 );
xor \U$39229 ( \46964 , \29849 , \46963 );
buf \U$39230 ( \46965 , \46964 );
buf \U$39232 ( \46966 , \46965 );
xor \U$39233 ( \46967 , \46960 , \46966 );
buf \U$39234 ( \46968 , \46967 );
and \U$39235 ( \46969 , \24792 , \42848_nG9b54 );
and \U$39236 ( \46970 , \24789 , \43179_nG9b51 );
or \U$39237 ( \46971 , \46969 , \46970 );
xor \U$39238 ( \46972 , \24788 , \46971 );
buf \U$39239 ( \46973 , \46972 );
buf \U$39241 ( \46974 , \46973 );
xor \U$39245 ( \46975 , \23197 , 1'b0 );
not \U$39246 ( \46976 , \46975 );
buf \U$39247 ( \46977 , \46976 );
buf \U$39249 ( \46978 , \46977 );
xor \U$39250 ( \46979 , \46974 , \46978 );
and \U$39251 ( \46980 , \28118 , \41963_nG9b60 );
and \U$39252 ( \46981 , \28115 , \42201_nG9b5d );
or \U$39253 ( \46982 , \46980 , \46981 );
xor \U$39254 ( \46983 , \28114 , \46982 );
buf \U$39255 ( \46984 , \46983 );
buf \U$39257 ( \46985 , \46984 );
xor \U$39258 ( \46986 , \46979 , \46985 );
buf \U$39259 ( \46987 , \46986 );
xor \U$39260 ( \46988 , \46968 , \46987 );
and \U$39261 ( \46989 , \46843 , \46849 );
and \U$39262 ( \46990 , \46843 , \46856 );
and \U$39263 ( \46991 , \46849 , \46856 );
or \U$39264 ( \46992 , \46989 , \46990 , \46991 );
buf \U$39265 ( \46993 , \46992 );
xor \U$39266 ( \46994 , \46988 , \46993 );
buf \U$39267 ( \46995 , \46994 );
xor \U$39268 ( \46996 , \46948 , \46995 );
and \U$39269 ( \46997 , \46914 , \46996 );
and \U$39271 ( \46998 , \46908 , \46913 );
or \U$39273 ( \46999 , 1'b0 , \46998 , 1'b0 );
xor \U$39274 ( \47000 , \46997 , \46999 );
and \U$39276 ( \47001 , \46901 , \46907 );
and \U$39277 ( \47002 , \46903 , \46907 );
or \U$39278 ( \47003 , 1'b0 , \47001 , \47002 );
xor \U$39279 ( \47004 , \47000 , \47003 );
xor \U$39286 ( \47005 , \47004 , 1'b0 );
and \U$39287 ( \47006 , \46919 , \46947 );
and \U$39288 ( \47007 , \46919 , \46995 );
and \U$39289 ( \47008 , \46947 , \46995 );
or \U$39290 ( \47009 , \47006 , \47007 , \47008 );
xor \U$39291 ( \47010 , \47005 , \47009 );
and \U$39292 ( \47011 , \46924 , \46929 );
and \U$39293 ( \47012 , \46924 , \46945 );
and \U$39294 ( \47013 , \46929 , \46945 );
or \U$39295 ( \47014 , \47011 , \47012 , \47013 );
buf \U$39296 ( \47015 , \47014 );
and \U$39297 ( \47016 , \46968 , \46987 );
and \U$39298 ( \47017 , \46968 , \46993 );
and \U$39299 ( \47018 , \46987 , \46993 );
or \U$39300 ( \47019 , \47016 , \47017 , \47018 );
buf \U$39301 ( \47020 , \47019 );
and \U$39302 ( \47021 , \46935 , \46936 );
and \U$39303 ( \47022 , \46935 , \46943 );
and \U$39304 ( \47023 , \46936 , \46943 );
or \U$39305 ( \47024 , \47021 , \47022 , \47023 );
buf \U$39306 ( \47025 , \47024 );
xor \U$39307 ( \47026 , \47020 , \47025 );
and \U$39308 ( \47027 , \29853 , \41685_nG9b63 );
and \U$39309 ( \47028 , \29850 , \41963_nG9b60 );
or \U$39310 ( \47029 , \47027 , \47028 );
xor \U$39311 ( \47030 , \29849 , \47029 );
buf \U$39312 ( \47031 , \47030 );
buf \U$39313 ( \47032 , \47031 );
not \U$39314 ( \47033 , \47032 );
and \U$39315 ( \47034 , \28118 , \42201_nG9b5d );
and \U$39316 ( \47035 , \28115 , \42433_nG9b5a );
or \U$39317 ( \47036 , \47034 , \47035 );
xor \U$39318 ( \47037 , \28114 , \47036 );
buf \U$39319 ( \47038 , \47037 );
buf \U$39321 ( \47039 , \47038 );
xor \U$39322 ( \47040 , \47033 , \47039 );
and \U$39323 ( \47041 , \26431 , \42766_nG9b57 );
and \U$39324 ( \47042 , \26428 , \42848_nG9b54 );
or \U$39325 ( \47043 , \47041 , \47042 );
xor \U$39326 ( \47044 , \26427 , \47043 );
buf \U$39327 ( \47045 , \47044 );
buf \U$39329 ( \47046 , \47045 );
xor \U$39330 ( \47047 , \47040 , \47046 );
buf \U$39331 ( \47048 , \47047 );
xor \U$39332 ( \47049 , \47026 , \47048 );
buf \U$39333 ( \47050 , \47049 );
xor \U$39334 ( \47051 , \47015 , \47050 );
and \U$39335 ( \47052 , \46974 , \46978 );
and \U$39336 ( \47053 , \46974 , \46985 );
and \U$39337 ( \47054 , \46978 , \46985 );
or \U$39338 ( \47055 , \47052 , \47053 , \47054 );
buf \U$39339 ( \47056 , \47055 );
and \U$39340 ( \47057 , \24792 , \43179_nG9b51 );
or \U$39342 ( \47058 , \47057 , 1'b0 );
xor \U$39343 ( \47059 , \24788 , \47058 );
buf \U$39344 ( \47060 , \47059 );
buf \U$39346 ( \47061 , \47060 );
and \U$39348 ( \47062 , \32916 , \40843_nG9b6c );
or \U$39349 ( \47063 , 1'b0 , \47062 );
xor \U$39350 ( \47064 , 1'b0 , \47063 );
buf \U$39351 ( \47065 , \47064 );
buf \U$39353 ( \47066 , \47065 );
xor \U$39354 ( \47067 , \47061 , \47066 );
and \U$39355 ( \47068 , \31636 , \41040_nG9b69 );
and \U$39356 ( \47069 , \31633 , \41381_nG9b66 );
or \U$39357 ( \47070 , \47068 , \47069 );
xor \U$39358 ( \47071 , \31632 , \47070 );
buf \U$39359 ( \47072 , \47071 );
buf \U$39361 ( \47073 , \47072 );
xor \U$39362 ( \47074 , \47067 , \47073 );
buf \U$39363 ( \47075 , \47074 );
xor \U$39364 ( \47076 , \47056 , \47075 );
and \U$39365 ( \47077 , \46953 , \46959 );
and \U$39366 ( \47078 , \46953 , \46966 );
and \U$39367 ( \47079 , \46959 , \46966 );
or \U$39368 ( \47080 , \47077 , \47078 , \47079 );
buf \U$39369 ( \47081 , \47080 );
xor \U$39370 ( \47082 , \47076 , \47081 );
buf \U$39371 ( \47083 , \47082 );
xor \U$39372 ( \47084 , \47051 , \47083 );
and \U$39373 ( \47085 , \47010 , \47084 );
and \U$39375 ( \47086 , \47004 , \47009 );
or \U$39377 ( \47087 , 1'b0 , \47086 , 1'b0 );
xor \U$39378 ( \47088 , \47085 , \47087 );
and \U$39380 ( \47089 , \46997 , \47003 );
and \U$39381 ( \47090 , \46999 , \47003 );
or \U$39382 ( \47091 , 1'b0 , \47089 , \47090 );
xor \U$39383 ( \47092 , \47088 , \47091 );
xor \U$39390 ( \47093 , \47092 , 1'b0 );
and \U$39391 ( \47094 , \26431 , \42848_nG9b54 );
and \U$39392 ( \47095 , \26428 , \43179_nG9b51 );
or \U$39393 ( \47096 , \47094 , \47095 );
xor \U$39394 ( \47097 , \26427 , \47096 );
buf \U$39395 ( \47098 , \47097 );
buf \U$39397 ( \47099 , \47098 );
xor \U$39401 ( \47100 , \24788 , 1'b0 );
not \U$39402 ( \47101 , \47100 );
buf \U$39403 ( \47102 , \47101 );
buf \U$39405 ( \47103 , \47102 );
xor \U$39406 ( \47104 , \47099 , \47103 );
and \U$39407 ( \47105 , \29853 , \41963_nG9b60 );
and \U$39408 ( \47106 , \29850 , \42201_nG9b5d );
or \U$39409 ( \47107 , \47105 , \47106 );
xor \U$39410 ( \47108 , \29849 , \47107 );
buf \U$39411 ( \47109 , \47108 );
buf \U$39413 ( \47110 , \47109 );
xor \U$39414 ( \47111 , \47104 , \47110 );
buf \U$39415 ( \47112 , \47111 );
and \U$39416 ( \47113 , \47033 , \47039 );
and \U$39417 ( \47114 , \47033 , \47046 );
and \U$39418 ( \47115 , \47039 , \47046 );
or \U$39419 ( \47116 , \47113 , \47114 , \47115 );
buf \U$39420 ( \47117 , \47116 );
xor \U$39421 ( \47118 , \47112 , \47117 );
and \U$39422 ( \47119 , \47061 , \47066 );
and \U$39423 ( \47120 , \47061 , \47073 );
and \U$39424 ( \47121 , \47066 , \47073 );
or \U$39425 ( \47122 , \47119 , \47120 , \47121 );
buf \U$39426 ( \47123 , \47122 );
and \U$39428 ( \47124 , \32916 , \41040_nG9b69 );
or \U$39429 ( \47125 , 1'b0 , \47124 );
xor \U$39430 ( \47126 , 1'b0 , \47125 );
buf \U$39431 ( \47127 , \47126 );
buf \U$39433 ( \47128 , \47127 );
and \U$39434 ( \47129 , \31636 , \41381_nG9b66 );
and \U$39435 ( \47130 , \31633 , \41685_nG9b63 );
or \U$39436 ( \47131 , \47129 , \47130 );
xor \U$39437 ( \47132 , \31632 , \47131 );
buf \U$39438 ( \47133 , \47132 );
buf \U$39440 ( \47134 , \47133 );
xor \U$39441 ( \47135 , \47128 , \47134 );
and \U$39442 ( \47136 , \28118 , \42433_nG9b5a );
and \U$39443 ( \47137 , \28115 , \42766_nG9b57 );
or \U$39444 ( \47138 , \47136 , \47137 );
xor \U$39445 ( \47139 , \28114 , \47138 );
buf \U$39446 ( \47140 , \47139 );
buf \U$39448 ( \47141 , \47140 );
xor \U$39449 ( \47142 , \47135 , \47141 );
buf \U$39450 ( \47143 , \47142 );
xor \U$39451 ( \47144 , \47123 , \47143 );
buf \U$39452 ( \47145 , \47032 );
xor \U$39453 ( \47146 , \47144 , \47145 );
buf \U$39454 ( \47147 , \47146 );
xor \U$39455 ( \47148 , \47118 , \47147 );
buf \U$39456 ( \47149 , \47148 );
and \U$39457 ( \47150 , \47020 , \47025 );
and \U$39458 ( \47151 , \47020 , \47048 );
and \U$39459 ( \47152 , \47025 , \47048 );
or \U$39460 ( \47153 , \47150 , \47151 , \47152 );
buf \U$39461 ( \47154 , \47153 );
xor \U$39462 ( \47155 , \47149 , \47154 );
and \U$39463 ( \47156 , \47056 , \47075 );
and \U$39464 ( \47157 , \47056 , \47081 );
and \U$39465 ( \47158 , \47075 , \47081 );
or \U$39466 ( \47159 , \47156 , \47157 , \47158 );
buf \U$39467 ( \47160 , \47159 );
xor \U$39468 ( \47161 , \47155 , \47160 );
xor \U$39469 ( \47162 , \47093 , \47161 );
and \U$39470 ( \47163 , \47015 , \47050 );
and \U$39471 ( \47164 , \47015 , \47083 );
and \U$39472 ( \47165 , \47050 , \47083 );
or \U$39473 ( \47166 , \47163 , \47164 , \47165 );
and \U$39474 ( \47167 , \47162 , \47166 );
and \U$39476 ( \47168 , \47092 , \47161 );
or \U$39478 ( \47169 , 1'b0 , \47168 , 1'b0 );
xor \U$39479 ( \47170 , \47167 , \47169 );
and \U$39481 ( \47171 , \47085 , \47091 );
and \U$39482 ( \47172 , \47087 , \47091 );
or \U$39483 ( \47173 , 1'b0 , \47171 , \47172 );
xor \U$39484 ( \47174 , \47170 , \47173 );
xor \U$39491 ( \47175 , \47174 , 1'b0 );
and \U$39492 ( \47176 , \47112 , \47117 );
and \U$39493 ( \47177 , \47112 , \47147 );
and \U$39494 ( \47178 , \47117 , \47147 );
or \U$39495 ( \47179 , \47176 , \47177 , \47178 );
buf \U$39496 ( \47180 , \47179 );
and \U$39497 ( \47181 , \47099 , \47103 );
and \U$39498 ( \47182 , \47099 , \47110 );
and \U$39499 ( \47183 , \47103 , \47110 );
or \U$39500 ( \47184 , \47181 , \47182 , \47183 );
buf \U$39501 ( \47185 , \47184 );
and \U$39502 ( \47186 , \31636 , \41685_nG9b63 );
and \U$39503 ( \47187 , \31633 , \41963_nG9b60 );
or \U$39504 ( \47188 , \47186 , \47187 );
xor \U$39505 ( \47189 , \31632 , \47188 );
buf \U$39506 ( \47190 , \47189 );
buf \U$39507 ( \47191 , \47190 );
not \U$39508 ( \47192 , \47191 );
xor \U$39509 ( \47193 , \47185 , \47192 );
and \U$39510 ( \47194 , \28118 , \42766_nG9b57 );
and \U$39511 ( \47195 , \28115 , \42848_nG9b54 );
or \U$39512 ( \47196 , \47194 , \47195 );
xor \U$39513 ( \47197 , \28114 , \47196 );
buf \U$39514 ( \47198 , \47197 );
buf \U$39516 ( \47199 , \47198 );
xor \U$39517 ( \47200 , \47193 , \47199 );
buf \U$39518 ( \47201 , \47200 );
and \U$39519 ( \47202 , \26431 , \43179_nG9b51 );
or \U$39521 ( \47203 , \47202 , 1'b0 );
xor \U$39522 ( \47204 , \26427 , \47203 );
buf \U$39523 ( \47205 , \47204 );
buf \U$39525 ( \47206 , \47205 );
and \U$39527 ( \47207 , \32916 , \41381_nG9b66 );
or \U$39528 ( \47208 , 1'b0 , \47207 );
xor \U$39529 ( \47209 , 1'b0 , \47208 );
buf \U$39530 ( \47210 , \47209 );
buf \U$39532 ( \47211 , \47210 );
xor \U$39533 ( \47212 , \47206 , \47211 );
and \U$39534 ( \47213 , \29853 , \42201_nG9b5d );
and \U$39535 ( \47214 , \29850 , \42433_nG9b5a );
or \U$39536 ( \47215 , \47213 , \47214 );
xor \U$39537 ( \47216 , \29849 , \47215 );
buf \U$39538 ( \47217 , \47216 );
buf \U$39540 ( \47218 , \47217 );
xor \U$39541 ( \47219 , \47212 , \47218 );
buf \U$39542 ( \47220 , \47219 );
xor \U$39543 ( \47221 , \47201 , \47220 );
and \U$39544 ( \47222 , \47128 , \47134 );
and \U$39545 ( \47223 , \47128 , \47141 );
and \U$39546 ( \47224 , \47134 , \47141 );
or \U$39547 ( \47225 , \47222 , \47223 , \47224 );
buf \U$39548 ( \47226 , \47225 );
xor \U$39549 ( \47227 , \47221 , \47226 );
buf \U$39550 ( \47228 , \47227 );
xor \U$39551 ( \47229 , \47180 , \47228 );
and \U$39552 ( \47230 , \47123 , \47143 );
and \U$39553 ( \47231 , \47123 , \47145 );
and \U$39554 ( \47232 , \47143 , \47145 );
or \U$39555 ( \47233 , \47230 , \47231 , \47232 );
buf \U$39556 ( \47234 , \47233 );
xor \U$39557 ( \47235 , \47229 , \47234 );
xor \U$39558 ( \47236 , \47175 , \47235 );
and \U$39559 ( \47237 , \47149 , \47154 );
and \U$39560 ( \47238 , \47149 , \47160 );
and \U$39561 ( \47239 , \47154 , \47160 );
or \U$39562 ( \47240 , \47237 , \47238 , \47239 );
and \U$39563 ( \47241 , \47236 , \47240 );
and \U$39565 ( \47242 , \47174 , \47235 );
or \U$39567 ( \47243 , 1'b0 , \47242 , 1'b0 );
xor \U$39568 ( \47244 , \47241 , \47243 );
and \U$39570 ( \47245 , \47167 , \47173 );
and \U$39571 ( \47246 , \47169 , \47173 );
or \U$39572 ( \47247 , 1'b0 , \47245 , \47246 );
xor \U$39573 ( \47248 , \47244 , \47247 );
xor \U$39580 ( \47249 , \47248 , 1'b0 );
and \U$39581 ( \47250 , \47180 , \47228 );
and \U$39582 ( \47251 , \47180 , \47234 );
and \U$39583 ( \47252 , \47228 , \47234 );
or \U$39584 ( \47253 , \47250 , \47251 , \47252 );
xor \U$39585 ( \47254 , \47249 , \47253 );
and \U$39586 ( \47255 , \47185 , \47192 );
and \U$39587 ( \47256 , \47185 , \47199 );
and \U$39588 ( \47257 , \47192 , \47199 );
or \U$39589 ( \47258 , \47255 , \47256 , \47257 );
buf \U$39590 ( \47259 , \47258 );
and \U$39592 ( \47260 , \32916 , \41685_nG9b63 );
or \U$39593 ( \47261 , 1'b0 , \47260 );
xor \U$39594 ( \47262 , 1'b0 , \47261 );
buf \U$39595 ( \47263 , \47262 );
buf \U$39597 ( \47264 , \47263 );
buf \U$39598 ( \47265 , \47191 );
xor \U$39599 ( \47266 , \47264 , \47265 );
and \U$39600 ( \47267 , \29853 , \42433_nG9b5a );
and \U$39601 ( \47268 , \29850 , \42766_nG9b57 );
or \U$39602 ( \47269 , \47267 , \47268 );
xor \U$39603 ( \47270 , \29849 , \47269 );
buf \U$39604 ( \47271 , \47270 );
buf \U$39606 ( \47272 , \47271 );
xor \U$39607 ( \47273 , \47266 , \47272 );
buf \U$39608 ( \47274 , \47273 );
and \U$39609 ( \47275 , \28118 , \42848_nG9b54 );
and \U$39610 ( \47276 , \28115 , \43179_nG9b51 );
or \U$39611 ( \47277 , \47275 , \47276 );
xor \U$39612 ( \47278 , \28114 , \47277 );
buf \U$39613 ( \47279 , \47278 );
buf \U$39615 ( \47280 , \47279 );
xor \U$39619 ( \47281 , \26427 , 1'b0 );
not \U$39620 ( \47282 , \47281 );
buf \U$39621 ( \47283 , \47282 );
buf \U$39623 ( \47284 , \47283 );
xor \U$39624 ( \47285 , \47280 , \47284 );
and \U$39625 ( \47286 , \31636 , \41963_nG9b60 );
and \U$39626 ( \47287 , \31633 , \42201_nG9b5d );
or \U$39627 ( \47288 , \47286 , \47287 );
xor \U$39628 ( \47289 , \31632 , \47288 );
buf \U$39629 ( \47290 , \47289 );
buf \U$39631 ( \47291 , \47290 );
xor \U$39632 ( \47292 , \47285 , \47291 );
buf \U$39633 ( \47293 , \47292 );
xor \U$39634 ( \47294 , \47274 , \47293 );
and \U$39635 ( \47295 , \47206 , \47211 );
and \U$39636 ( \47296 , \47206 , \47218 );
and \U$39637 ( \47297 , \47211 , \47218 );
or \U$39638 ( \47298 , \47295 , \47296 , \47297 );
buf \U$39639 ( \47299 , \47298 );
xor \U$39640 ( \47300 , \47294 , \47299 );
buf \U$39641 ( \47301 , \47300 );
xor \U$39642 ( \47302 , \47259 , \47301 );
and \U$39643 ( \47303 , \47201 , \47220 );
and \U$39644 ( \47304 , \47201 , \47226 );
and \U$39645 ( \47305 , \47220 , \47226 );
or \U$39646 ( \47306 , \47303 , \47304 , \47305 );
buf \U$39647 ( \47307 , \47306 );
xor \U$39648 ( \47308 , \47302 , \47307 );
and \U$39649 ( \47309 , \47254 , \47308 );
and \U$39651 ( \47310 , \47248 , \47253 );
or \U$39653 ( \47311 , 1'b0 , \47310 , 1'b0 );
xor \U$39654 ( \47312 , \47309 , \47311 );
and \U$39656 ( \47313 , \47241 , \47247 );
and \U$39657 ( \47314 , \47243 , \47247 );
or \U$39658 ( \47315 , 1'b0 , \47313 , \47314 );
xor \U$39659 ( \47316 , \47312 , \47315 );
xor \U$39666 ( \47317 , \47316 , 1'b0 );
and \U$39667 ( \47318 , \47274 , \47293 );
and \U$39668 ( \47319 , \47274 , \47299 );
and \U$39669 ( \47320 , \47293 , \47299 );
or \U$39670 ( \47321 , \47318 , \47319 , \47320 );
buf \U$39671 ( \47322 , \47321 );
and \U$39672 ( \47323 , \47280 , \47284 );
and \U$39673 ( \47324 , \47280 , \47291 );
and \U$39674 ( \47325 , \47284 , \47291 );
or \U$39675 ( \47326 , \47323 , \47324 , \47325 );
buf \U$39676 ( \47327 , \47326 );
and \U$39678 ( \47328 , \32916 , \41963_nG9b60 );
or \U$39679 ( \47329 , 1'b0 , \47328 );
xor \U$39680 ( \47330 , 1'b0 , \47329 );
buf \U$39681 ( \47331 , \47330 );
buf \U$39683 ( \47332 , \47331 );
and \U$39684 ( \47333 , \31636 , \42201_nG9b5d );
and \U$39685 ( \47334 , \31633 , \42433_nG9b5a );
or \U$39686 ( \47335 , \47333 , \47334 );
xor \U$39687 ( \47336 , \31632 , \47335 );
buf \U$39688 ( \47337 , \47336 );
buf \U$39690 ( \47338 , \47337 );
xor \U$39691 ( \47339 , \47332 , \47338 );
and \U$39692 ( \47340 , \29853 , \42766_nG9b57 );
and \U$39693 ( \47341 , \29850 , \42848_nG9b54 );
or \U$39694 ( \47342 , \47340 , \47341 );
xor \U$39695 ( \47343 , \29849 , \47342 );
buf \U$39696 ( \47344 , \47343 );
buf \U$39698 ( \47345 , \47344 );
xor \U$39699 ( \47346 , \47339 , \47345 );
buf \U$39700 ( \47347 , \47346 );
xor \U$39701 ( \47348 , \47327 , \47347 );
and \U$39702 ( \47349 , \28118 , \43179_nG9b51 );
or \U$39704 ( \47350 , \47349 , 1'b0 );
xor \U$39705 ( \47351 , \28114 , \47350 );
buf \U$39706 ( \47352 , \47351 );
buf \U$39707 ( \47353 , \47352 );
not \U$39708 ( \47354 , \47353 );
xor \U$39709 ( \47355 , \47348 , \47354 );
buf \U$39710 ( \47356 , \47355 );
xor \U$39711 ( \47357 , \47322 , \47356 );
and \U$39712 ( \47358 , \47264 , \47265 );
and \U$39713 ( \47359 , \47264 , \47272 );
and \U$39714 ( \47360 , \47265 , \47272 );
or \U$39715 ( \47361 , \47358 , \47359 , \47360 );
buf \U$39716 ( \47362 , \47361 );
xor \U$39717 ( \47363 , \47357 , \47362 );
xor \U$39718 ( \47364 , \47317 , \47363 );
and \U$39719 ( \47365 , \47259 , \47301 );
and \U$39720 ( \47366 , \47259 , \47307 );
and \U$39721 ( \47367 , \47301 , \47307 );
or \U$39722 ( \47368 , \47365 , \47366 , \47367 );
and \U$39723 ( \47369 , \47364 , \47368 );
and \U$39725 ( \47370 , \47316 , \47363 );
or \U$39727 ( \47371 , 1'b0 , \47370 , 1'b0 );
xor \U$39728 ( \47372 , \47369 , \47371 );
and \U$39730 ( \47373 , \47309 , \47315 );
and \U$39731 ( \47374 , \47311 , \47315 );
or \U$39732 ( \47375 , 1'b0 , \47373 , \47374 );
xor \U$39733 ( \47376 , \47372 , \47375 );
xor \U$39740 ( \47377 , \47376 , 1'b0 );
and \U$39741 ( \47378 , \47322 , \47356 );
and \U$39742 ( \47379 , \47322 , \47362 );
and \U$39743 ( \47380 , \47356 , \47362 );
or \U$39744 ( \47381 , \47378 , \47379 , \47380 );
xor \U$39745 ( \47382 , \47377 , \47381 );
and \U$39746 ( \47383 , \47327 , \47347 );
and \U$39747 ( \47384 , \47327 , \47354 );
and \U$39748 ( \47385 , \47347 , \47354 );
or \U$39749 ( \47386 , \47383 , \47384 , \47385 );
buf \U$39750 ( \47387 , \47386 );
and \U$39751 ( \47388 , \29853 , \42848_nG9b54 );
and \U$39752 ( \47389 , \29850 , \43179_nG9b51 );
or \U$39753 ( \47390 , \47388 , \47389 );
xor \U$39754 ( \47391 , \29849 , \47390 );
buf \U$39755 ( \47392 , \47391 );
buf \U$39757 ( \47393 , \47392 );
xor \U$39761 ( \47394 , \28114 , 1'b0 );
not \U$39762 ( \47395 , \47394 );
buf \U$39763 ( \47396 , \47395 );
buf \U$39765 ( \47397 , \47396 );
xor \U$39766 ( \47398 , \47393 , \47397 );
and \U$39768 ( \47399 , \32916 , \42201_nG9b5d );
or \U$39769 ( \47400 , 1'b0 , \47399 );
xor \U$39770 ( \47401 , 1'b0 , \47400 );
buf \U$39771 ( \47402 , \47401 );
buf \U$39773 ( \47403 , \47402 );
xor \U$39774 ( \47404 , \47398 , \47403 );
buf \U$39775 ( \47405 , \47404 );
buf \U$39776 ( \47406 , \47353 );
xor \U$39777 ( \47407 , \47405 , \47406 );
and \U$39778 ( \47408 , \31636 , \42433_nG9b5a );
and \U$39779 ( \47409 , \31633 , \42766_nG9b57 );
or \U$39780 ( \47410 , \47408 , \47409 );
xor \U$39781 ( \47411 , \31632 , \47410 );
buf \U$39782 ( \47412 , \47411 );
buf \U$39784 ( \47413 , \47412 );
xor \U$39785 ( \47414 , \47407 , \47413 );
buf \U$39786 ( \47415 , \47414 );
xor \U$39787 ( \47416 , \47387 , \47415 );
and \U$39788 ( \47417 , \47332 , \47338 );
and \U$39789 ( \47418 , \47332 , \47345 );
and \U$39790 ( \47419 , \47338 , \47345 );
or \U$39791 ( \47420 , \47417 , \47418 , \47419 );
buf \U$39792 ( \47421 , \47420 );
xor \U$39793 ( \47422 , \47416 , \47421 );
and \U$39794 ( \47423 , \47382 , \47422 );
and \U$39796 ( \47424 , \47376 , \47381 );
or \U$39798 ( \47425 , 1'b0 , \47424 , 1'b0 );
xor \U$39799 ( \47426 , \47423 , \47425 );
and \U$39801 ( \47427 , \47369 , \47375 );
and \U$39802 ( \47428 , \47371 , \47375 );
or \U$39803 ( \47429 , 1'b0 , \47427 , \47428 );
xor \U$39804 ( \47430 , \47426 , \47429 );
xor \U$39811 ( \47431 , \47430 , 1'b0 );
and \U$39812 ( \47432 , \47405 , \47406 );
and \U$39813 ( \47433 , \47405 , \47413 );
and \U$39814 ( \47434 , \47406 , \47413 );
or \U$39815 ( \47435 , \47432 , \47433 , \47434 );
buf \U$39816 ( \47436 , \47435 );
and \U$39817 ( \47437 , \29853 , \43179_nG9b51 );
or \U$39819 ( \47438 , \47437 , 1'b0 );
xor \U$39820 ( \47439 , \29849 , \47438 );
buf \U$39821 ( \47440 , \47439 );
buf \U$39822 ( \47441 , \47440 );
not \U$39823 ( \47442 , \47441 );
and \U$39825 ( \47443 , \32916 , \42433_nG9b5a );
or \U$39826 ( \47444 , 1'b0 , \47443 );
xor \U$39827 ( \47445 , 1'b0 , \47444 );
buf \U$39828 ( \47446 , \47445 );
buf \U$39830 ( \47447 , \47446 );
xor \U$39831 ( \47448 , \47442 , \47447 );
and \U$39832 ( \47449 , \31636 , \42766_nG9b57 );
and \U$39833 ( \47450 , \31633 , \42848_nG9b54 );
or \U$39834 ( \47451 , \47449 , \47450 );
xor \U$39835 ( \47452 , \31632 , \47451 );
buf \U$39836 ( \47453 , \47452 );
buf \U$39838 ( \47454 , \47453 );
xor \U$39839 ( \47455 , \47448 , \47454 );
buf \U$39840 ( \47456 , \47455 );
xor \U$39841 ( \47457 , \47436 , \47456 );
and \U$39842 ( \47458 , \47393 , \47397 );
and \U$39843 ( \47459 , \47393 , \47403 );
and \U$39844 ( \47460 , \47397 , \47403 );
or \U$39845 ( \47461 , \47458 , \47459 , \47460 );
buf \U$39846 ( \47462 , \47461 );
xor \U$39847 ( \47463 , \47457 , \47462 );
xor \U$39848 ( \47464 , \47431 , \47463 );
and \U$39849 ( \47465 , \47387 , \47415 );
and \U$39850 ( \47466 , \47387 , \47421 );
and \U$39851 ( \47467 , \47415 , \47421 );
or \U$39852 ( \47468 , \47465 , \47466 , \47467 );
and \U$39853 ( \47469 , \47464 , \47468 );
and \U$39855 ( \47470 , \47430 , \47463 );
or \U$39857 ( \47471 , 1'b0 , \47470 , 1'b0 );
xor \U$39858 ( \47472 , \47469 , \47471 );
and \U$39860 ( \47473 , \47423 , \47429 );
and \U$39861 ( \47474 , \47425 , \47429 );
or \U$39862 ( \47475 , 1'b0 , \47473 , \47474 );
xor \U$39863 ( \47476 , \47472 , \47475 );
xor \U$39865 ( \47477 , \47476 , 1'b1 );
buf \U$39867 ( \47478 , \47441 );
xor \U$39868 ( \47479 , 1'b1 , \47478 );
and \U$39870 ( \47480 , \32916 , \42766_nG9b57 );
or \U$39871 ( \47481 , 1'b0 , \47480 );
xor \U$39872 ( \47482 , 1'b0 , \47481 );
buf \U$39873 ( \47483 , \47482 );
buf \U$39874 ( \47484 , \47483 );
not \U$39875 ( \47485 , \47484 );
xor \U$39876 ( \47486 , \47479 , \47485 );
buf \U$39877 ( \47487 , \47486 );
xor \U$39881 ( \47488 , \29849 , 1'b0 );
not \U$39882 ( \47489 , \47488 );
buf \U$39883 ( \47490 , \47489 );
buf \U$39885 ( \47491 , \47490 );
buf \U$39886 ( \47492 , \47484 );
xor \U$39887 ( \47493 , \47491 , \47492 );
buf \U$39888 ( \47494 , \47493 );
xor \U$39889 ( \47495 , \47487 , \47494 );
xor \U$39890 ( \47496 , \47477 , \47495 );
xor \U$39897 ( \47497 , \47496 , 1'b0 );
and \U$39898 ( \47498 , \47442 , \47447 );
and \U$39899 ( \47499 , \47442 , \47454 );
and \U$39900 ( \47500 , \47447 , \47454 );
or \U$39901 ( \47501 , \47498 , \47499 , \47500 );
buf \U$39902 ( \47502 , \47501 );
and \U$39903 ( \47503 , \31636 , \42848_nG9b54 );
and \U$39904 ( \47504 , \31633 , \43179_nG9b51 );
or \U$39905 ( \47505 , \47503 , \47504 );
xor \U$39906 ( \47506 , \31632 , \47505 );
buf \U$39907 ( \47507 , \47506 );
buf \U$39909 ( \47508 , \47507 );
not \U$39910 ( \47509 , \47441 );
xor \U$39911 ( \47510 , \47508 , \47509 );
buf \U$39912 ( \47511 , \47484 );
xor \U$39913 ( \47512 , \47510 , \47511 );
buf \U$39914 ( \47513 , \47512 );
xor \U$39915 ( \47514 , \47502 , \47513 );
buf \U$39916 ( \47515 , \47441 );
xor \U$39917 ( \47516 , \47514 , \47515 );
xor \U$39918 ( \47517 , \47497 , \47516 );
and \U$39919 ( \47518 , \47436 , \47456 );
and \U$39920 ( \47519 , \47436 , \47462 );
and \U$39921 ( \47520 , \47456 , \47462 );
or \U$39922 ( \47521 , \47518 , \47519 , \47520 );
and \U$39923 ( \47522 , \47517 , \47521 );
and \U$39925 ( \47523 , \47496 , \47516 );
or \U$39927 ( \47524 , 1'b0 , \47523 , 1'b0 );
xor \U$39928 ( \47525 , \47522 , \47524 );
and \U$39929 ( \47526 , \47476 , 1'b1 );
and \U$39930 ( \47527 , \47476 , \47495 );
and \U$39931 ( \47528 , 1'b1 , \47495 );
or \U$39932 ( \47529 , \47526 , \47527 , \47528 );
xor \U$39933 ( \47530 , \47525 , \47529 );
and \U$39935 ( \47531 , \47469 , \47475 );
and \U$39936 ( \47532 , \47471 , \47475 );
or \U$39937 ( \47533 , 1'b0 , \47531 , \47532 );
xor \U$39938 ( \47534 , \47530 , \47533 );
and \U$39939 ( \47535 , \47487 , \47494 );
xor \U$39940 ( \47536 , \47534 , \47535 );
xor \U$39947 ( \47537 , \47536 , 1'b0 );
and \U$39949 ( \47538 , \32916 , \42848_nG9b54 );
or \U$39950 ( \47539 , 1'b0 , \47538 );
xor \U$39951 ( \47540 , 1'b0 , \47539 );
buf \U$39952 ( \47541 , \47540 );
buf \U$39953 ( \47542 , \47541 );
xor \U$39954 ( \47543 , \47537 , \47542 );
and \U$39955 ( \47544 , \47508 , \47509 );
and \U$39956 ( \47545 , \47508 , \47511 );
and \U$39957 ( \47546 , \47509 , \47511 );
or \U$39958 ( \47547 , \47544 , \47545 , \47546 );
buf \U$39959 ( \47548 , \47547 );
and \U$39960 ( \47549 , 1'b1 , \47478 );
and \U$39961 ( \47550 , 1'b1 , \47485 );
and \U$39962 ( \47551 , \47478 , \47485 );
or \U$39963 ( \47552 , \47549 , \47550 , \47551 );
buf \U$39964 ( \47553 , \47552 );
xor \U$39965 ( \47554 , \47548 , \47553 );
and \U$39967 ( \47555 , \47491 , \47492 );
buf \U$39968 ( \47556 , \47555 );
xor \U$39969 ( \47557 , 1'b1 , \47556 );
and \U$39970 ( \47558 , \31636 , \43179_nG9b51 );
or \U$39972 ( \47559 , \47558 , 1'b0 );
xor \U$39973 ( \47560 , \31632 , \47559 );
buf \U$39974 ( \47561 , \47560 );
buf \U$39976 ( \47562 , \47561 );
xor \U$39977 ( \47563 , \47557 , \47562 );
xor \U$39978 ( \47564 , \47554 , \47563 );
and \U$39979 ( \47565 , \47543 , \47564 );
and \U$39980 ( \47566 , \47502 , \47513 );
and \U$39981 ( \47567 , \47502 , \47515 );
and \U$39982 ( \47568 , \47513 , \47515 );
or \U$39983 ( \47569 , \47566 , \47567 , \47568 );
and \U$39984 ( \47570 , \47543 , \47569 );
and \U$39985 ( \47571 , \47564 , \47569 );
or \U$39986 ( \47572 , \47565 , \47570 , \47571 );
and \U$39988 ( \47573 , \47536 , \47542 );
or \U$39990 ( \47574 , 1'b0 , \47573 , 1'b0 );
xor \U$39991 ( \47575 , \47572 , \47574 );
and \U$39992 ( \47576 , \47530 , \47533 );
and \U$39993 ( \47577 , \47530 , \47535 );
and \U$39994 ( \47578 , \47533 , \47535 );
or \U$39995 ( \47579 , \47576 , \47577 , \47578 );
xor \U$39996 ( \47580 , \47575 , \47579 );
and \U$39998 ( \47581 , \47522 , \47529 );
and \U$39999 ( \47582 , \47524 , \47529 );
or \U$40000 ( \47583 , 1'b0 , \47581 , \47582 );
xor \U$40001 ( \47584 , \47580 , \47583 );
xor \U$40003 ( \47585 , \47584 , 1'b1 );
xor \U$40010 ( \47586 , \47585 , 1'b0 );
and \U$40012 ( \47587 , \32916 , \43179_nG9b51 );
or \U$40013 ( \47588 , 1'b0 , \47587 );
xor \U$40014 ( \47589 , 1'b0 , \47588 );
buf \U$40015 ( \47590 , \47589 );
buf \U$40016 ( \47591 , \47590 );
xor \U$40017 ( \47592 , \47586 , \47591 );
and \U$40018 ( \47593 , \47548 , \47553 );
and \U$40019 ( \47594 , \47548 , \47563 );
and \U$40020 ( \47595 , \47553 , \47563 );
or \U$40021 ( \47596 , \47593 , \47594 , \47595 );
xor \U$40022 ( \47597 , \47592 , \47596 );
and \U$40023 ( \47598 , 1'b1 , \47556 );
and \U$40024 ( \47599 , 1'b1 , \47562 );
and \U$40025 ( \47600 , \47556 , \47562 );
or \U$40026 ( \47601 , \47598 , \47599 , \47600 );
xor \U$40027 ( \47602 , \47597 , \47601 );
xor \U$40031 ( \47603 , \31632 , 1'b0 );
not \U$40032 ( \47604 , \47603 );
buf \U$40033 ( \47605 , \47604 );
buf \U$40034 ( \47606 , \47605 );
xor \U$40035 ( \47607 , \47602 , \47606 );
buf gdf4e ( \47608_nGdf4e , \47607 );
buf \U$40036 ( \47609 , \47608_nGdf4e );
xor \U$40037 ( \47610 , \47543 , \47564 );
xor \U$40038 ( \47611 , \47610 , \47569 );
buf gdf51 ( \47612_nGdf51 , \47611 );
buf \U$40039 ( \47613 , \47612_nGdf51 );
xor \U$40040 ( \47614 , \47517 , \47521 );
buf gdf53 ( \47615_nGdf53 , \47614 );
buf \U$40041 ( \47616 , \47615_nGdf53 );
xor \U$40042 ( \47617 , \47464 , \47468 );
buf gdf55 ( \47618_nGdf55 , \47617 );
buf \U$40043 ( \47619 , \47618_nGdf55 );
xor \U$40044 ( \47620 , \47382 , \47422 );
buf gdf57 ( \47621_nGdf57 , \47620 );
buf \U$40045 ( \47622 , \47621_nGdf57 );
xor \U$40046 ( \47623 , \47364 , \47368 );
buf gdf59 ( \47624_nGdf59 , \47623 );
buf \U$40047 ( \47625 , \47624_nGdf59 );
xor \U$40048 ( \47626 , \47254 , \47308 );
buf gdf5b ( \47627_nGdf5b , \47626 );
buf \U$40049 ( \47628 , \47627_nGdf5b );
xor \U$40050 ( \47629 , \47236 , \47240 );
buf gdf5d ( \47630_nGdf5d , \47629 );
buf \U$40051 ( \47631 , \47630_nGdf5d );
xor \U$40052 ( \47632 , \47162 , \47166 );
buf gdf5f ( \47633_nGdf5f , \47632 );
buf \U$40053 ( \47634 , \47633_nGdf5f );
xor \U$40054 ( \47635 , \47010 , \47084 );
buf gdf61 ( \47636_nGdf61 , \47635 );
buf \U$40055 ( \47637 , \47636_nGdf61 );
xor \U$40056 ( \47638 , \46914 , \46996 );
buf gdf63 ( \47639_nGdf63 , \47638 );
buf \U$40057 ( \47640 , \47639_nGdf63 );
xor \U$40058 ( \47641 , \46812 , \46900 );
buf gdf65 ( \47642_nGdf65 , \47641 );
buf \U$40059 ( \47643 , \47642_nGdf65 );
xor \U$40060 ( \47644 , \46702 , \46798 );
buf gdf67 ( \47645_nGdf67 , \47644 );
buf \U$40061 ( \47646 , \47645_nGdf67 );
xor \U$40062 ( \47647 , \46586 , \46688 );
buf gdf69 ( \47648_nGdf69 , \47647 );
buf \U$40063 ( \47649 , \47648_nGdf69 );
xor \U$40064 ( \47650 , \46462 , \46572 );
buf gdf6b ( \47651_nGdf6b , \47650 );
buf \U$40065 ( \47652 , \47651_nGdf6b );
xor \U$40066 ( \47653 , \46332 , \46448 );
buf gdf6d ( \47654_nGdf6d , \47653 );
buf \U$40067 ( \47655 , \47654_nGdf6d );
xor \U$40068 ( \47656 , \46314 , \46318 );
buf gdf6f ( \47657_nGdf6f , \47656 );
buf \U$40069 ( \47658 , \47657_nGdf6f );
xor \U$40070 ( \47659 , \46176 , \46180 );
buf gdf71 ( \47660_nGdf71 , \47659 );
buf \U$40071 ( \47661 , \47660_nGdf71 );
xor \U$40072 ( \47662 , \45898 , \46036 );
buf gdf73 ( \47663_nGdf73 , \47662 );
buf \U$40073 ( \47664 , \47663_nGdf73 );
xor \U$40074 ( \47665 , \45740 , \45884 );
buf gdf75 ( \47666_nGdf75 , \47665 );
buf \U$40075 ( \47667 , \47666_nGdf75 );
xor \U$40076 ( \47668 , \45574 , \45726 );
buf gdf77 ( \47669_nGdf77 , \47668 );
buf \U$40077 ( \47670 , \47669_nGdf77 );
xor \U$40078 ( \47671 , \45402 , \45560 );
buf gdf79 ( \47672_nGdf79 , \47671 );
buf \U$40079 ( \47673 , \47672_nGdf79 );
xor \U$40080 ( \47674 , \45222 , \45388 );
buf gdf7b ( \47675_nGdf7b , \47674 );
buf \U$40081 ( \47676 , \47675_nGdf7b );
xor \U$40082 ( \47677 , \45036 , \45208 );
buf gdf7d ( \47678_nGdf7d , \47677 );
buf \U$40083 ( \47679 , \47678_nGdf7d );
xor \U$40084 ( \47680 , \45018 , \45022 );
buf gdf7f ( \47681_nGdf7f , \47680 );
buf \U$40085 ( \47682 , \47681_nGdf7f );
xor \U$40086 ( \47683 , \44642 , \44828 );
buf gdf81 ( \47684_nGdf81 , \47683 );
buf \U$40087 ( \47685 , \47684_nGdf81 );
xor \U$40088 ( \47686 , \44434 , \44628 );
buf gdf83 ( \47687_nGdf83 , \47686 );
buf \U$40089 ( \47688 , \47687_nGdf83 );
xor \U$40090 ( \47689 , \44220 , \44420 );
buf gdf85 ( \47690_nGdf85 , \47689 );
buf \U$40091 ( \47691 , \47690_nGdf85 );
xor \U$40092 ( \47692 , \43998 , \44206 );
buf gdf87 ( \47693_nGdf87 , \47692 );
buf \U$40093 ( \47694 , \47693_nGdf87 );
xor \U$40094 ( \47695 , \43770 , \43984 );
buf gdf89 ( \47696_nGdf89 , \47695 );
buf \U$40095 ( \47697 , \47696_nGdf89 );
xor \U$40096 ( \47698 , \43538 , \43756 );
buf gdf8b ( \47699_nGdf8b , \47698 );
buf \U$40097 ( \47700 , \47699_nGdf8b );
xor \U$40098 ( \47701 , \43306 , \43524 );
buf gdf8d ( \47702_nGdf8d , \47701 );
buf \U$40099 ( \47703 , \47702_nGdf8d );
xor \U$40100 ( \47704 , \43058 , \43292 );
buf gdf8f ( \47705_nGdf8f , \47704 );
buf \U$40101 ( \47706 , \47705_nGdf8f );
xor \U$40102 ( \47707 , \42804 , \43044 );
buf gdf91 ( \47708_nGdf91 , \47707 );
buf \U$40103 ( \47709 , \47708_nGdf91 );
xor \U$40104 ( \47710 , \42546 , \42790 );
buf gdf93 ( \47711_nGdf93 , \47710 );
buf \U$40105 ( \47712 , \47711_nGdf93 );
xor \U$40106 ( \47713 , \42282 , \42532 );
buf gdf95 ( \47714_nGdf95 , \47713 );
buf \U$40107 ( \47715 , \47714_nGdf95 );
xor \U$40108 ( \47716 , \42014 , \42268 );
buf gdf97 ( \47717_nGdf97 , \47716 );
buf \U$40109 ( \47718 , \47717_nGdf97 );
xor \U$40110 ( \47719 , \41740 , \42000 );
buf gdf99 ( \47720_nGdf99 , \47719 );
buf \U$40111 ( \47721 , \47720_nGdf99 );
xor \U$40112 ( \47722 , \41462 , \41726 );
buf gdf9b ( \47723_nGdf9b , \47722 );
buf \U$40113 ( \47724 , \47723_nGdf9b );
xor \U$40114 ( \47725 , \41178 , \41448 );
buf gdf9d ( \47726_nGdf9d , \47725 );
buf \U$40115 ( \47727 , \47726_nGdf9d );
xor \U$40116 ( \47728 , \40890 , \41164 );
buf gdf9f ( \47729_nGdf9f , \47728 );
buf \U$40117 ( \47730 , \47729_nGdf9f );
xor \U$40118 ( \47731 , \40596 , \40876 );
buf gdfa1 ( \47732_nGdfa1 , \47731 );
buf \U$40119 ( \47733 , \47732_nGdfa1 );
xor \U$40120 ( \47734 , \40298 , \40582 );
buf gdfa3 ( \47735_nGdfa3 , \47734 );
buf \U$40121 ( \47736 , \47735_nGdfa3 );
xor \U$40122 ( \47737 , \39994 , \40284 );
buf gdfa5 ( \47738_nGdfa5 , \47737 );
buf \U$40123 ( \47739 , \47738_nGdfa5 );
xor \U$40124 ( \47740 , \39976 , \39980 );
buf gdfa7 ( \47741_nGdfa7 , \47740 );
buf \U$40125 ( \47742 , \47741_nGdfa7 );
xor \U$40126 ( \47743 , \39372 , \39672 );
buf gdfa9 ( \47744_nGdfa9 , \47743 );
buf \U$40127 ( \47745 , \47744_nGdfa9 );
xor \U$40128 ( \47746 , \39054 , \39358 );
buf gdfab ( \47747_nGdfab , \47746 );
buf \U$40129 ( \47748 , \47747_nGdfab );
xor \U$40130 ( \47749 , \38730 , \39040 );
buf gdfad ( \47750_nGdfad , \47749 );
buf \U$40131 ( \47751 , \47750_nGdfad );
xor \U$40132 ( \47752 , \38712 , \38716 );
buf gdfaf ( \47753_nGdfaf , \47752 );
buf \U$40133 ( \47754 , \47753_nGdfaf );
xor \U$40134 ( \47755 , \38068 , \38388 );
buf gdfb1 ( \47756_nGdfb1 , \47755 );
buf \U$40135 ( \47757 , \47756_nGdfb1 );
xor \U$40136 ( \47758 , \37730 , \38054 );
buf gdfb3 ( \47759_nGdfb3 , \47758 );
buf \U$40137 ( \47760 , \47759_nGdfb3 );
xor \U$40138 ( \47761 , \37386 , \37716 );
buf gdfb5 ( \47762_nGdfb5 , \47761 );
buf \U$40139 ( \47763 , \47762_nGdfb5 );
xor \U$40140 ( \47764 , \37038 , \37372 );
buf gdfb7 ( \47765_nGdfb7 , \47764 );
buf \U$40141 ( \47766 , \47765_nGdfb7 );
xor \U$40142 ( \47767 , \36684 , \37024 );
buf gdfb9 ( \47768_nGdfb9 , \47767 );
buf \U$40143 ( \47769 , \47768_nGdfb9 );
xor \U$40144 ( \47770 , \36326 , \36670 );
buf gdfbb ( \47771_nGdfbb , \47770 );
buf \U$40145 ( \47772 , \47771_nGdfbb );
xor \U$40146 ( \47773 , \35962 , \36312 );
buf gdfbd ( \47774_nGdfbd , \47773 );
buf \U$40147 ( \47775 , \47774_nGdfbd );
xor \U$40148 ( \47776 , \35594 , \35948 );
buf gdfbf ( \47777_nGdfbf , \47776 );
buf \U$40149 ( \47778 , \47777_nGdfbf );
xor \U$40150 ( \47779 , \35220 , \35580 );
buf gdfc1 ( \47780_nGdfc1 , \47779 );
buf \U$40151 ( \47781 , \47780_nGdfc1 );
xor \U$40152 ( \47782 , \34842 , \35206 );
buf gdfc3 ( \47783_nGdfc3 , \47782 );
buf \U$40153 ( \47784 , \47783_nGdfc3 );
xor \U$40154 ( \47785 , \34459 , \34829 );
buf gdfc5 ( \47786_nGdfc5 , \47785 );
buf \U$40155 ( \47787 , \47786_nGdfc5 );
xor \U$40156 ( \47788 , \34075 , \34446 );
buf gdfc7 ( \47789_nGdfc7 , \47788 );
buf \U$40157 ( \47790 , \47789_nGdfc7 );
xor \U$40158 ( \47791 , \33682 , \33686 );
xor \U$40159 ( \47792 , \47791 , \34062 );
buf gdfca ( \47793_nGdfca , \47792 );
buf \U$40160 ( \47794 , \47793_nGdfca );
xor \U$40161 ( \47795 , \33301 , \33670 );
xor \U$40162 ( \47796 , \47795 , \33675 );
buf gdfcd ( \47797_nGdfcd , \47796 );
buf \U$40163 ( \47798 , \47797_nGdfcd );
xor \U$40164 ( \47799 , \32924 , \32928 );
xor \U$40165 ( \47800 , \47799 , \33292 );
buf gdfd0 ( \47801_nGdfd0 , \47800 );
buf \U$40166 ( \47802 , \47801_nGdfd0 );
xor \U$40167 ( \47803 , \32905 , \32909 );
buf gdfd2 ( \47804_nGdfd2 , \47803 );
buf \U$40168 ( \47805 , \47804_nGdfd2 );
xor \U$40169 ( \47806 , \31643 , \31647 );
xor \U$40170 ( \47807 , \47806 , \32259 );
buf gdfd5 ( \47808_nGdfd5 , \47807 );
buf \U$40171 ( \47809 , \47808_nGdfd5 );
xor \U$40172 ( \47810 , \30465 , \31078 );
buf gdfd7 ( \47811_nGdfd7 , \47810 );
buf \U$40173 ( \47812 , \47811_nGdfd7 );
xor \U$40174 ( \47813 , \29860 , \29864 );
xor \U$40175 ( \47814 , \47813 , \30452 );
buf gdfda ( \47815_nGdfda , \47814 );
buf \U$40176 ( \47816 , \47815_nGdfda );
xor \U$40177 ( \47817 , \28706 , \29295 );
buf gdfdc ( \47818_nGdfdc , \47817 );
buf \U$40178 ( \47819 , \47818_nGdfdc );
xor \U$40179 ( \47820 , \28125 , \28129 );
xor \U$40180 ( \47821 , \47820 , \28693 );
buf gdfdf ( \47822_nGdfdf , \47821 );
buf \U$40181 ( \47823 , \47822_nGdfdf );
xor \U$40182 ( \47824 , \26995 , \27560 );
buf gdfe1 ( \47825_nGdfe1 , \47824 );
buf \U$40183 ( \47826 , \47825_nGdfe1 );
xor \U$40184 ( \47827 , \26438 , \26442 );
xor \U$40185 ( \47828 , \47827 , \26982 );
buf gdfe4 ( \47829_nGdfe4 , \47828 );
buf \U$40186 ( \47830 , \47829_nGdfe4 );
xor \U$40187 ( \47831 , \25869 , \25873 );
buf gdfe6 ( \47832_nGdfe6 , \47831 );
buf \U$40188 ( \47833 , \47832_nGdfe6 );
xor \U$40189 ( \47834 , \24799 , \25314 );
xor \U$40190 ( \47835 , \47834 , \25319 );
buf gdfe9 ( \47836_nGdfe9 , \47835 );
buf \U$40191 ( \47837 , \47836_nGdfe9 );
xor \U$40192 ( \47838 , \23717 , \24234 );
buf gdfeb ( \47839_nGdfeb , \47838 );
buf \U$40193 ( \47840 , \47839_nGdfeb );
xor \U$40194 ( \47841 , \23208 , \23212 );
xor \U$40195 ( \47842 , \47841 , \23704 );
buf gdfee ( \47843_nGdfee , \47842 );
buf \U$40196 ( \47844 , \47843_nGdfee );
xor \U$40197 ( \47845 , \22150 , \22643 );
buf gdff0 ( \47846_nGdff0 , \47845 );
buf \U$40198 ( \47847 , \47846_nGdff0 );
xor \U$40199 ( \47848 , \21665 , \21669 );
xor \U$40200 ( \47849 , \47848 , \22137 );
buf gdff3 ( \47850_nGdff3 , \47849 );
buf \U$40201 ( \47851 , \47850_nGdff3 );
xor \U$40202 ( \47852 , \20631 , \21100 );
buf gdff5 ( \47853_nGdff5 , \47852 );
buf \U$40203 ( \47854 , \47853_nGdff5 );
xor \U$40204 ( \47855 , \19603 , \20161 );
xor \U$40205 ( \47856 , \47855 , \20618 );
buf gdff8 ( \47857_nGdff8 , \47856 );
buf \U$40206 ( \47858 , \47857_nGdff8 );
xor \U$40207 ( \47859 , \19144 , \19602 );
buf gdffa ( \47860_nGdffa , \47859 );
buf \U$40208 ( \47861 , \47860_nGdffa );
xor \U$40209 ( \47862 , \18150 , \18708 );
xor \U$40210 ( \47863 , \47862 , \19141 );
buf gdffd ( \47864_nGdffd , \47863 );
buf \U$40211 ( \47865 , \47864_nGdffd );
xor \U$40212 ( \47866 , \17715 , \18149 );
buf gdfff ( \47867_nGdfff , \47866 );
buf \U$40213 ( \47868 , \47867_nGdfff );
xor \U$40214 ( \47869 , \16745 , \17303 );
xor \U$40215 ( \47870 , \47869 , \17712 );
buf ge002 ( \47871_nGe002 , \47870 );
buf \U$40216 ( \47872 , \47871_nGe002 );
xor \U$40217 ( \47873 , \16334 , \16744 );
buf ge004 ( \47874_nGe004 , \47873 );
buf \U$40218 ( \47875 , \47874_nGe004 );
xor \U$40219 ( \47876 , \15388 , \15946 );
xor \U$40220 ( \47877 , \47876 , \16331 );
buf ge007 ( \47878_nGe007 , \47877 );
buf \U$40221 ( \47879 , \47878_nGe007 );
xor \U$40222 ( \47880 , \15001 , \15387 );
buf ge009 ( \47881_nGe009 , \47880 );
buf \U$40223 ( \47882 , \47881_nGe009 );
xor \U$40224 ( \47883 , \14079 , \14637 );
xor \U$40225 ( \47884 , \47883 , \14998 );
buf ge00c ( \47885_nGe00c , \47884 );
buf \U$40226 ( \47886 , \47885_nGe00c );
xor \U$40227 ( \47887 , \13716 , \14078 );
buf ge00e ( \47888_nGe00e , \47887 );
buf \U$40228 ( \47889 , \47888_nGe00e );
xor \U$40229 ( \47890 , \12818 , \13376 );
xor \U$40230 ( \47891 , \47890 , \13713 );
buf ge011 ( \47892_nGe011 , \47891 );
buf \U$40231 ( \47893 , \47892_nGe011 );
xor \U$40232 ( \47894 , \12479 , \12817 );
buf ge013 ( \47895_nGe013 , \47894 );
buf \U$40233 ( \47896 , \47895_nGe013 );
xor \U$40234 ( \47897 , \11605 , \12163 );
xor \U$40235 ( \47898 , \47897 , \12476 );
buf ge016 ( \47899_nGe016 , \47898 );
buf \U$40236 ( \47900 , \47899_nGe016 );
xor \U$40237 ( \47901 , \11290 , \11604 );
buf ge018 ( \47902_nGe018 , \47901 );
buf \U$40238 ( \47903 , \47902_nGe018 );
endmodule

