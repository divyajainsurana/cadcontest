//
// Conformal-LEC Version 20.10-d005 (29-Apr-2020)
//
module top(RIb4ca3e8_33,RIa167a08_1,RIa167990_2,RIb4c6c20_34,RIa167918_3,RIb4c6ba8_35,RIa1678a0_4,RIb4c6b30_36,RIa167828_5,
        RIb4c6ab8_37,RIa1677b0_6,RIb4c6a40_38,RIa167738_7,RIb4c69c8_39,RIa1676c0_8,RIb4c6950_40,RIa167648_9,RIb4c68d8_41,RIa1675d0_10,
        RIb4c6860_42,RIa167558_11,RIb4c67e8_43,RIa1674e0_12,RIb4c6770_44,RIa167468_13,RIb4c3368_45,RIa1673f0_14,RIb4c32f0_46,RIa167378_15,
        RIb4c3278_47,RIa167300_16,RIb4c3200_48,RIa167288_17,RIb4c3188_49,RIa167210_18,RIb4c3110_50,RIa167198_19,RIb4c3098_51,RIa167120_20,
        RIb4c3020_52,RIa1670a8_21,RIb4c2fa8_53,RIa167030_22,RIb4c2f30_54,RIa166fb8_23,RIb4c2eb8_55,RIa166f40_24,RIb4c2e40_56,RIa166ec8_25,
        RIb4c2dc8_57,RIa166e50_26,RIb4c2d50_58,RIa166dd8_27,RIb4c2cd8_59,RIa166d60_28,RIb4c2c60_60,RIa166ce8_29,RIb4c2be8_61,RIa166c70_30,
        RIb4c2b70_62,RIb4ca4d8_31,RIb4c2af8_63,RIb4ca460_32,RIb4bfab0_64,RIb4bfa38_65,RIb4bf948_67,RIb4bf9c0_66,RIb4bf858_69,RIb4bf8d0_68,
        RIb4bf768_71,RIb4bf7e0_70,RIb4bf678_73,RIb4bf6f0_72,RIb4bf588_75,RIb4bf600_74,RIb4bf498_77,RIb4bf510_76,RIb4bf3a8_79,RIb4bf420_78,
        RIb4bf2b8_81,RIb4bf330_80,RIb4bf1c8_83,RIb4bf240_82,RIb4bf0d8_85,RIb4bf150_84,RIb4befe8_87,RIb4bf060_86,RIb4beef8_89,RIb4bef70_88,
        RIb4bc1f8_91,RIb4bee80_90,RIb4bc108_93,RIb4bc180_92,RIb4bc018_95,RIb4bc090_94,RIb4bbfa0_96,R_61_85b54e8,R_62_85b5590,R_63_85b5638,
        R_64_85b56e0,R_65_85b5788,R_66_85b5830,R_67_85b58d8,R_68_85b5980,R_69_85b5a28,R_6a_85b5ad0,R_6b_85b5b78,R_6c_85b5c20,R_6d_85b5cc8,
        R_6e_85b5d70,R_6f_85b5e18,R_70_85b5ec0,R_71_85b5f68,R_72_85b6010,R_73_85b60b8,R_74_85b6160,R_75_85b6208,R_76_85b62b0,R_77_85b6358,
        R_78_85b6400,R_79_85b64a8,R_7a_85b6550,R_7b_85b65f8,R_7c_85b66a0,R_7d_85b6748,R_7e_85b67f0,R_7f_85b6898,R_80_85b6940,R_81_85b69e8,
        R_82_85b6a90,R_83_85b6b38,R_84_85b6be0,R_85_85b6c88,R_86_85b6d30,R_87_85b6dd8,R_88_85b6e80,R_89_85b6f28,R_8a_85b6fd0,R_8b_85b7078,
        R_8c_85b7120,R_8d_85b71c8,R_8e_85b7270,R_8f_85b7318,R_90_85b73c0,R_91_85b7468,R_92_85b7510,R_93_85b75b8,R_94_85b7660,R_95_85b7708,
        R_96_85b77b0,R_97_85b7858,R_98_85b7900,R_99_85b79a8,R_9a_85b7a50);
input RIb4ca3e8_33,RIa167a08_1,RIa167990_2,RIb4c6c20_34,RIa167918_3,RIb4c6ba8_35,RIa1678a0_4,RIb4c6b30_36,RIa167828_5,
        RIb4c6ab8_37,RIa1677b0_6,RIb4c6a40_38,RIa167738_7,RIb4c69c8_39,RIa1676c0_8,RIb4c6950_40,RIa167648_9,RIb4c68d8_41,RIa1675d0_10,
        RIb4c6860_42,RIa167558_11,RIb4c67e8_43,RIa1674e0_12,RIb4c6770_44,RIa167468_13,RIb4c3368_45,RIa1673f0_14,RIb4c32f0_46,RIa167378_15,
        RIb4c3278_47,RIa167300_16,RIb4c3200_48,RIa167288_17,RIb4c3188_49,RIa167210_18,RIb4c3110_50,RIa167198_19,RIb4c3098_51,RIa167120_20,
        RIb4c3020_52,RIa1670a8_21,RIb4c2fa8_53,RIa167030_22,RIb4c2f30_54,RIa166fb8_23,RIb4c2eb8_55,RIa166f40_24,RIb4c2e40_56,RIa166ec8_25,
        RIb4c2dc8_57,RIa166e50_26,RIb4c2d50_58,RIa166dd8_27,RIb4c2cd8_59,RIa166d60_28,RIb4c2c60_60,RIa166ce8_29,RIb4c2be8_61,RIa166c70_30,
        RIb4c2b70_62,RIb4ca4d8_31,RIb4c2af8_63,RIb4ca460_32,RIb4bfab0_64,RIb4bfa38_65,RIb4bf948_67,RIb4bf9c0_66,RIb4bf858_69,RIb4bf8d0_68,
        RIb4bf768_71,RIb4bf7e0_70,RIb4bf678_73,RIb4bf6f0_72,RIb4bf588_75,RIb4bf600_74,RIb4bf498_77,RIb4bf510_76,RIb4bf3a8_79,RIb4bf420_78,
        RIb4bf2b8_81,RIb4bf330_80,RIb4bf1c8_83,RIb4bf240_82,RIb4bf0d8_85,RIb4bf150_84,RIb4befe8_87,RIb4bf060_86,RIb4beef8_89,RIb4bef70_88,
        RIb4bc1f8_91,RIb4bee80_90,RIb4bc108_93,RIb4bc180_92,RIb4bc018_95,RIb4bc090_94,RIb4bbfa0_96;
output R_61_85b54e8,R_62_85b5590,R_63_85b5638,R_64_85b56e0,R_65_85b5788,R_66_85b5830,R_67_85b58d8,R_68_85b5980,R_69_85b5a28,
        R_6a_85b5ad0,R_6b_85b5b78,R_6c_85b5c20,R_6d_85b5cc8,R_6e_85b5d70,R_6f_85b5e18,R_70_85b5ec0,R_71_85b5f68,R_72_85b6010,R_73_85b60b8,
        R_74_85b6160,R_75_85b6208,R_76_85b62b0,R_77_85b6358,R_78_85b6400,R_79_85b64a8,R_7a_85b6550,R_7b_85b65f8,R_7c_85b66a0,R_7d_85b6748,
        R_7e_85b67f0,R_7f_85b6898,R_80_85b6940,R_81_85b69e8,R_82_85b6a90,R_83_85b6b38,R_84_85b6be0,R_85_85b6c88,R_86_85b6d30,R_87_85b6dd8,
        R_88_85b6e80,R_89_85b6f28,R_8a_85b6fd0,R_8b_85b7078,R_8c_85b7120,R_8d_85b71c8,R_8e_85b7270,R_8f_85b7318,R_90_85b73c0,R_91_85b7468,
        R_92_85b7510,R_93_85b75b8,R_94_85b7660,R_95_85b7708,R_96_85b77b0,R_97_85b7858,R_98_85b7900,R_99_85b79a8,R_9a_85b7a50;

wire \155_ZERO , \156 , \157_N$1 , \158_ONE , \159 , \160 , \161 , \162 , \163 ,
         \164 , \165 , \166 , \167 , \168 , \169 , \170 , \171 , \172 , \173 ,
         \174 , \175 , \176 , \177 , \178 , \179 , \180 , \181 , \182 , \183 ,
         \184 , \185 , \186 , \187 , \188 , \189 , \190 , \191 , \192 , \193 ,
         \194 , \195 , \196 , \197 , \198 , \199 , \200 , \201 , \202 , \203 ,
         \204 , \205 , \206 , \207 , \208 , \209 , \210 , \211 , \212 , \213 ,
         \214 , \215 , \216 , \217 , \218 , \219 , \220 , \221 , \222 , \223 ,
         \224 , \225 , \226 , \227 , \228 , \229 , \230 , \231 , \232 , \233 ,
         \234 , \235 , \236 , \237 , \238 , \239 , \240 , \241 , \242 , \243 ,
         \244 , \245 , \246 , \247 , \248 , \249 , \250 , \251 , \252 , \253 ,
         \254 , \255 , \256 , \257 , \258 , \259 , \260 , \261 , \262 , \263 ,
         \264 , \265 , \266 , \267 , \268 , \269 , \270 , \271 , \272 , \273 ,
         \274 , \275 , \276 , \277 , \278 , \279 , \280 , \281 , \282 , \283 ,
         \284 , \285 , \286 , \287 , \288_nG143 , \289 , \290 , \291 , \292 , \293 ,
         \294 , \295 , \296 , \297 , \298 , \299 , \300 , \301 , \302 , \303_nG141 ,
         \304 , \305 , \306 , \307 , \308 , \309 , \310 , \311 , \312_nG142 , \313 ,
         \314 , \315 , \316 , \317 , \318 , \319 , \320 , \321_nG13f , \322 , \323 ,
         \324 , \325 , \326 , \327 , \328 , \329 , \330_nG140 , \331 , \332 , \333 ,
         \334 , \335 , \336 , \337 , \338 , \339 , \340 , \341_nG13d , \342 , \343 ,
         \344 , \345 , \346 , \347 , \348 , \349 , \350_nG13e , \351 , \352 , \353 ,
         \354 , \355 , \356 , \357 , \358_nG13c , \359 , \360 , \361 , \362 , \363 ,
         \364 , \365 , \366 , \367 , \368 , \369 , \370 , \371 , \372 , \373 ,
         \374 , \375 , \376 , \377 , \378 , \379 , \380 , \381 , \382 , \383 ,
         \384 , \385 , \386 , \387 , \388 , \389 , \390 , \391 , \392 , \393 ,
         \394 , \395 , \396 , \397 , \398 , \399 , \400 , \401 , \402 , \403 ,
         \404 , \405 , \406 , \407 , \408 , \409 , \410 , \411 , \412 , \413 ,
         \414 , \415 , \416 , \417 , \418 , \419 , \420 , \421 , \422 , \423 ,
         \424 , \425 , \426 , \427 , \428 , \429 , \430 , \431 , \432 , \433 ,
         \434 , \435 , \436 , \437 , \438 , \439 , \440 , \441 , \442 , \443_nG13b ,
         \444 , \445 , \446 , \447 , \448 , \449 , \450 , \451 , \452 , \453 ,
         \454 , \455 , \456 , \457 , \458 , \459 , \460 , \461 , \462 , \463 ,
         \464 , \465 , \466 , \467 , \468 , \469 , \470 , \471 , \472 , \473 ,
         \474 , \475 , \476 , \477 , \478 , \479 , \480 , \481 , \482 , \483 ,
         \484 , \485 , \486 , \487 , \488 , \489 , \490 , \491 , \492 , \493_nG13a ,
         \494 , \495 , \496 , \497 , \498 , \499 , \500 , \501 , \502 , \503 ,
         \504 , \505 , \506 , \507 , \508 , \509 , \510 , \511 , \512 , \513 ,
         \514 , \515 , \516 , \517 , \518 , \519 , \520 , \521 , \522 , \523 ,
         \524 , \525 , \526 , \527 , \528 , \529 , \530 , \531 , \532 , \533 ,
         \534 , \535 , \536 , \537 , \538 , \539 , \540 , \541 , \542 , \543 ,
         \544 , \545 , \546 , \547 , \548 , \549 , \550 , \551 , \552 , \553 ,
         \554 , \555 , \556 , \557 , \558 , \559 , \560 , \561 , \562 , \563 ,
         \564 , \565 , \566 , \567 , \568 , \569 , \570 , \571 , \572 , \573 ,
         \574 , \575 , \576 , \577 , \578 , \579 , \580 , \581 , \582 , \583 ,
         \584 , \585 , \586 , \587 , \588 , \589 , \590_nG139 , \591 , \592 , \593 ,
         \594 , \595 , \596 , \597 , \598 , \599 , \600 , \601 , \602 , \603 ,
         \604 , \605 , \606 , \607 , \608 , \609 , \610 , \611 , \612 , \613 ,
         \614 , \615 , \616 , \617 , \618 , \619_nG138 , \620 , \621 , \622 , \623 ,
         \624 , \625 , \626 , \627 , \628 , \629 , \630 , \631 , \632 , \633 ,
         \634 , \635 , \636 , \637 , \638 , \639 , \640 , \641 , \642 , \643 ,
         \644 , \645 , \646 , \647 , \648 , \649 , \650 , \651 , \652 , \653 ,
         \654 , \655 , \656 , \657 , \658 , \659 , \660 , \661 , \662 , \663 ,
         \664 , \665 , \666 , \667 , \668 , \669 , \670 , \671 , \672 , \673 ,
         \674 , \675 , \676 , \677 , \678 , \679 , \680 , \681 , \682 , \683 ,
         \684 , \685 , \686 , \687 , \688 , \689 , \690 , \691 , \692 , \693 ,
         \694 , \695 , \696 , \697 , \698 , \699 , \700_nG137 , \701 , \702 , \703 ,
         \704 , \705 , \706 , \707 , \708 , \709 , \710 , \711 , \712 , \713 ,
         \714 , \715 , \716 , \717 , \718 , \719 , \720 , \721 , \722 , \723 ,
         \724 , \725 , \726 , \727 , \728 , \729 , \730 , \731 , \732 , \733 ,
         \734 , \735 , \736 , \737 , \738 , \739 , \740 , \741 , \742 , \743 ,
         \744 , \745 , \746 , \747 , \748 , \749 , \750 , \751 , \752 , \753 ,
         \754 , \755 , \756 , \757 , \758 , \759 , \760 , \761 , \762 , \763 ,
         \764 , \765 , \766 , \767 , \768 , \769 , \770 , \771 , \772 , \773 ,
         \774 , \775_nG136 , \776 , \777 , \778 , \779 , \780 , \781 , \782 , \783 ,
         \784 , \785 , \786 , \787 , \788 , \789 , \790 , \791 , \792 , \793 ,
         \794 , \795 , \796 , \797 , \798 , \799 , \800 , \801 , \802 , \803 ,
         \804 , \805 , \806 , \807 , \808 , \809 , \810 , \811 , \812 , \813 ,
         \814 , \815 , \816 , \817 , \818 , \819 , \820 , \821 , \822 , \823 ,
         \824 , \825 , \826 , \827 , \828 , \829 , \830 , \831 , \832 , \833 ,
         \834 , \835 , \836 , \837 , \838_nG135 , \839 , \840 , \841 , \842 , \843 ,
         \844 , \845 , \846 , \847 , \848 , \849 , \850 , \851 , \852 , \853 ,
         \854 , \855 , \856 , \857 , \858 , \859 , \860 , \861 , \862 , \863 ,
         \864 , \865 , \866 , \867 , \868 , \869 , \870 , \871 , \872 , \873 ,
         \874 , \875 , \876 , \877 , \878 , \879 , \880 , \881 , \882 , \883 ,
         \884 , \885 , \886 , \887 , \888 , \889 , \890 , \891 , \892 , \893 ,
         \894 , \895 , \896 , \897 , \898 , \899 , \900 , \901 , \902_nG134 , \903 ,
         \904 , \905 , \906 , \907 , \908 , \909 , \910 , \911 , \912 , \913 ,
         \914 , \915 , \916 , \917 , \918 , \919 , \920 , \921 , \922 , \923 ,
         \924 , \925 , \926 , \927 , \928 , \929 , \930 , \931 , \932 , \933 ,
         \934 , \935 , \936 , \937 , \938 , \939 , \940 , \941 , \942 , \943 ,
         \944 , \945 , \946 , \947 , \948 , \949 , \950 , \951 , \952 , \953 ,
         \954 , \955 , \956 , \957 , \958 , \959 , \960 , \961 , \962 , \963 ,
         \964 , \965 , \966 , \967 , \968 , \969 , \970 , \971 , \972 , \973 ,
         \974 , \975 , \976 , \977 , \978 , \979 , \980 , \981 , \982 , \983 ,
         \984 , \985 , \986 , \987 , \988 , \989 , \990 , \991 , \992 , \993 ,
         \994 , \995 , \996 , \997 , \998 , \999 , \1000 , \1001 , \1002 , \1003 ,
         \1004 , \1005 , \1006 , \1007 , \1008 , \1009 , \1010 , \1011 , \1012 , \1013 ,
         \1014 , \1015 , \1016 , \1017 , \1018 , \1019 , \1020 , \1021 , \1022 , \1023 ,
         \1024 , \1025 , \1026 , \1027 , \1028 , \1029 , \1030 , \1031 , \1032 , \1033 ,
         \1034 , \1035 , \1036 , \1037 , \1038 , \1039 , \1040 , \1041 , \1042 , \1043 ,
         \1044 , \1045 , \1046 , \1047 , \1048 , \1049 , \1050 , \1051 , \1052 , \1053 ,
         \1054 , \1055 , \1056 , \1057 , \1058 , \1059 , \1060 , \1061 , \1062 , \1063 ,
         \1064 , \1065 , \1066 , \1067 , \1068 , \1069 , \1070 , \1071 , \1072 , \1073 ,
         \1074 , \1075 , \1076 , \1077 , \1078 , \1079 , \1080 , \1081 , \1082 , \1083 ,
         \1084 , \1085 , \1086 , \1087 , \1088 , \1089 , \1090 , \1091 , \1092 , \1093 ,
         \1094 , \1095 , \1096 , \1097 , \1098 , \1099 , \1100 , \1101_nG133 , \1102 , \1103 ,
         \1104 , \1105 , \1106 , \1107 , \1108 , \1109 , \1110 , \1111 , \1112 , \1113 ,
         \1114 , \1115 , \1116 , \1117 , \1118 , \1119 , \1120 , \1121 , \1122 , \1123 ,
         \1124 , \1125 , \1126 , \1127 , \1128 , \1129 , \1130 , \1131 , \1132 , \1133 ,
         \1134 , \1135 , \1136 , \1137 , \1138 , \1139 , \1140 , \1141 , \1142 , \1143 ,
         \1144 , \1145 , \1146 , \1147 , \1148 , \1149 , \1150 , \1151 , \1152 , \1153 ,
         \1154 , \1155 , \1156 , \1157 , \1158 , \1159 , \1160 , \1161 , \1162 , \1163 ,
         \1164 , \1165 , \1166 , \1167 , \1168 , \1169 , \1170 , \1171 , \1172 , \1173 ,
         \1174 , \1175 , \1176 , \1177 , \1178 , \1179 , \1180 , \1181 , \1182 , \1183 ,
         \1184 , \1185 , \1186 , \1187 , \1188 , \1189 , \1190_nG132 , \1191 , \1192 , \1193 ,
         \1194 , \1195 , \1196 , \1197 , \1198 , \1199 , \1200 , \1201 , \1202 , \1203 ,
         \1204 , \1205 , \1206 , \1207 , \1208 , \1209 , \1210 , \1211 , \1212 , \1213 ,
         \1214 , \1215 , \1216 , \1217 , \1218 , \1219 , \1220 , \1221 , \1222 , \1223 ,
         \1224 , \1225 , \1226 , \1227 , \1228 , \1229 , \1230 , \1231 , \1232 , \1233 ,
         \1234 , \1235 , \1236 , \1237 , \1238 , \1239 , \1240 , \1241 , \1242 , \1243 ,
         \1244 , \1245 , \1246 , \1247 , \1248 , \1249 , \1250 , \1251 , \1252 , \1253 ,
         \1254 , \1255 , \1256 , \1257 , \1258 , \1259 , \1260 , \1261 , \1262 , \1263 ,
         \1264 , \1265 , \1266 , \1267 , \1268 , \1269 , \1270 , \1271 , \1272 , \1273 ,
         \1274 , \1275 , \1276 , \1277 , \1278 , \1279 , \1280 , \1281 , \1282 , \1283 ,
         \1284 , \1285 , \1286 , \1287 , \1288 , \1289 , \1290 , \1291 , \1292 , \1293 ,
         \1294 , \1295 , \1296_nG131 , \1297 , \1298 , \1299 , \1300 , \1301 , \1302_nG130 , \1303 ,
         \1304 , \1305 , \1306 , \1307 , \1308 , \1309 , \1310 , \1311 , \1312 , \1313 ,
         \1314 , \1315 , \1316 , \1317 , \1318 , \1319 , \1320 , \1321 , \1322 , \1323 ,
         \1324 , \1325 , \1326 , \1327 , \1328 , \1329 , \1330 , \1331 , \1332 , \1333 ,
         \1334 , \1335 , \1336 , \1337 , \1338 , \1339 , \1340 , \1341 , \1342 , \1343 ,
         \1344 , \1345 , \1346 , \1347 , \1348 , \1349 , \1350 , \1351 , \1352 , \1353 ,
         \1354 , \1355 , \1356 , \1357 , \1358 , \1359 , \1360 , \1361 , \1362 , \1363 ,
         \1364 , \1365 , \1366 , \1367 , \1368 , \1369 , \1370 , \1371 , \1372 , \1373 ,
         \1374 , \1375 , \1376 , \1377 , \1378 , \1379 , \1380 , \1381 , \1382 , \1383 ,
         \1384 , \1385 , \1386 , \1387 , \1388 , \1389 , \1390 , \1391 , \1392 , \1393 ,
         \1394 , \1395 , \1396 , \1397 , \1398 , \1399 , \1400 , \1401 , \1402 , \1403 ,
         \1404 , \1405 , \1406 , \1407 , \1408 , \1409 , \1410 , \1411 , \1412 , \1413 ,
         \1414 , \1415 , \1416 , \1417 , \1418 , \1419_nG12f , \1420 , \1421 , \1422 , \1423 ,
         \1424 , \1425 , \1426 , \1427 , \1428 , \1429 , \1430 , \1431 , \1432 , \1433 ,
         \1434 , \1435 , \1436 , \1437 , \1438 , \1439 , \1440 , \1441 , \1442 , \1443 ,
         \1444 , \1445 , \1446 , \1447 , \1448 , \1449 , \1450 , \1451 , \1452 , \1453 ,
         \1454 , \1455 , \1456 , \1457 , \1458 , \1459 , \1460 , \1461 , \1462 , \1463 ,
         \1464 , \1465 , \1466 , \1467 , \1468 , \1469 , \1470 , \1471 , \1472 , \1473 ,
         \1474 , \1475 , \1476 , \1477 , \1478 , \1479 , \1480 , \1481 , \1482 , \1483 ,
         \1484 , \1485 , \1486 , \1487 , \1488 , \1489 , \1490 , \1491 , \1492 , \1493 ,
         \1494 , \1495 , \1496 , \1497 , \1498 , \1499 , \1500 , \1501 , \1502 , \1503 ,
         \1504 , \1505 , \1506 , \1507 , \1508 , \1509 , \1510 , \1511 , \1512 , \1513 ,
         \1514 , \1515 , \1516 , \1517 , \1518 , \1519 , \1520 , \1521 , \1522 , \1523 ,
         \1524 , \1525 , \1526 , \1527 , \1528 , \1529 , \1530 , \1531 , \1532 , \1533 ,
         \1534 , \1535_nG12e , \1536 , \1537 , \1538 , \1539 , \1540 , \1541 , \1542 , \1543 ,
         \1544 , \1545 , \1546 , \1547 , \1548 , \1549 , \1550 , \1551 , \1552 , \1553 ,
         \1554 , \1555 , \1556 , \1557 , \1558 , \1559 , \1560 , \1561 , \1562 , \1563 ,
         \1564 , \1565 , \1566 , \1567 , \1568 , \1569 , \1570 , \1571 , \1572 , \1573 ,
         \1574 , \1575 , \1576 , \1577 , \1578 , \1579 , \1580 , \1581 , \1582 , \1583 ,
         \1584 , \1585 , \1586 , \1587 , \1588 , \1589 , \1590 , \1591 , \1592 , \1593 ,
         \1594 , \1595 , \1596 , \1597 , \1598 , \1599 , \1600 , \1601 , \1602 , \1603 ,
         \1604 , \1605 , \1606 , \1607 , \1608 , \1609 , \1610 , \1611 , \1612 , \1613 ,
         \1614 , \1615 , \1616 , \1617 , \1618 , \1619 , \1620 , \1621 , \1622 , \1623 ,
         \1624 , \1625 , \1626 , \1627 , \1628 , \1629 , \1630 , \1631 , \1632 , \1633 ,
         \1634 , \1635 , \1636 , \1637 , \1638 , \1639 , \1640 , \1641 , \1642 , \1643 ,
         \1644 , \1645 , \1646 , \1647 , \1648 , \1649 , \1650 , \1651 , \1652 , \1653 ,
         \1654 , \1655 , \1656 , \1657 , \1658 , \1659 , \1660 , \1661 , \1662 , \1663 ,
         \1664 , \1665 , \1666 , \1667 , \1668 , \1669 , \1670 , \1671 , \1672 , \1673 ,
         \1674 , \1675 , \1676 , \1677 , \1678 , \1679 , \1680 , \1681 , \1682 , \1683 ,
         \1684 , \1685 , \1686 , \1687 , \1688 , \1689 , \1690 , \1691 , \1692 , \1693 ,
         \1694 , \1695 , \1696 , \1697 , \1698 , \1699 , \1700 , \1701 , \1702 , \1703 ,
         \1704 , \1705 , \1706 , \1707 , \1708 , \1709 , \1710 , \1711 , \1712 , \1713 ,
         \1714 , \1715 , \1716 , \1717 , \1718 , \1719 , \1720 , \1721 , \1722 , \1723 ,
         \1724 , \1725 , \1726 , \1727 , \1728 , \1729 , \1730 , \1731 , \1732 , \1733 ,
         \1734 , \1735 , \1736 , \1737 , \1738 , \1739 , \1740 , \1741 , \1742 , \1743 ,
         \1744 , \1745 , \1746 , \1747 , \1748 , \1749 , \1750 , \1751 , \1752 , \1753 ,
         \1754 , \1755 , \1756 , \1757 , \1758 , \1759 , \1760 , \1761 , \1762 , \1763 ,
         \1764 , \1765 , \1766 , \1767_nG12d , \1768 , \1769 , \1770 , \1771 , \1772 , \1773 ,
         \1774 , \1775 , \1776_nG12c , \1777 , \1778 , \1779 , \1780 , \1781 , \1782 , \1783 ,
         \1784 , \1785 , \1786 , \1787 , \1788 , \1789 , \1790 , \1791 , \1792 , \1793 ,
         \1794 , \1795 , \1796 , \1797 , \1798 , \1799 , \1800 , \1801 , \1802 , \1803 ,
         \1804 , \1805 , \1806 , \1807 , \1808 , \1809 , \1810 , \1811 , \1812 , \1813 ,
         \1814 , \1815 , \1816 , \1817 , \1818 , \1819 , \1820 , \1821 , \1822 , \1823 ,
         \1824 , \1825 , \1826 , \1827 , \1828 , \1829 , \1830 , \1831 , \1832 , \1833 ,
         \1834 , \1835 , \1836 , \1837 , \1838 , \1839 , \1840 , \1841 , \1842 , \1843 ,
         \1844 , \1845 , \1846 , \1847 , \1848 , \1849 , \1850 , \1851 , \1852 , \1853 ,
         \1854 , \1855 , \1856 , \1857 , \1858 , \1859 , \1860 , \1861 , \1862 , \1863 ,
         \1864 , \1865 , \1866 , \1867 , \1868 , \1869 , \1870 , \1871 , \1872 , \1873 ,
         \1874 , \1875 , \1876 , \1877 , \1878 , \1879 , \1880 , \1881 , \1882 , \1883 ,
         \1884 , \1885 , \1886 , \1887 , \1888 , \1889 , \1890 , \1891 , \1892 , \1893 ,
         \1894 , \1895 , \1896 , \1897 , \1898 , \1899 , \1900 , \1901 , \1902 , \1903 ,
         \1904 , \1905 , \1906 , \1907 , \1908 , \1909 , \1910 , \1911 , \1912 , \1913 ,
         \1914 , \1915 , \1916 , \1917 , \1918 , \1919 , \1920 , \1921 , \1922 , \1923 ,
         \1924 , \1925 , \1926 , \1927 , \1928 , \1929 , \1930 , \1931 , \1932 , \1933 ,
         \1934 , \1935 , \1936 , \1937 , \1938 , \1939 , \1940 , \1941 , \1942 , \1943 ,
         \1944 , \1945 , \1946 , \1947 , \1948 , \1949 , \1950 , \1951 , \1952 , \1953 ,
         \1954 , \1955 , \1956 , \1957 , \1958 , \1959 , \1960 , \1961 , \1962 , \1963 ,
         \1964 , \1965 , \1966 , \1967 , \1968 , \1969 , \1970 , \1971 , \1972 , \1973 ,
         \1974 , \1975 , \1976 , \1977 , \1978 , \1979 , \1980 , \1981 , \1982 , \1983 ,
         \1984 , \1985 , \1986 , \1987 , \1988 , \1989 , \1990 , \1991 , \1992 , \1993 ,
         \1994 , \1995 , \1996 , \1997 , \1998 , \1999 , \2000 , \2001 , \2002 , \2003 ,
         \2004 , \2005 , \2006 , \2007 , \2008 , \2009 , \2010 , \2011 , \2012 , \2013 ,
         \2014 , \2015 , \2016 , \2017 , \2018 , \2019 , \2020_nG12b , \2021 , \2022 , \2023 ,
         \2024 , \2025 , \2026_nG12a , \2027 , \2028 , \2029 , \2030 , \2031 , \2032 , \2033 ,
         \2034 , \2035 , \2036 , \2037 , \2038 , \2039 , \2040 , \2041 , \2042 , \2043 ,
         \2044 , \2045 , \2046 , \2047 , \2048 , \2049 , \2050 , \2051 , \2052 , \2053 ,
         \2054 , \2055 , \2056 , \2057 , \2058 , \2059 , \2060 , \2061 , \2062 , \2063 ,
         \2064 , \2065 , \2066 , \2067 , \2068 , \2069 , \2070 , \2071 , \2072 , \2073 ,
         \2074 , \2075 , \2076 , \2077 , \2078 , \2079 , \2080 , \2081 , \2082 , \2083 ,
         \2084 , \2085 , \2086 , \2087 , \2088 , \2089 , \2090 , \2091 , \2092 , \2093 ,
         \2094 , \2095 , \2096 , \2097 , \2098 , \2099 , \2100 , \2101 , \2102 , \2103 ,
         \2104 , \2105 , \2106 , \2107 , \2108 , \2109 , \2110 , \2111 , \2112 , \2113 ,
         \2114 , \2115 , \2116 , \2117 , \2118 , \2119 , \2120 , \2121 , \2122 , \2123 ,
         \2124 , \2125 , \2126 , \2127 , \2128 , \2129 , \2130 , \2131 , \2132 , \2133 ,
         \2134 , \2135 , \2136 , \2137 , \2138 , \2139 , \2140 , \2141 , \2142 , \2143 ,
         \2144 , \2145 , \2146 , \2147 , \2148 , \2149 , \2150 , \2151 , \2152 , \2153 ,
         \2154 , \2155 , \2156 , \2157 , \2158_nG129 , \2159 , \2160 , \2161 , \2162 , \2163 ,
         \2164 , \2165 , \2166 , \2167 , \2168 , \2169 , \2170 , \2171 , \2172 , \2173 ,
         \2174 , \2175 , \2176 , \2177 , \2178 , \2179 , \2180 , \2181 , \2182 , \2183 ,
         \2184 , \2185 , \2186 , \2187 , \2188 , \2189 , \2190 , \2191 , \2192 , \2193 ,
         \2194 , \2195 , \2196 , \2197 , \2198 , \2199 , \2200 , \2201 , \2202 , \2203 ,
         \2204 , \2205 , \2206 , \2207 , \2208 , \2209 , \2210 , \2211 , \2212 , \2213 ,
         \2214 , \2215 , \2216 , \2217 , \2218 , \2219 , \2220 , \2221 , \2222 , \2223 ,
         \2224 , \2225 , \2226 , \2227 , \2228 , \2229 , \2230 , \2231 , \2232 , \2233 ,
         \2234 , \2235 , \2236 , \2237 , \2238 , \2239 , \2240 , \2241 , \2242 , \2243 ,
         \2244 , \2245 , \2246 , \2247 , \2248 , \2249 , \2250 , \2251 , \2252 , \2253 ,
         \2254 , \2255 , \2256 , \2257 , \2258 , \2259 , \2260 , \2261 , \2262 , \2263 ,
         \2264 , \2265 , \2266 , \2267 , \2268 , \2269 , \2270 , \2271 , \2272 , \2273 ,
         \2274 , \2275 , \2276 , \2277 , \2278 , \2279 , \2280 , \2281 , \2282 , \2283 ,
         \2284 , \2285 , \2286 , \2287 , \2288 , \2289 , \2290 , \2291 , \2292 , \2293 ,
         \2294 , \2295 , \2296 , \2297 , \2298 , \2299 , \2300 , \2301 , \2302 , \2303_nG128 ,
         \2304 , \2305 , \2306 , \2307 , \2308 , \2309 , \2310 , \2311 , \2312 , \2313 ,
         \2314 , \2315 , \2316 , \2317 , \2318 , \2319 , \2320 , \2321 , \2322 , \2323 ,
         \2324 , \2325 , \2326 , \2327 , \2328 , \2329 , \2330 , \2331 , \2332 , \2333 ,
         \2334 , \2335 , \2336 , \2337 , \2338 , \2339 , \2340 , \2341 , \2342 , \2343 ,
         \2344 , \2345 , \2346 , \2347 , \2348 , \2349 , \2350 , \2351 , \2352 , \2353 ,
         \2354 , \2355 , \2356 , \2357 , \2358 , \2359 , \2360 , \2361 , \2362 , \2363 ,
         \2364 , \2365 , \2366 , \2367 , \2368 , \2369 , \2370 , \2371 , \2372 , \2373 ,
         \2374 , \2375 , \2376 , \2377 , \2378 , \2379 , \2380 , \2381 , \2382 , \2383 ,
         \2384 , \2385 , \2386 , \2387 , \2388 , \2389 , \2390 , \2391 , \2392 , \2393 ,
         \2394 , \2395 , \2396 , \2397 , \2398 , \2399 , \2400 , \2401 , \2402 , \2403 ,
         \2404 , \2405 , \2406 , \2407 , \2408 , \2409 , \2410 , \2411 , \2412 , \2413 ,
         \2414 , \2415 , \2416 , \2417 , \2418 , \2419 , \2420 , \2421 , \2422 , \2423 ,
         \2424 , \2425 , \2426 , \2427 , \2428 , \2429 , \2430 , \2431 , \2432 , \2433 ,
         \2434 , \2435 , \2436 , \2437 , \2438 , \2439 , \2440 , \2441 , \2442 , \2443 ,
         \2444 , \2445 , \2446 , \2447 , \2448 , \2449 , \2450 , \2451 , \2452 , \2453 ,
         \2454 , \2455 , \2456 , \2457 , \2458 , \2459 , \2460 , \2461 , \2462 , \2463 ,
         \2464 , \2465 , \2466 , \2467 , \2468 , \2469 , \2470 , \2471 , \2472 , \2473 ,
         \2474 , \2475 , \2476 , \2477 , \2478 , \2479 , \2480 , \2481 , \2482 , \2483 ,
         \2484 , \2485 , \2486 , \2487 , \2488 , \2489 , \2490 , \2491 , \2492 , \2493 ,
         \2494 , \2495 , \2496 , \2497 , \2498 , \2499 , \2500 , \2501 , \2502 , \2503 ,
         \2504 , \2505 , \2506 , \2507 , \2508 , \2509 , \2510 , \2511 , \2512 , \2513 ,
         \2514 , \2515 , \2516 , \2517 , \2518 , \2519 , \2520 , \2521 , \2522 , \2523 ,
         \2524 , \2525 , \2526 , \2527 , \2528 , \2529_nG127 , \2530 , \2531 , \2532 , \2533 ,
         \2534 , \2535 , \2536 , \2537 , \2538 , \2539_nG126 , \2540 , \2541 , \2542 , \2543 ,
         \2544 , \2545 , \2546 , \2547 , \2548 , \2549 , \2550 , \2551 , \2552 , \2553 ,
         \2554 , \2555 , \2556 , \2557 , \2558 , \2559 , \2560 , \2561 , \2562 , \2563 ,
         \2564 , \2565 , \2566 , \2567 , \2568 , \2569 , \2570 , \2571 , \2572 , \2573 ,
         \2574 , \2575 , \2576 , \2577 , \2578 , \2579 , \2580 , \2581 , \2582 , \2583 ,
         \2584 , \2585 , \2586 , \2587 , \2588 , \2589 , \2590 , \2591 , \2592 , \2593 ,
         \2594 , \2595 , \2596 , \2597 , \2598 , \2599 , \2600 , \2601 , \2602 , \2603 ,
         \2604 , \2605 , \2606 , \2607 , \2608 , \2609 , \2610 , \2611 , \2612 , \2613 ,
         \2614 , \2615 , \2616 , \2617 , \2618 , \2619 , \2620 , \2621 , \2622 , \2623 ,
         \2624 , \2625 , \2626 , \2627 , \2628 , \2629 , \2630 , \2631 , \2632 , \2633 ,
         \2634 , \2635 , \2636 , \2637 , \2638 , \2639 , \2640 , \2641 , \2642 , \2643 ,
         \2644 , \2645 , \2646 , \2647 , \2648 , \2649 , \2650 , \2651 , \2652 , \2653 ,
         \2654 , \2655 , \2656 , \2657 , \2658 , \2659 , \2660 , \2661 , \2662 , \2663 ,
         \2664 , \2665 , \2666 , \2667 , \2668 , \2669 , \2670 , \2671 , \2672 , \2673 ,
         \2674 , \2675 , \2676 , \2677 , \2678 , \2679 , \2680 , \2681 , \2682 , \2683 ,
         \2684 , \2685 , \2686 , \2687 , \2688 , \2689 , \2690 , \2691 , \2692 , \2693 ,
         \2694 , \2695 , \2696 , \2697 , \2698 , \2699 , \2700 , \2701 , \2702 , \2703 ,
         \2704 , \2705 , \2706 , \2707 , \2708 , \2709 , \2710 , \2711 , \2712 , \2713 ,
         \2714 , \2715 , \2716 , \2717 , \2718 , \2719 , \2720 , \2721 , \2722 , \2723 ,
         \2724 , \2725 , \2726 , \2727 , \2728 , \2729 , \2730 , \2731 , \2732 , \2733 ,
         \2734 , \2735 , \2736 , \2737 , \2738 , \2739 , \2740 , \2741 , \2742 , \2743 ,
         \2744 , \2745 , \2746 , \2747 , \2748 , \2749 , \2750 , \2751 , \2752 , \2753 ,
         \2754 , \2755 , \2756 , \2757 , \2758 , \2759 , \2760 , \2761 , \2762_nG125 , \2763 ,
         \2764 , \2765 , \2766 , \2767 , \2768 , \2769 , \2770 , \2771 , \2772 , \2773 ,
         \2774 , \2775 , \2776 , \2777 , \2778 , \2779 , \2780 , \2781 , \2782 , \2783 ,
         \2784 , \2785 , \2786 , \2787 , \2788 , \2789 , \2790 , \2791 , \2792 , \2793 ,
         \2794 , \2795 , \2796 , \2797 , \2798 , \2799 , \2800 , \2801 , \2802 , \2803 ,
         \2804 , \2805 , \2806 , \2807 , \2808 , \2809 , \2810 , \2811 , \2812 , \2813 ,
         \2814 , \2815 , \2816 , \2817 , \2818 , \2819 , \2820 , \2821 , \2822 , \2823 ,
         \2824 , \2825 , \2826 , \2827 , \2828 , \2829 , \2830 , \2831 , \2832 , \2833 ,
         \2834 , \2835 , \2836 , \2837 , \2838 , \2839 , \2840 , \2841 , \2842 , \2843 ,
         \2844 , \2845 , \2846 , \2847 , \2848 , \2849 , \2850_nG124 , \2851 , \2852 , \2853 ,
         \2854 , \2855 , \2856 , \2857 , \2858 , \2859 , \2860 , \2861 , \2862 , \2863 ,
         \2864 , \2865 , \2866 , \2867 , \2868 , \2869 , \2870 , \2871 , \2872 , \2873 ,
         \2874 , \2875 , \2876 , \2877 , \2878 , \2879 , \2880 , \2881 , \2882 , \2883 ,
         \2884 , \2885 , \2886 , \2887 , \2888 , \2889 , \2890 , \2891 , \2892 , \2893 ,
         \2894 , \2895 , \2896 , \2897 , \2898 , \2899 , \2900 , \2901 , \2902 , \2903 ,
         \2904 , \2905 , \2906 , \2907 , \2908 , \2909 , \2910 , \2911 , \2912 , \2913 ,
         \2914 , \2915 , \2916 , \2917 , \2918 , \2919 , \2920 , \2921 , \2922 , \2923 ,
         \2924 , \2925 , \2926 , \2927 , \2928 , \2929 , \2930 , \2931 , \2932 , \2933 ,
         \2934 , \2935 , \2936 , \2937 , \2938 , \2939 , \2940 , \2941 , \2942 , \2943 ,
         \2944 , \2945 , \2946 , \2947 , \2948 , \2949 , \2950 , \2951 , \2952 , \2953 ,
         \2954 , \2955 , \2956 , \2957 , \2958 , \2959 , \2960 , \2961 , \2962 , \2963 ,
         \2964 , \2965 , \2966 , \2967 , \2968 , \2969 , \2970 , \2971 , \2972 , \2973 ,
         \2974 , \2975 , \2976 , \2977 , \2978 , \2979 , \2980 , \2981 , \2982 , \2983 ,
         \2984 , \2985 , \2986 , \2987 , \2988 , \2989 , \2990 , \2991 , \2992 , \2993 ,
         \2994 , \2995 , \2996 , \2997 , \2998 , \2999 , \3000 , \3001 , \3002 , \3003 ,
         \3004 , \3005 , \3006 , \3007 , \3008 , \3009 , \3010 , \3011 , \3012 , \3013 ,
         \3014 , \3015 , \3016 , \3017 , \3018 , \3019 , \3020 , \3021 , \3022 , \3023 ,
         \3024 , \3025 , \3026 , \3027 , \3028 , \3029 , \3030 , \3031 , \3032 , \3033 ,
         \3034 , \3035 , \3036 , \3037 , \3038 , \3039 , \3040 , \3041 , \3042 , \3043 ,
         \3044 , \3045 , \3046 , \3047 , \3048 , \3049 , \3050 , \3051 , \3052 , \3053 ,
         \3054 , \3055 , \3056 , \3057 , \3058 , \3059 , \3060 , \3061 , \3062 , \3063 ,
         \3064 , \3065 , \3066 , \3067 , \3068 , \3069 , \3070 , \3071 , \3072 , \3073 ,
         \3074 , \3075 , \3076 , \3077 , \3078 , \3079 , \3080 , \3081 , \3082 , \3083 ,
         \3084 , \3085 , \3086 , \3087 , \3088 , \3089 , \3090 , \3091 , \3092 , \3093 ,
         \3094 , \3095 , \3096 , \3097 , \3098 , \3099 , \3100 , \3101 , \3102 , \3103 ,
         \3104 , \3105 , \3106 , \3107 , \3108 , \3109 , \3110 , \3111 , \3112 , \3113 ,
         \3114 , \3115 , \3116 , \3117 , \3118 , \3119 , \3120 , \3121 , \3122 , \3123 ,
         \3124 , \3125 , \3126 , \3127 , \3128 , \3129 , \3130 , \3131 , \3132 , \3133 ,
         \3134 , \3135 , \3136 , \3137 , \3138 , \3139 , \3140 , \3141 , \3142 , \3143 ,
         \3144 , \3145 , \3146 , \3147 , \3148 , \3149 , \3150 , \3151 , \3152 , \3153 ,
         \3154 , \3155 , \3156 , \3157 , \3158 , \3159 , \3160 , \3161 , \3162 , \3163 ,
         \3164 , \3165 , \3166 , \3167 , \3168 , \3169 , \3170 , \3171 , \3172 , \3173 ,
         \3174 , \3175 , \3176 , \3177 , \3178 , \3179 , \3180 , \3181 , \3182 , \3183 ,
         \3184 , \3185 , \3186 , \3187 , \3188 , \3189 , \3190 , \3191 , \3192 , \3193 ,
         \3194 , \3195 , \3196 , \3197 , \3198 , \3199 , \3200 , \3201 , \3202 , \3203 ,
         \3204 , \3205 , \3206 , \3207 , \3208 , \3209 , \3210 , \3211 , \3212 , \3213 ,
         \3214 , \3215 , \3216 , \3217 , \3218 , \3219 , \3220 , \3221 , \3222 , \3223 ,
         \3224 , \3225 , \3226 , \3227 , \3228 , \3229 , \3230 , \3231 , \3232 , \3233 ,
         \3234 , \3235 , \3236 , \3237 , \3238 , \3239 , \3240 , \3241 , \3242 , \3243 ,
         \3244 , \3245 , \3246 , \3247 , \3248 , \3249 , \3250 , \3251 , \3252 , \3253 ,
         \3254 , \3255 , \3256 , \3257 , \3258 , \3259 , \3260 , \3261 , \3262 , \3263 ,
         \3264 , \3265 , \3266 , \3267 , \3268 , \3269 , \3270 , \3271 , \3272 , \3273 ,
         \3274 , \3275 , \3276 , \3277 , \3278 , \3279 , \3280 , \3281 , \3282 , \3283 ,
         \3284 , \3285 , \3286 , \3287 , \3288 , \3289 , \3290 , \3291 , \3292 , \3293 ,
         \3294 , \3295 , \3296 , \3297 , \3298 , \3299 , \3300 , \3301 , \3302 , \3303 ,
         \3304 , \3305 , \3306 , \3307 , \3308 , \3309 , \3310 , \3311 , \3312 , \3313 ,
         \3314 , \3315 , \3316 , \3317 , \3318 , \3319 , \3320 , \3321 , \3322 , \3323 ,
         \3324 , \3325 , \3326 , \3327 , \3328 , \3329 , \3330 , \3331 , \3332 , \3333 ,
         \3334 , \3335 , \3336 , \3337 , \3338 , \3339 , \3340 , \3341 , \3342 , \3343 ,
         \3344 , \3345 , \3346 , \3347 , \3348 , \3349 , \3350 , \3351 , \3352 , \3353 ,
         \3354 , \3355 , \3356 , \3357 , \3358 , \3359 , \3360 , \3361 , \3362 , \3363 ,
         \3364 , \3365 , \3366 , \3367 , \3368 , \3369 , \3370 , \3371 , \3372 , \3373 ,
         \3374 , \3375 , \3376 , \3377 , \3378 , \3379 , \3380 , \3381 , \3382 , \3383 ,
         \3384 , \3385 , \3386 , \3387 , \3388 , \3389 , \3390 , \3391 , \3392 , \3393 ,
         \3394 , \3395 , \3396 , \3397 , \3398 , \3399 , \3400 , \3401 , \3402 , \3403 ,
         \3404 , \3405 , \3406 , \3407 , \3408 , \3409 , \3410 , \3411 , \3412 , \3413 ,
         \3414 , \3415 , \3416 , \3417 , \3418 , \3419 , \3420 , \3421 , \3422 , \3423 ,
         \3424 , \3425 , \3426 , \3427 , \3428 , \3429 , \3430 , \3431 , \3432 , \3433 ,
         \3434 , \3435 , \3436 , \3437 , \3438 , \3439 , \3440 , \3441 , \3442 , \3443 ,
         \3444 , \3445 , \3446 , \3447 , \3448 , \3449 , \3450 , \3451 , \3452 , \3453 ,
         \3454 , \3455 , \3456 , \3457 , \3458 , \3459 , \3460 , \3461 , \3462 , \3463 ,
         \3464 , \3465 , \3466 , \3467 , \3468 , \3469 , \3470 , \3471 , \3472 , \3473 ,
         \3474 , \3475 , \3476 , \3477 , \3478 , \3479 , \3480 , \3481 , \3482 , \3483 ,
         \3484 , \3485 , \3486 , \3487 , \3488 , \3489 , \3490 , \3491 , \3492 , \3493 ,
         \3494 , \3495 , \3496 , \3497 , \3498 , \3499 , \3500 , \3501 , \3502 , \3503 ,
         \3504 , \3505 , \3506 , \3507 , \3508 , \3509 , \3510 , \3511 , \3512 , \3513 ,
         \3514 , \3515 , \3516 , \3517 , \3518 , \3519 , \3520 , \3521 , \3522 , \3523 ,
         \3524 , \3525 , \3526 , \3527 , \3528 , \3529 , \3530 , \3531 , \3532 , \3533 ,
         \3534 , \3535 , \3536 , \3537 , \3538 , \3539 , \3540 , \3541 , \3542 , \3543 ,
         \3544 , \3545 , \3546 , \3547 , \3548 , \3549 , \3550 , \3551 , \3552 , \3553 ,
         \3554 , \3555 , \3556 , \3557 , \3558 , \3559 , \3560 , \3561 , \3562 , \3563 ,
         \3564 , \3565 , \3566 , \3567 , \3568 , \3569 , \3570 , \3571 , \3572 , \3573 ,
         \3574 , \3575 , \3576 , \3577 , \3578 , \3579 , \3580 , \3581 , \3582 , \3583 ,
         \3584 , \3585 , \3586 , \3587 , \3588 , \3589 , \3590 , \3591 , \3592 , \3593 ,
         \3594 , \3595 , \3596 , \3597 , \3598 , \3599 , \3600 , \3601 , \3602 , \3603 ,
         \3604 , \3605 , \3606 , \3607 , \3608 , \3609 , \3610 , \3611 , \3612 , \3613 ,
         \3614 , \3615 , \3616 , \3617 , \3618 , \3619 , \3620 , \3621 , \3622 , \3623 ,
         \3624 , \3625 , \3626 , \3627 , \3628 , \3629 , \3630 , \3631 , \3632 , \3633 ,
         \3634 , \3635 , \3636 , \3637 , \3638 , \3639 , \3640 , \3641 , \3642 , \3643 ,
         \3644 , \3645 , \3646 , \3647 , \3648 , \3649 , \3650 , \3651 , \3652 , \3653 ,
         \3654 , \3655 , \3656 , \3657 , \3658 , \3659 , \3660 , \3661 , \3662 , \3663 ,
         \3664 , \3665 , \3666 , \3667 , \3668 , \3669 , \3670 , \3671 , \3672 , \3673 ,
         \3674 , \3675 , \3676 , \3677 , \3678 , \3679 , \3680 , \3681 , \3682 , \3683 ,
         \3684 , \3685 , \3686 , \3687 , \3688 , \3689 , \3690 , \3691 , \3692 , \3693 ,
         \3694 , \3695 , \3696 , \3697 , \3698 , \3699 , \3700 , \3701 , \3702 , \3703 ,
         \3704 , \3705 , \3706 , \3707 , \3708 , \3709 , \3710 , \3711 , \3712 , \3713 ,
         \3714 , \3715 , \3716 , \3717 , \3718 , \3719 , \3720 , \3721 , \3722 , \3723 ,
         \3724 , \3725 , \3726 , \3727 , \3728 , \3729 , \3730 , \3731 , \3732 , \3733 ,
         \3734 , \3735 , \3736 , \3737 , \3738 , \3739 , \3740 , \3741 , \3742 , \3743 ,
         \3744 , \3745 , \3746 , \3747 , \3748 , \3749 , \3750 , \3751 , \3752 , \3753 ,
         \3754 , \3755 , \3756 , \3757 , \3758 , \3759 , \3760 , \3761 , \3762 , \3763 ,
         \3764 , \3765 , \3766 , \3767 , \3768 , \3769 , \3770 , \3771 , \3772 , \3773 ,
         \3774 , \3775 , \3776 , \3777 , \3778 , \3779 , \3780 , \3781 , \3782 , \3783 ,
         \3784 , \3785 , \3786 , \3787 , \3788 , \3789 , \3790 , \3791 , \3792 , \3793 ,
         \3794 , \3795 , \3796 , \3797 , \3798 , \3799 , \3800 , \3801 , \3802 , \3803 ,
         \3804 , \3805 , \3806 , \3807 , \3808 , \3809 , \3810 , \3811 , \3812 , \3813 ,
         \3814 , \3815 , \3816 , \3817 , \3818 , \3819 , \3820 , \3821 , \3822 , \3823 ,
         \3824 , \3825 , \3826 , \3827 , \3828 , \3829 , \3830 , \3831 , \3832 , \3833 ,
         \3834 , \3835 , \3836 , \3837 , \3838 , \3839 , \3840 , \3841 , \3842 , \3843 ,
         \3844 , \3845 , \3846 , \3847 , \3848 , \3849 , \3850 , \3851 , \3852 , \3853 ,
         \3854 , \3855 , \3856 , \3857 , \3858 , \3859 , \3860 , \3861 , \3862 , \3863 ,
         \3864 , \3865 , \3866 , \3867 , \3868 , \3869 , \3870 , \3871 , \3872 , \3873 ,
         \3874 , \3875 , \3876 , \3877 , \3878 , \3879 , \3880 , \3881 , \3882 , \3883 ,
         \3884 , \3885 , \3886 , \3887 , \3888 , \3889 , \3890 , \3891 , \3892 , \3893 ,
         \3894 , \3895 , \3896 , \3897 , \3898 , \3899 , \3900 , \3901 , \3902 , \3903 ,
         \3904 , \3905 , \3906 , \3907 , \3908 , \3909 , \3910 , \3911 , \3912 , \3913 ,
         \3914 , \3915 , \3916 , \3917 , \3918 , \3919 , \3920 , \3921 , \3922 , \3923 ,
         \3924 , \3925 , \3926 , \3927 , \3928 , \3929 , \3930 , \3931 , \3932 , \3933 ,
         \3934 , \3935 , \3936 , \3937 , \3938 , \3939 , \3940 , \3941 , \3942 , \3943 ,
         \3944 , \3945 , \3946 , \3947 , \3948 , \3949 , \3950 , \3951 , \3952 , \3953 ,
         \3954 , \3955 , \3956 , \3957 , \3958 , \3959 , \3960 , \3961 , \3962 , \3963 ,
         \3964 , \3965 , \3966 , \3967 , \3968 , \3969 , \3970 , \3971 , \3972 , \3973 ,
         \3974 , \3975 , \3976 , \3977 , \3978 , \3979 , \3980 , \3981 , \3982 , \3983 ,
         \3984 , \3985 , \3986 , \3987 , \3988 , \3989 , \3990 , \3991 , \3992 , \3993 ,
         \3994 , \3995 , \3996 , \3997 , \3998 , \3999 , \4000 , \4001 , \4002 , \4003 ,
         \4004 , \4005 , \4006 , \4007 , \4008 , \4009 , \4010 , \4011 , \4012 , \4013 ,
         \4014 , \4015 , \4016 , \4017 , \4018 , \4019 , \4020 , \4021 , \4022 , \4023 ,
         \4024 , \4025 , \4026 , \4027 , \4028 , \4029 , \4030 , \4031 , \4032 , \4033 ,
         \4034 , \4035 , \4036 , \4037 , \4038 , \4039 , \4040 , \4041 , \4042 , \4043 ,
         \4044 , \4045 , \4046 , \4047 , \4048 , \4049 , \4050 , \4051 , \4052 , \4053 ,
         \4054 , \4055 , \4056 , \4057 , \4058 , \4059 , \4060 , \4061 , \4062 , \4063 ,
         \4064 , \4065 , \4066 , \4067 , \4068 , \4069 , \4070 , \4071 , \4072 , \4073 ,
         \4074 , \4075 , \4076 , \4077 , \4078 , \4079 , \4080 , \4081 , \4082 , \4083 ,
         \4084 , \4085 , \4086 , \4087 , \4088 , \4089 , \4090 , \4091 , \4092 , \4093 ,
         \4094 , \4095 , \4096 , \4097 , \4098 , \4099 , \4100 , \4101 , \4102 , \4103 ,
         \4104 , \4105 , \4106 , \4107 , \4108 , \4109 , \4110 , \4111 , \4112 , \4113 ,
         \4114 , \4115 , \4116 , \4117 , \4118 , \4119 , \4120 , \4121 , \4122 , \4123 ,
         \4124 , \4125 , \4126 , \4127 , \4128 , \4129 , \4130 , \4131 , \4132 , \4133 ,
         \4134 , \4135 , \4136 , \4137 , \4138 , \4139 , \4140 , \4141 , \4142 , \4143 ,
         \4144 , \4145 , \4146 , \4147 , \4148 , \4149 , \4150 , \4151 , \4152 , \4153 ,
         \4154 , \4155 , \4156 , \4157 , \4158 , \4159 , \4160 , \4161 , \4162 , \4163 ,
         \4164 , \4165 , \4166 , \4167 , \4168 , \4169 , \4170 , \4171 , \4172 , \4173 ,
         \4174 , \4175 , \4176 , \4177 , \4178 , \4179 , \4180 , \4181 , \4182 , \4183 ,
         \4184 , \4185 , \4186 , \4187 , \4188 , \4189 , \4190 , \4191 , \4192 , \4193 ,
         \4194 , \4195 , \4196 , \4197 , \4198 , \4199 , \4200 , \4201 , \4202 , \4203 ,
         \4204 , \4205 , \4206 , \4207 , \4208 , \4209 , \4210 , \4211 , \4212 , \4213 ,
         \4214 , \4215 , \4216 , \4217 , \4218 , \4219 , \4220 , \4221 , \4222 , \4223 ,
         \4224 , \4225 , \4226 , \4227 , \4228 , \4229 , \4230 , \4231 , \4232 , \4233 ,
         \4234 , \4235 , \4236 , \4237 , \4238 , \4239 , \4240 , \4241 , \4242 , \4243 ,
         \4244 , \4245 , \4246 , \4247 , \4248 , \4249 , \4250 , \4251 , \4252 , \4253 ,
         \4254 , \4255 , \4256 , \4257 , \4258 , \4259 , \4260 , \4261 , \4262 , \4263 ,
         \4264 , \4265 , \4266 , \4267 , \4268 , \4269 , \4270 , \4271 , \4272 , \4273 ,
         \4274 , \4275 , \4276 , \4277 , \4278 , \4279 , \4280 , \4281 , \4282 , \4283 ,
         \4284 , \4285 , \4286 , \4287 , \4288 , \4289 , \4290 , \4291 , \4292 , \4293 ,
         \4294 , \4295 , \4296 , \4297 , \4298 , \4299 , \4300 , \4301 , \4302 , \4303 ,
         \4304 , \4305 , \4306 , \4307 , \4308 , \4309 , \4310 , \4311 , \4312 , \4313 ,
         \4314 , \4315 , \4316 , \4317 , \4318 , \4319 , \4320 , \4321 , \4322 , \4323 ,
         \4324 , \4325 , \4326 , \4327 , \4328 , \4329 , \4330 , \4331 , \4332 , \4333 ,
         \4334 , \4335 , \4336 , \4337 , \4338 , \4339 , \4340 , \4341 , \4342 , \4343 ,
         \4344 , \4345 , \4346 , \4347 , \4348 , \4349 , \4350 , \4351 , \4352 , \4353 ,
         \4354 , \4355 , \4356 , \4357 , \4358 , \4359 , \4360 , \4361 , \4362 , \4363 ,
         \4364 , \4365 , \4366 , \4367 , \4368 , \4369 , \4370 , \4371 , \4372 , \4373 ,
         \4374 , \4375 , \4376 , \4377 , \4378 , \4379 , \4380 , \4381 , \4382 , \4383 ,
         \4384 , \4385 , \4386 , \4387 , \4388 , \4389 , \4390 , \4391 , \4392 , \4393 ,
         \4394 , \4395 , \4396 , \4397 , \4398 , \4399 , \4400 , \4401 , \4402 , \4403 ,
         \4404 , \4405 , \4406 , \4407 , \4408 , \4409 , \4410 , \4411 , \4412 , \4413 ,
         \4414 , \4415 , \4416 , \4417 , \4418 , \4419 , \4420 , \4421 , \4422 , \4423 ,
         \4424 , \4425 , \4426 , \4427 , \4428 , \4429 , \4430 , \4431 , \4432 , \4433 ,
         \4434 , \4435 , \4436 , \4437 , \4438 , \4439 , \4440 , \4441 , \4442 , \4443 ,
         \4444 , \4445 , \4446 , \4447 , \4448 , \4449 , \4450 , \4451 , \4452 , \4453 ,
         \4454 , \4455 , \4456 , \4457 , \4458 , \4459 , \4460 , \4461 , \4462 , \4463 ,
         \4464 , \4465 , \4466 , \4467 , \4468 , \4469 , \4470 , \4471 , \4472 , \4473 ,
         \4474 , \4475 , \4476 , \4477 , \4478 , \4479 , \4480 , \4481 , \4482 , \4483 ,
         \4484 , \4485 , \4486 , \4487 , \4488 , \4489 , \4490 , \4491 , \4492 , \4493 ,
         \4494 , \4495 , \4496 , \4497 , \4498 , \4499 , \4500 , \4501 , \4502 , \4503 ,
         \4504 , \4505 , \4506 , \4507 , \4508 , \4509 , \4510 , \4511 , \4512 , \4513 ,
         \4514 , \4515 , \4516 , \4517 , \4518 , \4519 , \4520 , \4521 , \4522 , \4523 ,
         \4524 , \4525 , \4526 , \4527 , \4528 , \4529 , \4530 , \4531 , \4532 , \4533 ,
         \4534 , \4535 , \4536 , \4537 , \4538 , \4539 , \4540 , \4541 , \4542 , \4543 ,
         \4544 , \4545 , \4546 , \4547 , \4548 , \4549 , \4550 , \4551 , \4552 , \4553 ,
         \4554 , \4555 , \4556 , \4557 , \4558 , \4559 , \4560 , \4561 , \4562 , \4563 ,
         \4564 , \4565 , \4566 , \4567 , \4568 , \4569 , \4570 , \4571 , \4572 , \4573 ,
         \4574 , \4575 , \4576 , \4577 , \4578 , \4579 , \4580 , \4581 , \4582 , \4583 ,
         \4584 , \4585 , \4586 , \4587 , \4588 , \4589 , \4590 , \4591 , \4592 , \4593 ,
         \4594 , \4595 , \4596 , \4597 , \4598 , \4599 , \4600 , \4601 , \4602 , \4603 ,
         \4604 , \4605 , \4606 , \4607 , \4608 , \4609 , \4610 , \4611 , \4612 , \4613 ,
         \4614 , \4615 , \4616 , \4617 , \4618 , \4619 , \4620 , \4621 , \4622 , \4623 ,
         \4624 , \4625 , \4626 , \4627 , \4628 , \4629 , \4630 , \4631 , \4632 , \4633 ,
         \4634 , \4635 , \4636 , \4637 , \4638 , \4639 , \4640 , \4641 , \4642 , \4643 ,
         \4644 , \4645 , \4646 , \4647 , \4648 , \4649 , \4650 , \4651 , \4652 , \4653 ,
         \4654 , \4655 , \4656 , \4657 , \4658 , \4659 , \4660 , \4661 , \4662 , \4663 ,
         \4664 , \4665 , \4666 , \4667 , \4668 , \4669 , \4670 , \4671 , \4672 , \4673 ,
         \4674 , \4675 , \4676 , \4677 , \4678 , \4679 , \4680 , \4681 , \4682 , \4683 ,
         \4684 , \4685 , \4686 , \4687 , \4688 , \4689 , \4690 , \4691 , \4692 , \4693 ,
         \4694 , \4695 , \4696 , \4697 , \4698 , \4699 , \4700 , \4701 , \4702 , \4703 ,
         \4704 , \4705 , \4706 , \4707 , \4708 , \4709 , \4710 , \4711 , \4712 , \4713 ,
         \4714 , \4715 , \4716 , \4717 , \4718 , \4719 , \4720 , \4721 , \4722 , \4723 ,
         \4724 , \4725 , \4726 , \4727 , \4728 , \4729 , \4730 , \4731 , \4732 , \4733 ,
         \4734 , \4735 , \4736 , \4737 , \4738 , \4739 , \4740 , \4741 , \4742 , \4743 ,
         \4744 , \4745 , \4746 , \4747 , \4748 , \4749 , \4750 , \4751 , \4752 , \4753 ,
         \4754 , \4755 , \4756 , \4757 , \4758 , \4759 , \4760 , \4761 , \4762 , \4763 ,
         \4764 , \4765 , \4766 , \4767 , \4768 , \4769 , \4770 , \4771 , \4772 , \4773 ,
         \4774 , \4775 , \4776 , \4777 , \4778 , \4779 , \4780 , \4781 , \4782 , \4783 ,
         \4784 , \4785 , \4786 , \4787 , \4788 , \4789 , \4790 , \4791 , \4792 , \4793 ,
         \4794 , \4795 , \4796 , \4797 , \4798 , \4799 , \4800 , \4801 , \4802 , \4803 ,
         \4804 , \4805 , \4806 , \4807 , \4808 , \4809 , \4810 , \4811 , \4812 , \4813 ,
         \4814 , \4815 , \4816 , \4817 , \4818 , \4819 , \4820 , \4821 , \4822 , \4823 ,
         \4824 , \4825 , \4826 , \4827 , \4828 , \4829 , \4830 , \4831 , \4832 , \4833 ,
         \4834 , \4835 , \4836 , \4837 , \4838 , \4839 , \4840 , \4841 , \4842 , \4843 ,
         \4844 , \4845 , \4846 , \4847 , \4848 , \4849 , \4850 , \4851 , \4852 , \4853 ,
         \4854 , \4855 , \4856 , \4857 , \4858 , \4859 , \4860 , \4861 , \4862 , \4863 ,
         \4864 , \4865 , \4866 , \4867 , \4868 , \4869 , \4870 , \4871 , \4872 , \4873 ,
         \4874 , \4875 , \4876 , \4877 , \4878 , \4879 , \4880 , \4881 , \4882 , \4883 ,
         \4884 , \4885 , \4886 , \4887 , \4888 , \4889 , \4890 , \4891 , \4892 , \4893 ,
         \4894 , \4895 , \4896 , \4897 , \4898 , \4899 , \4900 , \4901 , \4902 , \4903 ,
         \4904 , \4905 , \4906 , \4907 , \4908 , \4909 , \4910 , \4911 , \4912 , \4913 ,
         \4914 , \4915 , \4916 , \4917 , \4918 , \4919 , \4920 , \4921 , \4922 , \4923 ,
         \4924 , \4925 , \4926 , \4927 , \4928 , \4929 , \4930 , \4931 , \4932 , \4933 ,
         \4934 , \4935 , \4936 , \4937 , \4938 , \4939 , \4940 , \4941 , \4942 , \4943 ,
         \4944 , \4945 , \4946 , \4947 , \4948 , \4949 , \4950 , \4951 , \4952 , \4953 ,
         \4954 , \4955 , \4956 , \4957 , \4958 , \4959 , \4960 , \4961 , \4962 , \4963 ,
         \4964 , \4965 , \4966 , \4967 , \4968 , \4969 , \4970 , \4971 , \4972 , \4973 ,
         \4974 , \4975 , \4976 , \4977 , \4978 , \4979 , \4980 , \4981 , \4982 , \4983 ,
         \4984 , \4985 , \4986 , \4987 , \4988 , \4989 , \4990 , \4991 , \4992 , \4993 ,
         \4994 , \4995 , \4996 , \4997 , \4998 , \4999 , \5000 , \5001 , \5002 , \5003 ,
         \5004 , \5005 , \5006 , \5007 , \5008 , \5009 , \5010 , \5011 , \5012 , \5013 ,
         \5014 , \5015 , \5016 , \5017 , \5018 , \5019 , \5020 , \5021 , \5022 , \5023 ,
         \5024 , \5025 , \5026 , \5027 , \5028 , \5029 , \5030 , \5031 , \5032 , \5033 ,
         \5034 , \5035 , \5036 , \5037 , \5038 , \5039 , \5040 , \5041 , \5042 , \5043 ,
         \5044 , \5045 , \5046 , \5047 , \5048 , \5049 , \5050 , \5051 , \5052 , \5053 ,
         \5054 , \5055 , \5056 , \5057 , \5058 , \5059 , \5060 , \5061 , \5062 , \5063 ,
         \5064 , \5065 , \5066 , \5067 , \5068 , \5069 , \5070 , \5071 , \5072 , \5073 ,
         \5074 , \5075 , \5076 , \5077 , \5078 , \5079 , \5080 , \5081 , \5082 , \5083 ,
         \5084 , \5085 , \5086 , \5087 , \5088 , \5089 , \5090 , \5091 , \5092 , \5093 ,
         \5094 , \5095 , \5096 , \5097 , \5098 , \5099 , \5100 , \5101 , \5102 , \5103 ,
         \5104 , \5105 , \5106 , \5107 , \5108 , \5109 , \5110 , \5111 , \5112 , \5113 ,
         \5114 , \5115 , \5116 , \5117 , \5118 , \5119 , \5120 , \5121 , \5122 , \5123 ,
         \5124 , \5125 , \5126 , \5127 , \5128 , \5129 , \5130 , \5131 , \5132 , \5133 ,
         \5134 , \5135 , \5136 , \5137 , \5138 , \5139 , \5140 , \5141 , \5142 , \5143 ,
         \5144 , \5145 , \5146 , \5147 , \5148 , \5149 , \5150 , \5151 , \5152 , \5153 ,
         \5154 , \5155 , \5156 , \5157 , \5158 , \5159 , \5160 , \5161 , \5162 , \5163 ,
         \5164 , \5165 , \5166 , \5167 , \5168 , \5169 , \5170 , \5171 , \5172 , \5173 ,
         \5174 , \5175 , \5176 , \5177 , \5178 , \5179 , \5180 , \5181 , \5182 , \5183 ,
         \5184 , \5185 , \5186 , \5187 , \5188 , \5189 , \5190 , \5191 , \5192 , \5193 ,
         \5194 , \5195 , \5196 , \5197 , \5198 , \5199 , \5200 , \5201 , \5202 , \5203 ,
         \5204 , \5205 , \5206 , \5207 , \5208 , \5209 , \5210 , \5211 , \5212 , \5213 ,
         \5214 , \5215 , \5216 , \5217 , \5218 , \5219 , \5220 , \5221 , \5222 , \5223 ,
         \5224 , \5225 , \5226 , \5227 , \5228 , \5229 , \5230 , \5231 , \5232 , \5233 ,
         \5234 , \5235 , \5236 , \5237 , \5238 , \5239 , \5240 , \5241 , \5242 , \5243 ,
         \5244 , \5245 , \5246 , \5247 , \5248 , \5249 , \5250 , \5251 , \5252 , \5253 ,
         \5254 , \5255 , \5256 , \5257 , \5258 , \5259 , \5260 , \5261 , \5262 , \5263 ,
         \5264 , \5265 , \5266 , \5267 , \5268 , \5269 , \5270 , \5271 , \5272 , \5273 ,
         \5274 , \5275 , \5276 , \5277 , \5278 , \5279 , \5280 , \5281 , \5282 , \5283 ,
         \5284 , \5285 , \5286 , \5287 , \5288 , \5289 , \5290 , \5291 , \5292 , \5293 ,
         \5294 , \5295 , \5296 , \5297 , \5298 , \5299 , \5300 , \5301 , \5302 , \5303 ,
         \5304 , \5305 , \5306 , \5307 , \5308 , \5309 , \5310 , \5311 , \5312 , \5313 ,
         \5314 , \5315 , \5316 , \5317 , \5318 , \5319 , \5320 , \5321 , \5322 , \5323 ,
         \5324 , \5325 , \5326 , \5327 , \5328 , \5329 , \5330 , \5331 , \5332 , \5333 ,
         \5334 , \5335 , \5336 , \5337 , \5338 , \5339 , \5340 , \5341 , \5342 , \5343 ,
         \5344 , \5345 , \5346 , \5347 , \5348 , \5349 , \5350 , \5351 , \5352 , \5353 ,
         \5354 , \5355 , \5356 , \5357 , \5358 , \5359 , \5360 , \5361 , \5362 , \5363 ,
         \5364 , \5365 , \5366 , \5367 , \5368 , \5369 , \5370 , \5371 , \5372 , \5373 ,
         \5374 , \5375 , \5376 , \5377 , \5378 , \5379 , \5380 , \5381 , \5382 , \5383 ,
         \5384 , \5385 , \5386 , \5387 , \5388 , \5389 , \5390 , \5391 , \5392 , \5393 ,
         \5394 , \5395 , \5396 , \5397 , \5398 , \5399 , \5400 , \5401 , \5402 , \5403 ,
         \5404 , \5405 , \5406 , \5407 , \5408 , \5409 , \5410 , \5411 , \5412 , \5413 ,
         \5414 , \5415 , \5416 , \5417 , \5418 , \5419 , \5420 , \5421 , \5422 , \5423 ,
         \5424 , \5425 , \5426 , \5427 , \5428 , \5429 , \5430 , \5431 , \5432 , \5433 ,
         \5434 , \5435 , \5436 , \5437 , \5438 , \5439 , \5440 , \5441 , \5442 , \5443 ,
         \5444 , \5445 , \5446 , \5447 , \5448 , \5449 , \5450 , \5451 , \5452 , \5453 ,
         \5454 , \5455 , \5456 , \5457 , \5458 , \5459 , \5460 , \5461 , \5462 , \5463 ,
         \5464 , \5465 , \5466 , \5467 , \5468 , \5469 , \5470 , \5471 , \5472 , \5473 ,
         \5474 , \5475 , \5476 , \5477 , \5478 , \5479 , \5480 , \5481 , \5482 , \5483 ,
         \5484 , \5485 , \5486 , \5487 , \5488 , \5489 , \5490 , \5491 , \5492 , \5493 ,
         \5494 , \5495 , \5496 , \5497 , \5498 , \5499 , \5500 , \5501 , \5502 , \5503 ,
         \5504 , \5505 , \5506 , \5507 , \5508 , \5509 , \5510 , \5511 , \5512 , \5513 ,
         \5514 , \5515 , \5516 , \5517 , \5518 , \5519 , \5520 , \5521 , \5522 , \5523 ,
         \5524 , \5525 , \5526 , \5527 , \5528 , \5529 , \5530 , \5531 , \5532 , \5533 ,
         \5534 , \5535 , \5536 , \5537 , \5538 , \5539 , \5540 , \5541 , \5542 , \5543 ,
         \5544 , \5545 , \5546 , \5547 , \5548 , \5549 , \5550 , \5551 , \5552 , \5553 ,
         \5554 , \5555 , \5556 , \5557 , \5558 , \5559 , \5560 , \5561 , \5562 , \5563 ,
         \5564 , \5565 , \5566 , \5567 , \5568 , \5569 , \5570 , \5571 , \5572 , \5573 ,
         \5574 , \5575 , \5576 , \5577 , \5578 , \5579 , \5580 , \5581 , \5582 , \5583 ,
         \5584 , \5585 , \5586 , \5587 , \5588 , \5589 , \5590 , \5591 , \5592 , \5593 ,
         \5594 , \5595 , \5596 , \5597 , \5598 , \5599 , \5600 , \5601 , \5602 , \5603 ,
         \5604 , \5605 , \5606 , \5607 , \5608 , \5609 , \5610 , \5611 , \5612 , \5613 ,
         \5614 , \5615 , \5616 , \5617 , \5618 , \5619 , \5620 , \5621 , \5622 , \5623 ,
         \5624 , \5625 , \5626 , \5627 , \5628 , \5629 , \5630 , \5631 , \5632 , \5633 ,
         \5634 , \5635 , \5636 , \5637 , \5638 , \5639 , \5640 , \5641 , \5642 , \5643 ,
         \5644 , \5645 , \5646 , \5647 , \5648 , \5649 , \5650 , \5651 , \5652 , \5653 ,
         \5654 , \5655 , \5656 , \5657 , \5658 , \5659 , \5660 , \5661 , \5662 , \5663 ,
         \5664 , \5665 , \5666 , \5667 , \5668 , \5669 , \5670 , \5671 , \5672 , \5673 ,
         \5674 , \5675 , \5676 , \5677 , \5678 , \5679 , \5680 , \5681 , \5682 , \5683 ,
         \5684 , \5685 , \5686 , \5687 , \5688 , \5689 , \5690 , \5691 , \5692 , \5693 ,
         \5694 , \5695 , \5696 , \5697 , \5698 , \5699 , \5700 , \5701 , \5702 , \5703 ,
         \5704 , \5705 , \5706 , \5707 , \5708 , \5709 , \5710 , \5711 , \5712 , \5713 ,
         \5714 , \5715 , \5716 , \5717 , \5718 , \5719 , \5720 , \5721 , \5722 , \5723 ,
         \5724 , \5725 , \5726_nG16bf , \5727 , \5728 , \5729_nG16c2 , \5730 , \5731 , \5732_nG16c5 , \5733 ,
         \5734 , \5735 , \5736 , \5737 , \5738 , \5739_nG171f , \5740 , \5741 , \5742_nG1722 , \5743 ,
         \5744 , \5745 , \5746_nG1725 , \5747 , \5748 , \5749 , \5750 , \5751 , \5752 , \5753 ,
         \5754 , \5755 , \5756 , \5757 , \5758 , \5759 , \5760_nG1719 , \5761 , \5762 , \5763_nG171c ,
         \5764 , \5765 , \5766 , \5767 , \5768 , \5769 , \5770 , \5771 , \5772 , \5773 ,
         \5774 , \5775 , \5776 , \5777 , \5778 , \5779 , \5780 , \5781 , \5782_nG1713 , \5783 ,
         \5784 , \5785_nG1716 , \5786 , \5787 , \5788 , \5789 , \5790 , \5791 , \5792 , \5793 ,
         \5794 , \5795 , \5796 , \5797 , \5798 , \5799 , \5800 , \5801_nG170d , \5802 , \5803 ,
         \5804_nG1710 , \5805 , \5806 , \5807 , \5808 , \5809 , \5810 , \5811 , \5812 , \5813 ,
         \5814 , \5815 , \5816 , \5817 , \5818 , \5819 , \5820 , \5821_nG1707 , \5822 , \5823 ,
         \5824_nG170a , \5825 , \5826 , \5827 , \5828 , \5829 , \5830 , \5831 , \5832 , \5833 ,
         \5834 , \5835 , \5836 , \5837 , \5838 , \5839 , \5840 , \5841 , \5842 , \5843 ,
         \5844_nG1701 , \5845 , \5846 , \5847_nG1704 , \5848 , \5849 , \5850 , \5851 , \5852 , \5853 ,
         \5854 , \5855 , \5856 , \5857 , \5858 , \5859 , \5860 , \5861 , \5862 , \5863_nG16fb ,
         \5864 , \5865 , \5866_nG16fe , \5867 , \5868 , \5869 , \5870 , \5871 , \5872 , \5873 ,
         \5874 , \5875 , \5876 , \5877 , \5878 , \5879 , \5880 , \5881 , \5882 , \5883_nG16f5 ,
         \5884 , \5885 , \5886_nG16f8 , \5887 , \5888 , \5889 , \5890 , \5891 , \5892 , \5893 ,
         \5894 , \5895 , \5896 , \5897 , \5898 , \5899 , \5900 , \5901 , \5902 , \5903 ,
         \5904 , \5905 , \5906 , \5907 , \5908_nG16ef , \5909 , \5910 , \5911_nG16f2 , \5912 , \5913 ,
         \5914 , \5915 , \5916 , \5917 , \5918 , \5919 , \5920 , \5921 , \5922 , \5923 ,
         \5924 , \5925 , \5926 , \5927_nG16e9 , \5928 , \5929 , \5930_nG16ec , \5931 , \5932 , \5933 ,
         \5934 , \5935 , \5936 , \5937 , \5938 , \5939 , \5940 , \5941 , \5942 , \5943 ,
         \5944 , \5945 , \5946 , \5947_nG16e3 , \5948 , \5949 , \5950_nG16e6 , \5951 , \5952 , \5953 ,
         \5954 , \5955 , \5956 , \5957 , \5958 , \5959 , \5960 , \5961 , \5962 , \5963 ,
         \5964 , \5965 , \5966 , \5967 , \5968 , \5969_nG16dd , \5970 , \5971 , \5972_nG16e0 , \5973 ,
         \5974 , \5975 , \5976 , \5977 , \5978 , \5979 , \5980 , \5981 , \5982 , \5983 ,
         \5984 , \5985 , \5986 , \5987 , \5988_nG16d7 , \5989 , \5990 , \5991_nG16da , \5992 , \5993 ,
         \5994 , \5995 , \5996 , \5997 , \5998 , \5999 , \6000 , \6001 , \6002 , \6003 ,
         \6004 , \6005 , \6006 , \6007 , \6008_nG16d1 , \6009 , \6010 , \6011_nG16d4 , \6012 , \6013 ,
         \6014 , \6015 , \6016 , \6017 , \6018 , \6019 , \6020 , \6021 , \6022 , \6023 ,
         \6024 , \6025 , \6026 , \6027 , \6028 , \6029 , \6030 , \6031_nG16cb , \6032 , \6033 ,
         \6034_nG16ce , \6035 , \6036 , \6037 , \6038 , \6039 , \6040 , \6041 , \6042 , \6043 ,
         \6044 , \6045 , \6046 , \6047 , \6048 , \6049 , \6050_nG16c8 , \6051 , \6052 , \6053 ,
         \6054 , \6055 , \6056 , \6057 , \6058 , \6059 , \6060 , \6061 , \6062 , \6063 ,
         \6064 , \6065 , \6066 , \6067 , \6068 , \6069 , \6070 , \6071 , \6072 , \6073 ,
         \6074 , \6075 , \6076 , \6077 , \6078 , \6079 , \6080 , \6081 , \6082 , \6083 ,
         \6084 , \6085 , \6086 , \6087 , \6088 , \6089 , \6090 , \6091 , \6092 , \6093 ,
         \6094 , \6095 , \6096 , \6097 , \6098 , \6099 , \6100 , \6101 , \6102 , \6103 ,
         \6104 , \6105 , \6106 , \6107 , \6108 , \6109 , \6110 , \6111 , \6112 , \6113 ,
         \6114 , \6115 , \6116 , \6117 , \6118 , \6119 , \6120 , \6121 , \6122 , \6123 ,
         \6124 , \6125 , \6126 , \6127 , \6128 , \6129 , \6130 , \6131 , \6132 , \6133 ,
         \6134 , \6135 , \6136 , \6137 , \6138 , \6139 , \6140 , \6141 , \6142 , \6143 ,
         \6144 , \6145 , \6146 , \6147 , \6148 , \6149 , \6150 , \6151 , \6152 , \6153 ,
         \6154 , \6155 , \6156 , \6157 , \6158 , \6159 , \6160 , \6161 , \6162 , \6163 ,
         \6164 , \6165 , \6166 , \6167 , \6168 , \6169 , \6170 , \6171 , \6172 , \6173 ,
         \6174 , \6175 , \6176 , \6177 , \6178 , \6179 , \6180 , \6181 , \6182 , \6183 ,
         \6184 , \6185 , \6186 , \6187 , \6188 , \6189 , \6190 , \6191 , \6192 , \6193 ,
         \6194 , \6195 , \6196 , \6197 , \6198 , \6199 , \6200 , \6201 , \6202 , \6203 ,
         \6204 , \6205 , \6206 , \6207 , \6208 , \6209 , \6210 , \6211 , \6212 , \6213 ,
         \6214 , \6215 , \6216 , \6217 , \6218 , \6219 , \6220_nG16b9 , \6221 , \6222 , \6223_nG16bc ,
         \6224 , \6225 , \6226 , \6227 , \6228 , \6229 , \6230 , \6231 , \6232 , \6233 ,
         \6234 , \6235 , \6236 , \6237 , \6238 , \6239 , \6240 , \6241 , \6242 , \6243 ,
         \6244 , \6245 , \6246 , \6247 , \6248 , \6249 , \6250 , \6251 , \6252 , \6253 ,
         \6254 , \6255 , \6256 , \6257 , \6258 , \6259 , \6260 , \6261 , \6262 , \6263 ,
         \6264 , \6265 , \6266 , \6267 , \6268 , \6269 , \6270 , \6271 , \6272 , \6273 ,
         \6274 , \6275 , \6276 , \6277 , \6278 , \6279 , \6280 , \6281 , \6282 , \6283 ,
         \6284 , \6285 , \6286 , \6287 , \6288 , \6289 , \6290 , \6291 , \6292 , \6293 ,
         \6294 , \6295 , \6296 , \6297 , \6298 , \6299 , \6300 , \6301 , \6302 , \6303 ,
         \6304 , \6305 , \6306 , \6307 , \6308 , \6309 , \6310 , \6311 , \6312 , \6313 ,
         \6314 , \6315 , \6316 , \6317 , \6318 , \6319 , \6320 , \6321 , \6322 , \6323 ,
         \6324 , \6325 , \6326 , \6327 , \6328 , \6329 , \6330 , \6331 , \6332 , \6333 ,
         \6334 , \6335 , \6336 , \6337 , \6338 , \6339 , \6340 , \6341 , \6342 , \6343 ,
         \6344 , \6345 , \6346 , \6347 , \6348 , \6349 , \6350 , \6351 , \6352 , \6353 ,
         \6354 , \6355 , \6356 , \6357 , \6358 , \6359 , \6360 , \6361 , \6362 , \6363 ,
         \6364 , \6365 , \6366 , \6367 , \6368 , \6369 , \6370 , \6371 , \6372 , \6373 ,
         \6374 , \6375 , \6376 , \6377 , \6378 , \6379 , \6380 , \6381 , \6382 , \6383 ,
         \6384 , \6385 , \6386 , \6387 , \6388 , \6389 , \6390 , \6391 , \6392 , \6393 ,
         \6394 , \6395 , \6396 , \6397 , \6398 , \6399 , \6400 , \6401 , \6402 , \6403 ,
         \6404 , \6405 , \6406 , \6407 , \6408 , \6409 , \6410 , \6411 , \6412 , \6413 ,
         \6414 , \6415 , \6416 , \6417 , \6418 , \6419 , \6420 , \6421 , \6422 , \6423 ,
         \6424 , \6425 , \6426 , \6427 , \6428 , \6429 , \6430 , \6431 , \6432 , \6433 ,
         \6434 , \6435 , \6436 , \6437 , \6438 , \6439 , \6440 , \6441 , \6442 , \6443 ,
         \6444 , \6445 , \6446 , \6447 , \6448 , \6449 , \6450 , \6451 , \6452 , \6453 ,
         \6454 , \6455 , \6456 , \6457 , \6458 , \6459 , \6460 , \6461 , \6462 , \6463 ,
         \6464 , \6465 , \6466 , \6467 , \6468 , \6469 , \6470 , \6471 , \6472 , \6473 ,
         \6474 , \6475 , \6476 , \6477 , \6478 , \6479 , \6480 , \6481 , \6482 , \6483 ,
         \6484 , \6485 , \6486 , \6487 , \6488 , \6489 , \6490 , \6491 , \6492 , \6493 ,
         \6494 , \6495 , \6496 , \6497 , \6498 , \6499 , \6500 , \6501 , \6502 , \6503 ,
         \6504 , \6505 , \6506 , \6507 , \6508_nG16b6 , \6509 , \6510 , \6511 , \6512 , \6513 ,
         \6514 , \6515 , \6516 , \6517 , \6518 , \6519 , \6520 , \6521 , \6522 , \6523_nG16b3 ,
         \6524 , \6525 , \6526 , \6527 , \6528 , \6529 , \6530 , \6531 , \6532 , \6533 ,
         \6534 , \6535 , \6536 , \6537 , \6538 , \6539 , \6540 , \6541 , \6542 , \6543 ,
         \6544 , \6545 , \6546 , \6547 , \6548 , \6549 , \6550 , \6551 , \6552 , \6553 ,
         \6554 , \6555 , \6556 , \6557 , \6558 , \6559 , \6560 , \6561 , \6562 , \6563 ,
         \6564 , \6565 , \6566 , \6567 , \6568 , \6569 , \6570 , \6571 , \6572 , \6573 ,
         \6574 , \6575 , \6576 , \6577 , \6578 , \6579 , \6580 , \6581 , \6582 , \6583 ,
         \6584 , \6585 , \6586 , \6587 , \6588 , \6589 , \6590 , \6591 , \6592 , \6593 ,
         \6594 , \6595 , \6596 , \6597 , \6598 , \6599 , \6600 , \6601 , \6602 , \6603 ,
         \6604 , \6605 , \6606 , \6607 , \6608 , \6609 , \6610 , \6611 , \6612 , \6613 ,
         \6614 , \6615 , \6616 , \6617 , \6618 , \6619 , \6620 , \6621 , \6622 , \6623 ,
         \6624 , \6625 , \6626 , \6627 , \6628 , \6629 , \6630 , \6631 , \6632 , \6633 ,
         \6634 , \6635 , \6636 , \6637 , \6638 , \6639 , \6640 , \6641 , \6642 , \6643 ,
         \6644 , \6645 , \6646 , \6647 , \6648 , \6649 , \6650 , \6651 , \6652 , \6653 ,
         \6654 , \6655 , \6656 , \6657 , \6658 , \6659 , \6660 , \6661 , \6662 , \6663 ,
         \6664 , \6665 , \6666 , \6667 , \6668 , \6669 , \6670 , \6671 , \6672 , \6673 ,
         \6674 , \6675 , \6676 , \6677 , \6678 , \6679 , \6680 , \6681 , \6682 , \6683 ,
         \6684 , \6685 , \6686 , \6687 , \6688 , \6689 , \6690 , \6691 , \6692 , \6693 ,
         \6694 , \6695 , \6696 , \6697 , \6698 , \6699 , \6700 , \6701 , \6702 , \6703 ,
         \6704 , \6705 , \6706 , \6707 , \6708 , \6709 , \6710 , \6711 , \6712 , \6713 ,
         \6714 , \6715 , \6716 , \6717 , \6718 , \6719 , \6720 , \6721 , \6722 , \6723 ,
         \6724 , \6725 , \6726 , \6727 , \6728 , \6729 , \6730 , \6731 , \6732 , \6733 ,
         \6734 , \6735 , \6736 , \6737 , \6738 , \6739 , \6740 , \6741 , \6742 , \6743 ,
         \6744 , \6745 , \6746 , \6747 , \6748 , \6749 , \6750 , \6751 , \6752 , \6753 ,
         \6754 , \6755 , \6756 , \6757 , \6758 , \6759 , \6760 , \6761 , \6762 , \6763 ,
         \6764 , \6765 , \6766 , \6767 , \6768 , \6769 , \6770 , \6771 , \6772 , \6773 ,
         \6774 , \6775 , \6776 , \6777 , \6778 , \6779 , \6780 , \6781 , \6782 , \6783 ,
         \6784 , \6785 , \6786 , \6787 , \6788 , \6789 , \6790 , \6791 , \6792 , \6793 ,
         \6794 , \6795 , \6796 , \6797 , \6798 , \6799 , \6800 , \6801 , \6802 , \6803 ,
         \6804 , \6805 , \6806 , \6807 , \6808 , \6809 , \6810 , \6811 , \6812 , \6813 ,
         \6814 , \6815 , \6816 , \6817_nG1728 , \6818 , \6819 , \6820_nG172b , \6821 , \6822 , \6823 ,
         \6824 , \6825 , \6826 , \6827 , \6828 , \6829 , \6830 , \6831 , \6832 , \6833 ,
         \6834 , \6835 , \6836 , \6837 , \6838 , \6839 , \6840 , \6841 , \6842 , \6843 ,
         \6844 , \6845 , \6846 , \6847 , \6848 , \6849 , \6850 , \6851 , \6852 , \6853 ,
         \6854 , \6855 , \6856 , \6857 , \6858 , \6859 , \6860 , \6861 , \6862 , \6863 ,
         \6864 , \6865 , \6866 , \6867 , \6868 , \6869 , \6870 , \6871 , \6872 , \6873 ,
         \6874 , \6875 , \6876 , \6877 , \6878 , \6879 , \6880 , \6881 , \6882 , \6883 ,
         \6884 , \6885 , \6886 , \6887 , \6888 , \6889 , \6890 , \6891 , \6892 , \6893 ,
         \6894 , \6895 , \6896 , \6897 , \6898 , \6899 , \6900 , \6901 , \6902 , \6903 ,
         \6904 , \6905 , \6906 , \6907 , \6908 , \6909 , \6910 , \6911 , \6912 , \6913 ,
         \6914 , \6915 , \6916 , \6917 , \6918 , \6919 , \6920 , \6921 , \6922 , \6923 ,
         \6924 , \6925 , \6926 , \6927 , \6928 , \6929 , \6930 , \6931 , \6932 , \6933 ,
         \6934 , \6935 , \6936 , \6937 , \6938 , \6939 , \6940 , \6941 , \6942 , \6943 ,
         \6944 , \6945 , \6946 , \6947 , \6948 , \6949 , \6950 , \6951 , \6952 , \6953 ,
         \6954 , \6955 , \6956 , \6957 , \6958 , \6959 , \6960 , \6961 , \6962 , \6963 ,
         \6964 , \6965 , \6966 , \6967 , \6968 , \6969 , \6970 , \6971 , \6972 , \6973 ,
         \6974 , \6975 , \6976 , \6977 , \6978 , \6979 , \6980 , \6981 , \6982 , \6983 ,
         \6984_nG176d , \6985 , \6986 , \6987_nG1770 , \6988 , \6989 , \6990 , \6991 , \6992 , \6993 ,
         \6994 , \6995 , \6996 , \6997 , \6998_nG1767 , \6999 , \7000 , \7001_nG176a , \7002 , \7003 ,
         \7004 , \7005 , \7006 , \7007 , \7008 , \7009 , \7010 , \7011 , \7012 , \7013 ,
         \7014 , \7015 , \7016 , \7017 , \7018_nG1761 , \7019 , \7020 , \7021_nG1764 , \7022 , \7023 ,
         \7024 , \7025 , \7026 , \7027 , \7028 , \7029 , \7030 , \7031 , \7032 , \7033 ,
         \7034 , \7035_nG175b , \7036 , \7037 , \7038_nG175e , \7039 , \7040 , \7041 , \7042 , \7043 ,
         \7044 , \7045 , \7046 , \7047 , \7048 , \7049 , \7050 , \7051 , \7052 , \7053_nG1755 ,
         \7054 , \7055 , \7056_nG1758 , \7057 , \7058 , \7059 , \7060 , \7061 , \7062 , \7063 ,
         \7064 , \7065 , \7066 , \7067 , \7068 , \7069 , \7070 , \7071 , \7072 , \7073 ,
         \7074_nG174f , \7075 , \7076 , \7077_nG1752 , \7078 , \7079 , \7080 , \7081 , \7082 , \7083 ,
         \7084 , \7085 , \7086 , \7087 , \7088 , \7089 , \7090 , \7091_nG1749 , \7092 , \7093 ,
         \7094_nG174c , \7095 , \7096 , \7097 , \7098 , \7099 , \7100 , \7101 , \7102 , \7103 ,
         \7104 , \7105 , \7106 , \7107 , \7108 , \7109_nG1743 , \7110 , \7111 , \7112_nG1746 , \7113 ,
         \7114 , \7115 , \7116 , \7117 , \7118 , \7119 , \7120 , \7121 , \7122 , \7123 ,
         \7124 , \7125 , \7126 , \7127 , \7128 , \7129 , \7130 , \7131 , \7132_nG173d , \7133 ,
         \7134 , \7135_nG1740 , \7136 , \7137 , \7138 , \7139 , \7140 , \7141 , \7142 , \7143 ,
         \7144 , \7145 , \7146 , \7147 , \7148 , \7149_nG1737 , \7150 , \7151 , \7152_nG173a , \7153 ,
         \7154 , \7155 , \7156 , \7157 , \7158 , \7159 , \7160 , \7161 , \7162 , \7163 ,
         \7164 , \7165 , \7166 , \7167_nG1731 , \7168 , \7169 , \7170_nG1734 , \7171 , \7172 , \7173 ,
         \7174 , \7175 , \7176 , \7177 , \7178 , \7179 , \7180 , \7181 , \7182 , \7183 ,
         \7184 , \7185 , \7186 , \7187_nG172e , \7188 , \7189 , \7190 , \7191 , \7192 , \7193 ,
         \7194 , \7195 , \7196 , \7197 , \7198 , \7199 , \7200 , \7201 , \7202 , \7203 ,
         \7204 , \7205 , \7206 , \7207 , \7208 , \7209 , \7210 , \7211 , \7212 , \7213 ,
         \7214 , \7215 , \7216 , \7217 , \7218 , \7219 , \7220 , \7221 , \7222 , \7223 ,
         \7224 , \7225 , \7226 , \7227 , \7228 , \7229 , \7230 , \7231 , \7232 , \7233 ,
         \7234 , \7235 , \7236 , \7237 , \7238 , \7239 , \7240 , \7241 , \7242 , \7243 ,
         \7244 , \7245 , \7246 , \7247 , \7248 , \7249 , \7250 , \7251 , \7252 , \7253 ,
         \7254 , \7255 , \7256 , \7257 , \7258 , \7259 , \7260 , \7261 , \7262 , \7263 ,
         \7264 , \7265 , \7266 , \7267 , \7268 , \7269 , \7270 , \7271 , \7272 , \7273 ,
         \7274 , \7275 , \7276 , \7277 , \7278 , \7279 , \7280 , \7281 , \7282 , \7283 ,
         \7284 , \7285 , \7286 , \7287 , \7288 , \7289 , \7290 , \7291 , \7292 , \7293 ,
         \7294 , \7295 , \7296 , \7297 , \7298 , \7299 , \7300 , \7301 , \7302 , \7303 ,
         \7304 , \7305 , \7306 , \7307 , \7308 , \7309 , \7310 , \7311 , \7312 , \7313 ,
         \7314 , \7315 , \7316 , \7317 , \7318 , \7319 , \7320 , \7321 , \7322 , \7323 ,
         \7324 , \7325 , \7326 , \7327 , \7328 , \7329 , \7330 , \7331 , \7332 , \7333 ,
         \7334 , \7335 , \7336 , \7337 , \7338 , \7339 , \7340 , \7341 , \7342 , \7343 ,
         \7344 , \7345 , \7346 , \7347 , \7348 , \7349 , \7350 , \7351 , \7352 , \7353 ,
         \7354 , \7355 , \7356 , \7357 , \7358 , \7359 , \7360 , \7361 , \7362 , \7363 ,
         \7364 , \7365 , \7366 , \7367 , \7368 , \7369 , \7370 , \7371 , \7372 , \7373 ,
         \7374 , \7375 , \7376 , \7377 , \7378 , \7379 , \7380 , \7381 , \7382 , \7383 ,
         \7384 , \7385 , \7386 , \7387 , \7388 , \7389 , \7390 , \7391 , \7392 , \7393 ,
         \7394 , \7395 , \7396 , \7397 , \7398 , \7399 , \7400 , \7401 , \7402 , \7403 ,
         \7404 , \7405 , \7406 , \7407 , \7408 , \7409 , \7410 , \7411 , \7412 , \7413 ,
         \7414 , \7415 , \7416 , \7417 , \7418 , \7419 , \7420 , \7421 , \7422 , \7423 ,
         \7424 , \7425 , \7426 , \7427 , \7428 , \7429 , \7430 , \7431 , \7432 , \7433 ,
         \7434 , \7435 , \7436 , \7437 , \7438 , \7439 , \7440 , \7441 , \7442 , \7443 ,
         \7444 , \7445 , \7446 , \7447 , \7448 , \7449 , \7450 , \7451 , \7452 , \7453 ,
         \7454 , \7455 , \7456 , \7457 , \7458 , \7459 , \7460 , \7461 , \7462 , \7463 ,
         \7464 , \7465 , \7466 , \7467 , \7468 , \7469 , \7470 , \7471 , \7472 , \7473 ,
         \7474 , \7475 , \7476 , \7477 , \7478 , \7479 , \7480 , \7481 , \7482 , \7483 ,
         \7484 , \7485 , \7486 , \7487 , \7488 , \7489 , \7490 , \7491 , \7492 , \7493 ,
         \7494 , \7495 , \7496 , \7497 , \7498 , \7499 , \7500 , \7501 , \7502 , \7503 ,
         \7504 , \7505 , \7506 , \7507 , \7508 , \7509 , \7510 , \7511 , \7512 , \7513 ,
         \7514 , \7515 , \7516 , \7517 , \7518 , \7519 , \7520 , \7521 , \7522 , \7523 ,
         \7524 , \7525 , \7526 , \7527 , \7528 , \7529 , \7530 , \7531 , \7532 , \7533 ,
         \7534 , \7535 , \7536 , \7537 , \7538 , \7539 , \7540 , \7541 , \7542 , \7543 ,
         \7544 , \7545 , \7546 , \7547 , \7548 , \7549 , \7550 , \7551 , \7552 , \7553 ,
         \7554 , \7555 , \7556 , \7557 , \7558 , \7559 , \7560 , \7561 , \7562 , \7563 ,
         \7564 , \7565 , \7566 , \7567 , \7568 , \7569 , \7570 , \7571 , \7572 , \7573 ,
         \7574 , \7575 , \7576 , \7577 , \7578 , \7579 , \7580 , \7581 , \7582 , \7583 ,
         \7584 , \7585 , \7586 , \7587 , \7588 , \7589 , \7590 , \7591 , \7592 , \7593 ,
         \7594 , \7595 , \7596 , \7597 , \7598 , \7599 , \7600 , \7601 , \7602 , \7603 ,
         \7604 , \7605 , \7606 , \7607 , \7608 , \7609 , \7610 , \7611 , \7612 , \7613 ,
         \7614 , \7615 , \7616 , \7617 , \7618 , \7619 , \7620 , \7621 , \7622 , \7623 ,
         \7624 , \7625 , \7626 , \7627 , \7628 , \7629 , \7630 , \7631 , \7632 , \7633 ,
         \7634 , \7635 , \7636 , \7637 , \7638 , \7639 , \7640 , \7641 , \7642 , \7643 ,
         \7644 , \7645 , \7646 , \7647 , \7648 , \7649 , \7650 , \7651 , \7652 , \7653 ,
         \7654 , \7655 , \7656 , \7657 , \7658 , \7659 , \7660 , \7661 , \7662 , \7663 ,
         \7664 , \7665 , \7666 , \7667 , \7668 , \7669 , \7670 , \7671 , \7672 , \7673 ,
         \7674 , \7675 , \7676 , \7677 , \7678 , \7679 , \7680 , \7681 , \7682 , \7683 ,
         \7684 , \7685 , \7686 , \7687 , \7688 , \7689 , \7690 , \7691 , \7692 , \7693 ,
         \7694 , \7695 , \7696 , \7697 , \7698 , \7699 , \7700 , \7701 , \7702 , \7703 ,
         \7704 , \7705 , \7706 , \7707 , \7708 , \7709 , \7710 , \7711 , \7712 , \7713 ,
         \7714 , \7715 , \7716 , \7717 , \7718 , \7719 , \7720 , \7721 , \7722 , \7723 ,
         \7724 , \7725 , \7726 , \7727 , \7728 , \7729 , \7730 , \7731 , \7732 , \7733 ,
         \7734 , \7735 , \7736 , \7737 , \7738 , \7739 , \7740 , \7741 , \7742 , \7743 ,
         \7744 , \7745 , \7746 , \7747 , \7748 , \7749 , \7750 , \7751 , \7752 , \7753 ,
         \7754 , \7755 , \7756 , \7757 , \7758 , \7759 , \7760 , \7761 , \7762 , \7763 ,
         \7764 , \7765 , \7766 , \7767 , \7768 , \7769 , \7770 , \7771 , \7772 , \7773 ,
         \7774 , \7775 , \7776 , \7777 , \7778 , \7779 , \7780 , \7781 , \7782 , \7783 ,
         \7784 , \7785 , \7786 , \7787 , \7788 , \7789 , \7790 , \7791 , \7792 , \7793 ,
         \7794 , \7795 , \7796 , \7797 , \7798 , \7799 , \7800 , \7801 , \7802 , \7803 ,
         \7804 , \7805 , \7806 , \7807 , \7808 , \7809 , \7810 , \7811 , \7812 , \7813 ,
         \7814 , \7815 , \7816 , \7817 , \7818 , \7819 , \7820 , \7821 , \7822 , \7823 ,
         \7824 , \7825 , \7826 , \7827 , \7828 , \7829 , \7830 , \7831 , \7832 , \7833 ,
         \7834 , \7835 , \7836 , \7837 , \7838 , \7839 , \7840 , \7841 , \7842 , \7843 ,
         \7844 , \7845 , \7846 , \7847 , \7848 , \7849 , \7850 , \7851 , \7852 , \7853 ,
         \7854 , \7855 , \7856 , \7857 , \7858 , \7859 , \7860 , \7861 , \7862 , \7863 ,
         \7864 , \7865 , \7866 , \7867 , \7868 , \7869 , \7870 , \7871 , \7872 , \7873 ,
         \7874 , \7875 , \7876 , \7877 , \7878 , \7879 , \7880 , \7881 , \7882 , \7883 ,
         \7884 , \7885 , \7886 , \7887 , \7888 , \7889 , \7890 , \7891 , \7892 , \7893 ,
         \7894 , \7895 , \7896 , \7897 , \7898 , \7899 , \7900 , \7901 , \7902 , \7903 ,
         \7904 , \7905 , \7906 , \7907 , \7908 , \7909 , \7910 , \7911 , \7912 , \7913 ,
         \7914 , \7915 , \7916 , \7917 , \7918 , \7919 , \7920 , \7921 , \7922 , \7923 ,
         \7924 , \7925 , \7926 , \7927 , \7928 , \7929 , \7930 , \7931 , \7932 , \7933 ,
         \7934 , \7935 , \7936 , \7937 , \7938 , \7939 , \7940 , \7941 , \7942 , \7943 ,
         \7944 , \7945 , \7946 , \7947 , \7948 , \7949 , \7950 , \7951 , \7952 , \7953 ,
         \7954 , \7955 , \7956 , \7957 , \7958 , \7959 , \7960 , \7961 , \7962 , \7963 ,
         \7964 , \7965 , \7966 , \7967 , \7968 , \7969 , \7970 , \7971 , \7972 , \7973 ,
         \7974 , \7975 , \7976 , \7977 , \7978 , \7979 , \7980 , \7981 , \7982 , \7983 ,
         \7984 , \7985 , \7986 , \7987 , \7988 , \7989 , \7990 , \7991 , \7992 , \7993 ,
         \7994 , \7995 , \7996 , \7997 , \7998 , \7999 , \8000 , \8001 , \8002 , \8003 ,
         \8004 , \8005 , \8006 , \8007 , \8008 , \8009 , \8010 , \8011 , \8012 , \8013 ,
         \8014 , \8015 , \8016 , \8017 , \8018 , \8019 , \8020 , \8021 , \8022 , \8023 ,
         \8024 , \8025 , \8026 , \8027 , \8028 , \8029 , \8030 , \8031 , \8032 , \8033 ,
         \8034 , \8035 , \8036 , \8037 , \8038 , \8039 , \8040 , \8041 , \8042 , \8043 ,
         \8044 , \8045 , \8046 , \8047 , \8048 , \8049 , \8050 , \8051 , \8052 , \8053 ,
         \8054 , \8055 , \8056 , \8057 , \8058 , \8059 , \8060 , \8061 , \8062 , \8063 ,
         \8064 , \8065 , \8066 , \8067 , \8068 , \8069 , \8070 , \8071 , \8072 , \8073 ,
         \8074 , \8075 , \8076 , \8077 , \8078 , \8079 , \8080 , \8081 , \8082 , \8083 ,
         \8084 , \8085 , \8086 , \8087 , \8088 , \8089 , \8090 , \8091 , \8092 , \8093 ,
         \8094 , \8095 , \8096 , \8097 , \8098 , \8099 , \8100 , \8101 , \8102 , \8103 ,
         \8104 , \8105 , \8106 , \8107 , \8108 , \8109 , \8110 , \8111 , \8112 , \8113 ,
         \8114 , \8115 , \8116 , \8117 , \8118 , \8119 , \8120 , \8121 , \8122 , \8123 ,
         \8124 , \8125 , \8126 , \8127 , \8128 , \8129 , \8130 , \8131 , \8132 , \8133 ,
         \8134 , \8135 , \8136 , \8137 , \8138 , \8139 , \8140 , \8141 , \8142 , \8143 ,
         \8144 , \8145 , \8146 , \8147 , \8148 , \8149 , \8150 , \8151 , \8152 , \8153 ,
         \8154 , \8155 , \8156 , \8157 , \8158 , \8159 , \8160 , \8161 , \8162 , \8163 ,
         \8164 , \8165 , \8166 , \8167 , \8168 , \8169 , \8170 , \8171 , \8172 , \8173 ,
         \8174 , \8175 , \8176 , \8177 , \8178 , \8179 , \8180 , \8181 , \8182 , \8183 ,
         \8184 , \8185 , \8186 , \8187 , \8188 , \8189 , \8190 , \8191 , \8192 , \8193 ,
         \8194 , \8195 , \8196 , \8197 , \8198 , \8199 , \8200 , \8201 , \8202 , \8203 ,
         \8204 , \8205 , \8206 , \8207 , \8208 , \8209 , \8210 , \8211 , \8212 , \8213 ,
         \8214 , \8215 , \8216 , \8217 , \8218 , \8219 , \8220 , \8221 , \8222 , \8223 ,
         \8224 , \8225 , \8226 , \8227 , \8228 , \8229 , \8230 , \8231 , \8232 , \8233 ,
         \8234 , \8235 , \8236 , \8237 , \8238 , \8239 , \8240 , \8241 , \8242 , \8243 ,
         \8244 , \8245 , \8246 , \8247 , \8248 , \8249 , \8250 , \8251 , \8252 , \8253 ,
         \8254 , \8255 , \8256 , \8257 , \8258 , \8259 , \8260 , \8261 , \8262 , \8263 ,
         \8264 , \8265 , \8266 , \8267 , \8268 , \8269 , \8270 , \8271 , \8272 , \8273 ,
         \8274 , \8275 , \8276 , \8277 , \8278 , \8279 , \8280 , \8281 , \8282 , \8283 ,
         \8284 , \8285 , \8286 , \8287 , \8288 , \8289 , \8290 , \8291 , \8292 , \8293 ,
         \8294 , \8295 , \8296 , \8297 , \8298 , \8299 , \8300 , \8301 , \8302 , \8303 ,
         \8304 , \8305 , \8306 , \8307 , \8308 , \8309 , \8310 , \8311 , \8312 , \8313 ,
         \8314 , \8315 , \8316 , \8317 , \8318 , \8319 , \8320 , \8321 , \8322 , \8323 ,
         \8324 , \8325 , \8326 , \8327 , \8328 , \8329 , \8330 , \8331 , \8332 , \8333 ,
         \8334 , \8335 , \8336 , \8337 , \8338 , \8339 , \8340 , \8341 , \8342 , \8343 ,
         \8344 , \8345 , \8346 , \8347 , \8348 , \8349 , \8350 , \8351 , \8352 , \8353 ,
         \8354 , \8355 , \8356 , \8357 , \8358 , \8359 , \8360 , \8361 , \8362 , \8363 ,
         \8364 , \8365 , \8366 , \8367 , \8368 , \8369 , \8370 , \8371 , \8372 , \8373 ,
         \8374 , \8375 , \8376 , \8377 , \8378 , \8379 , \8380 , \8381 , \8382 , \8383 ,
         \8384 , \8385 , \8386 , \8387 , \8388 , \8389 , \8390 , \8391 , \8392 , \8393 ,
         \8394 , \8395 , \8396 , \8397 , \8398 , \8399 , \8400 , \8401 , \8402 , \8403 ,
         \8404 , \8405 , \8406 , \8407 , \8408 , \8409 , \8410 , \8411 , \8412 , \8413 ,
         \8414 , \8415 , \8416 , \8417 , \8418 , \8419 , \8420 , \8421 , \8422 , \8423 ,
         \8424 , \8425 , \8426 , \8427 , \8428 , \8429 , \8430 , \8431 , \8432 , \8433 ,
         \8434 , \8435 , \8436 , \8437 , \8438 , \8439 , \8440 , \8441 , \8442 , \8443 ,
         \8444 , \8445 , \8446 , \8447 , \8448 , \8449 , \8450 , \8451 , \8452 , \8453 ,
         \8454 , \8455 , \8456 , \8457 , \8458 , \8459 , \8460 , \8461 , \8462 , \8463 ,
         \8464 , \8465 , \8466 , \8467 , \8468 , \8469 , \8470 , \8471 , \8472 , \8473 ,
         \8474 , \8475 , \8476 , \8477 , \8478 , \8479 , \8480 , \8481 , \8482 , \8483 ,
         \8484 , \8485 , \8486 , \8487 , \8488 , \8489 , \8490 , \8491 , \8492 , \8493 ,
         \8494 , \8495 , \8496 , \8497 , \8498 , \8499 , \8500 , \8501 , \8502 , \8503 ,
         \8504 , \8505 , \8506 , \8507 , \8508 , \8509 , \8510 , \8511 , \8512 , \8513 ,
         \8514 , \8515 , \8516 , \8517 , \8518 , \8519 , \8520 , \8521 , \8522 , \8523 ,
         \8524 , \8525 , \8526 , \8527 , \8528 , \8529 , \8530 , \8531 , \8532 , \8533 ,
         \8534 , \8535 , \8536 , \8537 , \8538 , \8539 , \8540 , \8541 , \8542 , \8543 ,
         \8544 , \8545 , \8546 , \8547 , \8548 , \8549 , \8550 , \8551 , \8552 , \8553 ,
         \8554 , \8555 , \8556 , \8557 , \8558 , \8559 , \8560 , \8561 , \8562 , \8563 ,
         \8564 , \8565 , \8566 , \8567 , \8568 , \8569 , \8570 , \8571 , \8572 , \8573 ,
         \8574 , \8575 , \8576 , \8577 , \8578 , \8579 , \8580 , \8581 , \8582 , \8583 ,
         \8584 , \8585 , \8586 , \8587 , \8588 , \8589 , \8590 , \8591 , \8592 , \8593 ,
         \8594 , \8595 , \8596 , \8597 , \8598 , \8599 , \8600 , \8601 , \8602 , \8603 ,
         \8604 , \8605 , \8606 , \8607 , \8608 , \8609 , \8610 , \8611 , \8612 , \8613 ,
         \8614 , \8615 , \8616 , \8617 , \8618 , \8619 , \8620 , \8621 , \8622 , \8623 ,
         \8624 , \8625 , \8626 , \8627 , \8628 , \8629 , \8630 , \8631 , \8632 , \8633 ,
         \8634 , \8635 , \8636 , \8637 , \8638 , \8639 , \8640 , \8641 , \8642 , \8643 ,
         \8644 , \8645 , \8646 , \8647 , \8648 , \8649 , \8650 , \8651 , \8652 , \8653 ,
         \8654 , \8655 , \8656 , \8657 , \8658 , \8659 , \8660 , \8661 , \8662 , \8663 ,
         \8664 , \8665 , \8666 , \8667 , \8668 , \8669 , \8670 , \8671 , \8672 , \8673 ,
         \8674 , \8675 , \8676 , \8677 , \8678 , \8679 , \8680 , \8681 , \8682 , \8683 ,
         \8684 , \8685 , \8686 , \8687 , \8688 , \8689 , \8690 , \8691 , \8692 , \8693 ,
         \8694 , \8695 , \8696 , \8697 , \8698 , \8699 , \8700 , \8701 , \8702 , \8703 ,
         \8704 , \8705 , \8706 , \8707 , \8708 , \8709 , \8710 , \8711 , \8712 , \8713 ,
         \8714 , \8715 , \8716 , \8717 , \8718 , \8719 , \8720 , \8721 , \8722 , \8723 ,
         \8724 , \8725 , \8726 , \8727 , \8728 , \8729 , \8730 , \8731 , \8732 , \8733 ,
         \8734 , \8735 , \8736 , \8737 , \8738 , \8739 , \8740 , \8741 , \8742 , \8743 ,
         \8744 , \8745 , \8746 , \8747 , \8748 , \8749 , \8750 , \8751 , \8752 , \8753 ,
         \8754 , \8755 , \8756 , \8757 , \8758 , \8759 , \8760 , \8761 , \8762 , \8763 ,
         \8764 , \8765 , \8766 , \8767 , \8768 , \8769 , \8770 , \8771 , \8772 , \8773 ,
         \8774 , \8775 , \8776 , \8777 , \8778 , \8779 , \8780 , \8781 , \8782 , \8783 ,
         \8784 , \8785 , \8786 , \8787 , \8788 , \8789 , \8790 , \8791 , \8792 , \8793 ,
         \8794 , \8795 , \8796 , \8797 , \8798 , \8799 , \8800 , \8801 , \8802 , \8803 ,
         \8804 , \8805 , \8806 , \8807 , \8808 , \8809 , \8810 , \8811 , \8812 , \8813 ,
         \8814 , \8815 , \8816 , \8817 , \8818 , \8819 , \8820 , \8821 , \8822 , \8823 ,
         \8824 , \8825 , \8826 , \8827 , \8828 , \8829 , \8830 , \8831 , \8832 , \8833 ,
         \8834 , \8835 , \8836 , \8837 , \8838 , \8839 , \8840 , \8841 , \8842 , \8843 ,
         \8844 , \8845 , \8846 , \8847 , \8848 , \8849 , \8850 , \8851 , \8852 , \8853 ,
         \8854 , \8855 , \8856 , \8857 , \8858 , \8859 , \8860 , \8861 , \8862 , \8863 ,
         \8864 , \8865 , \8866 , \8867 , \8868 , \8869 , \8870 , \8871 , \8872 , \8873 ,
         \8874 , \8875 , \8876 , \8877 , \8878 , \8879 , \8880 , \8881 , \8882 , \8883 ,
         \8884 , \8885 , \8886 , \8887 , \8888 , \8889 , \8890 , \8891 , \8892 , \8893 ,
         \8894 , \8895 , \8896 , \8897 , \8898 , \8899 , \8900 , \8901 , \8902 , \8903 ,
         \8904 , \8905 , \8906 , \8907 , \8908 , \8909 , \8910 , \8911 , \8912 , \8913 ,
         \8914 , \8915 , \8916 , \8917 , \8918 , \8919 , \8920 , \8921 , \8922 , \8923 ,
         \8924 , \8925 , \8926 , \8927 , \8928 , \8929 , \8930 , \8931 , \8932 , \8933 ,
         \8934 , \8935 , \8936 , \8937 , \8938 , \8939 , \8940 , \8941 , \8942 , \8943 ,
         \8944 , \8945 , \8946 , \8947 , \8948 , \8949 , \8950 , \8951 , \8952 , \8953 ,
         \8954 , \8955 , \8956 , \8957 , \8958 , \8959 , \8960 , \8961 , \8962 , \8963 ,
         \8964 , \8965 , \8966 , \8967 , \8968 , \8969 , \8970 , \8971 , \8972 , \8973 ,
         \8974 , \8975 , \8976 , \8977 , \8978 , \8979 , \8980 , \8981 , \8982 , \8983 ,
         \8984 , \8985 , \8986 , \8987 , \8988 , \8989 , \8990 , \8991 , \8992 , \8993 ,
         \8994 , \8995 , \8996 , \8997 , \8998 , \8999 , \9000 , \9001 , \9002 , \9003 ,
         \9004 , \9005 , \9006 , \9007 , \9008 , \9009 , \9010 , \9011 , \9012 , \9013 ,
         \9014 , \9015 , \9016 , \9017 , \9018 , \9019 , \9020 , \9021 , \9022 , \9023 ,
         \9024 , \9025 , \9026 , \9027 , \9028 , \9029 , \9030 , \9031 , \9032 , \9033 ,
         \9034 , \9035 , \9036 , \9037 , \9038 , \9039 , \9040 , \9041 , \9042 , \9043 ,
         \9044 , \9045 , \9046 , \9047 , \9048 , \9049 , \9050 , \9051 , \9052 , \9053 ,
         \9054 , \9055 , \9056 , \9057 , \9058 , \9059 , \9060 , \9061 , \9062 , \9063 ,
         \9064 , \9065 , \9066 , \9067 , \9068 , \9069 , \9070 , \9071 , \9072 , \9073 ,
         \9074 , \9075 , \9076 , \9077 , \9078 , \9079 , \9080 , \9081 , \9082 , \9083 ,
         \9084 , \9085 , \9086 , \9087 , \9088 , \9089 , \9090 , \9091 , \9092 , \9093 ,
         \9094 , \9095 , \9096 , \9097 , \9098 , \9099 , \9100 , \9101 , \9102 , \9103 ,
         \9104 , \9105 , \9106 , \9107 , \9108 , \9109 , \9110 , \9111 , \9112 , \9113 ,
         \9114 , \9115 , \9116 , \9117 , \9118 , \9119 , \9120 , \9121 , \9122 , \9123 ,
         \9124 , \9125 , \9126 , \9127 , \9128 , \9129 , \9130 , \9131 , \9132 , \9133 ,
         \9134 , \9135 , \9136 , \9137 , \9138 , \9139 , \9140 , \9141 , \9142 , \9143 ,
         \9144 , \9145 , \9146 , \9147 , \9148 , \9149 , \9150 , \9151 , \9152 , \9153 ,
         \9154 , \9155 , \9156 , \9157 , \9158 , \9159 , \9160 , \9161 , \9162 , \9163 ,
         \9164 , \9165 , \9166 , \9167 , \9168 , \9169 , \9170 , \9171 , \9172 , \9173 ,
         \9174 , \9175 , \9176 , \9177 , \9178 , \9179 , \9180 , \9181 , \9182 , \9183 ,
         \9184 , \9185 , \9186 , \9187 , \9188 , \9189 , \9190 , \9191 , \9192 , \9193 ,
         \9194 , \9195 , \9196 , \9197 , \9198 , \9199 , \9200 , \9201 , \9202 , \9203 ,
         \9204 , \9205 , \9206 , \9207 , \9208 , \9209 , \9210 , \9211 , \9212 , \9213 ,
         \9214 , \9215 , \9216 , \9217 , \9218 , \9219 , \9220 , \9221 , \9222 , \9223 ,
         \9224 , \9225 , \9226 , \9227 , \9228 , \9229 , \9230 , \9231 , \9232 , \9233 ,
         \9234 , \9235 , \9236 , \9237 , \9238 , \9239 , \9240 , \9241 , \9242 , \9243 ,
         \9244 , \9245 , \9246 , \9247 , \9248 , \9249 , \9250 , \9251 , \9252 , \9253 ,
         \9254 , \9255 , \9256 , \9257 , \9258 , \9259 , \9260 , \9261 , \9262 , \9263 ,
         \9264 , \9265 , \9266 , \9267 , \9268 , \9269 , \9270 , \9271 , \9272 , \9273 ,
         \9274 , \9275 , \9276 , \9277 , \9278 , \9279 , \9280 , \9281 , \9282 , \9283 ,
         \9284 , \9285 , \9286 , \9287 , \9288 , \9289 , \9290 , \9291 , \9292 , \9293 ,
         \9294 , \9295 , \9296 , \9297 , \9298 , \9299 , \9300 , \9301 , \9302 , \9303 ,
         \9304 , \9305 , \9306 , \9307 , \9308 , \9309 , \9310 , \9311 , \9312 , \9313 ,
         \9314 , \9315 , \9316 , \9317 , \9318 , \9319 , \9320 , \9321 , \9322 , \9323 ,
         \9324 , \9325 , \9326 , \9327 , \9328 , \9329 , \9330 , \9331 , \9332 , \9333 ,
         \9334 , \9335 , \9336 , \9337 , \9338 , \9339 , \9340 , \9341 , \9342 , \9343 ,
         \9344 , \9345 , \9346 , \9347 , \9348 , \9349 , \9350 , \9351 , \9352 , \9353 ,
         \9354 , \9355 , \9356 , \9357 , \9358 , \9359 , \9360 , \9361 , \9362 , \9363 ,
         \9364 , \9365 , \9366 , \9367 , \9368 , \9369 , \9370 , \9371 , \9372 , \9373 ,
         \9374 , \9375 , \9376 , \9377 , \9378 , \9379 , \9380 , \9381 , \9382 , \9383 ,
         \9384 , \9385 , \9386 , \9387 , \9388 , \9389 , \9390 , \9391 , \9392 , \9393 ,
         \9394 , \9395 , \9396 , \9397 , \9398 , \9399 , \9400 , \9401 , \9402 , \9403 ,
         \9404 , \9405 , \9406 , \9407 , \9408 , \9409 , \9410 , \9411 , \9412 , \9413 ,
         \9414 , \9415 , \9416 , \9417 , \9418 , \9419 , \9420 , \9421 , \9422 , \9423 ,
         \9424 , \9425 , \9426 , \9427 , \9428 , \9429 , \9430 , \9431 , \9432 , \9433 ,
         \9434 , \9435 , \9436 , \9437 , \9438 , \9439 , \9440 , \9441 , \9442 , \9443 ,
         \9444 , \9445 , \9446 , \9447 , \9448 , \9449 , \9450 , \9451 , \9452 , \9453 ,
         \9454 , \9455 , \9456 , \9457 , \9458 , \9459 , \9460 , \9461 , \9462 , \9463 ,
         \9464 , \9465 , \9466 , \9467 , \9468 , \9469 , \9470 , \9471 , \9472 , \9473 ,
         \9474 , \9475 , \9476 , \9477 , \9478 , \9479 , \9480 , \9481 , \9482 , \9483 ,
         \9484 , \9485 , \9486 , \9487 , \9488 , \9489 , \9490 , \9491 , \9492 , \9493 ,
         \9494 , \9495 , \9496 , \9497 , \9498 , \9499 , \9500 , \9501 , \9502 , \9503 ,
         \9504 , \9505 , \9506 , \9507 , \9508 , \9509 , \9510 , \9511 , \9512 , \9513 ,
         \9514 , \9515 , \9516 , \9517 , \9518 , \9519 , \9520 , \9521 , \9522 , \9523 ,
         \9524 , \9525 , \9526 , \9527 , \9528 , \9529 , \9530 , \9531 , \9532 , \9533 ,
         \9534 , \9535 , \9536 , \9537 , \9538 , \9539 , \9540 , \9541 , \9542 , \9543 ,
         \9544 , \9545 , \9546 , \9547 , \9548 , \9549 , \9550 , \9551 , \9552 , \9553 ,
         \9554 , \9555 , \9556 , \9557 , \9558 , \9559 , \9560 , \9561 , \9562 , \9563 ,
         \9564 , \9565 , \9566 , \9567 , \9568 , \9569 , \9570 , \9571 , \9572 , \9573 ,
         \9574 , \9575 , \9576 , \9577 , \9578 , \9579 , \9580 , \9581 , \9582 , \9583 ,
         \9584 , \9585 , \9586 , \9587 , \9588 , \9589 , \9590 , \9591 , \9592 , \9593 ,
         \9594 , \9595 , \9596 , \9597 , \9598 , \9599 , \9600 , \9601 , \9602 , \9603 ,
         \9604 , \9605 , \9606 , \9607 , \9608 , \9609 , \9610 , \9611 , \9612 , \9613 ,
         \9614 , \9615 , \9616 , \9617 , \9618 , \9619 , \9620 , \9621 , \9622 , \9623 ,
         \9624 , \9625 , \9626 , \9627 , \9628 , \9629 , \9630 , \9631 , \9632 , \9633 ,
         \9634 , \9635 , \9636 , \9637 , \9638 , \9639 , \9640 , \9641 , \9642 , \9643 ,
         \9644 , \9645 , \9646 , \9647 , \9648 , \9649 , \9650 , \9651 , \9652 , \9653 ,
         \9654 , \9655 , \9656 , \9657 , \9658 , \9659 , \9660 , \9661 , \9662 , \9663 ,
         \9664 , \9665 , \9666 , \9667 , \9668 , \9669 , \9670 , \9671 , \9672 , \9673 ,
         \9674 , \9675 , \9676 , \9677 , \9678 , \9679 , \9680 , \9681 , \9682 , \9683 ,
         \9684 , \9685 , \9686 , \9687 , \9688 , \9689 , \9690 , \9691 , \9692 , \9693 ,
         \9694 , \9695 , \9696 , \9697 , \9698 , \9699 , \9700 , \9701 , \9702 , \9703 ,
         \9704 , \9705 , \9706 , \9707 , \9708 , \9709 , \9710 , \9711 , \9712 , \9713 ,
         \9714 , \9715 , \9716 , \9717 , \9718 , \9719 , \9720 , \9721 , \9722 , \9723 ,
         \9724 , \9725 , \9726 , \9727 , \9728 , \9729 , \9730 , \9731 , \9732 , \9733 ,
         \9734 , \9735 , \9736 , \9737 , \9738 , \9739 , \9740 , \9741 , \9742 , \9743 ,
         \9744 , \9745 , \9746 , \9747 , \9748 , \9749 , \9750 , \9751 , \9752 , \9753 ,
         \9754 , \9755 , \9756 , \9757 , \9758 , \9759 , \9760 , \9761 , \9762 , \9763 ,
         \9764 , \9765 , \9766 , \9767 , \9768 , \9769 , \9770 , \9771 , \9772 , \9773 ,
         \9774 , \9775 , \9776 , \9777 , \9778 , \9779 , \9780 , \9781 , \9782 , \9783 ,
         \9784 , \9785 , \9786 , \9787 , \9788 , \9789 , \9790 , \9791 , \9792 , \9793 ,
         \9794 , \9795 , \9796 , \9797 , \9798 , \9799 , \9800 , \9801 , \9802 , \9803 ,
         \9804 , \9805 , \9806 , \9807 , \9808 , \9809 , \9810 , \9811 , \9812 , \9813 ,
         \9814 , \9815 , \9816 , \9817 , \9818 , \9819 , \9820 , \9821 , \9822 , \9823 ,
         \9824 , \9825 , \9826 , \9827 , \9828 , \9829 , \9830 , \9831 , \9832 , \9833 ,
         \9834 , \9835 , \9836 , \9837 , \9838 , \9839 , \9840 , \9841 , \9842 , \9843 ,
         \9844 , \9845 , \9846 , \9847 , \9848 , \9849 , \9850 , \9851 , \9852 , \9853 ,
         \9854 , \9855 , \9856 , \9857 , \9858 , \9859 , \9860 , \9861 , \9862 , \9863 ,
         \9864 , \9865 , \9866 , \9867 , \9868 , \9869 , \9870 , \9871 , \9872 , \9873 ,
         \9874 , \9875 , \9876 , \9877 , \9878 , \9879 , \9880 , \9881 , \9882 , \9883 ,
         \9884 , \9885 , \9886 , \9887 , \9888 , \9889 , \9890 , \9891 , \9892 , \9893 ,
         \9894 , \9895 , \9896 , \9897 , \9898 , \9899 , \9900 , \9901 , \9902 , \9903 ,
         \9904 , \9905 , \9906 , \9907 , \9908 , \9909 , \9910 , \9911 , \9912 , \9913 ,
         \9914 , \9915 , \9916 , \9917 , \9918 , \9919 , \9920 , \9921 , \9922 , \9923 ,
         \9924 , \9925 , \9926 , \9927 , \9928 , \9929 , \9930 , \9931 , \9932 , \9933 ,
         \9934 , \9935 , \9936 , \9937 , \9938 , \9939 , \9940 , \9941 , \9942 , \9943 ,
         \9944 , \9945 , \9946 , \9947 , \9948 , \9949 , \9950 , \9951 , \9952 , \9953 ,
         \9954 , \9955 , \9956 , \9957 , \9958 , \9959 , \9960 , \9961 , \9962 , \9963 ,
         \9964 , \9965 , \9966 , \9967 , \9968 , \9969 , \9970 , \9971 , \9972 , \9973 ,
         \9974 , \9975 , \9976 , \9977 , \9978 , \9979 , \9980 , \9981 , \9982 , \9983 ,
         \9984 , \9985 , \9986 , \9987 , \9988 , \9989 , \9990 , \9991 , \9992 , \9993 ,
         \9994 , \9995 , \9996 , \9997 , \9998 , \9999 , \10000 , \10001 , \10002 , \10003 ,
         \10004 , \10005 , \10006 , \10007 , \10008 , \10009 , \10010 , \10011 , \10012 , \10013 ,
         \10014 , \10015 , \10016 , \10017 , \10018 , \10019 , \10020 , \10021 , \10022 , \10023 ,
         \10024 , \10025 , \10026 , \10027 , \10028 , \10029 , \10030 , \10031 , \10032 , \10033 ,
         \10034 , \10035 , \10036 , \10037 , \10038 , \10039 , \10040 , \10041 , \10042 , \10043 ,
         \10044 , \10045 , \10046 , \10047 , \10048 , \10049 , \10050 , \10051 , \10052 , \10053 ,
         \10054 , \10055 , \10056 , \10057 , \10058 , \10059 , \10060 , \10061 , \10062 , \10063 ,
         \10064 , \10065 , \10066 , \10067 , \10068 , \10069 , \10070 , \10071 , \10072 , \10073 ,
         \10074 , \10075 , \10076 , \10077 , \10078 , \10079 , \10080 , \10081 , \10082 , \10083 ,
         \10084 , \10085 , \10086 , \10087 , \10088 , \10089 , \10090 , \10091 , \10092 , \10093 ,
         \10094 , \10095 , \10096 , \10097 , \10098 , \10099 , \10100 , \10101 , \10102 , \10103 ,
         \10104 , \10105 , \10106 , \10107 , \10108 , \10109 , \10110 , \10111 , \10112 , \10113 ,
         \10114 , \10115 , \10116 , \10117 , \10118 , \10119 , \10120 , \10121 , \10122 , \10123 ,
         \10124 , \10125 , \10126 , \10127 , \10128 , \10129 , \10130 , \10131 , \10132 , \10133 ,
         \10134 , \10135 , \10136 , \10137 , \10138 , \10139 , \10140 , \10141 , \10142 , \10143 ,
         \10144 , \10145 , \10146 , \10147 , \10148 , \10149 , \10150 , \10151 , \10152 , \10153 ,
         \10154 , \10155 , \10156 , \10157 , \10158 , \10159 , \10160 , \10161 , \10162 , \10163 ,
         \10164 , \10165 , \10166 , \10167 , \10168 , \10169 , \10170 , \10171 , \10172 , \10173 ,
         \10174 , \10175 , \10176 , \10177 , \10178 , \10179 , \10180 , \10181 , \10182 , \10183 ,
         \10184 , \10185 , \10186 , \10187 , \10188 , \10189 , \10190 , \10191 , \10192 , \10193 ,
         \10194 , \10195 , \10196 , \10197 , \10198 , \10199 , \10200 , \10201 , \10202 , \10203 ,
         \10204 , \10205 , \10206 , \10207 , \10208 , \10209 , \10210 , \10211 , \10212 , \10213 ,
         \10214 , \10215 , \10216 , \10217 , \10218 , \10219 , \10220 , \10221 , \10222 , \10223 ,
         \10224 , \10225 , \10226 , \10227 , \10228 , \10229 , \10230 , \10231 , \10232 , \10233 ,
         \10234 , \10235 , \10236 , \10237 , \10238 , \10239 , \10240 , \10241 , \10242 , \10243 ,
         \10244 , \10245 , \10246 , \10247 , \10248 , \10249 , \10250 , \10251 , \10252 , \10253 ,
         \10254 , \10255 , \10256 , \10257 , \10258 , \10259 , \10260 , \10261 , \10262 , \10263 ,
         \10264 , \10265 , \10266 , \10267 , \10268 , \10269 , \10270 , \10271 , \10272 , \10273 ,
         \10274 , \10275 , \10276 , \10277 , \10278 , \10279 , \10280 , \10281 , \10282 , \10283 ,
         \10284 , \10285 , \10286 , \10287 , \10288 , \10289 , \10290 , \10291 , \10292 , \10293 ,
         \10294 , \10295 , \10296 , \10297 , \10298 , \10299 , \10300 , \10301 , \10302 , \10303 ,
         \10304 , \10305 , \10306 , \10307 , \10308 , \10309 , \10310 , \10311 , \10312 , \10313 ,
         \10314 , \10315 , \10316 , \10317 , \10318 , \10319 , \10320 , \10321 , \10322 , \10323 ,
         \10324 , \10325 , \10326 , \10327 , \10328 , \10329 , \10330 , \10331 , \10332 , \10333 ,
         \10334 , \10335 , \10336 , \10337 , \10338 , \10339 , \10340 , \10341 , \10342 , \10343 ,
         \10344 , \10345 , \10346 , \10347 , \10348 , \10349 , \10350 , \10351 , \10352 , \10353 ,
         \10354 , \10355 , \10356 , \10357 , \10358 , \10359 , \10360 , \10361 , \10362 , \10363 ,
         \10364 , \10365 , \10366 , \10367 , \10368 , \10369 , \10370 , \10371 , \10372 , \10373 ,
         \10374 , \10375 , \10376 , \10377 , \10378 , \10379 , \10380 , \10381 , \10382 , \10383 ,
         \10384 , \10385 , \10386 , \10387 , \10388 , \10389 , \10390 , \10391 , \10392 , \10393 ,
         \10394 , \10395 , \10396 , \10397 , \10398 , \10399 , \10400 , \10401 , \10402 , \10403 ,
         \10404 , \10405 , \10406 , \10407 , \10408 , \10409 , \10410 , \10411 , \10412 , \10413 ,
         \10414 , \10415 , \10416 , \10417 , \10418 , \10419 , \10420 , \10421 , \10422 , \10423 ,
         \10424 , \10425 , \10426 , \10427 , \10428 , \10429 , \10430 , \10431 , \10432 , \10433 ,
         \10434 , \10435 , \10436 , \10437 , \10438 , \10439 , \10440 , \10441 , \10442 , \10443 ,
         \10444 , \10445 , \10446 , \10447 , \10448 , \10449 , \10450 , \10451 , \10452 , \10453 ,
         \10454 , \10455 , \10456 , \10457 , \10458 , \10459 , \10460 , \10461 , \10462 , \10463 ,
         \10464 , \10465 , \10466 , \10467 , \10468 , \10469 , \10470 , \10471 , \10472 , \10473 ,
         \10474 , \10475 , \10476 , \10477 , \10478 , \10479 , \10480 , \10481 , \10482 , \10483 ,
         \10484 , \10485 , \10486 , \10487 , \10488 , \10489 , \10490 , \10491 , \10492 , \10493 ,
         \10494 , \10495 , \10496 , \10497 , \10498 , \10499 , \10500 , \10501 , \10502 , \10503 ,
         \10504 , \10505 , \10506 , \10507 , \10508 , \10509 , \10510 , \10511 , \10512 , \10513 ,
         \10514 , \10515 , \10516 , \10517 , \10518 , \10519 , \10520 , \10521 , \10522 , \10523 ,
         \10524 , \10525 , \10526 , \10527 , \10528 , \10529 , \10530 , \10531 , \10532 , \10533 ,
         \10534 , \10535 , \10536 , \10537 , \10538 , \10539 , \10540 , \10541 , \10542 , \10543 ,
         \10544 , \10545 , \10546 , \10547 , \10548 , \10549 , \10550 , \10551 , \10552 , \10553 ,
         \10554 , \10555 , \10556 , \10557 , \10558 , \10559 , \10560 , \10561 , \10562 , \10563 ,
         \10564 , \10565 , \10566 , \10567 , \10568 , \10569 , \10570 , \10571 , \10572 , \10573 ,
         \10574 , \10575 , \10576 , \10577 , \10578 , \10579 , \10580 , \10581 , \10582 , \10583 ,
         \10584 , \10585 , \10586 , \10587 , \10588 , \10589 , \10590 , \10591 , \10592 , \10593 ,
         \10594 , \10595 , \10596 , \10597 , \10598 , \10599 , \10600 , \10601 , \10602 , \10603 ,
         \10604 , \10605 , \10606 , \10607 , \10608 , \10609 , \10610 , \10611 , \10612 , \10613 ,
         \10614 , \10615 , \10616 , \10617 , \10618 , \10619 , \10620 , \10621 , \10622 , \10623 ,
         \10624 , \10625 , \10626 , \10627 , \10628 , \10629 , \10630 , \10631 , \10632 , \10633 ,
         \10634 , \10635 , \10636 , \10637 , \10638 , \10639 , \10640 , \10641 , \10642 , \10643 ,
         \10644 , \10645 , \10646 , \10647 , \10648 , \10649 , \10650 , \10651 , \10652 , \10653 ,
         \10654 , \10655 , \10656 , \10657 , \10658 , \10659 , \10660 , \10661 , \10662 , \10663 ,
         \10664 , \10665 , \10666 , \10667 , \10668 , \10669 , \10670 , \10671 , \10672 , \10673 ,
         \10674 , \10675 , \10676 , \10677 , \10678 , \10679 , \10680 , \10681 , \10682 , \10683 ,
         \10684 , \10685 , \10686 , \10687 , \10688 , \10689 , \10690 , \10691 , \10692 , \10693 ,
         \10694 , \10695 , \10696 , \10697 , \10698 , \10699 , \10700 , \10701 , \10702 , \10703 ,
         \10704 , \10705 , \10706 , \10707 , \10708 , \10709 , \10710 , \10711 , \10712 , \10713 ,
         \10714 , \10715 , \10716 , \10717 , \10718 , \10719 , \10720 , \10721 , \10722 , \10723 ,
         \10724 , \10725 , \10726 , \10727 , \10728 , \10729 , \10730 , \10731 , \10732 , \10733 ,
         \10734 , \10735 , \10736 , \10737 , \10738 , \10739 , \10740 , \10741 , \10742 , \10743 ,
         \10744 , \10745 , \10746 , \10747 , \10748 , \10749 , \10750 , \10751 , \10752 , \10753 ,
         \10754 , \10755 , \10756 , \10757 , \10758 , \10759 , \10760 , \10761 , \10762 , \10763 ,
         \10764 , \10765 , \10766 , \10767 , \10768 , \10769 , \10770 , \10771 , \10772 , \10773 ,
         \10774 , \10775 , \10776 , \10777 , \10778 , \10779 , \10780 , \10781 , \10782 , \10783 ,
         \10784 , \10785 , \10786 , \10787 , \10788 , \10789 , \10790 , \10791 , \10792 , \10793 ,
         \10794 , \10795 , \10796 , \10797 , \10798 , \10799 , \10800 , \10801 , \10802 , \10803 ,
         \10804 , \10805 , \10806 , \10807 , \10808 , \10809 , \10810 , \10811 , \10812 , \10813 ,
         \10814 , \10815 , \10816 , \10817 , \10818 , \10819 , \10820 , \10821 , \10822 , \10823 ,
         \10824 , \10825 , \10826 , \10827 , \10828 , \10829 , \10830 , \10831 , \10832 , \10833 ,
         \10834 , \10835 , \10836 , \10837 , \10838 , \10839 , \10840 , \10841 , \10842 , \10843 ,
         \10844 , \10845 , \10846 , \10847 , \10848 , \10849 , \10850 , \10851 , \10852 , \10853 ,
         \10854 , \10855 , \10856 , \10857 , \10858 , \10859 , \10860 , \10861 , \10862 , \10863 ,
         \10864 , \10865 , \10866 , \10867 , \10868 , \10869 , \10870 , \10871 , \10872 , \10873 ,
         \10874 , \10875 , \10876 , \10877 , \10878 , \10879 , \10880 , \10881 , \10882 , \10883 ,
         \10884 , \10885 , \10886 , \10887 , \10888 , \10889 , \10890 , \10891 , \10892 , \10893 ,
         \10894 , \10895 , \10896 , \10897 , \10898 , \10899 , \10900 , \10901 , \10902 , \10903 ,
         \10904 , \10905 , \10906 , \10907 , \10908 , \10909 , \10910 , \10911 , \10912 , \10913 ,
         \10914 , \10915 , \10916 , \10917 , \10918 , \10919 , \10920 , \10921 , \10922 , \10923 ,
         \10924 , \10925 , \10926 , \10927 , \10928 , \10929 , \10930 , \10931 , \10932 , \10933 ,
         \10934 , \10935 , \10936 , \10937 , \10938 , \10939 , \10940 , \10941 , \10942 , \10943 ,
         \10944 , \10945 , \10946 , \10947 , \10948 , \10949 , \10950 , \10951 , \10952 , \10953 ,
         \10954 , \10955 , \10956 , \10957 , \10958 , \10959 , \10960 , \10961 , \10962 , \10963 ,
         \10964 , \10965 , \10966 , \10967 , \10968 , \10969 , \10970 , \10971 , \10972 , \10973 ,
         \10974 , \10975 , \10976 , \10977 , \10978 , \10979 , \10980 , \10981 , \10982 , \10983 ,
         \10984 , \10985 , \10986 , \10987 , \10988 , \10989 , \10990 , \10991 , \10992 , \10993 ,
         \10994 , \10995 , \10996 , \10997 , \10998 , \10999 , \11000 , \11001 , \11002 , \11003 ,
         \11004 , \11005 , \11006 , \11007 , \11008 , \11009 , \11010 , \11011 , \11012 , \11013 ,
         \11014 , \11015 , \11016 , \11017 , \11018 , \11019 , \11020 , \11021 , \11022 , \11023 ,
         \11024 , \11025 , \11026 , \11027 , \11028 , \11029 , \11030 , \11031 , \11032 , \11033 ,
         \11034 , \11035 , \11036 , \11037 , \11038 , \11039 , \11040 , \11041 , \11042 , \11043 ,
         \11044 , \11045 , \11046 , \11047 , \11048 , \11049 , \11050 , \11051 , \11052 , \11053 ,
         \11054 , \11055 , \11056 , \11057 , \11058 , \11059 , \11060 , \11061 , \11062 , \11063 ,
         \11064 , \11065 , \11066 , \11067 , \11068 , \11069 , \11070 , \11071 , \11072 , \11073 ,
         \11074 , \11075 , \11076 , \11077 , \11078 , \11079 , \11080 , \11081 , \11082 , \11083 ,
         \11084 , \11085 , \11086 , \11087 , \11088 , \11089 , \11090 , \11091 , \11092 , \11093 ,
         \11094 , \11095 , \11096 , \11097 , \11098 , \11099 , \11100 , \11101 , \11102 , \11103 ,
         \11104 , \11105 , \11106 , \11107 , \11108 , \11109 , \11110 , \11111 , \11112 , \11113 ,
         \11114 , \11115 , \11116 , \11117 , \11118 , \11119 , \11120 , \11121 , \11122 , \11123 ,
         \11124 , \11125 , \11126 , \11127 , \11128 , \11129 , \11130 , \11131 , \11132 , \11133 ,
         \11134 , \11135 , \11136 , \11137 , \11138 , \11139 , \11140 , \11141 , \11142 , \11143 ,
         \11144 , \11145 , \11146 , \11147 , \11148 , \11149 , \11150 , \11151 , \11152 , \11153 ,
         \11154 , \11155 , \11156 , \11157 , \11158 , \11159 , \11160 , \11161 , \11162 , \11163 ,
         \11164 , \11165 , \11166 , \11167 , \11168 , \11169 , \11170 , \11171 , \11172 , \11173 ,
         \11174 , \11175 , \11176 , \11177 , \11178 , \11179 , \11180 , \11181 , \11182 , \11183 ,
         \11184 , \11185 , \11186 , \11187 , \11188 , \11189 , \11190 , \11191 , \11192 , \11193 ,
         \11194 , \11195 , \11196 , \11197 , \11198 , \11199 , \11200 , \11201 , \11202 , \11203 ,
         \11204 , \11205 , \11206 , \11207 , \11208 , \11209 , \11210 , \11211 , \11212 , \11213 ,
         \11214 , \11215 , \11216 , \11217 , \11218 , \11219 , \11220 , \11221 , \11222 , \11223 ,
         \11224 , \11225 , \11226 , \11227 , \11228 , \11229 , \11230 , \11231 , \11232 , \11233 ,
         \11234 , \11235 , \11236 , \11237 , \11238 , \11239 , \11240 , \11241 , \11242 , \11243 ,
         \11244 , \11245 , \11246 , \11247 , \11248 , \11249 , \11250 , \11251 , \11252 , \11253 ,
         \11254 , \11255 , \11256 , \11257 , \11258 , \11259 , \11260 , \11261 , \11262 , \11263 ,
         \11264 , \11265 , \11266 , \11267 , \11268 , \11269 , \11270 , \11271 , \11272 , \11273 ,
         \11274 , \11275 , \11276 , \11277 , \11278 , \11279 , \11280 , \11281 , \11282 , \11283 ,
         \11284 , \11285 , \11286 , \11287 , \11288 , \11289 , \11290 , \11291 , \11292 , \11293 ,
         \11294 , \11295 , \11296 , \11297 , \11298 , \11299 , \11300 , \11301 , \11302 , \11303 ,
         \11304 , \11305 , \11306 , \11307 , \11308 , \11309 , \11310 , \11311 , \11312 , \11313 ,
         \11314 , \11315 , \11316 , \11317 , \11318 , \11319 , \11320 , \11321 , \11322 , \11323 ,
         \11324 , \11325 , \11326 , \11327 , \11328 , \11329 , \11330 , \11331 , \11332 , \11333 ,
         \11334 , \11335 , \11336 , \11337 , \11338 , \11339 , \11340 , \11341 , \11342 , \11343 ,
         \11344 , \11345 , \11346 , \11347 , \11348 , \11349 , \11350 , \11351 , \11352 , \11353 ,
         \11354 , \11355 , \11356 , \11357 , \11358 , \11359 , \11360 , \11361 , \11362 , \11363 ,
         \11364 , \11365 , \11366 , \11367 , \11368 , \11369 , \11370 , \11371 , \11372 , \11373 ,
         \11374 , \11375 , \11376 , \11377 , \11378 , \11379 , \11380 , \11381 , \11382 , \11383 ,
         \11384 , \11385 , \11386 , \11387 , \11388 , \11389 , \11390 , \11391 , \11392 , \11393 ,
         \11394 , \11395 , \11396 , \11397 , \11398 , \11399 , \11400 , \11401 , \11402 , \11403 ,
         \11404 , \11405 , \11406 , \11407 , \11408 , \11409 , \11410 , \11411 , \11412 , \11413 ,
         \11414 , \11415 , \11416 , \11417 , \11418 , \11419 , \11420 , \11421 , \11422 , \11423 ,
         \11424 , \11425 , \11426 , \11427 , \11428 , \11429 , \11430 , \11431 , \11432 , \11433 ,
         \11434 , \11435 , \11436 , \11437 , \11438 , \11439 , \11440 , \11441 , \11442 , \11443 ,
         \11444 , \11445 , \11446 , \11447 , \11448 , \11449 , \11450 , \11451 , \11452 , \11453 ,
         \11454 , \11455 , \11456 , \11457 , \11458 , \11459 , \11460 , \11461 , \11462 , \11463 ,
         \11464 , \11465 , \11466 , \11467 , \11468 , \11469 , \11470 , \11471 , \11472 , \11473 ,
         \11474 , \11475 , \11476 , \11477 , \11478 , \11479 , \11480 , \11481 , \11482 , \11483 ,
         \11484 , \11485 , \11486 , \11487 , \11488 , \11489 , \11490 , \11491 , \11492 , \11493 ,
         \11494 , \11495 , \11496 , \11497 , \11498 , \11499 , \11500 , \11501 , \11502 , \11503 ,
         \11504 , \11505 , \11506 , \11507 , \11508 , \11509 , \11510 , \11511 , \11512 , \11513 ,
         \11514 , \11515 , \11516 , \11517 , \11518 , \11519 , \11520 , \11521 , \11522 , \11523 ,
         \11524 , \11525 , \11526 , \11527 , \11528 , \11529 , \11530 , \11531 , \11532 , \11533 ,
         \11534 , \11535 , \11536 , \11537 , \11538 , \11539 , \11540 , \11541 , \11542 , \11543 ,
         \11544 , \11545 , \11546 , \11547 , \11548 , \11549 , \11550 , \11551 , \11552 , \11553 ,
         \11554 , \11555 , \11556 , \11557 , \11558 , \11559 , \11560 , \11561 , \11562 , \11563 ,
         \11564 , \11565 , \11566 , \11567 , \11568 , \11569 , \11570 , \11571 , \11572 , \11573 ,
         \11574 , \11575 , \11576 , \11577 , \11578 , \11579 , \11580 , \11581 , \11582 , \11583 ,
         \11584 , \11585 , \11586 , \11587 , \11588 , \11589 , \11590 , \11591 , \11592 , \11593 ,
         \11594 , \11595 , \11596 , \11597 , \11598 , \11599 , \11600 , \11601 , \11602 , \11603 ,
         \11604 , \11605 , \11606 , \11607 , \11608 , \11609 , \11610 , \11611 , \11612 , \11613 ,
         \11614 , \11615 , \11616 , \11617 , \11618 , \11619 , \11620 , \11621 , \11622 , \11623 ,
         \11624 , \11625 , \11626 , \11627 , \11628 , \11629 , \11630 , \11631 , \11632 , \11633 ,
         \11634 , \11635 , \11636 , \11637 , \11638 , \11639 , \11640 , \11641 , \11642 , \11643 ,
         \11644 , \11645 , \11646 , \11647 , \11648 , \11649 , \11650 , \11651 , \11652 , \11653 ,
         \11654 , \11655 , \11656 , \11657 , \11658 , \11659 , \11660 , \11661 , \11662 , \11663 ,
         \11664 , \11665 , \11666 , \11667 , \11668 , \11669 , \11670 , \11671 , \11672 , \11673 ,
         \11674 , \11675 , \11676 , \11677 , \11678 , \11679 , \11680 , \11681 , \11682 , \11683 ,
         \11684 , \11685 , \11686 , \11687 , \11688 , \11689 , \11690 , \11691 , \11692 , \11693 ,
         \11694 , \11695 , \11696 , \11697 , \11698 , \11699 , \11700 , \11701 , \11702 , \11703 ,
         \11704 , \11705 , \11706 , \11707 , \11708 , \11709 , \11710 , \11711 , \11712 , \11713 ,
         \11714 , \11715 , \11716 , \11717 , \11718 , \11719 , \11720 , \11721 , \11722 , \11723 ,
         \11724 , \11725 , \11726 , \11727 , \11728 , \11729 , \11730 , \11731 , \11732 , \11733 ,
         \11734 , \11735 , \11736 , \11737 , \11738 , \11739 , \11740 , \11741 , \11742 , \11743 ,
         \11744 , \11745 , \11746 , \11747 , \11748 , \11749 , \11750 , \11751 , \11752 , \11753 ,
         \11754 , \11755 , \11756 , \11757 , \11758 , \11759 , \11760 , \11761 , \11762 , \11763 ,
         \11764 , \11765 , \11766 , \11767 , \11768 , \11769 , \11770 , \11771 , \11772 , \11773 ,
         \11774 , \11775 , \11776 , \11777 , \11778 , \11779 , \11780 , \11781 , \11782 , \11783 ,
         \11784 , \11785 , \11786 , \11787 , \11788 , \11789 , \11790 , \11791 , \11792 , \11793 ,
         \11794 , \11795 , \11796 , \11797 , \11798 , \11799 , \11800 , \11801 , \11802 , \11803 ,
         \11804 , \11805 , \11806 , \11807 , \11808 , \11809 , \11810 , \11811 , \11812 , \11813 ,
         \11814 , \11815 , \11816 , \11817 , \11818 , \11819 , \11820 , \11821 , \11822 , \11823 ,
         \11824 , \11825 , \11826 , \11827 , \11828 , \11829 , \11830 , \11831 , \11832 , \11833 ,
         \11834 , \11835 , \11836 , \11837 , \11838 , \11839 , \11840 , \11841 , \11842 , \11843 ,
         \11844 , \11845 , \11846 , \11847 , \11848 , \11849 , \11850 , \11851 , \11852 , \11853 ,
         \11854 , \11855 , \11856 , \11857 , \11858 , \11859 , \11860 , \11861 , \11862 , \11863 ,
         \11864 , \11865 , \11866 , \11867 , \11868 , \11869 , \11870 , \11871 , \11872 , \11873 ,
         \11874 , \11875 , \11876 , \11877 , \11878 , \11879 , \11880 , \11881 , \11882 , \11883 ,
         \11884 , \11885 , \11886 , \11887 , \11888 , \11889 , \11890 , \11891 , \11892 , \11893 ,
         \11894 , \11895 , \11896 , \11897 , \11898 , \11899 , \11900 , \11901 , \11902 , \11903 ,
         \11904 , \11905 , \11906 , \11907 , \11908 , \11909 , \11910 , \11911 , \11912 , \11913 ,
         \11914 , \11915 , \11916 , \11917 , \11918 , \11919 , \11920 , \11921 , \11922 , \11923 ,
         \11924 , \11925 , \11926 , \11927 , \11928 , \11929 , \11930 , \11931 , \11932 , \11933 ,
         \11934 , \11935 , \11936 , \11937 , \11938 , \11939 , \11940 , \11941 , \11942 , \11943 ,
         \11944 , \11945 , \11946 , \11947 , \11948 , \11949 , \11950 , \11951 , \11952 , \11953 ,
         \11954 , \11955 , \11956 , \11957 , \11958 , \11959 , \11960 , \11961 , \11962 , \11963 ,
         \11964 , \11965 , \11966 , \11967 , \11968 , \11969 , \11970 , \11971 , \11972 , \11973 ,
         \11974 , \11975 , \11976 , \11977 , \11978 , \11979 , \11980 , \11981 , \11982 , \11983 ,
         \11984 , \11985 , \11986 , \11987 , \11988 , \11989 , \11990 , \11991 , \11992 , \11993 ,
         \11994 , \11995 , \11996 , \11997 , \11998 , \11999 , \12000 , \12001 , \12002 , \12003 ,
         \12004 , \12005 , \12006 , \12007 , \12008 , \12009 , \12010 , \12011 , \12012 , \12013 ,
         \12014 , \12015 , \12016 , \12017 , \12018 , \12019 , \12020 , \12021 , \12022 , \12023 ,
         \12024 , \12025 , \12026 , \12027 , \12028 , \12029 , \12030 , \12031 , \12032 , \12033 ,
         \12034 , \12035 , \12036 , \12037 , \12038 , \12039 , \12040 , \12041 , \12042 , \12043 ,
         \12044 , \12045 , \12046 , \12047 , \12048 , \12049 , \12050 , \12051 , \12052 , \12053 ,
         \12054 , \12055 , \12056 , \12057 , \12058 , \12059 , \12060 , \12061 , \12062 , \12063 ,
         \12064 , \12065 , \12066 , \12067 , \12068 , \12069 , \12070 , \12071 , \12072 , \12073 ,
         \12074 , \12075 , \12076 , \12077 , \12078 , \12079 , \12080 , \12081 , \12082 , \12083 ,
         \12084 , \12085 , \12086 , \12087 , \12088 , \12089 , \12090 , \12091 , \12092 , \12093 ,
         \12094 , \12095 , \12096 , \12097 , \12098 , \12099 , \12100 , \12101 , \12102 , \12103 ,
         \12104 , \12105 , \12106 , \12107 , \12108 , \12109 , \12110 , \12111 , \12112 , \12113 ,
         \12114 , \12115 , \12116 , \12117 , \12118 , \12119 , \12120 , \12121 , \12122 , \12123 ,
         \12124 , \12125 , \12126 , \12127 , \12128 , \12129 , \12130 , \12131 , \12132 , \12133 ,
         \12134 , \12135 , \12136 , \12137 , \12138 , \12139 , \12140 , \12141 , \12142 , \12143 ,
         \12144 , \12145 , \12146 , \12147 , \12148 , \12149 , \12150 , \12151 , \12152 , \12153 ,
         \12154 , \12155 , \12156 , \12157 , \12158 , \12159 , \12160 , \12161 , \12162 , \12163 ,
         \12164 , \12165 , \12166 , \12167 , \12168 , \12169 , \12170 , \12171 , \12172 , \12173 ,
         \12174 , \12175 , \12176 , \12177 , \12178 , \12179 , \12180 , \12181 , \12182 , \12183 ,
         \12184 , \12185 , \12186 , \12187 , \12188 , \12189 , \12190 , \12191 , \12192 , \12193 ,
         \12194 , \12195 , \12196 , \12197 , \12198 , \12199 , \12200 , \12201 , \12202 , \12203 ,
         \12204 , \12205 , \12206 , \12207 , \12208 , \12209 , \12210 , \12211 , \12212 , \12213 ,
         \12214 , \12215 , \12216 , \12217 , \12218 , \12219 , \12220 , \12221 , \12222 , \12223 ,
         \12224 , \12225 , \12226 , \12227 , \12228 , \12229 , \12230 , \12231 , \12232 , \12233 ,
         \12234 , \12235 , \12236 , \12237 , \12238 , \12239 , \12240 , \12241 , \12242 , \12243 ,
         \12244 , \12245 , \12246 , \12247 , \12248 , \12249 , \12250 , \12251 , \12252 , \12253 ,
         \12254 , \12255 , \12256 , \12257 , \12258 , \12259 , \12260 , \12261 , \12262 , \12263 ,
         \12264 , \12265 , \12266 , \12267 , \12268 , \12269 , \12270 , \12271 , \12272 , \12273 ,
         \12274 , \12275 , \12276 , \12277 , \12278 , \12279 , \12280 , \12281 , \12282 , \12283 ,
         \12284 , \12285 , \12286 , \12287 , \12288 , \12289 , \12290 , \12291 , \12292 , \12293 ,
         \12294 , \12295 , \12296 , \12297 , \12298 , \12299 , \12300 , \12301 , \12302 , \12303 ,
         \12304 , \12305 , \12306 , \12307 , \12308 , \12309 , \12310 , \12311 , \12312 , \12313 ,
         \12314 , \12315 , \12316 , \12317 , \12318 , \12319 , \12320 , \12321 , \12322 , \12323 ,
         \12324 , \12325 , \12326 , \12327 , \12328 , \12329 , \12330 , \12331 , \12332 , \12333 ,
         \12334 , \12335 , \12336 , \12337 , \12338 , \12339 , \12340 , \12341 , \12342 , \12343 ,
         \12344 , \12345 , \12346 , \12347 , \12348 , \12349 , \12350 , \12351 , \12352 , \12353 ,
         \12354 , \12355 , \12356 , \12357 , \12358 , \12359 , \12360 , \12361 , \12362 , \12363 ,
         \12364 , \12365 , \12366 , \12367 , \12368 , \12369 , \12370 , \12371 , \12372 , \12373 ,
         \12374 , \12375 , \12376 , \12377 , \12378 , \12379 , \12380 , \12381 , \12382 , \12383 ,
         \12384 , \12385 , \12386 , \12387 , \12388 , \12389 , \12390 , \12391 , \12392 , \12393 ,
         \12394 , \12395 , \12396 , \12397 , \12398 , \12399 , \12400 , \12401 , \12402 , \12403 ,
         \12404 , \12405 , \12406 , \12407 , \12408 , \12409 , \12410 , \12411 , \12412 , \12413 ,
         \12414 , \12415 , \12416 , \12417 , \12418 , \12419 , \12420 , \12421 , \12422 , \12423 ,
         \12424 , \12425 , \12426 , \12427 , \12428 , \12429 , \12430 , \12431 , \12432 , \12433 ,
         \12434 , \12435 , \12436 , \12437 , \12438 , \12439 , \12440 , \12441 , \12442 , \12443 ,
         \12444 , \12445 , \12446 , \12447 , \12448 , \12449 , \12450 , \12451 , \12452 , \12453 ,
         \12454 , \12455 , \12456 , \12457 , \12458 , \12459 , \12460 , \12461 , \12462 , \12463 ,
         \12464 , \12465 , \12466 , \12467 , \12468 , \12469 , \12470 , \12471 , \12472 , \12473 ,
         \12474 , \12475 , \12476 , \12477 , \12478 , \12479 , \12480 , \12481 , \12482 , \12483 ,
         \12484 , \12485 , \12486 , \12487 , \12488 , \12489 , \12490 , \12491 , \12492 , \12493 ,
         \12494 , \12495 , \12496 , \12497 , \12498 , \12499 , \12500 , \12501 , \12502 , \12503 ,
         \12504 , \12505 , \12506 , \12507 , \12508 , \12509 , \12510 , \12511 , \12512 , \12513 ,
         \12514 , \12515 , \12516 , \12517 , \12518 , \12519 , \12520 , \12521 , \12522 , \12523 ,
         \12524 , \12525 , \12526 , \12527 , \12528 , \12529 , \12530 , \12531 , \12532 , \12533 ,
         \12534 , \12535 , \12536 , \12537 , \12538 , \12539 , \12540 , \12541 , \12542 , \12543 ,
         \12544 , \12545 , \12546 , \12547 , \12548 , \12549 , \12550 , \12551 , \12552 , \12553 ,
         \12554 , \12555 , \12556 , \12557 , \12558 , \12559 , \12560 , \12561 , \12562 , \12563 ,
         \12564 , \12565 , \12566 , \12567 , \12568 , \12569 , \12570 , \12571 , \12572 , \12573 ,
         \12574 , \12575 , \12576 , \12577 , \12578 , \12579 , \12580 , \12581 , \12582 , \12583 ,
         \12584 , \12585 , \12586 , \12587 , \12588 , \12589 , \12590 , \12591 , \12592 , \12593 ,
         \12594 , \12595 , \12596 , \12597 , \12598 , \12599 , \12600 , \12601 , \12602 , \12603 ,
         \12604 , \12605 , \12606 , \12607 , \12608 , \12609 , \12610 , \12611 , \12612 , \12613 ,
         \12614 , \12615 , \12616 , \12617 , \12618 , \12619 , \12620 , \12621 , \12622 , \12623 ,
         \12624 , \12625 , \12626 , \12627 , \12628 , \12629 , \12630 , \12631 , \12632 , \12633 ,
         \12634 , \12635 , \12636 , \12637 , \12638 , \12639 , \12640 , \12641 , \12642 , \12643 ,
         \12644 , \12645 , \12646 , \12647 , \12648 , \12649 , \12650 , \12651 , \12652 , \12653 ,
         \12654 , \12655 , \12656 , \12657 , \12658 , \12659 , \12660 , \12661 , \12662 , \12663 ,
         \12664 , \12665 , \12666 , \12667 , \12668 , \12669 , \12670 , \12671 , \12672 , \12673 ,
         \12674 , \12675 , \12676 , \12677 , \12678 , \12679 , \12680 , \12681 , \12682 , \12683 ,
         \12684 , \12685 , \12686 , \12687 , \12688 , \12689 , \12690 , \12691 , \12692 , \12693 ,
         \12694 , \12695 , \12696 , \12697 , \12698 , \12699 , \12700 , \12701 , \12702 , \12703 ,
         \12704 , \12705 , \12706 , \12707 , \12708 , \12709 , \12710 , \12711 , \12712 , \12713 ,
         \12714 , \12715 , \12716 , \12717 , \12718 , \12719 , \12720 , \12721 , \12722 , \12723 ,
         \12724 , \12725 , \12726 , \12727 , \12728 , \12729 , \12730 , \12731 , \12732 , \12733 ,
         \12734 , \12735 , \12736 , \12737 , \12738 , \12739 , \12740 , \12741 , \12742 , \12743 ,
         \12744 , \12745 , \12746 , \12747 , \12748 , \12749 , \12750 , \12751 , \12752 , \12753 ,
         \12754 , \12755 , \12756 , \12757 , \12758 , \12759 , \12760 , \12761 , \12762 , \12763 ,
         \12764 , \12765 , \12766 , \12767 , \12768 , \12769 , \12770 , \12771 , \12772 , \12773 ,
         \12774 , \12775 , \12776 , \12777 , \12778 , \12779 , \12780 , \12781 , \12782 , \12783 ,
         \12784 , \12785 , \12786 , \12787 , \12788 , \12789 , \12790 , \12791 , \12792 , \12793 ,
         \12794 , \12795 , \12796 , \12797 , \12798 , \12799 , \12800 , \12801 , \12802 , \12803 ,
         \12804 , \12805 , \12806 , \12807 , \12808 , \12809 , \12810 , \12811 , \12812 , \12813 ,
         \12814 , \12815 , \12816 , \12817 , \12818 , \12819 , \12820 , \12821 , \12822 , \12823 ,
         \12824 , \12825 , \12826 , \12827 , \12828 , \12829 , \12830 , \12831 , \12832 , \12833 ,
         \12834 , \12835 , \12836 , \12837 , \12838 , \12839 , \12840 , \12841 , \12842 , \12843 ,
         \12844 , \12845 , \12846 , \12847 , \12848 , \12849 , \12850 , \12851 , \12852 , \12853 ,
         \12854 , \12855 , \12856 , \12857 , \12858 , \12859 , \12860 , \12861 , \12862 , \12863 ,
         \12864 , \12865 , \12866 , \12867 , \12868 , \12869 , \12870 , \12871 , \12872 , \12873 ,
         \12874 , \12875 , \12876 , \12877 , \12878 , \12879 , \12880 , \12881 , \12882 , \12883 ,
         \12884 , \12885 , \12886 , \12887 , \12888 , \12889 , \12890 , \12891 , \12892 , \12893 ,
         \12894 , \12895 , \12896 , \12897 , \12898 , \12899 , \12900 , \12901 , \12902 , \12903 ,
         \12904 , \12905 , \12906 , \12907 , \12908 , \12909 , \12910 , \12911 , \12912 , \12913 ,
         \12914 , \12915 , \12916 , \12917 , \12918 , \12919 , \12920 , \12921 , \12922 , \12923 ,
         \12924 , \12925 , \12926 , \12927 , \12928 , \12929 , \12930 , \12931 , \12932 , \12933 ,
         \12934 , \12935 , \12936 , \12937 , \12938 , \12939 , \12940 , \12941 , \12942 , \12943 ,
         \12944 , \12945 , \12946 , \12947 , \12948 , \12949 , \12950 , \12951 , \12952 , \12953 ,
         \12954 , \12955 , \12956 , \12957 , \12958 , \12959 , \12960 , \12961 , \12962 , \12963 ,
         \12964 , \12965 , \12966 , \12967 , \12968 , \12969 , \12970 , \12971 , \12972 , \12973 ,
         \12974 , \12975 , \12976 , \12977 , \12978 , \12979 , \12980 , \12981 , \12982 , \12983 ,
         \12984 , \12985 , \12986 , \12987 , \12988 , \12989 , \12990 , \12991 , \12992 , \12993 ,
         \12994 , \12995 , \12996 , \12997 , \12998 , \12999 , \13000 , \13001 , \13002 , \13003 ,
         \13004 , \13005 , \13006 , \13007 , \13008 , \13009 , \13010 , \13011 , \13012 , \13013 ,
         \13014 , \13015 , \13016 , \13017 , \13018 , \13019 , \13020 , \13021 , \13022 , \13023 ,
         \13024 , \13025 , \13026 , \13027 , \13028 , \13029 , \13030 , \13031 , \13032 , \13033 ,
         \13034 , \13035 , \13036 , \13037 , \13038 , \13039 , \13040 , \13041 , \13042 , \13043 ,
         \13044 , \13045 , \13046 , \13047 , \13048 , \13049 , \13050 , \13051 , \13052 , \13053 ,
         \13054 , \13055 , \13056 , \13057 , \13058 , \13059 , \13060 , \13061 , \13062 , \13063 ,
         \13064 , \13065 , \13066 , \13067 , \13068 , \13069 , \13070 , \13071 , \13072 , \13073 ,
         \13074 , \13075 , \13076 , \13077 , \13078 , \13079 , \13080 , \13081 , \13082 , \13083 ,
         \13084 , \13085 , \13086 , \13087 , \13088 , \13089 , \13090 , \13091 , \13092 , \13093 ,
         \13094 , \13095 , \13096 , \13097 , \13098 , \13099 , \13100 , \13101 , \13102 , \13103 ,
         \13104 , \13105 , \13106 , \13107 , \13108 , \13109 , \13110 , \13111 , \13112 , \13113 ,
         \13114 , \13115 , \13116 , \13117 , \13118 , \13119 , \13120 , \13121 , \13122 , \13123 ,
         \13124 , \13125 , \13126 , \13127 , \13128 , \13129 , \13130 , \13131 , \13132 , \13133 ,
         \13134 , \13135 , \13136 , \13137 , \13138 , \13139 , \13140 , \13141 , \13142 , \13143 ,
         \13144 , \13145 , \13146 , \13147 , \13148 , \13149 , \13150 , \13151 , \13152 , \13153 ,
         \13154 , \13155 , \13156 , \13157 , \13158 , \13159 , \13160 , \13161 , \13162 , \13163 ,
         \13164 , \13165 , \13166 , \13167 , \13168 , \13169 , \13170 , \13171 , \13172 , \13173 ,
         \13174 , \13175 , \13176 , \13177 , \13178 , \13179 , \13180 , \13181 , \13182 , \13183 ,
         \13184 , \13185 , \13186 , \13187 , \13188 , \13189 , \13190 , \13191 , \13192 , \13193 ,
         \13194 , \13195 , \13196 , \13197 , \13198 , \13199 , \13200 , \13201 , \13202 , \13203 ,
         \13204 , \13205 , \13206 , \13207 , \13208 , \13209 , \13210 , \13211 , \13212 , \13213 ,
         \13214 , \13215 , \13216 , \13217 , \13218 , \13219 , \13220 , \13221 , \13222 , \13223 ,
         \13224 , \13225 , \13226 , \13227 , \13228 , \13229 , \13230 , \13231 , \13232 , \13233 ,
         \13234 , \13235 , \13236 , \13237 , \13238 , \13239 , \13240 , \13241 , \13242 , \13243 ,
         \13244 , \13245 , \13246 , \13247 , \13248 , \13249 , \13250 , \13251 , \13252 , \13253 ,
         \13254 , \13255 , \13256 , \13257 , \13258 , \13259 , \13260 , \13261 , \13262 , \13263 ,
         \13264 , \13265 , \13266 , \13267 , \13268 , \13269 , \13270 , \13271 , \13272 , \13273 ,
         \13274 , \13275 , \13276 , \13277 , \13278 , \13279 , \13280 , \13281 , \13282 , \13283 ,
         \13284 , \13285 , \13286 , \13287 , \13288 , \13289 , \13290 , \13291 , \13292 , \13293 ,
         \13294 , \13295 , \13296 , \13297 , \13298 , \13299 , \13300 , \13301 , \13302 , \13303 ,
         \13304 , \13305 , \13306 , \13307 , \13308 , \13309 , \13310 , \13311 , \13312 , \13313 ,
         \13314 , \13315 , \13316 , \13317 , \13318 , \13319 , \13320 , \13321 , \13322 , \13323 ,
         \13324 , \13325 , \13326 , \13327 , \13328 , \13329 , \13330 , \13331 , \13332 , \13333 ,
         \13334 , \13335 , \13336 , \13337 , \13338 , \13339 , \13340 , \13341 , \13342 , \13343 ,
         \13344 , \13345 , \13346 , \13347 , \13348 , \13349 , \13350 , \13351 , \13352 , \13353 ,
         \13354 , \13355 , \13356 , \13357 , \13358 , \13359 , \13360 , \13361 , \13362 , \13363 ,
         \13364 , \13365 , \13366 , \13367 , \13368 , \13369 , \13370 , \13371 , \13372 , \13373 ,
         \13374 , \13375 , \13376 , \13377 , \13378 , \13379 , \13380 , \13381 , \13382 , \13383 ,
         \13384 , \13385 , \13386 , \13387 , \13388 , \13389 , \13390 , \13391 , \13392 , \13393 ,
         \13394 , \13395 , \13396 , \13397 , \13398 , \13399 , \13400 , \13401 , \13402 , \13403 ,
         \13404 , \13405 , \13406 , \13407 , \13408 , \13409 , \13410 , \13411 , \13412 , \13413 ,
         \13414 , \13415 , \13416 , \13417 , \13418 , \13419 , \13420 , \13421 , \13422 , \13423 ,
         \13424 , \13425 , \13426 , \13427 , \13428 , \13429 , \13430 , \13431 , \13432 , \13433 ,
         \13434 , \13435 , \13436 , \13437 , \13438 , \13439 , \13440 , \13441 , \13442 , \13443 ,
         \13444 , \13445 , \13446 , \13447 , \13448 , \13449 , \13450 , \13451 , \13452 , \13453 ,
         \13454 , \13455 , \13456 , \13457 , \13458 , \13459 , \13460 , \13461 , \13462 , \13463 ,
         \13464 , \13465 , \13466 , \13467 , \13468 , \13469 , \13470 , \13471 , \13472 , \13473 ,
         \13474 , \13475 , \13476 , \13477 , \13478 , \13479 , \13480 , \13481 , \13482 , \13483 ,
         \13484 , \13485 , \13486 , \13487 , \13488 , \13489 , \13490 , \13491 , \13492 , \13493 ,
         \13494 , \13495 , \13496 , \13497 , \13498 , \13499 , \13500 , \13501 , \13502 , \13503 ,
         \13504 , \13505 , \13506 , \13507 , \13508 , \13509 , \13510 , \13511 , \13512 , \13513 ,
         \13514 , \13515 , \13516 , \13517 , \13518 , \13519 , \13520 , \13521 , \13522 , \13523 ,
         \13524 , \13525 , \13526 , \13527 , \13528 , \13529 , \13530 , \13531 , \13532 , \13533 ,
         \13534 , \13535 , \13536 , \13537 , \13538 , \13539 , \13540 , \13541 , \13542 , \13543 ,
         \13544 , \13545 , \13546 , \13547 , \13548 , \13549 , \13550 , \13551 , \13552 , \13553 ,
         \13554 , \13555 , \13556 , \13557 , \13558 , \13559 , \13560 , \13561 , \13562 , \13563 ,
         \13564 , \13565 , \13566 , \13567 , \13568 , \13569 , \13570 , \13571 , \13572 , \13573 ,
         \13574 , \13575 , \13576 , \13577 , \13578 , \13579 , \13580 , \13581 , \13582 , \13583 ,
         \13584 , \13585 , \13586 , \13587 , \13588 , \13589 , \13590 , \13591 , \13592 , \13593 ,
         \13594 , \13595 , \13596 , \13597 , \13598 , \13599 , \13600 , \13601 , \13602 , \13603 ,
         \13604 , \13605 , \13606 , \13607 , \13608 , \13609 , \13610 , \13611 , \13612 , \13613 ,
         \13614 , \13615 , \13616 , \13617 , \13618 , \13619 , \13620 , \13621 , \13622 , \13623 ,
         \13624 , \13625 , \13626 , \13627 , \13628 , \13629 , \13630 , \13631 , \13632 , \13633 ,
         \13634 , \13635 , \13636 , \13637 , \13638 , \13639 , \13640 , \13641 , \13642 , \13643 ,
         \13644 , \13645 , \13646 , \13647 , \13648 , \13649 , \13650 , \13651 , \13652 , \13653 ,
         \13654 , \13655 , \13656 , \13657 , \13658 , \13659 , \13660 , \13661 , \13662 , \13663 ,
         \13664 , \13665 , \13666 , \13667 , \13668 , \13669 , \13670 , \13671 , \13672 , \13673 ,
         \13674 , \13675 , \13676 , \13677 , \13678 , \13679 , \13680 , \13681 , \13682 , \13683 ,
         \13684 , \13685 , \13686 , \13687 , \13688 , \13689 , \13690 , \13691 , \13692 , \13693 ,
         \13694 , \13695 , \13696 , \13697 , \13698 , \13699 , \13700 , \13701 , \13702 , \13703 ,
         \13704 , \13705 , \13706 , \13707 , \13708 , \13709 , \13710 , \13711 , \13712 , \13713 ,
         \13714 , \13715 , \13716 , \13717 , \13718 , \13719 , \13720 , \13721 , \13722 , \13723 ,
         \13724 , \13725 , \13726 , \13727 , \13728 , \13729 , \13730 , \13731 , \13732 , \13733 ,
         \13734 , \13735 , \13736 , \13737 , \13738 , \13739 , \13740 , \13741 , \13742 , \13743 ,
         \13744 , \13745 , \13746 , \13747 , \13748 , \13749 , \13750 , \13751 , \13752 , \13753 ,
         \13754 , \13755 , \13756 , \13757 , \13758 , \13759 , \13760 , \13761 , \13762 , \13763 ,
         \13764 , \13765 , \13766 , \13767 , \13768 , \13769 , \13770 , \13771 , \13772 , \13773 ,
         \13774 , \13775 , \13776 , \13777 , \13778 , \13779 , \13780 , \13781 , \13782 , \13783 ,
         \13784 , \13785 , \13786 , \13787 , \13788 , \13789 , \13790 , \13791 , \13792 , \13793 ,
         \13794 , \13795 , \13796 , \13797 , \13798 , \13799 , \13800 , \13801 , \13802 , \13803 ,
         \13804 , \13805 , \13806 , \13807 , \13808 , \13809 , \13810 , \13811 , \13812 , \13813 ,
         \13814 , \13815 , \13816 , \13817 , \13818 , \13819 , \13820 , \13821 , \13822 , \13823 ,
         \13824 , \13825 , \13826 , \13827 , \13828 , \13829 , \13830 , \13831 , \13832 , \13833 ,
         \13834 , \13835 , \13836 , \13837 , \13838 , \13839 , \13840 , \13841 , \13842 , \13843 ,
         \13844 , \13845 , \13846 , \13847 , \13848 , \13849 , \13850 , \13851 , \13852 , \13853 ,
         \13854 , \13855 , \13856 , \13857 , \13858 , \13859 , \13860 , \13861 , \13862 , \13863 ,
         \13864 , \13865 , \13866 , \13867 , \13868 , \13869 , \13870 , \13871 , \13872 , \13873 ,
         \13874 , \13875 , \13876 , \13877 , \13878 , \13879 , \13880 , \13881 , \13882 , \13883 ,
         \13884 , \13885 , \13886 , \13887 , \13888 , \13889 , \13890 , \13891 , \13892 , \13893 ,
         \13894 , \13895 , \13896 , \13897 , \13898 , \13899 , \13900 , \13901 , \13902 , \13903 ,
         \13904 , \13905 , \13906 , \13907 , \13908 , \13909 , \13910 , \13911 , \13912 , \13913 ,
         \13914 , \13915 , \13916 , \13917 , \13918 , \13919 , \13920 , \13921 , \13922 , \13923 ,
         \13924 , \13925 , \13926 , \13927 , \13928 , \13929 , \13930 , \13931 , \13932 , \13933 ,
         \13934 , \13935 , \13936 , \13937 , \13938 , \13939 , \13940 , \13941 , \13942 , \13943 ,
         \13944 , \13945 , \13946 , \13947 , \13948 , \13949 , \13950 , \13951 , \13952 , \13953 ,
         \13954 , \13955 , \13956 , \13957 , \13958 , \13959 , \13960 , \13961 , \13962 , \13963 ,
         \13964 , \13965 , \13966 , \13967 , \13968 , \13969 , \13970 , \13971 , \13972 , \13973 ,
         \13974 , \13975 , \13976 , \13977 , \13978 , \13979 , \13980 , \13981 , \13982 , \13983 ,
         \13984 , \13985 , \13986 , \13987 , \13988 , \13989 , \13990 , \13991 , \13992 , \13993 ,
         \13994 , \13995 , \13996 , \13997 , \13998 , \13999 , \14000 , \14001 , \14002 , \14003 ,
         \14004 , \14005 , \14006 , \14007 , \14008 , \14009 , \14010 , \14011 , \14012 , \14013_nG36c1 ,
         \14014 , \14015 , \14016 , \14017 , \14018 , \14019 , \14020 , \14021 , \14022 , \14023 ,
         \14024 , \14025 , \14026 , \14027 , \14028 , \14029 , \14030 , \14031 , \14032 , \14033 ,
         \14034 , \14035 , \14036 , \14037 , \14038 , \14039 , \14040 , \14041 , \14042 , \14043 ,
         \14044 , \14045 , \14046 , \14047 , \14048 , \14049 , \14050 , \14051 , \14052 , \14053 ,
         \14054 , \14055 , \14056 , \14057 , \14058 , \14059 , \14060 , \14061 , \14062 , \14063 ,
         \14064 , \14065 , \14066 , \14067 , \14068 , \14069 , \14070 , \14071 , \14072 , \14073 ,
         \14074 , \14075 , \14076 , \14077 , \14078 , \14079 , \14080 , \14081 , \14082 , \14083 ,
         \14084 , \14085 , \14086 , \14087 , \14088 , \14089 , \14090 , \14091 , \14092 , \14093 ,
         \14094 , \14095 , \14096 , \14097 , \14098 , \14099 , \14100 , \14101 , \14102 , \14103 ,
         \14104 , \14105 , \14106 , \14107 , \14108 , \14109 , \14110 , \14111 , \14112 , \14113 ,
         \14114 , \14115 , \14116 , \14117 , \14118 , \14119 , \14120 , \14121 , \14122 , \14123 ,
         \14124 , \14125 , \14126 , \14127 , \14128 , \14129 , \14130 , \14131 , \14132 , \14133 ,
         \14134 , \14135 , \14136 , \14137 , \14138 , \14139 , \14140 , \14141 , \14142 , \14143 ,
         \14144 , \14145 , \14146 , \14147 , \14148 , \14149 , \14150 , \14151 , \14152 , \14153 ,
         \14154 , \14155 , \14156 , \14157 , \14158 , \14159 , \14160 , \14161 , \14162 , \14163 ,
         \14164 , \14165 , \14166 , \14167 , \14168 , \14169 , \14170 , \14171 , \14172 , \14173 ,
         \14174 , \14175 , \14176 , \14177 , \14178 , \14179 , \14180 , \14181 , \14182 , \14183 ,
         \14184 , \14185 , \14186 , \14187 , \14188 , \14189 , \14190 , \14191 , \14192 , \14193 ,
         \14194 , \14195_nG3776 , \14196 , \14197 , \14198 , \14199 , \14200 , \14201 , \14202 , \14203 ,
         \14204 , \14205 , \14206 , \14207 , \14208 , \14209 , \14210 , \14211 , \14212 , \14213 ,
         \14214 , \14215 , \14216 , \14217 , \14218 , \14219 , \14220 , \14221 , \14222 , \14223 ,
         \14224 , \14225 , \14226 , \14227 , \14228 , \14229 , \14230 , \14231 , \14232 , \14233 ,
         \14234 , \14235 , \14236 , \14237 , \14238 , \14239 , \14240 , \14241 , \14242 , \14243 ,
         \14244 , \14245 , \14246 , \14247 , \14248 , \14249 , \14250 , \14251 , \14252 , \14253 ,
         \14254 , \14255 , \14256 , \14257 , \14258 , \14259 , \14260 , \14261 , \14262 , \14263 ,
         \14264 , \14265 , \14266 , \14267 , \14268 , \14269 , \14270 , \14271 , \14272 , \14273 ,
         \14274 , \14275 , \14276 , \14277 , \14278 , \14279 , \14280 , \14281 , \14282 , \14283 ,
         \14284 , \14285_nG37cf , \14286 , \14287 , \14288 , \14289 , \14290 , \14291 , \14292 , \14293 ,
         \14294 , \14295 , \14296 , \14297 , \14298 , \14299 , \14300 , \14301 , \14302 , \14303 ,
         \14304 , \14305 , \14306 , \14307 , \14308 , \14309 , \14310 , \14311 , \14312 , \14313 ,
         \14314 , \14315 , \14316 , \14317 , \14318 , \14319 , \14320 , \14321 , \14322 , \14323 ,
         \14324 , \14325 , \14326 , \14327 , \14328 , \14329 , \14330 , \14331 , \14332 , \14333 ,
         \14334 , \14335 , \14336 , \14337 , \14338 , \14339 , \14340 , \14341 , \14342 , \14343 ,
         \14344 , \14345 , \14346 , \14347 , \14348 , \14349 , \14350 , \14351 , \14352 , \14353 ,
         \14354 , \14355 , \14356 , \14357 , \14358 , \14359 , \14360 , \14361 , \14362 , \14363 ,
         \14364 , \14365 , \14366 , \14367 , \14368 , \14369 , \14370 , \14371 , \14372 , \14373 ,
         \14374 , \14375 , \14376_nG3829 , \14377 , \14378 , \14379 , \14380 , \14381 , \14382 , \14383 ,
         \14384 , \14385 , \14386 , \14387 , \14388 , \14389 , \14390 , \14391 , \14392 , \14393 ,
         \14394 , \14395 , \14396 , \14397 , \14398 , \14399 , \14400 , \14401 , \14402 , \14403 ,
         \14404 , \14405 , \14406 , \14407 , \14408 , \14409 , \14410 , \14411 , \14412 , \14413 ,
         \14414 , \14415 , \14416 , \14417 , \14418 , \14419 , \14420 , \14421_nG3855 , \14422 , \14423 ,
         \14424 , \14425 , \14426 , \14427 , \14428 , \14429 , \14430 , \14431 , \14432 , \14433 ,
         \14434 , \14435 , \14436 , \14437 , \14438 , \14439 , \14440 , \14441 , \14442 , \14443 ,
         \14444 , \14445 , \14446 , \14447 , \14448 , \14449 , \14450 , \14451 , \14452 , \14453 ,
         \14454 , \14455 , \14456 , \14457 , \14458 , \14459 , \14460 , \14461 , \14462 , \14463 ,
         \14464 , \14465 , \14466_nG3881 , \14467 , \14468 , \14469 , \14470 , \14471 , \14472 , \14473 ,
         \14474 , \14475 , \14476 , \14477 , \14478 , \14479 , \14480 , \14481 , \14482 , \14483 ,
         \14484 , \14485 , \14486 , \14487 , \14488 , \14489 , \14490 , \14491 , \14492 , \14493 ,
         \14494 , \14495 , \14496 , \14497 , \14498 , \14499 , \14500 , \14501 , \14502 , \14503 ,
         \14504 , \14505 , \14506 , \14507 , \14508 , \14509_nG38ab , \14510 , \14511 , \14512 , \14513 ,
         \14514 , \14515 , \14516 , \14517 , \14518 , \14519 , \14520 , \14521 , \14522 , \14523 ,
         \14524 , \14525 , \14526 , \14527 , \14528 , \14529 , \14530 , \14531 , \14532 , \14533 ,
         \14534 , \14535 , \14536 , \14537 , \14538 , \14539 , \14540 , \14541 , \14542 , \14543 ,
         \14544 , \14545 , \14546 , \14547 , \14548 , \14549 , \14550 , \14551 , \14552_nG38d5 , \14553 ,
         \14554 , \14555 , \14556 , \14557 , \14558 , \14559 , \14560 , \14561 , \14562 , \14563 ,
         \14564 , \14565 , \14566 , \14567 , \14568 , \14569 , \14570 , \14571 , \14572 , \14573 ,
         \14574 , \14575_nG38eb , \14576 , \14577 , \14578 , \14579 , \14580 , \14581 , \14582 , \14583 ,
         \14584 , \14585 , \14586 , \14587 , \14588 , \14589 , \14590 , \14591 , \14592 , \14593 ,
         \14594 , \14595 , \14596 , \14597 , \14598_nG3901 , \14599 , \14600 , \14601 , \14602 , \14603 ,
         \14604 , \14605 , \14606 , \14607 , \14608 , \14609 , \14610 , \14611 , \14612 , \14613 ,
         \14614 , \14615 , \14616 , \14617 , \14618 , \14619 , \14620_nG3916 , \14621 , \14622 , \14623 ,
         \14624 , \14625 , \14626 , \14627 , \14628 , \14629 , \14630 , \14631 , \14632 , \14633 ,
         \14634 , \14635 , \14636 , \14637 , \14638 , \14639 , \14640 , \14641 , \14642_nG392b , \14643 ,
         \14644 , \14645 , \14646 , \14647 , \14648 , \14649 , \14650 , \14651 , \14652 , \14653 ,
         \14654 , \14655 , \14656 , \14657 , \14658 , \14659 , \14660 , \14661 , \14662 , \14663 ,
         \14664_nG3940 , \14665 , \14666 , \14667 , \14668 , \14669 , \14670 , \14671 , \14672 , \14673 ,
         \14674 , \14675 , \14676 , \14677 , \14678 , \14679 , \14680 , \14681 , \14682 , \14683 ,
         \14684 , \14685 , \14686_nG3955 , \14687 , \14688 , \14689 , \14690 , \14691 , \14692 , \14693 ,
         \14694 , \14695 , \14696 , \14697 , \14698 , \14699 , \14700 , \14701 , \14702 , \14703 ,
         \14704 , \14705 , \14706_nG3968 , \14707 , \14708 , \14709 , \14710 , \14711 , \14712 , \14713 ,
         \14714 , \14715 , \14716 , \14717 , \14718 , \14719 , \14720 , \14721 , \14722 , \14723 ,
         \14724 , \14725 , \14726_nG397b , \14727 , \14728 , \14729 , \14730 , \14731 , \14732 , \14733 ,
         \14734 , \14735 , \14736 , \14737 , \14738_nG3986 , \14739 , \14740 , \14741 , \14742 , \14743 ,
         \14744 , \14745 , \14746 , \14747 , \14748 , \14749 , \14750_nG3991 , \14751 , \14752 , \14753 ,
         \14754 , \14755 , \14756 , \14757 , \14758 , \14759 , \14760 , \14761 , \14762_nG399c , \14763 ,
         \14764 , \14765 , \14766 , \14767 , \14768 , \14769 , \14770 , \14771 , \14772 , \14773 ,
         \14774_nG39a7 , \14775 , \14776 , \14777 , \14778 , \14779 , \14780 , \14781 , \14782 , \14783 ,
         \14784 , \14785 , \14786_nG39b2 , \14787 , \14788 , \14789 , \14790 , \14791 , \14792 , \14793 ,
         \14794 , \14795 , \14796 , \14797 , \14798_nG39bd , \14799 , \14800 , \14801 , \14802 , \14803 ,
         \14804 , \14805 , \14806 , \14807 , \14808 , \14809_nG39c7 , \14810 , \14811 , \14812 , \14813 ,
         \14814 , \14815 , \14816 , \14817 , \14818 , \14819 , \14820_nG39d1 , \14821 , \14822 , \14823 ,
         \14824 , \14825 , \14826 , \14827 , \14828 , \14829 , \14830 , \14831_nG39db , \14832 , \14833 ,
         \14834 , \14835 , \14836 , \14837 , \14838 , \14839 , \14840 , \14841 , \14842_nG39e5 , \14843 ,
         \14844 , \14845 , \14846 , \14847 , \14848 , \14849 , \14850 , \14851 , \14852 , \14853_nG39ef ,
         \14854 , \14855 , \14856 , \14857 , \14858 , \14859 , \14860 , \14861 , \14862 , \14863 ,
         \14864_nG39f9 , \14865 , \14866 , \14867 , \14868 , \14869 , \14870 , \14871 , \14872 , \14873 ,
         \14874 , \14875_nG3a03 , \14876 , \14877 , \14878 , \14879 , \14880 , \14881 , \14882 , \14883 ,
         \14884 , \14885 , \14886_nG3a0d , \14887 , \14888 , \14889 , \14890 , \14891 , \14892 , \14893_nG3a13 ,
         \14894 , \14895 , \14896 , \14897 , \14898 , \14899 , \14900_nG3a19 , \14901 , \14902 , \14903 ,
         \14904 , \14905_nG3a1d , \14906 , \14907 , \14908 , \14909 , \14910_nG3a21 , \14911 , \14912 , \14913 ,
         \14914 , \14915_nG3a25 , \14916 , \14917 , \14918 , \14919 , \14920_nG3a29 , \14921 , \14922 , \14923 ,
         \14924 , \14925_nG3a2d , \14926 , \14927 , \14928 , \14929 , \14930_nG3a31 , \14931 , \14932 , \14933 ,
         \14934 , \14935_nG3a35 , \14936 , \14937 , \14938 , \14939 , \14940_nG3a39 , \14941 , \14942 , \14943 ,
         \14944 , \14945_nG3a3d , \14946 , \14947 , \14948 , \14949 , \14950_nG3a41 , \14951 , \14952 , \14953 ,
         \14954 , \14955_nG3a45 , \14956 , \14957 , \14958 , \14959 , \14960_nG3a49 , \14961 , \14962 , \14963 ,
         \14964 , \14965_nG3a4d , \14966 , \14967 , \14968 , \14969 , \14970_nG3a51 , \14971 , \14972 , \14973 ,
         \14974 , \14975_nG3a55 , \14976 , \14977 , \14978 , \14979 , \14980_nG3a59 , \14981 , \14982 , \14983 ,
         \14984 , \14985_nG3a5d , \14986 , \14987 , \14988 , \14989 , \14990_nG3a61 , \14991 , \14992 , \14993 ,
         \14994 , \14995_nG3a65 , \14996 , \14997 , \14998 , \14999 , \15000_nG3a69 , \15001 , \15002 , \15003 ,
         \15004 , \15005_nG3a6d , \15006 , \15007 , \15008 , \15009 , \15010_nG3a71 , \15011 , \15012 , \15013 ,
         \15014 , \15015_nG3a75 , \15016 , \15017 , \15018 , \15019 , \15020_nG3a79 , \15021 , \15022 , \15023 ,
         \15024 , \15025_nG3a7d , \15026 , \15027 , \15028 , \15029 , \15030_nG3a81 , \15031 ;
buf \U$labaj1525 ( R_61_85b54e8, \14014 );
buf \U$labaj1526 ( R_62_85b5590, \14196 );
buf \U$labaj1527 ( R_63_85b5638, \14286 );
buf \U$labaj1528 ( R_64_85b56e0, \14377 );
buf \U$labaj1529 ( R_65_85b5788, \14422 );
buf \U$labaj1530 ( R_66_85b5830, \14467 );
buf \U$labaj1531 ( R_67_85b58d8, \14510 );
buf \U$labaj1532 ( R_68_85b5980, \14553 );
buf \U$labaj1533 ( R_69_85b5a28, \14576 );
buf \U$labaj1534 ( R_6a_85b5ad0, \14599 );
buf \U$labaj1535 ( R_6b_85b5b78, \14621 );
buf \U$labaj1536 ( R_6c_85b5c20, \14643 );
buf \U$labaj1537 ( R_6d_85b5cc8, \14665 );
buf \U$labaj1538 ( R_6e_85b5d70, \14687 );
buf \U$labaj1539 ( R_6f_85b5e18, \14707 );
buf \U$labaj1540 ( R_70_85b5ec0, \14727 );
buf \U$labaj1541 ( R_71_85b5f68, \14739 );
buf \U$labaj1542 ( R_72_85b6010, \14751 );
buf \U$labaj1543 ( R_73_85b60b8, \14763 );
buf \U$labaj1544 ( R_74_85b6160, \14775 );
buf \U$labaj1545 ( R_75_85b6208, \14787 );
buf \U$labaj1546 ( R_76_85b62b0, \14799 );
buf \U$labaj1547 ( R_77_85b6358, \14810 );
buf \U$labaj1548 ( R_78_85b6400, \14821 );
buf \U$labaj1549 ( R_79_85b64a8, \14832 );
buf \U$labaj1550 ( R_7a_85b6550, \14843 );
buf \U$labaj1551 ( R_7b_85b65f8, \14854 );
buf \U$labaj1552 ( R_7c_85b66a0, \14865 );
buf \U$labaj1553 ( R_7d_85b6748, \14876 );
buf \U$labaj1554 ( R_7e_85b67f0, \14887 );
buf \U$labaj1555 ( R_7f_85b6898, \14894 );
buf \U$labaj1556 ( R_80_85b6940, \14901 );
buf \U$labaj1557 ( R_81_85b69e8, \14906 );
buf \U$labaj1558 ( R_82_85b6a90, \14911 );
buf \U$labaj1559 ( R_83_85b6b38, \14916 );
buf \U$labaj1560 ( R_84_85b6be0, \14921 );
buf \U$labaj1561 ( R_85_85b6c88, \14926 );
buf \U$labaj1562 ( R_86_85b6d30, \14931 );
buf \U$labaj1563 ( R_87_85b6dd8, \14936 );
buf \U$labaj1564 ( R_88_85b6e80, \14941 );
buf \U$labaj1565 ( R_89_85b6f28, \14946 );
buf \U$labaj1566 ( R_8a_85b6fd0, \14951 );
buf \U$labaj1567 ( R_8b_85b7078, \14956 );
buf \U$labaj1568 ( R_8c_85b7120, \14961 );
buf \U$labaj1569 ( R_8d_85b71c8, \14966 );
buf \U$labaj1570 ( R_8e_85b7270, \14971 );
buf \U$labaj1571 ( R_8f_85b7318, \14976 );
buf \U$labaj1572 ( R_90_85b73c0, \14981 );
buf \U$labaj1573 ( R_91_85b7468, \14986 );
buf \U$labaj1574 ( R_92_85b7510, \14991 );
buf \U$labaj1575 ( R_93_85b75b8, \14996 );
buf \U$labaj1576 ( R_94_85b7660, \15001 );
buf \U$labaj1577 ( R_95_85b7708, \15006 );
buf \U$labaj1578 ( R_96_85b77b0, \15011 );
buf \U$labaj1579 ( R_97_85b7858, \15016 );
buf \U$labaj1580 ( R_98_85b7900, \15021 );
buf \U$labaj1581 ( R_99_85b79a8, \15026 );
buf \U$labaj1582 ( R_9a_85b7a50, \15031 );
buf \U$1 ( \159 , RIa167a08_1);
buf \U$2 ( \160 , RIb4ca3e8_33);
xor \U$3 ( \161 , \159 , \160 );
buf \U$4 ( \162 , RIa167990_2);
buf \U$5 ( \163 , RIb4c6c20_34);
xor \U$6 ( \164 , \162 , \163 );
or \U$7 ( \165 , \161 , \164 );
buf \U$8 ( \166 , RIa167918_3);
buf \U$9 ( \167 , RIb4c6ba8_35);
xor \U$10 ( \168 , \166 , \167 );
or \U$11 ( \169 , \165 , \168 );
buf \U$12 ( \170 , RIa1678a0_4);
buf \U$13 ( \171 , RIb4c6b30_36);
xor \U$14 ( \172 , \170 , \171 );
or \U$15 ( \173 , \169 , \172 );
buf \U$16 ( \174 , RIa167828_5);
buf \U$17 ( \175 , RIb4c6ab8_37);
xor \U$18 ( \176 , \174 , \175 );
or \U$19 ( \177 , \173 , \176 );
buf \U$20 ( \178 , RIa1677b0_6);
buf \U$21 ( \179 , RIb4c6a40_38);
xor \U$22 ( \180 , \178 , \179 );
or \U$23 ( \181 , \177 , \180 );
buf \U$24 ( \182 , RIa167738_7);
buf \U$25 ( \183 , RIb4c69c8_39);
xor \U$26 ( \184 , \182 , \183 );
or \U$27 ( \185 , \181 , \184 );
buf \U$28 ( \186 , RIa1676c0_8);
buf \U$29 ( \187 , RIb4c6950_40);
xor \U$30 ( \188 , \186 , \187 );
or \U$31 ( \189 , \185 , \188 );
buf \U$32 ( \190 , RIa167648_9);
buf \U$33 ( \191 , RIb4c68d8_41);
xor \U$34 ( \192 , \190 , \191 );
or \U$35 ( \193 , \189 , \192 );
buf \U$36 ( \194 , RIa1675d0_10);
buf \U$37 ( \195 , RIb4c6860_42);
xor \U$38 ( \196 , \194 , \195 );
or \U$39 ( \197 , \193 , \196 );
buf \U$40 ( \198 , RIa167558_11);
buf \U$41 ( \199 , RIb4c67e8_43);
xor \U$42 ( \200 , \198 , \199 );
or \U$43 ( \201 , \197 , \200 );
buf \U$44 ( \202 , RIa1674e0_12);
buf \U$45 ( \203 , RIb4c6770_44);
xor \U$46 ( \204 , \202 , \203 );
or \U$47 ( \205 , \201 , \204 );
buf \U$48 ( \206 , RIa167468_13);
buf \U$49 ( \207 , RIb4c3368_45);
xor \U$50 ( \208 , \206 , \207 );
or \U$51 ( \209 , \205 , \208 );
buf \U$52 ( \210 , RIa1673f0_14);
buf \U$53 ( \211 , RIb4c32f0_46);
xor \U$54 ( \212 , \210 , \211 );
or \U$55 ( \213 , \209 , \212 );
buf \U$56 ( \214 , RIa167378_15);
buf \U$57 ( \215 , RIb4c3278_47);
xor \U$58 ( \216 , \214 , \215 );
or \U$59 ( \217 , \213 , \216 );
buf \U$60 ( \218 , RIa167300_16);
buf \U$61 ( \219 , RIb4c3200_48);
xor \U$62 ( \220 , \218 , \219 );
or \U$63 ( \221 , \217 , \220 );
buf \U$64 ( \222 , RIa167288_17);
buf \U$65 ( \223 , RIb4c3188_49);
xor \U$66 ( \224 , \222 , \223 );
or \U$67 ( \225 , \221 , \224 );
buf \U$68 ( \226 , RIa167210_18);
buf \U$69 ( \227 , RIb4c3110_50);
xor \U$70 ( \228 , \226 , \227 );
or \U$71 ( \229 , \225 , \228 );
buf \U$72 ( \230 , RIa167198_19);
buf \U$73 ( \231 , RIb4c3098_51);
xor \U$74 ( \232 , \230 , \231 );
or \U$75 ( \233 , \229 , \232 );
buf \U$76 ( \234 , RIa167120_20);
buf \U$77 ( \235 , RIb4c3020_52);
xor \U$78 ( \236 , \234 , \235 );
or \U$79 ( \237 , \233 , \236 );
buf \U$80 ( \238 , RIa1670a8_21);
buf \U$81 ( \239 , RIb4c2fa8_53);
xor \U$82 ( \240 , \238 , \239 );
or \U$83 ( \241 , \237 , \240 );
buf \U$84 ( \242 , RIa167030_22);
buf \U$85 ( \243 , RIb4c2f30_54);
xor \U$86 ( \244 , \242 , \243 );
or \U$87 ( \245 , \241 , \244 );
buf \U$88 ( \246 , RIa166fb8_23);
buf \U$89 ( \247 , RIb4c2eb8_55);
xor \U$90 ( \248 , \246 , \247 );
or \U$91 ( \249 , \245 , \248 );
buf \U$92 ( \250 , RIa166f40_24);
buf \U$93 ( \251 , RIb4c2e40_56);
xor \U$94 ( \252 , \250 , \251 );
or \U$95 ( \253 , \249 , \252 );
buf \U$96 ( \254 , RIa166ec8_25);
buf \U$97 ( \255 , RIb4c2dc8_57);
xor \U$98 ( \256 , \254 , \255 );
or \U$99 ( \257 , \253 , \256 );
buf \U$100 ( \258 , RIa166e50_26);
buf \U$101 ( \259 , RIb4c2d50_58);
xor \U$102 ( \260 , \258 , \259 );
or \U$103 ( \261 , \257 , \260 );
buf \U$104 ( \262 , RIa166dd8_27);
buf \U$105 ( \263 , RIb4c2cd8_59);
xor \U$106 ( \264 , \262 , \263 );
or \U$107 ( \265 , \261 , \264 );
buf \U$108 ( \266 , RIa166d60_28);
buf \U$109 ( \267 , RIb4c2c60_60);
xor \U$110 ( \268 , \266 , \267 );
or \U$111 ( \269 , \265 , \268 );
buf \U$112 ( \270 , RIa166ce8_29);
buf \U$113 ( \271 , RIb4c2be8_61);
xor \U$114 ( \272 , \270 , \271 );
or \U$115 ( \273 , \269 , \272 );
buf \U$116 ( \274 , RIa166c70_30);
buf \U$117 ( \275 , RIb4c2b70_62);
xor \U$118 ( \276 , \274 , \275 );
or \U$119 ( \277 , \273 , \276 );
buf \U$120 ( \278 , RIb4ca4d8_31);
buf \U$121 ( \279 , RIb4c2af8_63);
xor \U$122 ( \280 , \278 , \279 );
or \U$123 ( \281 , \277 , \280 );
buf \U$124 ( \282 , RIb4ca460_32);
buf \U$125 ( \283 , RIb4bfab0_64);
xor \U$126 ( \284 , \282 , \283 );
or \U$127 ( \285 , \281 , \284 );
not \U$128 ( \286 , \285 );
buf \U$129 ( \287 , \286 );
_DC g143 ( \288_nG143 , RIb4ca3e8_33 , \287 );
buf \U$130 ( \289 , \288_nG143 );
buf \U$131 ( \290 , RIa167738_7);
buf \U$132 ( \291 , RIa1676c0_8);
xor \U$133 ( \292 , \290 , \291 );
buf \U$134 ( \293 , RIa167648_9);
xor \U$135 ( \294 , \291 , \293 );
not \U$136 ( \295 , \294 );
and \U$137 ( \296 , \292 , \295 );
and \U$138 ( \297 , \289 , \296 );
not \U$139 ( \298 , \297 );
and \U$140 ( \299 , \291 , \293 );
not \U$141 ( \300 , \299 );
and \U$142 ( \301 , \290 , \300 );
xnor \U$143 ( \302 , \298 , \301 );
_DC g141 ( \303_nG141 , RIb4c6ba8_35 , \287 );
buf \U$144 ( \304 , \303_nG141 );
buf \U$145 ( \305 , RIa167828_5);
buf \U$146 ( \306 , RIa1677b0_6);
xor \U$147 ( \307 , \305 , \306 );
xor \U$148 ( \308 , \306 , \290 );
not \U$149 ( \309 , \308 );
and \U$150 ( \310 , \307 , \309 );
and \U$151 ( \311 , \304 , \310 );
_DC g142 ( \312_nG142 , RIb4c6c20_34 , \287 );
buf \U$152 ( \313 , \312_nG142 );
and \U$153 ( \314 , \313 , \308 );
nor \U$154 ( \315 , \311 , \314 );
and \U$155 ( \316 , \306 , \290 );
not \U$156 ( \317 , \316 );
and \U$157 ( \318 , \305 , \317 );
xnor \U$158 ( \319 , \315 , \318 );
and \U$159 ( \320 , \302 , \319 );
_DC g13f ( \321_nG13f , RIb4c6ab8_37 , \287 );
buf \U$160 ( \322 , \321_nG13f );
buf \U$161 ( \323 , RIa167918_3);
buf \U$162 ( \324 , RIa1678a0_4);
xor \U$163 ( \325 , \323 , \324 );
xor \U$164 ( \326 , \324 , \305 );
not \U$165 ( \327 , \326 );
and \U$166 ( \328 , \325 , \327 );
and \U$167 ( \329 , \322 , \328 );
_DC g140 ( \330_nG140 , RIb4c6b30_36 , \287 );
buf \U$168 ( \331 , \330_nG140 );
and \U$169 ( \332 , \331 , \326 );
nor \U$170 ( \333 , \329 , \332 );
and \U$171 ( \334 , \324 , \305 );
not \U$172 ( \335 , \334 );
and \U$173 ( \336 , \323 , \335 );
xnor \U$174 ( \337 , \333 , \336 );
and \U$175 ( \338 , \319 , \337 );
and \U$176 ( \339 , \302 , \337 );
or \U$177 ( \340 , \320 , \338 , \339 );
_DC g13d ( \341_nG13d , RIb4c69c8_39 , \287 );
buf \U$178 ( \342 , \341_nG13d );
buf \U$179 ( \343 , RIa167a08_1);
buf \U$180 ( \344 , RIa167990_2);
xor \U$181 ( \345 , \343 , \344 );
xor \U$182 ( \346 , \344 , \323 );
not \U$183 ( \347 , \346 );
and \U$184 ( \348 , \345 , \347 );
and \U$185 ( \349 , \342 , \348 );
_DC g13e ( \350_nG13e , RIb4c6a40_38 , \287 );
buf \U$186 ( \351 , \350_nG13e );
and \U$187 ( \352 , \351 , \346 );
nor \U$188 ( \353 , \349 , \352 );
and \U$189 ( \354 , \344 , \323 );
not \U$190 ( \355 , \354 );
and \U$191 ( \356 , \343 , \355 );
xnor \U$192 ( \357 , \353 , \356 );
_DC g13c ( \358_nG13c , RIb4c6950_40 , \287 );
buf \U$193 ( \359 , \358_nG13c );
and \U$194 ( \360 , \359 , \343 );
or \U$195 ( \361 , \357 , \360 );
and \U$196 ( \362 , \340 , \361 );
and \U$197 ( \363 , \351 , \348 );
and \U$198 ( \364 , \322 , \346 );
nor \U$199 ( \365 , \363 , \364 );
xnor \U$200 ( \366 , \365 , \356 );
and \U$201 ( \367 , \361 , \366 );
and \U$202 ( \368 , \340 , \366 );
or \U$203 ( \369 , \362 , \367 , \368 );
and \U$204 ( \370 , \342 , \343 );
not \U$205 ( \371 , \301 );
and \U$206 ( \372 , \313 , \310 );
and \U$207 ( \373 , \289 , \308 );
nor \U$208 ( \374 , \372 , \373 );
xnor \U$209 ( \375 , \374 , \318 );
xor \U$210 ( \376 , \371 , \375 );
and \U$211 ( \377 , \331 , \328 );
and \U$212 ( \378 , \304 , \326 );
nor \U$213 ( \379 , \377 , \378 );
xnor \U$214 ( \380 , \379 , \336 );
xor \U$215 ( \381 , \376 , \380 );
and \U$216 ( \382 , \370 , \381 );
and \U$217 ( \383 , \369 , \382 );
and \U$218 ( \384 , \371 , \375 );
and \U$219 ( \385 , \375 , \380 );
and \U$220 ( \386 , \371 , \380 );
or \U$221 ( \387 , \384 , \385 , \386 );
and \U$222 ( \388 , \289 , \310 );
not \U$223 ( \389 , \388 );
xnor \U$224 ( \390 , \389 , \318 );
and \U$225 ( \391 , \304 , \328 );
and \U$226 ( \392 , \313 , \326 );
nor \U$227 ( \393 , \391 , \392 );
xnor \U$228 ( \394 , \393 , \336 );
xor \U$229 ( \395 , \390 , \394 );
and \U$230 ( \396 , \322 , \348 );
and \U$231 ( \397 , \331 , \346 );
nor \U$232 ( \398 , \396 , \397 );
xnor \U$233 ( \399 , \398 , \356 );
xor \U$234 ( \400 , \395 , \399 );
xor \U$235 ( \401 , \387 , \400 );
and \U$236 ( \402 , \351 , \343 );
not \U$237 ( \403 , \402 );
xor \U$238 ( \404 , \401 , \403 );
and \U$239 ( \405 , \382 , \404 );
and \U$240 ( \406 , \369 , \404 );
or \U$241 ( \407 , \383 , \405 , \406 );
and \U$242 ( \408 , \387 , \400 );
and \U$243 ( \409 , \400 , \403 );
and \U$244 ( \410 , \387 , \403 );
or \U$245 ( \411 , \408 , \409 , \410 );
not \U$246 ( \412 , \318 );
and \U$247 ( \413 , \313 , \328 );
and \U$248 ( \414 , \289 , \326 );
nor \U$249 ( \415 , \413 , \414 );
xnor \U$250 ( \416 , \415 , \336 );
xor \U$251 ( \417 , \412 , \416 );
and \U$252 ( \418 , \331 , \348 );
and \U$253 ( \419 , \304 , \346 );
nor \U$254 ( \420 , \418 , \419 );
xnor \U$255 ( \421 , \420 , \356 );
xor \U$256 ( \422 , \417 , \421 );
xor \U$257 ( \423 , \411 , \422 );
and \U$258 ( \424 , \390 , \394 );
and \U$259 ( \425 , \394 , \399 );
and \U$260 ( \426 , \390 , \399 );
or \U$261 ( \427 , \424 , \425 , \426 );
buf \U$262 ( \428 , \402 );
xor \U$263 ( \429 , \427 , \428 );
and \U$264 ( \430 , \322 , \343 );
xor \U$265 ( \431 , \429 , \430 );
xor \U$266 ( \432 , \423 , \431 );
xor \U$267 ( \433 , \407 , \432 );
and \U$268 ( \434 , \351 , \328 );
and \U$269 ( \435 , \322 , \326 );
nor \U$270 ( \436 , \434 , \435 );
xnor \U$271 ( \437 , \436 , \336 );
and \U$272 ( \438 , \359 , \348 );
and \U$273 ( \439 , \342 , \346 );
nor \U$274 ( \440 , \438 , \439 );
xnor \U$275 ( \441 , \440 , \356 );
and \U$276 ( \442 , \437 , \441 );
_DC g13b ( \443_nG13b , RIb4c68d8_41 , \287 );
buf \U$277 ( \444 , \443_nG13b );
and \U$278 ( \445 , \444 , \343 );
and \U$279 ( \446 , \441 , \445 );
and \U$280 ( \447 , \437 , \445 );
or \U$281 ( \448 , \442 , \446 , \447 );
buf \U$282 ( \449 , RIa1675d0_10);
buf \U$283 ( \450 , RIa167558_11);
and \U$284 ( \451 , \449 , \450 );
not \U$285 ( \452 , \451 );
and \U$286 ( \453 , \293 , \452 );
not \U$287 ( \454 , \453 );
and \U$288 ( \455 , \313 , \296 );
and \U$289 ( \456 , \289 , \294 );
nor \U$290 ( \457 , \455 , \456 );
xnor \U$291 ( \458 , \457 , \301 );
and \U$292 ( \459 , \454 , \458 );
and \U$293 ( \460 , \331 , \310 );
and \U$294 ( \461 , \304 , \308 );
nor \U$295 ( \462 , \460 , \461 );
xnor \U$296 ( \463 , \462 , \318 );
and \U$297 ( \464 , \458 , \463 );
and \U$298 ( \465 , \454 , \463 );
or \U$299 ( \466 , \459 , \464 , \465 );
and \U$300 ( \467 , \448 , \466 );
xnor \U$301 ( \468 , \357 , \360 );
and \U$302 ( \469 , \466 , \468 );
and \U$303 ( \470 , \448 , \468 );
or \U$304 ( \471 , \467 , \469 , \470 );
xor \U$305 ( \472 , \340 , \361 );
xor \U$306 ( \473 , \472 , \366 );
and \U$307 ( \474 , \471 , \473 );
xor \U$308 ( \475 , \370 , \381 );
and \U$309 ( \476 , \473 , \475 );
and \U$310 ( \477 , \471 , \475 );
or \U$311 ( \478 , \474 , \476 , \477 );
xor \U$312 ( \479 , \369 , \382 );
xor \U$313 ( \480 , \479 , \404 );
and \U$314 ( \481 , \478 , \480 );
xor \U$315 ( \482 , \433 , \481 );
xor \U$316 ( \483 , \478 , \480 );
and \U$317 ( \484 , \342 , \328 );
and \U$318 ( \485 , \351 , \326 );
nor \U$319 ( \486 , \484 , \485 );
xnor \U$320 ( \487 , \486 , \336 );
and \U$321 ( \488 , \444 , \348 );
and \U$322 ( \489 , \359 , \346 );
nor \U$323 ( \490 , \488 , \489 );
xnor \U$324 ( \491 , \490 , \356 );
and \U$325 ( \492 , \487 , \491 );
_DC g13a ( \493_nG13a , RIb4c6860_42 , \287 );
buf \U$326 ( \494 , \493_nG13a );
and \U$327 ( \495 , \494 , \343 );
and \U$328 ( \496 , \491 , \495 );
and \U$329 ( \497 , \487 , \495 );
or \U$330 ( \498 , \492 , \496 , \497 );
xor \U$331 ( \499 , \293 , \449 );
xor \U$332 ( \500 , \449 , \450 );
not \U$333 ( \501 , \500 );
and \U$334 ( \502 , \499 , \501 );
and \U$335 ( \503 , \289 , \502 );
not \U$336 ( \504 , \503 );
xnor \U$337 ( \505 , \504 , \453 );
and \U$338 ( \506 , \304 , \296 );
and \U$339 ( \507 , \313 , \294 );
nor \U$340 ( \508 , \506 , \507 );
xnor \U$341 ( \509 , \508 , \301 );
and \U$342 ( \510 , \505 , \509 );
and \U$343 ( \511 , \322 , \310 );
and \U$344 ( \512 , \331 , \308 );
nor \U$345 ( \513 , \511 , \512 );
xnor \U$346 ( \514 , \513 , \318 );
and \U$347 ( \515 , \509 , \514 );
and \U$348 ( \516 , \505 , \514 );
or \U$349 ( \517 , \510 , \515 , \516 );
and \U$350 ( \518 , \498 , \517 );
xor \U$351 ( \519 , \437 , \441 );
xor \U$352 ( \520 , \519 , \445 );
and \U$353 ( \521 , \517 , \520 );
and \U$354 ( \522 , \498 , \520 );
or \U$355 ( \523 , \518 , \521 , \522 );
xor \U$356 ( \524 , \302 , \319 );
xor \U$357 ( \525 , \524 , \337 );
and \U$358 ( \526 , \523 , \525 );
xor \U$359 ( \527 , \448 , \466 );
xor \U$360 ( \528 , \527 , \468 );
and \U$361 ( \529 , \525 , \528 );
and \U$362 ( \530 , \523 , \528 );
or \U$363 ( \531 , \526 , \529 , \530 );
xor \U$364 ( \532 , \471 , \473 );
xor \U$365 ( \533 , \532 , \475 );
and \U$366 ( \534 , \531 , \533 );
and \U$367 ( \535 , \483 , \534 );
xor \U$368 ( \536 , \483 , \534 );
xor \U$369 ( \537 , \531 , \533 );
and \U$370 ( \538 , \351 , \310 );
and \U$371 ( \539 , \322 , \308 );
nor \U$372 ( \540 , \538 , \539 );
xnor \U$373 ( \541 , \540 , \318 );
and \U$374 ( \542 , \359 , \328 );
and \U$375 ( \543 , \342 , \326 );
nor \U$376 ( \544 , \542 , \543 );
xnor \U$377 ( \545 , \544 , \336 );
and \U$378 ( \546 , \541 , \545 );
and \U$379 ( \547 , \494 , \348 );
and \U$380 ( \548 , \444 , \346 );
nor \U$381 ( \549 , \547 , \548 );
xnor \U$382 ( \550 , \549 , \356 );
and \U$383 ( \551 , \545 , \550 );
and \U$384 ( \552 , \541 , \550 );
or \U$385 ( \553 , \546 , \551 , \552 );
buf \U$386 ( \554 , RIa1674e0_12);
buf \U$387 ( \555 , RIa167468_13);
and \U$388 ( \556 , \554 , \555 );
not \U$389 ( \557 , \556 );
and \U$390 ( \558 , \450 , \557 );
not \U$391 ( \559 , \558 );
and \U$392 ( \560 , \313 , \502 );
and \U$393 ( \561 , \289 , \500 );
nor \U$394 ( \562 , \560 , \561 );
xnor \U$395 ( \563 , \562 , \453 );
and \U$396 ( \564 , \559 , \563 );
and \U$397 ( \565 , \331 , \296 );
and \U$398 ( \566 , \304 , \294 );
nor \U$399 ( \567 , \565 , \566 );
xnor \U$400 ( \568 , \567 , \301 );
and \U$401 ( \569 , \563 , \568 );
and \U$402 ( \570 , \559 , \568 );
or \U$403 ( \571 , \564 , \569 , \570 );
or \U$404 ( \572 , \553 , \571 );
xor \U$405 ( \573 , \454 , \458 );
xor \U$406 ( \574 , \573 , \463 );
and \U$407 ( \575 , \572 , \574 );
xor \U$408 ( \576 , \498 , \517 );
xor \U$409 ( \577 , \576 , \520 );
and \U$410 ( \578 , \574 , \577 );
and \U$411 ( \579 , \572 , \577 );
or \U$412 ( \580 , \575 , \578 , \579 );
and \U$413 ( \581 , \342 , \310 );
and \U$414 ( \582 , \351 , \308 );
nor \U$415 ( \583 , \581 , \582 );
xnor \U$416 ( \584 , \583 , \318 );
and \U$417 ( \585 , \444 , \328 );
and \U$418 ( \586 , \359 , \326 );
nor \U$419 ( \587 , \585 , \586 );
xnor \U$420 ( \588 , \587 , \336 );
and \U$421 ( \589 , \584 , \588 );
_DC g139 ( \590_nG139 , RIb4c67e8_43 , \287 );
buf \U$422 ( \591 , \590_nG139 );
and \U$423 ( \592 , \591 , \348 );
and \U$424 ( \593 , \494 , \346 );
nor \U$425 ( \594 , \592 , \593 );
xnor \U$426 ( \595 , \594 , \356 );
and \U$427 ( \596 , \588 , \595 );
and \U$428 ( \597 , \584 , \595 );
or \U$429 ( \598 , \589 , \596 , \597 );
xor \U$430 ( \599 , \450 , \554 );
xor \U$431 ( \600 , \554 , \555 );
not \U$432 ( \601 , \600 );
and \U$433 ( \602 , \599 , \601 );
and \U$434 ( \603 , \289 , \602 );
not \U$435 ( \604 , \603 );
xnor \U$436 ( \605 , \604 , \558 );
and \U$437 ( \606 , \304 , \502 );
and \U$438 ( \607 , \313 , \500 );
nor \U$439 ( \608 , \606 , \607 );
xnor \U$440 ( \609 , \608 , \453 );
and \U$441 ( \610 , \605 , \609 );
and \U$442 ( \611 , \322 , \296 );
and \U$443 ( \612 , \331 , \294 );
nor \U$444 ( \613 , \611 , \612 );
xnor \U$445 ( \614 , \613 , \301 );
and \U$446 ( \615 , \609 , \614 );
and \U$447 ( \616 , \605 , \614 );
or \U$448 ( \617 , \610 , \615 , \616 );
and \U$449 ( \618 , \598 , \617 );
_DC g138 ( \619_nG138 , RIb4c6770_44 , \287 );
buf \U$450 ( \620 , \619_nG138 );
and \U$451 ( \621 , \620 , \343 );
buf \U$452 ( \622 , \621 );
and \U$453 ( \623 , \617 , \622 );
and \U$454 ( \624 , \598 , \622 );
or \U$455 ( \625 , \618 , \623 , \624 );
and \U$456 ( \626 , \591 , \343 );
xor \U$457 ( \627 , \541 , \545 );
xor \U$458 ( \628 , \627 , \550 );
and \U$459 ( \629 , \626 , \628 );
xor \U$460 ( \630 , \559 , \563 );
xor \U$461 ( \631 , \630 , \568 );
and \U$462 ( \632 , \628 , \631 );
and \U$463 ( \633 , \626 , \631 );
or \U$464 ( \634 , \629 , \632 , \633 );
and \U$465 ( \635 , \625 , \634 );
xor \U$466 ( \636 , \487 , \491 );
xor \U$467 ( \637 , \636 , \495 );
and \U$468 ( \638 , \634 , \637 );
and \U$469 ( \639 , \625 , \637 );
or \U$470 ( \640 , \635 , \638 , \639 );
xor \U$471 ( \641 , \505 , \509 );
xor \U$472 ( \642 , \641 , \514 );
xnor \U$473 ( \643 , \553 , \571 );
and \U$474 ( \644 , \642 , \643 );
and \U$475 ( \645 , \640 , \644 );
xor \U$476 ( \646 , \572 , \574 );
xor \U$477 ( \647 , \646 , \577 );
and \U$478 ( \648 , \644 , \647 );
and \U$479 ( \649 , \640 , \647 );
or \U$480 ( \650 , \645 , \648 , \649 );
and \U$481 ( \651 , \580 , \650 );
xor \U$482 ( \652 , \523 , \525 );
xor \U$483 ( \653 , \652 , \528 );
and \U$484 ( \654 , \650 , \653 );
and \U$485 ( \655 , \580 , \653 );
or \U$486 ( \656 , \651 , \654 , \655 );
and \U$487 ( \657 , \537 , \656 );
xor \U$488 ( \658 , \537 , \656 );
xor \U$489 ( \659 , \580 , \650 );
xor \U$490 ( \660 , \659 , \653 );
buf \U$491 ( \661 , RIa1673f0_14);
buf \U$492 ( \662 , RIa167378_15);
and \U$493 ( \663 , \661 , \662 );
not \U$494 ( \664 , \663 );
and \U$495 ( \665 , \555 , \664 );
not \U$496 ( \666 , \665 );
and \U$497 ( \667 , \313 , \602 );
and \U$498 ( \668 , \289 , \600 );
nor \U$499 ( \669 , \667 , \668 );
xnor \U$500 ( \670 , \669 , \558 );
and \U$501 ( \671 , \666 , \670 );
and \U$502 ( \672 , \331 , \502 );
and \U$503 ( \673 , \304 , \500 );
nor \U$504 ( \674 , \672 , \673 );
xnor \U$505 ( \675 , \674 , \453 );
and \U$506 ( \676 , \670 , \675 );
and \U$507 ( \677 , \666 , \675 );
or \U$508 ( \678 , \671 , \676 , \677 );
and \U$509 ( \679 , \351 , \296 );
and \U$510 ( \680 , \322 , \294 );
nor \U$511 ( \681 , \679 , \680 );
xnor \U$512 ( \682 , \681 , \301 );
and \U$513 ( \683 , \359 , \310 );
and \U$514 ( \684 , \342 , \308 );
nor \U$515 ( \685 , \683 , \684 );
xnor \U$516 ( \686 , \685 , \318 );
and \U$517 ( \687 , \682 , \686 );
and \U$518 ( \688 , \494 , \328 );
and \U$519 ( \689 , \444 , \326 );
nor \U$520 ( \690 , \688 , \689 );
xnor \U$521 ( \691 , \690 , \336 );
and \U$522 ( \692 , \686 , \691 );
and \U$523 ( \693 , \682 , \691 );
or \U$524 ( \694 , \687 , \692 , \693 );
and \U$525 ( \695 , \678 , \694 );
and \U$526 ( \696 , \620 , \348 );
and \U$527 ( \697 , \591 , \346 );
nor \U$528 ( \698 , \696 , \697 );
xnor \U$529 ( \699 , \698 , \356 );
_DC g137 ( \700_nG137 , RIb4c3368_45 , \287 );
buf \U$530 ( \701 , \700_nG137 );
and \U$531 ( \702 , \701 , \343 );
and \U$532 ( \703 , \699 , \702 );
and \U$533 ( \704 , \694 , \703 );
and \U$534 ( \705 , \678 , \703 );
or \U$535 ( \706 , \695 , \704 , \705 );
xor \U$536 ( \707 , \584 , \588 );
xor \U$537 ( \708 , \707 , \595 );
xor \U$538 ( \709 , \605 , \609 );
xor \U$539 ( \710 , \709 , \614 );
and \U$540 ( \711 , \708 , \710 );
not \U$541 ( \712 , \621 );
and \U$542 ( \713 , \710 , \712 );
and \U$543 ( \714 , \708 , \712 );
or \U$544 ( \715 , \711 , \713 , \714 );
and \U$545 ( \716 , \706 , \715 );
xor \U$546 ( \717 , \626 , \628 );
xor \U$547 ( \718 , \717 , \631 );
and \U$548 ( \719 , \715 , \718 );
and \U$549 ( \720 , \706 , \718 );
or \U$550 ( \721 , \716 , \719 , \720 );
xor \U$551 ( \722 , \625 , \634 );
xor \U$552 ( \723 , \722 , \637 );
and \U$553 ( \724 , \721 , \723 );
xor \U$554 ( \725 , \642 , \643 );
and \U$555 ( \726 , \723 , \725 );
and \U$556 ( \727 , \721 , \725 );
or \U$557 ( \728 , \724 , \726 , \727 );
xor \U$558 ( \729 , \640 , \644 );
xor \U$559 ( \730 , \729 , \647 );
and \U$560 ( \731 , \728 , \730 );
and \U$561 ( \732 , \660 , \731 );
xor \U$562 ( \733 , \660 , \731 );
xor \U$563 ( \734 , \728 , \730 );
xor \U$564 ( \735 , \555 , \661 );
xor \U$565 ( \736 , \661 , \662 );
not \U$566 ( \737 , \736 );
and \U$567 ( \738 , \735 , \737 );
and \U$568 ( \739 , \289 , \738 );
not \U$569 ( \740 , \739 );
xnor \U$570 ( \741 , \740 , \665 );
and \U$571 ( \742 , \304 , \602 );
and \U$572 ( \743 , \313 , \600 );
nor \U$573 ( \744 , \742 , \743 );
xnor \U$574 ( \745 , \744 , \558 );
and \U$575 ( \746 , \741 , \745 );
and \U$576 ( \747 , \322 , \502 );
and \U$577 ( \748 , \331 , \500 );
nor \U$578 ( \749 , \747 , \748 );
xnor \U$579 ( \750 , \749 , \453 );
and \U$580 ( \751 , \745 , \750 );
and \U$581 ( \752 , \741 , \750 );
or \U$582 ( \753 , \746 , \751 , \752 );
and \U$583 ( \754 , \342 , \296 );
and \U$584 ( \755 , \351 , \294 );
nor \U$585 ( \756 , \754 , \755 );
xnor \U$586 ( \757 , \756 , \301 );
and \U$587 ( \758 , \444 , \310 );
and \U$588 ( \759 , \359 , \308 );
nor \U$589 ( \760 , \758 , \759 );
xnor \U$590 ( \761 , \760 , \318 );
and \U$591 ( \762 , \757 , \761 );
and \U$592 ( \763 , \591 , \328 );
and \U$593 ( \764 , \494 , \326 );
nor \U$594 ( \765 , \763 , \764 );
xnor \U$595 ( \766 , \765 , \336 );
and \U$596 ( \767 , \761 , \766 );
and \U$597 ( \768 , \757 , \766 );
or \U$598 ( \769 , \762 , \767 , \768 );
and \U$599 ( \770 , \753 , \769 );
and \U$600 ( \771 , \701 , \348 );
and \U$601 ( \772 , \620 , \346 );
nor \U$602 ( \773 , \771 , \772 );
xnor \U$603 ( \774 , \773 , \356 );
_DC g136 ( \775_nG136 , RIb4c32f0_46 , \287 );
buf \U$604 ( \776 , \775_nG136 );
and \U$605 ( \777 , \776 , \343 );
or \U$606 ( \778 , \774 , \777 );
and \U$607 ( \779 , \769 , \778 );
and \U$608 ( \780 , \753 , \778 );
or \U$609 ( \781 , \770 , \779 , \780 );
xor \U$610 ( \782 , \666 , \670 );
xor \U$611 ( \783 , \782 , \675 );
xor \U$612 ( \784 , \682 , \686 );
xor \U$613 ( \785 , \784 , \691 );
and \U$614 ( \786 , \783 , \785 );
xor \U$615 ( \787 , \699 , \702 );
and \U$616 ( \788 , \785 , \787 );
and \U$617 ( \789 , \783 , \787 );
or \U$618 ( \790 , \786 , \788 , \789 );
and \U$619 ( \791 , \781 , \790 );
xor \U$620 ( \792 , \708 , \710 );
xor \U$621 ( \793 , \792 , \712 );
and \U$622 ( \794 , \790 , \793 );
and \U$623 ( \795 , \781 , \793 );
or \U$624 ( \796 , \791 , \794 , \795 );
xor \U$625 ( \797 , \598 , \617 );
xor \U$626 ( \798 , \797 , \622 );
and \U$627 ( \799 , \796 , \798 );
xor \U$628 ( \800 , \706 , \715 );
xor \U$629 ( \801 , \800 , \718 );
and \U$630 ( \802 , \798 , \801 );
and \U$631 ( \803 , \796 , \801 );
or \U$632 ( \804 , \799 , \802 , \803 );
xor \U$633 ( \805 , \721 , \723 );
xor \U$634 ( \806 , \805 , \725 );
and \U$635 ( \807 , \804 , \806 );
and \U$636 ( \808 , \734 , \807 );
xor \U$637 ( \809 , \734 , \807 );
xor \U$638 ( \810 , \804 , \806 );
buf \U$639 ( \811 , RIa167300_16);
buf \U$640 ( \812 , RIa167288_17);
and \U$641 ( \813 , \811 , \812 );
not \U$642 ( \814 , \813 );
and \U$643 ( \815 , \662 , \814 );
not \U$644 ( \816 , \815 );
and \U$645 ( \817 , \313 , \738 );
and \U$646 ( \818 , \289 , \736 );
nor \U$647 ( \819 , \817 , \818 );
xnor \U$648 ( \820 , \819 , \665 );
and \U$649 ( \821 , \816 , \820 );
and \U$650 ( \822 , \331 , \602 );
and \U$651 ( \823 , \304 , \600 );
nor \U$652 ( \824 , \822 , \823 );
xnor \U$653 ( \825 , \824 , \558 );
and \U$654 ( \826 , \820 , \825 );
and \U$655 ( \827 , \816 , \825 );
or \U$656 ( \828 , \821 , \826 , \827 );
and \U$657 ( \829 , \620 , \328 );
and \U$658 ( \830 , \591 , \326 );
nor \U$659 ( \831 , \829 , \830 );
xnor \U$660 ( \832 , \831 , \336 );
and \U$661 ( \833 , \776 , \348 );
and \U$662 ( \834 , \701 , \346 );
nor \U$663 ( \835 , \833 , \834 );
xnor \U$664 ( \836 , \835 , \356 );
and \U$665 ( \837 , \832 , \836 );
_DC g135 ( \838_nG135 , RIb4c3278_47 , \287 );
buf \U$666 ( \839 , \838_nG135 );
and \U$667 ( \840 , \839 , \343 );
and \U$668 ( \841 , \836 , \840 );
and \U$669 ( \842 , \832 , \840 );
or \U$670 ( \843 , \837 , \841 , \842 );
and \U$671 ( \844 , \828 , \843 );
and \U$672 ( \845 , \351 , \502 );
and \U$673 ( \846 , \322 , \500 );
nor \U$674 ( \847 , \845 , \846 );
xnor \U$675 ( \848 , \847 , \453 );
and \U$676 ( \849 , \359 , \296 );
and \U$677 ( \850 , \342 , \294 );
nor \U$678 ( \851 , \849 , \850 );
xnor \U$679 ( \852 , \851 , \301 );
and \U$680 ( \853 , \848 , \852 );
and \U$681 ( \854 , \494 , \310 );
and \U$682 ( \855 , \444 , \308 );
nor \U$683 ( \856 , \854 , \855 );
xnor \U$684 ( \857 , \856 , \318 );
and \U$685 ( \858 , \852 , \857 );
and \U$686 ( \859 , \848 , \857 );
or \U$687 ( \860 , \853 , \858 , \859 );
and \U$688 ( \861 , \843 , \860 );
and \U$689 ( \862 , \828 , \860 );
or \U$690 ( \863 , \844 , \861 , \862 );
xor \U$691 ( \864 , \741 , \745 );
xor \U$692 ( \865 , \864 , \750 );
xor \U$693 ( \866 , \757 , \761 );
xor \U$694 ( \867 , \866 , \766 );
and \U$695 ( \868 , \865 , \867 );
xnor \U$696 ( \869 , \774 , \777 );
and \U$697 ( \870 , \867 , \869 );
and \U$698 ( \871 , \865 , \869 );
or \U$699 ( \872 , \868 , \870 , \871 );
and \U$700 ( \873 , \863 , \872 );
xor \U$701 ( \874 , \783 , \785 );
xor \U$702 ( \875 , \874 , \787 );
and \U$703 ( \876 , \872 , \875 );
and \U$704 ( \877 , \863 , \875 );
or \U$705 ( \878 , \873 , \876 , \877 );
xor \U$706 ( \879 , \678 , \694 );
xor \U$707 ( \880 , \879 , \703 );
and \U$708 ( \881 , \878 , \880 );
xor \U$709 ( \882 , \781 , \790 );
xor \U$710 ( \883 , \882 , \793 );
and \U$711 ( \884 , \880 , \883 );
and \U$712 ( \885 , \878 , \883 );
or \U$713 ( \886 , \881 , \884 , \885 );
xor \U$714 ( \887 , \796 , \798 );
xor \U$715 ( \888 , \887 , \801 );
and \U$716 ( \889 , \886 , \888 );
and \U$717 ( \890 , \810 , \889 );
xor \U$718 ( \891 , \810 , \889 );
xor \U$719 ( \892 , \886 , \888 );
and \U$720 ( \893 , \701 , \328 );
and \U$721 ( \894 , \620 , \326 );
nor \U$722 ( \895 , \893 , \894 );
xnor \U$723 ( \896 , \895 , \336 );
and \U$724 ( \897 , \839 , \348 );
and \U$725 ( \898 , \776 , \346 );
nor \U$726 ( \899 , \897 , \898 );
xnor \U$727 ( \900 , \899 , \356 );
and \U$728 ( \901 , \896 , \900 );
_DC g134 ( \902_nG134 , RIb4c3200_48 , \287 );
buf \U$729 ( \903 , \902_nG134 );
and \U$730 ( \904 , \903 , \343 );
and \U$731 ( \905 , \900 , \904 );
and \U$732 ( \906 , \896 , \904 );
or \U$733 ( \907 , \901 , \905 , \906 );
xor \U$734 ( \908 , \662 , \811 );
xor \U$735 ( \909 , \811 , \812 );
not \U$736 ( \910 , \909 );
and \U$737 ( \911 , \908 , \910 );
and \U$738 ( \912 , \289 , \911 );
not \U$739 ( \913 , \912 );
xnor \U$740 ( \914 , \913 , \815 );
and \U$741 ( \915 , \304 , \738 );
and \U$742 ( \916 , \313 , \736 );
nor \U$743 ( \917 , \915 , \916 );
xnor \U$744 ( \918 , \917 , \665 );
and \U$745 ( \919 , \914 , \918 );
and \U$746 ( \920 , \322 , \602 );
and \U$747 ( \921 , \331 , \600 );
nor \U$748 ( \922 , \920 , \921 );
xnor \U$749 ( \923 , \922 , \558 );
and \U$750 ( \924 , \918 , \923 );
and \U$751 ( \925 , \914 , \923 );
or \U$752 ( \926 , \919 , \924 , \925 );
and \U$753 ( \927 , \907 , \926 );
and \U$754 ( \928 , \342 , \502 );
and \U$755 ( \929 , \351 , \500 );
nor \U$756 ( \930 , \928 , \929 );
xnor \U$757 ( \931 , \930 , \453 );
and \U$758 ( \932 , \444 , \296 );
and \U$759 ( \933 , \359 , \294 );
nor \U$760 ( \934 , \932 , \933 );
xnor \U$761 ( \935 , \934 , \301 );
and \U$762 ( \936 , \931 , \935 );
and \U$763 ( \937 , \591 , \310 );
and \U$764 ( \938 , \494 , \308 );
nor \U$765 ( \939 , \937 , \938 );
xnor \U$766 ( \940 , \939 , \318 );
and \U$767 ( \941 , \935 , \940 );
and \U$768 ( \942 , \931 , \940 );
or \U$769 ( \943 , \936 , \941 , \942 );
and \U$770 ( \944 , \926 , \943 );
and \U$771 ( \945 , \907 , \943 );
or \U$772 ( \946 , \927 , \944 , \945 );
xor \U$773 ( \947 , \816 , \820 );
xor \U$774 ( \948 , \947 , \825 );
xor \U$775 ( \949 , \832 , \836 );
xor \U$776 ( \950 , \949 , \840 );
and \U$777 ( \951 , \948 , \950 );
xor \U$778 ( \952 , \848 , \852 );
xor \U$779 ( \953 , \952 , \857 );
and \U$780 ( \954 , \950 , \953 );
and \U$781 ( \955 , \948 , \953 );
or \U$782 ( \956 , \951 , \954 , \955 );
and \U$783 ( \957 , \946 , \956 );
xor \U$784 ( \958 , \865 , \867 );
xor \U$785 ( \959 , \958 , \869 );
and \U$786 ( \960 , \956 , \959 );
and \U$787 ( \961 , \946 , \959 );
or \U$788 ( \962 , \957 , \960 , \961 );
xor \U$789 ( \963 , \753 , \769 );
xor \U$790 ( \964 , \963 , \778 );
and \U$791 ( \965 , \962 , \964 );
xor \U$792 ( \966 , \863 , \872 );
xor \U$793 ( \967 , \966 , \875 );
and \U$794 ( \968 , \964 , \967 );
and \U$795 ( \969 , \962 , \967 );
or \U$796 ( \970 , \965 , \968 , \969 );
xor \U$797 ( \971 , \878 , \880 );
xor \U$798 ( \972 , \971 , \883 );
and \U$799 ( \973 , \970 , \972 );
and \U$800 ( \974 , \892 , \973 );
xor \U$801 ( \975 , \892 , \973 );
xor \U$802 ( \976 , \970 , \972 );
buf \U$803 ( \977 , RIa167210_18);
buf \U$804 ( \978 , RIa167198_19);
and \U$805 ( \979 , \977 , \978 );
not \U$806 ( \980 , \979 );
and \U$807 ( \981 , \812 , \980 );
not \U$808 ( \982 , \981 );
and \U$809 ( \983 , \313 , \911 );
and \U$810 ( \984 , \289 , \909 );
nor \U$811 ( \985 , \983 , \984 );
xnor \U$812 ( \986 , \985 , \815 );
and \U$813 ( \987 , \982 , \986 );
and \U$814 ( \988 , \331 , \738 );
and \U$815 ( \989 , \304 , \736 );
nor \U$816 ( \990 , \988 , \989 );
xnor \U$817 ( \991 , \990 , \665 );
and \U$818 ( \992 , \986 , \991 );
and \U$819 ( \993 , \982 , \991 );
or \U$820 ( \994 , \987 , \992 , \993 );
and \U$821 ( \995 , \351 , \602 );
and \U$822 ( \996 , \322 , \600 );
nor \U$823 ( \997 , \995 , \996 );
xnor \U$824 ( \998 , \997 , \558 );
and \U$825 ( \999 , \359 , \502 );
and \U$826 ( \1000 , \342 , \500 );
nor \U$827 ( \1001 , \999 , \1000 );
xnor \U$828 ( \1002 , \1001 , \453 );
and \U$829 ( \1003 , \998 , \1002 );
and \U$830 ( \1004 , \494 , \296 );
and \U$831 ( \1005 , \444 , \294 );
nor \U$832 ( \1006 , \1004 , \1005 );
xnor \U$833 ( \1007 , \1006 , \301 );
and \U$834 ( \1008 , \1002 , \1007 );
and \U$835 ( \1009 , \998 , \1007 );
or \U$836 ( \1010 , \1003 , \1008 , \1009 );
and \U$837 ( \1011 , \994 , \1010 );
and \U$838 ( \1012 , \620 , \310 );
and \U$839 ( \1013 , \591 , \308 );
nor \U$840 ( \1014 , \1012 , \1013 );
xnor \U$841 ( \1015 , \1014 , \318 );
and \U$842 ( \1016 , \776 , \328 );
and \U$843 ( \1017 , \701 , \326 );
nor \U$844 ( \1018 , \1016 , \1017 );
xnor \U$845 ( \1019 , \1018 , \336 );
and \U$846 ( \1020 , \1015 , \1019 );
and \U$847 ( \1021 , \903 , \348 );
and \U$848 ( \1022 , \839 , \346 );
nor \U$849 ( \1023 , \1021 , \1022 );
xnor \U$850 ( \1024 , \1023 , \356 );
and \U$851 ( \1025 , \1019 , \1024 );
and \U$852 ( \1026 , \1015 , \1024 );
or \U$853 ( \1027 , \1020 , \1025 , \1026 );
and \U$854 ( \1028 , \1010 , \1027 );
and \U$855 ( \1029 , \994 , \1027 );
or \U$856 ( \1030 , \1011 , \1028 , \1029 );
xor \U$857 ( \1031 , \896 , \900 );
xor \U$858 ( \1032 , \1031 , \904 );
xor \U$859 ( \1033 , \931 , \935 );
xor \U$860 ( \1034 , \1033 , \940 );
or \U$861 ( \1035 , \1032 , \1034 );
and \U$862 ( \1036 , \1030 , \1035 );
xor \U$863 ( \1037 , \948 , \950 );
xor \U$864 ( \1038 , \1037 , \953 );
and \U$865 ( \1039 , \1035 , \1038 );
and \U$866 ( \1040 , \1030 , \1038 );
or \U$867 ( \1041 , \1036 , \1039 , \1040 );
xor \U$868 ( \1042 , \828 , \843 );
xor \U$869 ( \1043 , \1042 , \860 );
and \U$870 ( \1044 , \1041 , \1043 );
xor \U$871 ( \1045 , \946 , \956 );
xor \U$872 ( \1046 , \1045 , \959 );
and \U$873 ( \1047 , \1043 , \1046 );
and \U$874 ( \1048 , \1041 , \1046 );
or \U$875 ( \1049 , \1044 , \1047 , \1048 );
xor \U$876 ( \1050 , \962 , \964 );
xor \U$877 ( \1051 , \1050 , \967 );
and \U$878 ( \1052 , \1049 , \1051 );
and \U$879 ( \1053 , \976 , \1052 );
xor \U$880 ( \1054 , \976 , \1052 );
xor \U$881 ( \1055 , \1049 , \1051 );
xor \U$882 ( \1056 , \812 , \977 );
xor \U$883 ( \1057 , \977 , \978 );
not \U$884 ( \1058 , \1057 );
and \U$885 ( \1059 , \1056 , \1058 );
and \U$886 ( \1060 , \289 , \1059 );
not \U$887 ( \1061 , \1060 );
xnor \U$888 ( \1062 , \1061 , \981 );
and \U$889 ( \1063 , \304 , \911 );
and \U$890 ( \1064 , \313 , \909 );
nor \U$891 ( \1065 , \1063 , \1064 );
xnor \U$892 ( \1066 , \1065 , \815 );
and \U$893 ( \1067 , \1062 , \1066 );
and \U$894 ( \1068 , \322 , \738 );
and \U$895 ( \1069 , \331 , \736 );
nor \U$896 ( \1070 , \1068 , \1069 );
xnor \U$897 ( \1071 , \1070 , \665 );
and \U$898 ( \1072 , \1066 , \1071 );
and \U$899 ( \1073 , \1062 , \1071 );
or \U$900 ( \1074 , \1067 , \1072 , \1073 );
and \U$901 ( \1075 , \342 , \602 );
and \U$902 ( \1076 , \351 , \600 );
nor \U$903 ( \1077 , \1075 , \1076 );
xnor \U$904 ( \1078 , \1077 , \558 );
and \U$905 ( \1079 , \444 , \502 );
and \U$906 ( \1080 , \359 , \500 );
nor \U$907 ( \1081 , \1079 , \1080 );
xnor \U$908 ( \1082 , \1081 , \453 );
and \U$909 ( \1083 , \1078 , \1082 );
and \U$910 ( \1084 , \591 , \296 );
and \U$911 ( \1085 , \494 , \294 );
nor \U$912 ( \1086 , \1084 , \1085 );
xnor \U$913 ( \1087 , \1086 , \301 );
and \U$914 ( \1088 , \1082 , \1087 );
and \U$915 ( \1089 , \1078 , \1087 );
or \U$916 ( \1090 , \1083 , \1088 , \1089 );
and \U$917 ( \1091 , \1074 , \1090 );
and \U$918 ( \1092 , \701 , \310 );
and \U$919 ( \1093 , \620 , \308 );
nor \U$920 ( \1094 , \1092 , \1093 );
xnor \U$921 ( \1095 , \1094 , \318 );
and \U$922 ( \1096 , \839 , \328 );
and \U$923 ( \1097 , \776 , \326 );
nor \U$924 ( \1098 , \1096 , \1097 );
xnor \U$925 ( \1099 , \1098 , \336 );
and \U$926 ( \1100 , \1095 , \1099 );
_DC g133 ( \1101_nG133 , RIb4c3188_49 , \287 );
buf \U$927 ( \1102 , \1101_nG133 );
and \U$928 ( \1103 , \1102 , \348 );
and \U$929 ( \1104 , \903 , \346 );
nor \U$930 ( \1105 , \1103 , \1104 );
xnor \U$931 ( \1106 , \1105 , \356 );
and \U$932 ( \1107 , \1099 , \1106 );
and \U$933 ( \1108 , \1095 , \1106 );
or \U$934 ( \1109 , \1100 , \1107 , \1108 );
and \U$935 ( \1110 , \1090 , \1109 );
and \U$936 ( \1111 , \1074 , \1109 );
or \U$937 ( \1112 , \1091 , \1110 , \1111 );
and \U$938 ( \1113 , \1102 , \343 );
xor \U$939 ( \1114 , \998 , \1002 );
xor \U$940 ( \1115 , \1114 , \1007 );
and \U$941 ( \1116 , \1113 , \1115 );
xor \U$942 ( \1117 , \1015 , \1019 );
xor \U$943 ( \1118 , \1117 , \1024 );
and \U$944 ( \1119 , \1115 , \1118 );
and \U$945 ( \1120 , \1113 , \1118 );
or \U$946 ( \1121 , \1116 , \1119 , \1120 );
and \U$947 ( \1122 , \1112 , \1121 );
xor \U$948 ( \1123 , \914 , \918 );
xor \U$949 ( \1124 , \1123 , \923 );
and \U$950 ( \1125 , \1121 , \1124 );
and \U$951 ( \1126 , \1112 , \1124 );
or \U$952 ( \1127 , \1122 , \1125 , \1126 );
xor \U$953 ( \1128 , \907 , \926 );
xor \U$954 ( \1129 , \1128 , \943 );
and \U$955 ( \1130 , \1127 , \1129 );
xor \U$956 ( \1131 , \1030 , \1035 );
xor \U$957 ( \1132 , \1131 , \1038 );
and \U$958 ( \1133 , \1129 , \1132 );
and \U$959 ( \1134 , \1127 , \1132 );
or \U$960 ( \1135 , \1130 , \1133 , \1134 );
and \U$961 ( \1136 , \351 , \738 );
and \U$962 ( \1137 , \322 , \736 );
nor \U$963 ( \1138 , \1136 , \1137 );
xnor \U$964 ( \1139 , \1138 , \665 );
and \U$965 ( \1140 , \359 , \602 );
and \U$966 ( \1141 , \342 , \600 );
nor \U$967 ( \1142 , \1140 , \1141 );
xnor \U$968 ( \1143 , \1142 , \558 );
and \U$969 ( \1144 , \1139 , \1143 );
and \U$970 ( \1145 , \494 , \502 );
and \U$971 ( \1146 , \444 , \500 );
nor \U$972 ( \1147 , \1145 , \1146 );
xnor \U$973 ( \1148 , \1147 , \453 );
and \U$974 ( \1149 , \1143 , \1148 );
and \U$975 ( \1150 , \1139 , \1148 );
or \U$976 ( \1151 , \1144 , \1149 , \1150 );
and \U$977 ( \1152 , \620 , \296 );
and \U$978 ( \1153 , \591 , \294 );
nor \U$979 ( \1154 , \1152 , \1153 );
xnor \U$980 ( \1155 , \1154 , \301 );
and \U$981 ( \1156 , \776 , \310 );
and \U$982 ( \1157 , \701 , \308 );
nor \U$983 ( \1158 , \1156 , \1157 );
xnor \U$984 ( \1159 , \1158 , \318 );
and \U$985 ( \1160 , \1155 , \1159 );
and \U$986 ( \1161 , \903 , \328 );
and \U$987 ( \1162 , \839 , \326 );
nor \U$988 ( \1163 , \1161 , \1162 );
xnor \U$989 ( \1164 , \1163 , \336 );
and \U$990 ( \1165 , \1159 , \1164 );
and \U$991 ( \1166 , \1155 , \1164 );
or \U$992 ( \1167 , \1160 , \1165 , \1166 );
and \U$993 ( \1168 , \1151 , \1167 );
buf \U$994 ( \1169 , RIa167120_20);
buf \U$995 ( \1170 , RIa1670a8_21);
and \U$996 ( \1171 , \1169 , \1170 );
not \U$997 ( \1172 , \1171 );
and \U$998 ( \1173 , \978 , \1172 );
not \U$999 ( \1174 , \1173 );
and \U$1000 ( \1175 , \313 , \1059 );
and \U$1001 ( \1176 , \289 , \1057 );
nor \U$1002 ( \1177 , \1175 , \1176 );
xnor \U$1003 ( \1178 , \1177 , \981 );
and \U$1004 ( \1179 , \1174 , \1178 );
and \U$1005 ( \1180 , \331 , \911 );
and \U$1006 ( \1181 , \304 , \909 );
nor \U$1007 ( \1182 , \1180 , \1181 );
xnor \U$1008 ( \1183 , \1182 , \815 );
and \U$1009 ( \1184 , \1178 , \1183 );
and \U$1010 ( \1185 , \1174 , \1183 );
or \U$1011 ( \1186 , \1179 , \1184 , \1185 );
and \U$1012 ( \1187 , \1167 , \1186 );
and \U$1013 ( \1188 , \1151 , \1186 );
or \U$1014 ( \1189 , \1168 , \1187 , \1188 );
_DC g132 ( \1190_nG132 , RIb4c3110_50 , \287 );
buf \U$1015 ( \1191 , \1190_nG132 );
and \U$1016 ( \1192 , \1191 , \343 );
xor \U$1017 ( \1193 , \1095 , \1099 );
xor \U$1018 ( \1194 , \1193 , \1106 );
or \U$1019 ( \1195 , \1192 , \1194 );
and \U$1020 ( \1196 , \1189 , \1195 );
xor \U$1021 ( \1197 , \1062 , \1066 );
xor \U$1022 ( \1198 , \1197 , \1071 );
xor \U$1023 ( \1199 , \1078 , \1082 );
xor \U$1024 ( \1200 , \1199 , \1087 );
and \U$1025 ( \1201 , \1198 , \1200 );
and \U$1026 ( \1202 , \1195 , \1201 );
and \U$1027 ( \1203 , \1189 , \1201 );
or \U$1028 ( \1204 , \1196 , \1202 , \1203 );
xor \U$1029 ( \1205 , \982 , \986 );
xor \U$1030 ( \1206 , \1205 , \991 );
xor \U$1031 ( \1207 , \1074 , \1090 );
xor \U$1032 ( \1208 , \1207 , \1109 );
and \U$1033 ( \1209 , \1206 , \1208 );
xor \U$1034 ( \1210 , \1113 , \1115 );
xor \U$1035 ( \1211 , \1210 , \1118 );
and \U$1036 ( \1212 , \1208 , \1211 );
and \U$1037 ( \1213 , \1206 , \1211 );
or \U$1038 ( \1214 , \1209 , \1212 , \1213 );
and \U$1039 ( \1215 , \1204 , \1214 );
xnor \U$1040 ( \1216 , \1032 , \1034 );
and \U$1041 ( \1217 , \1214 , \1216 );
and \U$1042 ( \1218 , \1204 , \1216 );
or \U$1043 ( \1219 , \1215 , \1217 , \1218 );
xor \U$1044 ( \1220 , \994 , \1010 );
xor \U$1045 ( \1221 , \1220 , \1027 );
xor \U$1046 ( \1222 , \1112 , \1121 );
xor \U$1047 ( \1223 , \1222 , \1124 );
and \U$1048 ( \1224 , \1221 , \1223 );
and \U$1049 ( \1225 , \1219 , \1224 );
xor \U$1050 ( \1226 , \1127 , \1129 );
xor \U$1051 ( \1227 , \1226 , \1132 );
and \U$1052 ( \1228 , \1224 , \1227 );
and \U$1053 ( \1229 , \1219 , \1227 );
or \U$1054 ( \1230 , \1225 , \1228 , \1229 );
and \U$1055 ( \1231 , \1135 , \1230 );
xor \U$1056 ( \1232 , \1041 , \1043 );
xor \U$1057 ( \1233 , \1232 , \1046 );
and \U$1058 ( \1234 , \1230 , \1233 );
and \U$1059 ( \1235 , \1135 , \1233 );
or \U$1060 ( \1236 , \1231 , \1234 , \1235 );
and \U$1061 ( \1237 , \1055 , \1236 );
xor \U$1062 ( \1238 , \1055 , \1236 );
xor \U$1063 ( \1239 , \1135 , \1230 );
xor \U$1064 ( \1240 , \1239 , \1233 );
and \U$1065 ( \1241 , \342 , \738 );
and \U$1066 ( \1242 , \351 , \736 );
nor \U$1067 ( \1243 , \1241 , \1242 );
xnor \U$1068 ( \1244 , \1243 , \665 );
and \U$1069 ( \1245 , \444 , \602 );
and \U$1070 ( \1246 , \359 , \600 );
nor \U$1071 ( \1247 , \1245 , \1246 );
xnor \U$1072 ( \1248 , \1247 , \558 );
and \U$1073 ( \1249 , \1244 , \1248 );
and \U$1074 ( \1250 , \591 , \502 );
and \U$1075 ( \1251 , \494 , \500 );
nor \U$1076 ( \1252 , \1250 , \1251 );
xnor \U$1077 ( \1253 , \1252 , \453 );
and \U$1078 ( \1254 , \1248 , \1253 );
and \U$1079 ( \1255 , \1244 , \1253 );
or \U$1080 ( \1256 , \1249 , \1254 , \1255 );
and \U$1081 ( \1257 , \701 , \296 );
and \U$1082 ( \1258 , \620 , \294 );
nor \U$1083 ( \1259 , \1257 , \1258 );
xnor \U$1084 ( \1260 , \1259 , \301 );
and \U$1085 ( \1261 , \839 , \310 );
and \U$1086 ( \1262 , \776 , \308 );
nor \U$1087 ( \1263 , \1261 , \1262 );
xnor \U$1088 ( \1264 , \1263 , \318 );
and \U$1089 ( \1265 , \1260 , \1264 );
and \U$1090 ( \1266 , \1102 , \328 );
and \U$1091 ( \1267 , \903 , \326 );
nor \U$1092 ( \1268 , \1266 , \1267 );
xnor \U$1093 ( \1269 , \1268 , \336 );
and \U$1094 ( \1270 , \1264 , \1269 );
and \U$1095 ( \1271 , \1260 , \1269 );
or \U$1096 ( \1272 , \1265 , \1270 , \1271 );
and \U$1097 ( \1273 , \1256 , \1272 );
xor \U$1098 ( \1274 , \978 , \1169 );
xor \U$1099 ( \1275 , \1169 , \1170 );
not \U$1100 ( \1276 , \1275 );
and \U$1101 ( \1277 , \1274 , \1276 );
and \U$1102 ( \1278 , \289 , \1277 );
not \U$1103 ( \1279 , \1278 );
xnor \U$1104 ( \1280 , \1279 , \1173 );
and \U$1105 ( \1281 , \304 , \1059 );
and \U$1106 ( \1282 , \313 , \1057 );
nor \U$1107 ( \1283 , \1281 , \1282 );
xnor \U$1108 ( \1284 , \1283 , \981 );
and \U$1109 ( \1285 , \1280 , \1284 );
and \U$1110 ( \1286 , \322 , \911 );
and \U$1111 ( \1287 , \331 , \909 );
nor \U$1112 ( \1288 , \1286 , \1287 );
xnor \U$1113 ( \1289 , \1288 , \815 );
and \U$1114 ( \1290 , \1284 , \1289 );
and \U$1115 ( \1291 , \1280 , \1289 );
or \U$1116 ( \1292 , \1285 , \1290 , \1291 );
and \U$1117 ( \1293 , \1272 , \1292 );
and \U$1118 ( \1294 , \1256 , \1292 );
or \U$1119 ( \1295 , \1273 , \1293 , \1294 );
_DC g131 ( \1296_nG131 , RIb4c3098_51 , \287 );
buf \U$1120 ( \1297 , \1296_nG131 );
and \U$1121 ( \1298 , \1297 , \348 );
and \U$1122 ( \1299 , \1191 , \346 );
nor \U$1123 ( \1300 , \1298 , \1299 );
xnor \U$1124 ( \1301 , \1300 , \356 );
_DC g130 ( \1302_nG130 , RIb4c3020_52 , \287 );
buf \U$1125 ( \1303 , \1302_nG130 );
and \U$1126 ( \1304 , \1303 , \343 );
or \U$1127 ( \1305 , \1301 , \1304 );
and \U$1128 ( \1306 , \1191 , \348 );
and \U$1129 ( \1307 , \1102 , \346 );
nor \U$1130 ( \1308 , \1306 , \1307 );
xnor \U$1131 ( \1309 , \1308 , \356 );
and \U$1132 ( \1310 , \1305 , \1309 );
and \U$1133 ( \1311 , \1297 , \343 );
and \U$1134 ( \1312 , \1309 , \1311 );
and \U$1135 ( \1313 , \1305 , \1311 );
or \U$1136 ( \1314 , \1310 , \1312 , \1313 );
and \U$1137 ( \1315 , \1295 , \1314 );
xor \U$1138 ( \1316 , \1139 , \1143 );
xor \U$1139 ( \1317 , \1316 , \1148 );
xor \U$1140 ( \1318 , \1155 , \1159 );
xor \U$1141 ( \1319 , \1318 , \1164 );
and \U$1142 ( \1320 , \1317 , \1319 );
xor \U$1143 ( \1321 , \1174 , \1178 );
xor \U$1144 ( \1322 , \1321 , \1183 );
and \U$1145 ( \1323 , \1319 , \1322 );
and \U$1146 ( \1324 , \1317 , \1322 );
or \U$1147 ( \1325 , \1320 , \1323 , \1324 );
and \U$1148 ( \1326 , \1314 , \1325 );
and \U$1149 ( \1327 , \1295 , \1325 );
or \U$1150 ( \1328 , \1315 , \1326 , \1327 );
xor \U$1151 ( \1329 , \1151 , \1167 );
xor \U$1152 ( \1330 , \1329 , \1186 );
xnor \U$1153 ( \1331 , \1192 , \1194 );
and \U$1154 ( \1332 , \1330 , \1331 );
xor \U$1155 ( \1333 , \1198 , \1200 );
and \U$1156 ( \1334 , \1331 , \1333 );
and \U$1157 ( \1335 , \1330 , \1333 );
or \U$1158 ( \1336 , \1332 , \1334 , \1335 );
and \U$1159 ( \1337 , \1328 , \1336 );
xor \U$1160 ( \1338 , \1206 , \1208 );
xor \U$1161 ( \1339 , \1338 , \1211 );
and \U$1162 ( \1340 , \1336 , \1339 );
and \U$1163 ( \1341 , \1328 , \1339 );
or \U$1164 ( \1342 , \1337 , \1340 , \1341 );
xor \U$1165 ( \1343 , \1204 , \1214 );
xor \U$1166 ( \1344 , \1343 , \1216 );
and \U$1167 ( \1345 , \1342 , \1344 );
xor \U$1168 ( \1346 , \1221 , \1223 );
and \U$1169 ( \1347 , \1344 , \1346 );
and \U$1170 ( \1348 , \1342 , \1346 );
or \U$1171 ( \1349 , \1345 , \1347 , \1348 );
xor \U$1172 ( \1350 , \1219 , \1224 );
xor \U$1173 ( \1351 , \1350 , \1227 );
and \U$1174 ( \1352 , \1349 , \1351 );
and \U$1175 ( \1353 , \1240 , \1352 );
xor \U$1176 ( \1354 , \1240 , \1352 );
xor \U$1177 ( \1355 , \1349 , \1351 );
buf \U$1178 ( \1356 , RIa167030_22);
buf \U$1179 ( \1357 , RIa166fb8_23);
and \U$1180 ( \1358 , \1356 , \1357 );
not \U$1181 ( \1359 , \1358 );
and \U$1182 ( \1360 , \1170 , \1359 );
not \U$1183 ( \1361 , \1360 );
and \U$1184 ( \1362 , \313 , \1277 );
and \U$1185 ( \1363 , \289 , \1275 );
nor \U$1186 ( \1364 , \1362 , \1363 );
xnor \U$1187 ( \1365 , \1364 , \1173 );
and \U$1188 ( \1366 , \1361 , \1365 );
and \U$1189 ( \1367 , \331 , \1059 );
and \U$1190 ( \1368 , \304 , \1057 );
nor \U$1191 ( \1369 , \1367 , \1368 );
xnor \U$1192 ( \1370 , \1369 , \981 );
and \U$1193 ( \1371 , \1365 , \1370 );
and \U$1194 ( \1372 , \1361 , \1370 );
or \U$1195 ( \1373 , \1366 , \1371 , \1372 );
and \U$1196 ( \1374 , \351 , \911 );
and \U$1197 ( \1375 , \322 , \909 );
nor \U$1198 ( \1376 , \1374 , \1375 );
xnor \U$1199 ( \1377 , \1376 , \815 );
and \U$1200 ( \1378 , \359 , \738 );
and \U$1201 ( \1379 , \342 , \736 );
nor \U$1202 ( \1380 , \1378 , \1379 );
xnor \U$1203 ( \1381 , \1380 , \665 );
and \U$1204 ( \1382 , \1377 , \1381 );
and \U$1205 ( \1383 , \494 , \602 );
and \U$1206 ( \1384 , \444 , \600 );
nor \U$1207 ( \1385 , \1383 , \1384 );
xnor \U$1208 ( \1386 , \1385 , \558 );
and \U$1209 ( \1387 , \1381 , \1386 );
and \U$1210 ( \1388 , \1377 , \1386 );
or \U$1211 ( \1389 , \1382 , \1387 , \1388 );
and \U$1212 ( \1390 , \1373 , \1389 );
and \U$1213 ( \1391 , \620 , \502 );
and \U$1214 ( \1392 , \591 , \500 );
nor \U$1215 ( \1393 , \1391 , \1392 );
xnor \U$1216 ( \1394 , \1393 , \453 );
and \U$1217 ( \1395 , \776 , \296 );
and \U$1218 ( \1396 , \701 , \294 );
nor \U$1219 ( \1397 , \1395 , \1396 );
xnor \U$1220 ( \1398 , \1397 , \301 );
and \U$1221 ( \1399 , \1394 , \1398 );
and \U$1222 ( \1400 , \903 , \310 );
and \U$1223 ( \1401 , \839 , \308 );
nor \U$1224 ( \1402 , \1400 , \1401 );
xnor \U$1225 ( \1403 , \1402 , \318 );
and \U$1226 ( \1404 , \1398 , \1403 );
and \U$1227 ( \1405 , \1394 , \1403 );
or \U$1228 ( \1406 , \1399 , \1404 , \1405 );
and \U$1229 ( \1407 , \1389 , \1406 );
and \U$1230 ( \1408 , \1373 , \1406 );
or \U$1231 ( \1409 , \1390 , \1407 , \1408 );
and \U$1232 ( \1410 , \1191 , \328 );
and \U$1233 ( \1411 , \1102 , \326 );
nor \U$1234 ( \1412 , \1410 , \1411 );
xnor \U$1235 ( \1413 , \1412 , \336 );
and \U$1236 ( \1414 , \1303 , \348 );
and \U$1237 ( \1415 , \1297 , \346 );
nor \U$1238 ( \1416 , \1414 , \1415 );
xnor \U$1239 ( \1417 , \1416 , \356 );
and \U$1240 ( \1418 , \1413 , \1417 );
_DC g12f ( \1419_nG12f , RIb4c2fa8_53 , \287 );
buf \U$1241 ( \1420 , \1419_nG12f );
and \U$1242 ( \1421 , \1420 , \343 );
and \U$1243 ( \1422 , \1417 , \1421 );
and \U$1244 ( \1423 , \1413 , \1421 );
or \U$1245 ( \1424 , \1418 , \1422 , \1423 );
xor \U$1246 ( \1425 , \1260 , \1264 );
xor \U$1247 ( \1426 , \1425 , \1269 );
and \U$1248 ( \1427 , \1424 , \1426 );
xnor \U$1249 ( \1428 , \1301 , \1304 );
and \U$1250 ( \1429 , \1426 , \1428 );
and \U$1251 ( \1430 , \1424 , \1428 );
or \U$1252 ( \1431 , \1427 , \1429 , \1430 );
and \U$1253 ( \1432 , \1409 , \1431 );
xor \U$1254 ( \1433 , \1244 , \1248 );
xor \U$1255 ( \1434 , \1433 , \1253 );
xor \U$1256 ( \1435 , \1280 , \1284 );
xor \U$1257 ( \1436 , \1435 , \1289 );
and \U$1258 ( \1437 , \1434 , \1436 );
and \U$1259 ( \1438 , \1431 , \1437 );
and \U$1260 ( \1439 , \1409 , \1437 );
or \U$1261 ( \1440 , \1432 , \1438 , \1439 );
xor \U$1262 ( \1441 , \1256 , \1272 );
xor \U$1263 ( \1442 , \1441 , \1292 );
xor \U$1264 ( \1443 , \1305 , \1309 );
xor \U$1265 ( \1444 , \1443 , \1311 );
and \U$1266 ( \1445 , \1442 , \1444 );
xor \U$1267 ( \1446 , \1317 , \1319 );
xor \U$1268 ( \1447 , \1446 , \1322 );
and \U$1269 ( \1448 , \1444 , \1447 );
and \U$1270 ( \1449 , \1442 , \1447 );
or \U$1271 ( \1450 , \1445 , \1448 , \1449 );
and \U$1272 ( \1451 , \1440 , \1450 );
xor \U$1273 ( \1452 , \1330 , \1331 );
xor \U$1274 ( \1453 , \1452 , \1333 );
and \U$1275 ( \1454 , \1450 , \1453 );
and \U$1276 ( \1455 , \1440 , \1453 );
or \U$1277 ( \1456 , \1451 , \1454 , \1455 );
xor \U$1278 ( \1457 , \1189 , \1195 );
xor \U$1279 ( \1458 , \1457 , \1201 );
and \U$1280 ( \1459 , \1456 , \1458 );
xor \U$1281 ( \1460 , \1328 , \1336 );
xor \U$1282 ( \1461 , \1460 , \1339 );
and \U$1283 ( \1462 , \1458 , \1461 );
and \U$1284 ( \1463 , \1456 , \1461 );
or \U$1285 ( \1464 , \1459 , \1462 , \1463 );
xor \U$1286 ( \1465 , \1342 , \1344 );
xor \U$1287 ( \1466 , \1465 , \1346 );
and \U$1288 ( \1467 , \1464 , \1466 );
and \U$1289 ( \1468 , \1355 , \1467 );
xor \U$1290 ( \1469 , \1355 , \1467 );
xor \U$1291 ( \1470 , \1464 , \1466 );
xor \U$1292 ( \1471 , \1170 , \1356 );
xor \U$1293 ( \1472 , \1356 , \1357 );
not \U$1294 ( \1473 , \1472 );
and \U$1295 ( \1474 , \1471 , \1473 );
and \U$1296 ( \1475 , \289 , \1474 );
not \U$1297 ( \1476 , \1475 );
xnor \U$1298 ( \1477 , \1476 , \1360 );
and \U$1299 ( \1478 , \304 , \1277 );
and \U$1300 ( \1479 , \313 , \1275 );
nor \U$1301 ( \1480 , \1478 , \1479 );
xnor \U$1302 ( \1481 , \1480 , \1173 );
and \U$1303 ( \1482 , \1477 , \1481 );
and \U$1304 ( \1483 , \322 , \1059 );
and \U$1305 ( \1484 , \331 , \1057 );
nor \U$1306 ( \1485 , \1483 , \1484 );
xnor \U$1307 ( \1486 , \1485 , \981 );
and \U$1308 ( \1487 , \1481 , \1486 );
and \U$1309 ( \1488 , \1477 , \1486 );
or \U$1310 ( \1489 , \1482 , \1487 , \1488 );
and \U$1311 ( \1490 , \342 , \911 );
and \U$1312 ( \1491 , \351 , \909 );
nor \U$1313 ( \1492 , \1490 , \1491 );
xnor \U$1314 ( \1493 , \1492 , \815 );
and \U$1315 ( \1494 , \444 , \738 );
and \U$1316 ( \1495 , \359 , \736 );
nor \U$1317 ( \1496 , \1494 , \1495 );
xnor \U$1318 ( \1497 , \1496 , \665 );
and \U$1319 ( \1498 , \1493 , \1497 );
and \U$1320 ( \1499 , \591 , \602 );
and \U$1321 ( \1500 , \494 , \600 );
nor \U$1322 ( \1501 , \1499 , \1500 );
xnor \U$1323 ( \1502 , \1501 , \558 );
and \U$1324 ( \1503 , \1497 , \1502 );
and \U$1325 ( \1504 , \1493 , \1502 );
or \U$1326 ( \1505 , \1498 , \1503 , \1504 );
and \U$1327 ( \1506 , \1489 , \1505 );
and \U$1328 ( \1507 , \701 , \502 );
and \U$1329 ( \1508 , \620 , \500 );
nor \U$1330 ( \1509 , \1507 , \1508 );
xnor \U$1331 ( \1510 , \1509 , \453 );
and \U$1332 ( \1511 , \839 , \296 );
and \U$1333 ( \1512 , \776 , \294 );
nor \U$1334 ( \1513 , \1511 , \1512 );
xnor \U$1335 ( \1514 , \1513 , \301 );
and \U$1336 ( \1515 , \1510 , \1514 );
and \U$1337 ( \1516 , \1102 , \310 );
and \U$1338 ( \1517 , \903 , \308 );
nor \U$1339 ( \1518 , \1516 , \1517 );
xnor \U$1340 ( \1519 , \1518 , \318 );
and \U$1341 ( \1520 , \1514 , \1519 );
and \U$1342 ( \1521 , \1510 , \1519 );
or \U$1343 ( \1522 , \1515 , \1520 , \1521 );
and \U$1344 ( \1523 , \1505 , \1522 );
and \U$1345 ( \1524 , \1489 , \1522 );
or \U$1346 ( \1525 , \1506 , \1523 , \1524 );
and \U$1347 ( \1526 , \1297 , \328 );
and \U$1348 ( \1527 , \1191 , \326 );
nor \U$1349 ( \1528 , \1526 , \1527 );
xnor \U$1350 ( \1529 , \1528 , \336 );
and \U$1351 ( \1530 , \1420 , \348 );
and \U$1352 ( \1531 , \1303 , \346 );
nor \U$1353 ( \1532 , \1530 , \1531 );
xnor \U$1354 ( \1533 , \1532 , \356 );
and \U$1355 ( \1534 , \1529 , \1533 );
_DC g12e ( \1535_nG12e , RIb4c2f30_54 , \287 );
buf \U$1356 ( \1536 , \1535_nG12e );
and \U$1357 ( \1537 , \1536 , \343 );
and \U$1358 ( \1538 , \1533 , \1537 );
and \U$1359 ( \1539 , \1529 , \1537 );
or \U$1360 ( \1540 , \1534 , \1538 , \1539 );
xor \U$1361 ( \1541 , \1413 , \1417 );
xor \U$1362 ( \1542 , \1541 , \1421 );
and \U$1363 ( \1543 , \1540 , \1542 );
xor \U$1364 ( \1544 , \1394 , \1398 );
xor \U$1365 ( \1545 , \1544 , \1403 );
and \U$1366 ( \1546 , \1542 , \1545 );
and \U$1367 ( \1547 , \1540 , \1545 );
or \U$1368 ( \1548 , \1543 , \1546 , \1547 );
and \U$1369 ( \1549 , \1525 , \1548 );
xor \U$1370 ( \1550 , \1361 , \1365 );
xor \U$1371 ( \1551 , \1550 , \1370 );
xor \U$1372 ( \1552 , \1377 , \1381 );
xor \U$1373 ( \1553 , \1552 , \1386 );
and \U$1374 ( \1554 , \1551 , \1553 );
and \U$1375 ( \1555 , \1548 , \1554 );
and \U$1376 ( \1556 , \1525 , \1554 );
or \U$1377 ( \1557 , \1549 , \1555 , \1556 );
xor \U$1378 ( \1558 , \1373 , \1389 );
xor \U$1379 ( \1559 , \1558 , \1406 );
xor \U$1380 ( \1560 , \1424 , \1426 );
xor \U$1381 ( \1561 , \1560 , \1428 );
and \U$1382 ( \1562 , \1559 , \1561 );
xor \U$1383 ( \1563 , \1434 , \1436 );
and \U$1384 ( \1564 , \1561 , \1563 );
and \U$1385 ( \1565 , \1559 , \1563 );
or \U$1386 ( \1566 , \1562 , \1564 , \1565 );
and \U$1387 ( \1567 , \1557 , \1566 );
xor \U$1388 ( \1568 , \1442 , \1444 );
xor \U$1389 ( \1569 , \1568 , \1447 );
and \U$1390 ( \1570 , \1566 , \1569 );
and \U$1391 ( \1571 , \1557 , \1569 );
or \U$1392 ( \1572 , \1567 , \1570 , \1571 );
xor \U$1393 ( \1573 , \1295 , \1314 );
xor \U$1394 ( \1574 , \1573 , \1325 );
and \U$1395 ( \1575 , \1572 , \1574 );
xor \U$1396 ( \1576 , \1440 , \1450 );
xor \U$1397 ( \1577 , \1576 , \1453 );
and \U$1398 ( \1578 , \1574 , \1577 );
and \U$1399 ( \1579 , \1572 , \1577 );
or \U$1400 ( \1580 , \1575 , \1578 , \1579 );
xor \U$1401 ( \1581 , \1456 , \1458 );
xor \U$1402 ( \1582 , \1581 , \1461 );
and \U$1403 ( \1583 , \1580 , \1582 );
and \U$1404 ( \1584 , \1470 , \1583 );
xor \U$1405 ( \1585 , \1470 , \1583 );
xor \U$1406 ( \1586 , \1580 , \1582 );
and \U$1407 ( \1587 , \620 , \602 );
and \U$1408 ( \1588 , \591 , \600 );
nor \U$1409 ( \1589 , \1587 , \1588 );
xnor \U$1410 ( \1590 , \1589 , \558 );
and \U$1411 ( \1591 , \776 , \502 );
and \U$1412 ( \1592 , \701 , \500 );
nor \U$1413 ( \1593 , \1591 , \1592 );
xnor \U$1414 ( \1594 , \1593 , \453 );
and \U$1415 ( \1595 , \1590 , \1594 );
and \U$1416 ( \1596 , \903 , \296 );
and \U$1417 ( \1597 , \839 , \294 );
nor \U$1418 ( \1598 , \1596 , \1597 );
xnor \U$1419 ( \1599 , \1598 , \301 );
and \U$1420 ( \1600 , \1594 , \1599 );
and \U$1421 ( \1601 , \1590 , \1599 );
or \U$1422 ( \1602 , \1595 , \1600 , \1601 );
buf \U$1423 ( \1603 , RIa166f40_24);
buf \U$1424 ( \1604 , RIa166ec8_25);
and \U$1425 ( \1605 , \1603 , \1604 );
not \U$1426 ( \1606 , \1605 );
and \U$1427 ( \1607 , \1357 , \1606 );
not \U$1428 ( \1608 , \1607 );
and \U$1429 ( \1609 , \313 , \1474 );
and \U$1430 ( \1610 , \289 , \1472 );
nor \U$1431 ( \1611 , \1609 , \1610 );
xnor \U$1432 ( \1612 , \1611 , \1360 );
and \U$1433 ( \1613 , \1608 , \1612 );
and \U$1434 ( \1614 , \331 , \1277 );
and \U$1435 ( \1615 , \304 , \1275 );
nor \U$1436 ( \1616 , \1614 , \1615 );
xnor \U$1437 ( \1617 , \1616 , \1173 );
and \U$1438 ( \1618 , \1612 , \1617 );
and \U$1439 ( \1619 , \1608 , \1617 );
or \U$1440 ( \1620 , \1613 , \1618 , \1619 );
and \U$1441 ( \1621 , \1602 , \1620 );
and \U$1442 ( \1622 , \351 , \1059 );
and \U$1443 ( \1623 , \322 , \1057 );
nor \U$1444 ( \1624 , \1622 , \1623 );
xnor \U$1445 ( \1625 , \1624 , \981 );
and \U$1446 ( \1626 , \359 , \911 );
and \U$1447 ( \1627 , \342 , \909 );
nor \U$1448 ( \1628 , \1626 , \1627 );
xnor \U$1449 ( \1629 , \1628 , \815 );
and \U$1450 ( \1630 , \1625 , \1629 );
and \U$1451 ( \1631 , \494 , \738 );
and \U$1452 ( \1632 , \444 , \736 );
nor \U$1453 ( \1633 , \1631 , \1632 );
xnor \U$1454 ( \1634 , \1633 , \665 );
and \U$1455 ( \1635 , \1629 , \1634 );
and \U$1456 ( \1636 , \1625 , \1634 );
or \U$1457 ( \1637 , \1630 , \1635 , \1636 );
and \U$1458 ( \1638 , \1620 , \1637 );
and \U$1459 ( \1639 , \1602 , \1637 );
or \U$1460 ( \1640 , \1621 , \1638 , \1639 );
xor \U$1461 ( \1641 , \1477 , \1481 );
xor \U$1462 ( \1642 , \1641 , \1486 );
xor \U$1463 ( \1643 , \1493 , \1497 );
xor \U$1464 ( \1644 , \1643 , \1502 );
and \U$1465 ( \1645 , \1642 , \1644 );
xor \U$1466 ( \1646 , \1510 , \1514 );
xor \U$1467 ( \1647 , \1646 , \1519 );
and \U$1468 ( \1648 , \1644 , \1647 );
and \U$1469 ( \1649 , \1642 , \1647 );
or \U$1470 ( \1650 , \1645 , \1648 , \1649 );
and \U$1471 ( \1651 , \1640 , \1650 );
and \U$1472 ( \1652 , \1191 , \310 );
and \U$1473 ( \1653 , \1102 , \308 );
nor \U$1474 ( \1654 , \1652 , \1653 );
xnor \U$1475 ( \1655 , \1654 , \318 );
and \U$1476 ( \1656 , \1303 , \328 );
and \U$1477 ( \1657 , \1297 , \326 );
nor \U$1478 ( \1658 , \1656 , \1657 );
xnor \U$1479 ( \1659 , \1658 , \336 );
and \U$1480 ( \1660 , \1655 , \1659 );
and \U$1481 ( \1661 , \1536 , \348 );
and \U$1482 ( \1662 , \1420 , \346 );
nor \U$1483 ( \1663 , \1661 , \1662 );
xnor \U$1484 ( \1664 , \1663 , \356 );
and \U$1485 ( \1665 , \1659 , \1664 );
and \U$1486 ( \1666 , \1655 , \1664 );
or \U$1487 ( \1667 , \1660 , \1665 , \1666 );
xor \U$1488 ( \1668 , \1529 , \1533 );
xor \U$1489 ( \1669 , \1668 , \1537 );
or \U$1490 ( \1670 , \1667 , \1669 );
and \U$1491 ( \1671 , \1650 , \1670 );
and \U$1492 ( \1672 , \1640 , \1670 );
or \U$1493 ( \1673 , \1651 , \1671 , \1672 );
xor \U$1494 ( \1674 , \1489 , \1505 );
xor \U$1495 ( \1675 , \1674 , \1522 );
xor \U$1496 ( \1676 , \1540 , \1542 );
xor \U$1497 ( \1677 , \1676 , \1545 );
and \U$1498 ( \1678 , \1675 , \1677 );
xor \U$1499 ( \1679 , \1551 , \1553 );
and \U$1500 ( \1680 , \1677 , \1679 );
and \U$1501 ( \1681 , \1675 , \1679 );
or \U$1502 ( \1682 , \1678 , \1680 , \1681 );
and \U$1503 ( \1683 , \1673 , \1682 );
xor \U$1504 ( \1684 , \1559 , \1561 );
xor \U$1505 ( \1685 , \1684 , \1563 );
and \U$1506 ( \1686 , \1682 , \1685 );
and \U$1507 ( \1687 , \1673 , \1685 );
or \U$1508 ( \1688 , \1683 , \1686 , \1687 );
xor \U$1509 ( \1689 , \1409 , \1431 );
xor \U$1510 ( \1690 , \1689 , \1437 );
and \U$1511 ( \1691 , \1688 , \1690 );
xor \U$1512 ( \1692 , \1557 , \1566 );
xor \U$1513 ( \1693 , \1692 , \1569 );
and \U$1514 ( \1694 , \1690 , \1693 );
and \U$1515 ( \1695 , \1688 , \1693 );
or \U$1516 ( \1696 , \1691 , \1694 , \1695 );
xor \U$1517 ( \1697 , \1572 , \1574 );
xor \U$1518 ( \1698 , \1697 , \1577 );
and \U$1519 ( \1699 , \1696 , \1698 );
and \U$1520 ( \1700 , \1586 , \1699 );
xor \U$1521 ( \1701 , \1586 , \1699 );
xor \U$1522 ( \1702 , \1696 , \1698 );
and \U$1523 ( \1703 , \701 , \602 );
and \U$1524 ( \1704 , \620 , \600 );
nor \U$1525 ( \1705 , \1703 , \1704 );
xnor \U$1526 ( \1706 , \1705 , \558 );
and \U$1527 ( \1707 , \839 , \502 );
and \U$1528 ( \1708 , \776 , \500 );
nor \U$1529 ( \1709 , \1707 , \1708 );
xnor \U$1530 ( \1710 , \1709 , \453 );
and \U$1531 ( \1711 , \1706 , \1710 );
and \U$1532 ( \1712 , \1102 , \296 );
and \U$1533 ( \1713 , \903 , \294 );
nor \U$1534 ( \1714 , \1712 , \1713 );
xnor \U$1535 ( \1715 , \1714 , \301 );
and \U$1536 ( \1716 , \1710 , \1715 );
and \U$1537 ( \1717 , \1706 , \1715 );
or \U$1538 ( \1718 , \1711 , \1716 , \1717 );
and \U$1539 ( \1719 , \342 , \1059 );
and \U$1540 ( \1720 , \351 , \1057 );
nor \U$1541 ( \1721 , \1719 , \1720 );
xnor \U$1542 ( \1722 , \1721 , \981 );
and \U$1543 ( \1723 , \444 , \911 );
and \U$1544 ( \1724 , \359 , \909 );
nor \U$1545 ( \1725 , \1723 , \1724 );
xnor \U$1546 ( \1726 , \1725 , \815 );
and \U$1547 ( \1727 , \1722 , \1726 );
and \U$1548 ( \1728 , \591 , \738 );
and \U$1549 ( \1729 , \494 , \736 );
nor \U$1550 ( \1730 , \1728 , \1729 );
xnor \U$1551 ( \1731 , \1730 , \665 );
and \U$1552 ( \1732 , \1726 , \1731 );
and \U$1553 ( \1733 , \1722 , \1731 );
or \U$1554 ( \1734 , \1727 , \1732 , \1733 );
and \U$1555 ( \1735 , \1718 , \1734 );
xor \U$1556 ( \1736 , \1357 , \1603 );
xor \U$1557 ( \1737 , \1603 , \1604 );
not \U$1558 ( \1738 , \1737 );
and \U$1559 ( \1739 , \1736 , \1738 );
and \U$1560 ( \1740 , \289 , \1739 );
not \U$1561 ( \1741 , \1740 );
xnor \U$1562 ( \1742 , \1741 , \1607 );
and \U$1563 ( \1743 , \304 , \1474 );
and \U$1564 ( \1744 , \313 , \1472 );
nor \U$1565 ( \1745 , \1743 , \1744 );
xnor \U$1566 ( \1746 , \1745 , \1360 );
and \U$1567 ( \1747 , \1742 , \1746 );
and \U$1568 ( \1748 , \322 , \1277 );
and \U$1569 ( \1749 , \331 , \1275 );
nor \U$1570 ( \1750 , \1748 , \1749 );
xnor \U$1571 ( \1751 , \1750 , \1173 );
and \U$1572 ( \1752 , \1746 , \1751 );
and \U$1573 ( \1753 , \1742 , \1751 );
or \U$1574 ( \1754 , \1747 , \1752 , \1753 );
and \U$1575 ( \1755 , \1734 , \1754 );
and \U$1576 ( \1756 , \1718 , \1754 );
or \U$1577 ( \1757 , \1735 , \1755 , \1756 );
and \U$1578 ( \1758 , \1297 , \310 );
and \U$1579 ( \1759 , \1191 , \308 );
nor \U$1580 ( \1760 , \1758 , \1759 );
xnor \U$1581 ( \1761 , \1760 , \318 );
and \U$1582 ( \1762 , \1420 , \328 );
and \U$1583 ( \1763 , \1303 , \326 );
nor \U$1584 ( \1764 , \1762 , \1763 );
xnor \U$1585 ( \1765 , \1764 , \336 );
and \U$1586 ( \1766 , \1761 , \1765 );
_DC g12d ( \1767_nG12d , RIb4c2eb8_55 , \287 );
buf \U$1587 ( \1768 , \1767_nG12d );
and \U$1588 ( \1769 , \1768 , \348 );
and \U$1589 ( \1770 , \1536 , \346 );
nor \U$1590 ( \1771 , \1769 , \1770 );
xnor \U$1591 ( \1772 , \1771 , \356 );
and \U$1592 ( \1773 , \1765 , \1772 );
and \U$1593 ( \1774 , \1761 , \1772 );
or \U$1594 ( \1775 , \1766 , \1773 , \1774 );
_DC g12c ( \1776_nG12c , RIb4c2e40_56 , \287 );
buf \U$1595 ( \1777 , \1776_nG12c );
and \U$1596 ( \1778 , \1777 , \343 );
buf \U$1597 ( \1779 , \1778 );
and \U$1598 ( \1780 , \1775 , \1779 );
and \U$1599 ( \1781 , \1768 , \343 );
and \U$1600 ( \1782 , \1779 , \1781 );
and \U$1601 ( \1783 , \1775 , \1781 );
or \U$1602 ( \1784 , \1780 , \1782 , \1783 );
and \U$1603 ( \1785 , \1757 , \1784 );
xor \U$1604 ( \1786 , \1655 , \1659 );
xor \U$1605 ( \1787 , \1786 , \1664 );
xor \U$1606 ( \1788 , \1590 , \1594 );
xor \U$1607 ( \1789 , \1788 , \1599 );
and \U$1608 ( \1790 , \1787 , \1789 );
xor \U$1609 ( \1791 , \1625 , \1629 );
xor \U$1610 ( \1792 , \1791 , \1634 );
and \U$1611 ( \1793 , \1789 , \1792 );
and \U$1612 ( \1794 , \1787 , \1792 );
or \U$1613 ( \1795 , \1790 , \1793 , \1794 );
and \U$1614 ( \1796 , \1784 , \1795 );
and \U$1615 ( \1797 , \1757 , \1795 );
or \U$1616 ( \1798 , \1785 , \1796 , \1797 );
xor \U$1617 ( \1799 , \1602 , \1620 );
xor \U$1618 ( \1800 , \1799 , \1637 );
xor \U$1619 ( \1801 , \1642 , \1644 );
xor \U$1620 ( \1802 , \1801 , \1647 );
and \U$1621 ( \1803 , \1800 , \1802 );
xnor \U$1622 ( \1804 , \1667 , \1669 );
and \U$1623 ( \1805 , \1802 , \1804 );
and \U$1624 ( \1806 , \1800 , \1804 );
or \U$1625 ( \1807 , \1803 , \1805 , \1806 );
and \U$1626 ( \1808 , \1798 , \1807 );
xor \U$1627 ( \1809 , \1675 , \1677 );
xor \U$1628 ( \1810 , \1809 , \1679 );
and \U$1629 ( \1811 , \1807 , \1810 );
and \U$1630 ( \1812 , \1798 , \1810 );
or \U$1631 ( \1813 , \1808 , \1811 , \1812 );
xor \U$1632 ( \1814 , \1525 , \1548 );
xor \U$1633 ( \1815 , \1814 , \1554 );
and \U$1634 ( \1816 , \1813 , \1815 );
xor \U$1635 ( \1817 , \1673 , \1682 );
xor \U$1636 ( \1818 , \1817 , \1685 );
and \U$1637 ( \1819 , \1815 , \1818 );
and \U$1638 ( \1820 , \1813 , \1818 );
or \U$1639 ( \1821 , \1816 , \1819 , \1820 );
xor \U$1640 ( \1822 , \1688 , \1690 );
xor \U$1641 ( \1823 , \1822 , \1693 );
and \U$1642 ( \1824 , \1821 , \1823 );
and \U$1643 ( \1825 , \1702 , \1824 );
xor \U$1644 ( \1826 , \1702 , \1824 );
xor \U$1645 ( \1827 , \1821 , \1823 );
buf \U$1646 ( \1828 , RIa166e50_26);
buf \U$1647 ( \1829 , RIa166dd8_27);
and \U$1648 ( \1830 , \1828 , \1829 );
not \U$1649 ( \1831 , \1830 );
and \U$1650 ( \1832 , \1604 , \1831 );
not \U$1651 ( \1833 , \1832 );
and \U$1652 ( \1834 , \313 , \1739 );
and \U$1653 ( \1835 , \289 , \1737 );
nor \U$1654 ( \1836 , \1834 , \1835 );
xnor \U$1655 ( \1837 , \1836 , \1607 );
and \U$1656 ( \1838 , \1833 , \1837 );
and \U$1657 ( \1839 , \331 , \1474 );
and \U$1658 ( \1840 , \304 , \1472 );
nor \U$1659 ( \1841 , \1839 , \1840 );
xnor \U$1660 ( \1842 , \1841 , \1360 );
and \U$1661 ( \1843 , \1837 , \1842 );
and \U$1662 ( \1844 , \1833 , \1842 );
or \U$1663 ( \1845 , \1838 , \1843 , \1844 );
and \U$1664 ( \1846 , \351 , \1277 );
and \U$1665 ( \1847 , \322 , \1275 );
nor \U$1666 ( \1848 , \1846 , \1847 );
xnor \U$1667 ( \1849 , \1848 , \1173 );
and \U$1668 ( \1850 , \359 , \1059 );
and \U$1669 ( \1851 , \342 , \1057 );
nor \U$1670 ( \1852 , \1850 , \1851 );
xnor \U$1671 ( \1853 , \1852 , \981 );
and \U$1672 ( \1854 , \1849 , \1853 );
and \U$1673 ( \1855 , \494 , \911 );
and \U$1674 ( \1856 , \444 , \909 );
nor \U$1675 ( \1857 , \1855 , \1856 );
xnor \U$1676 ( \1858 , \1857 , \815 );
and \U$1677 ( \1859 , \1853 , \1858 );
and \U$1678 ( \1860 , \1849 , \1858 );
or \U$1679 ( \1861 , \1854 , \1859 , \1860 );
and \U$1680 ( \1862 , \1845 , \1861 );
and \U$1681 ( \1863 , \620 , \738 );
and \U$1682 ( \1864 , \591 , \736 );
nor \U$1683 ( \1865 , \1863 , \1864 );
xnor \U$1684 ( \1866 , \1865 , \665 );
and \U$1685 ( \1867 , \776 , \602 );
and \U$1686 ( \1868 , \701 , \600 );
nor \U$1687 ( \1869 , \1867 , \1868 );
xnor \U$1688 ( \1870 , \1869 , \558 );
and \U$1689 ( \1871 , \1866 , \1870 );
and \U$1690 ( \1872 , \903 , \502 );
and \U$1691 ( \1873 , \839 , \500 );
nor \U$1692 ( \1874 , \1872 , \1873 );
xnor \U$1693 ( \1875 , \1874 , \453 );
and \U$1694 ( \1876 , \1870 , \1875 );
and \U$1695 ( \1877 , \1866 , \1875 );
or \U$1696 ( \1878 , \1871 , \1876 , \1877 );
and \U$1697 ( \1879 , \1861 , \1878 );
and \U$1698 ( \1880 , \1845 , \1878 );
or \U$1699 ( \1881 , \1862 , \1879 , \1880 );
xor \U$1700 ( \1882 , \1706 , \1710 );
xor \U$1701 ( \1883 , \1882 , \1715 );
xor \U$1702 ( \1884 , \1722 , \1726 );
xor \U$1703 ( \1885 , \1884 , \1731 );
and \U$1704 ( \1886 , \1883 , \1885 );
xor \U$1705 ( \1887 , \1742 , \1746 );
xor \U$1706 ( \1888 , \1887 , \1751 );
and \U$1707 ( \1889 , \1885 , \1888 );
and \U$1708 ( \1890 , \1883 , \1888 );
or \U$1709 ( \1891 , \1886 , \1889 , \1890 );
and \U$1710 ( \1892 , \1881 , \1891 );
and \U$1711 ( \1893 , \1191 , \296 );
and \U$1712 ( \1894 , \1102 , \294 );
nor \U$1713 ( \1895 , \1893 , \1894 );
xnor \U$1714 ( \1896 , \1895 , \301 );
and \U$1715 ( \1897 , \1303 , \310 );
and \U$1716 ( \1898 , \1297 , \308 );
nor \U$1717 ( \1899 , \1897 , \1898 );
xnor \U$1718 ( \1900 , \1899 , \318 );
and \U$1719 ( \1901 , \1896 , \1900 );
and \U$1720 ( \1902 , \1536 , \328 );
and \U$1721 ( \1903 , \1420 , \326 );
nor \U$1722 ( \1904 , \1902 , \1903 );
xnor \U$1723 ( \1905 , \1904 , \336 );
and \U$1724 ( \1906 , \1900 , \1905 );
and \U$1725 ( \1907 , \1896 , \1905 );
or \U$1726 ( \1908 , \1901 , \1906 , \1907 );
xor \U$1727 ( \1909 , \1761 , \1765 );
xor \U$1728 ( \1910 , \1909 , \1772 );
and \U$1729 ( \1911 , \1908 , \1910 );
not \U$1730 ( \1912 , \1778 );
and \U$1731 ( \1913 , \1910 , \1912 );
and \U$1732 ( \1914 , \1908 , \1912 );
or \U$1733 ( \1915 , \1911 , \1913 , \1914 );
and \U$1734 ( \1916 , \1891 , \1915 );
and \U$1735 ( \1917 , \1881 , \1915 );
or \U$1736 ( \1918 , \1892 , \1916 , \1917 );
xor \U$1737 ( \1919 , \1608 , \1612 );
xor \U$1738 ( \1920 , \1919 , \1617 );
xor \U$1739 ( \1921 , \1775 , \1779 );
xor \U$1740 ( \1922 , \1921 , \1781 );
and \U$1741 ( \1923 , \1920 , \1922 );
xor \U$1742 ( \1924 , \1787 , \1789 );
xor \U$1743 ( \1925 , \1924 , \1792 );
and \U$1744 ( \1926 , \1922 , \1925 );
and \U$1745 ( \1927 , \1920 , \1925 );
or \U$1746 ( \1928 , \1923 , \1926 , \1927 );
and \U$1747 ( \1929 , \1918 , \1928 );
xor \U$1748 ( \1930 , \1800 , \1802 );
xor \U$1749 ( \1931 , \1930 , \1804 );
and \U$1750 ( \1932 , \1928 , \1931 );
and \U$1751 ( \1933 , \1918 , \1931 );
or \U$1752 ( \1934 , \1929 , \1932 , \1933 );
xor \U$1753 ( \1935 , \1640 , \1650 );
xor \U$1754 ( \1936 , \1935 , \1670 );
and \U$1755 ( \1937 , \1934 , \1936 );
xor \U$1756 ( \1938 , \1798 , \1807 );
xor \U$1757 ( \1939 , \1938 , \1810 );
and \U$1758 ( \1940 , \1936 , \1939 );
and \U$1759 ( \1941 , \1934 , \1939 );
or \U$1760 ( \1942 , \1937 , \1940 , \1941 );
xor \U$1761 ( \1943 , \1813 , \1815 );
xor \U$1762 ( \1944 , \1943 , \1818 );
and \U$1763 ( \1945 , \1942 , \1944 );
and \U$1764 ( \1946 , \1827 , \1945 );
xor \U$1765 ( \1947 , \1827 , \1945 );
xor \U$1766 ( \1948 , \1942 , \1944 );
xor \U$1767 ( \1949 , \1604 , \1828 );
xor \U$1768 ( \1950 , \1828 , \1829 );
not \U$1769 ( \1951 , \1950 );
and \U$1770 ( \1952 , \1949 , \1951 );
and \U$1771 ( \1953 , \289 , \1952 );
not \U$1772 ( \1954 , \1953 );
xnor \U$1773 ( \1955 , \1954 , \1832 );
and \U$1774 ( \1956 , \304 , \1739 );
and \U$1775 ( \1957 , \313 , \1737 );
nor \U$1776 ( \1958 , \1956 , \1957 );
xnor \U$1777 ( \1959 , \1958 , \1607 );
and \U$1778 ( \1960 , \1955 , \1959 );
and \U$1779 ( \1961 , \322 , \1474 );
and \U$1780 ( \1962 , \331 , \1472 );
nor \U$1781 ( \1963 , \1961 , \1962 );
xnor \U$1782 ( \1964 , \1963 , \1360 );
and \U$1783 ( \1965 , \1959 , \1964 );
and \U$1784 ( \1966 , \1955 , \1964 );
or \U$1785 ( \1967 , \1960 , \1965 , \1966 );
and \U$1786 ( \1968 , \342 , \1277 );
and \U$1787 ( \1969 , \351 , \1275 );
nor \U$1788 ( \1970 , \1968 , \1969 );
xnor \U$1789 ( \1971 , \1970 , \1173 );
and \U$1790 ( \1972 , \444 , \1059 );
and \U$1791 ( \1973 , \359 , \1057 );
nor \U$1792 ( \1974 , \1972 , \1973 );
xnor \U$1793 ( \1975 , \1974 , \981 );
and \U$1794 ( \1976 , \1971 , \1975 );
and \U$1795 ( \1977 , \591 , \911 );
and \U$1796 ( \1978 , \494 , \909 );
nor \U$1797 ( \1979 , \1977 , \1978 );
xnor \U$1798 ( \1980 , \1979 , \815 );
and \U$1799 ( \1981 , \1975 , \1980 );
and \U$1800 ( \1982 , \1971 , \1980 );
or \U$1801 ( \1983 , \1976 , \1981 , \1982 );
and \U$1802 ( \1984 , \1967 , \1983 );
and \U$1803 ( \1985 , \701 , \738 );
and \U$1804 ( \1986 , \620 , \736 );
nor \U$1805 ( \1987 , \1985 , \1986 );
xnor \U$1806 ( \1988 , \1987 , \665 );
and \U$1807 ( \1989 , \839 , \602 );
and \U$1808 ( \1990 , \776 , \600 );
nor \U$1809 ( \1991 , \1989 , \1990 );
xnor \U$1810 ( \1992 , \1991 , \558 );
and \U$1811 ( \1993 , \1988 , \1992 );
and \U$1812 ( \1994 , \1102 , \502 );
and \U$1813 ( \1995 , \903 , \500 );
nor \U$1814 ( \1996 , \1994 , \1995 );
xnor \U$1815 ( \1997 , \1996 , \453 );
and \U$1816 ( \1998 , \1992 , \1997 );
and \U$1817 ( \1999 , \1988 , \1997 );
or \U$1818 ( \2000 , \1993 , \1998 , \1999 );
and \U$1819 ( \2001 , \1983 , \2000 );
and \U$1820 ( \2002 , \1967 , \2000 );
or \U$1821 ( \2003 , \1984 , \2001 , \2002 );
and \U$1822 ( \2004 , \1297 , \296 );
and \U$1823 ( \2005 , \1191 , \294 );
nor \U$1824 ( \2006 , \2004 , \2005 );
xnor \U$1825 ( \2007 , \2006 , \301 );
and \U$1826 ( \2008 , \1420 , \310 );
and \U$1827 ( \2009 , \1303 , \308 );
nor \U$1828 ( \2010 , \2008 , \2009 );
xnor \U$1829 ( \2011 , \2010 , \318 );
and \U$1830 ( \2012 , \2007 , \2011 );
and \U$1831 ( \2013 , \1768 , \328 );
and \U$1832 ( \2014 , \1536 , \326 );
nor \U$1833 ( \2015 , \2013 , \2014 );
xnor \U$1834 ( \2016 , \2015 , \336 );
and \U$1835 ( \2017 , \2011 , \2016 );
and \U$1836 ( \2018 , \2007 , \2016 );
or \U$1837 ( \2019 , \2012 , \2017 , \2018 );
_DC g12b ( \2020_nG12b , RIb4c2dc8_57 , \287 );
buf \U$1838 ( \2021 , \2020_nG12b );
and \U$1839 ( \2022 , \2021 , \348 );
and \U$1840 ( \2023 , \1777 , \346 );
nor \U$1841 ( \2024 , \2022 , \2023 );
xnor \U$1842 ( \2025 , \2024 , \356 );
_DC g12a ( \2026_nG12a , RIb4c2d50_58 , \287 );
buf \U$1843 ( \2027 , \2026_nG12a );
and \U$1844 ( \2028 , \2027 , \343 );
or \U$1845 ( \2029 , \2025 , \2028 );
and \U$1846 ( \2030 , \2019 , \2029 );
and \U$1847 ( \2031 , \1777 , \348 );
and \U$1848 ( \2032 , \1768 , \346 );
nor \U$1849 ( \2033 , \2031 , \2032 );
xnor \U$1850 ( \2034 , \2033 , \356 );
and \U$1851 ( \2035 , \2029 , \2034 );
and \U$1852 ( \2036 , \2019 , \2034 );
or \U$1853 ( \2037 , \2030 , \2035 , \2036 );
and \U$1854 ( \2038 , \2003 , \2037 );
and \U$1855 ( \2039 , \2021 , \343 );
xor \U$1856 ( \2040 , \1896 , \1900 );
xor \U$1857 ( \2041 , \2040 , \1905 );
and \U$1858 ( \2042 , \2039 , \2041 );
xor \U$1859 ( \2043 , \1866 , \1870 );
xor \U$1860 ( \2044 , \2043 , \1875 );
and \U$1861 ( \2045 , \2041 , \2044 );
and \U$1862 ( \2046 , \2039 , \2044 );
or \U$1863 ( \2047 , \2042 , \2045 , \2046 );
and \U$1864 ( \2048 , \2037 , \2047 );
and \U$1865 ( \2049 , \2003 , \2047 );
or \U$1866 ( \2050 , \2038 , \2048 , \2049 );
xor \U$1867 ( \2051 , \1845 , \1861 );
xor \U$1868 ( \2052 , \2051 , \1878 );
xor \U$1869 ( \2053 , \1883 , \1885 );
xor \U$1870 ( \2054 , \2053 , \1888 );
and \U$1871 ( \2055 , \2052 , \2054 );
xor \U$1872 ( \2056 , \1908 , \1910 );
xor \U$1873 ( \2057 , \2056 , \1912 );
and \U$1874 ( \2058 , \2054 , \2057 );
and \U$1875 ( \2059 , \2052 , \2057 );
or \U$1876 ( \2060 , \2055 , \2058 , \2059 );
and \U$1877 ( \2061 , \2050 , \2060 );
xor \U$1878 ( \2062 , \1718 , \1734 );
xor \U$1879 ( \2063 , \2062 , \1754 );
and \U$1880 ( \2064 , \2060 , \2063 );
and \U$1881 ( \2065 , \2050 , \2063 );
or \U$1882 ( \2066 , \2061 , \2064 , \2065 );
xor \U$1883 ( \2067 , \1881 , \1891 );
xor \U$1884 ( \2068 , \2067 , \1915 );
xor \U$1885 ( \2069 , \1920 , \1922 );
xor \U$1886 ( \2070 , \2069 , \1925 );
and \U$1887 ( \2071 , \2068 , \2070 );
and \U$1888 ( \2072 , \2066 , \2071 );
xor \U$1889 ( \2073 , \1757 , \1784 );
xor \U$1890 ( \2074 , \2073 , \1795 );
and \U$1891 ( \2075 , \2071 , \2074 );
and \U$1892 ( \2076 , \2066 , \2074 );
or \U$1893 ( \2077 , \2072 , \2075 , \2076 );
xor \U$1894 ( \2078 , \1934 , \1936 );
xor \U$1895 ( \2079 , \2078 , \1939 );
and \U$1896 ( \2080 , \2077 , \2079 );
and \U$1897 ( \2081 , \1948 , \2080 );
xor \U$1898 ( \2082 , \1948 , \2080 );
xor \U$1899 ( \2083 , \2077 , \2079 );
and \U$1900 ( \2084 , \620 , \911 );
and \U$1901 ( \2085 , \591 , \909 );
nor \U$1902 ( \2086 , \2084 , \2085 );
xnor \U$1903 ( \2087 , \2086 , \815 );
and \U$1904 ( \2088 , \776 , \738 );
and \U$1905 ( \2089 , \701 , \736 );
nor \U$1906 ( \2090 , \2088 , \2089 );
xnor \U$1907 ( \2091 , \2090 , \665 );
and \U$1908 ( \2092 , \2087 , \2091 );
and \U$1909 ( \2093 , \903 , \602 );
and \U$1910 ( \2094 , \839 , \600 );
nor \U$1911 ( \2095 , \2093 , \2094 );
xnor \U$1912 ( \2096 , \2095 , \558 );
and \U$1913 ( \2097 , \2091 , \2096 );
and \U$1914 ( \2098 , \2087 , \2096 );
or \U$1915 ( \2099 , \2092 , \2097 , \2098 );
and \U$1916 ( \2100 , \351 , \1474 );
and \U$1917 ( \2101 , \322 , \1472 );
nor \U$1918 ( \2102 , \2100 , \2101 );
xnor \U$1919 ( \2103 , \2102 , \1360 );
and \U$1920 ( \2104 , \359 , \1277 );
and \U$1921 ( \2105 , \342 , \1275 );
nor \U$1922 ( \2106 , \2104 , \2105 );
xnor \U$1923 ( \2107 , \2106 , \1173 );
and \U$1924 ( \2108 , \2103 , \2107 );
and \U$1925 ( \2109 , \494 , \1059 );
and \U$1926 ( \2110 , \444 , \1057 );
nor \U$1927 ( \2111 , \2109 , \2110 );
xnor \U$1928 ( \2112 , \2111 , \981 );
and \U$1929 ( \2113 , \2107 , \2112 );
and \U$1930 ( \2114 , \2103 , \2112 );
or \U$1931 ( \2115 , \2108 , \2113 , \2114 );
and \U$1932 ( \2116 , \2099 , \2115 );
buf \U$1933 ( \2117 , RIa166d60_28);
buf \U$1934 ( \2118 , RIa166ce8_29);
and \U$1935 ( \2119 , \2117 , \2118 );
not \U$1936 ( \2120 , \2119 );
and \U$1937 ( \2121 , \1829 , \2120 );
not \U$1938 ( \2122 , \2121 );
and \U$1939 ( \2123 , \313 , \1952 );
and \U$1940 ( \2124 , \289 , \1950 );
nor \U$1941 ( \2125 , \2123 , \2124 );
xnor \U$1942 ( \2126 , \2125 , \1832 );
and \U$1943 ( \2127 , \2122 , \2126 );
and \U$1944 ( \2128 , \331 , \1739 );
and \U$1945 ( \2129 , \304 , \1737 );
nor \U$1946 ( \2130 , \2128 , \2129 );
xnor \U$1947 ( \2131 , \2130 , \1607 );
and \U$1948 ( \2132 , \2126 , \2131 );
and \U$1949 ( \2133 , \2122 , \2131 );
or \U$1950 ( \2134 , \2127 , \2132 , \2133 );
and \U$1951 ( \2135 , \2115 , \2134 );
and \U$1952 ( \2136 , \2099 , \2134 );
or \U$1953 ( \2137 , \2116 , \2135 , \2136 );
xor \U$1954 ( \2138 , \2007 , \2011 );
xor \U$1955 ( \2139 , \2138 , \2016 );
xor \U$1956 ( \2140 , \1971 , \1975 );
xor \U$1957 ( \2141 , \2140 , \1980 );
and \U$1958 ( \2142 , \2139 , \2141 );
xor \U$1959 ( \2143 , \1988 , \1992 );
xor \U$1960 ( \2144 , \2143 , \1997 );
and \U$1961 ( \2145 , \2141 , \2144 );
and \U$1962 ( \2146 , \2139 , \2144 );
or \U$1963 ( \2147 , \2142 , \2145 , \2146 );
and \U$1964 ( \2148 , \2137 , \2147 );
and \U$1965 ( \2149 , \1777 , \328 );
and \U$1966 ( \2150 , \1768 , \326 );
nor \U$1967 ( \2151 , \2149 , \2150 );
xnor \U$1968 ( \2152 , \2151 , \336 );
and \U$1969 ( \2153 , \2027 , \348 );
and \U$1970 ( \2154 , \2021 , \346 );
nor \U$1971 ( \2155 , \2153 , \2154 );
xnor \U$1972 ( \2156 , \2155 , \356 );
and \U$1973 ( \2157 , \2152 , \2156 );
_DC g129 ( \2158_nG129 , RIb4c2cd8_59 , \287 );
buf \U$1974 ( \2159 , \2158_nG129 );
and \U$1975 ( \2160 , \2159 , \343 );
and \U$1976 ( \2161 , \2156 , \2160 );
and \U$1977 ( \2162 , \2152 , \2160 );
or \U$1978 ( \2163 , \2157 , \2161 , \2162 );
and \U$1979 ( \2164 , \1191 , \502 );
and \U$1980 ( \2165 , \1102 , \500 );
nor \U$1981 ( \2166 , \2164 , \2165 );
xnor \U$1982 ( \2167 , \2166 , \453 );
and \U$1983 ( \2168 , \1303 , \296 );
and \U$1984 ( \2169 , \1297 , \294 );
nor \U$1985 ( \2170 , \2168 , \2169 );
xnor \U$1986 ( \2171 , \2170 , \301 );
and \U$1987 ( \2172 , \2167 , \2171 );
and \U$1988 ( \2173 , \1536 , \310 );
and \U$1989 ( \2174 , \1420 , \308 );
nor \U$1990 ( \2175 , \2173 , \2174 );
xnor \U$1991 ( \2176 , \2175 , \318 );
and \U$1992 ( \2177 , \2171 , \2176 );
and \U$1993 ( \2178 , \2167 , \2176 );
or \U$1994 ( \2179 , \2172 , \2177 , \2178 );
and \U$1995 ( \2180 , \2163 , \2179 );
xnor \U$1996 ( \2181 , \2025 , \2028 );
and \U$1997 ( \2182 , \2179 , \2181 );
and \U$1998 ( \2183 , \2163 , \2181 );
or \U$1999 ( \2184 , \2180 , \2182 , \2183 );
and \U$2000 ( \2185 , \2147 , \2184 );
and \U$2001 ( \2186 , \2137 , \2184 );
or \U$2002 ( \2187 , \2148 , \2185 , \2186 );
xor \U$2003 ( \2188 , \1833 , \1837 );
xor \U$2004 ( \2189 , \2188 , \1842 );
xor \U$2005 ( \2190 , \1849 , \1853 );
xor \U$2006 ( \2191 , \2190 , \1858 );
and \U$2007 ( \2192 , \2189 , \2191 );
xor \U$2008 ( \2193 , \2039 , \2041 );
xor \U$2009 ( \2194 , \2193 , \2044 );
and \U$2010 ( \2195 , \2191 , \2194 );
and \U$2011 ( \2196 , \2189 , \2194 );
or \U$2012 ( \2197 , \2192 , \2195 , \2196 );
and \U$2013 ( \2198 , \2187 , \2197 );
xor \U$2014 ( \2199 , \2052 , \2054 );
xor \U$2015 ( \2200 , \2199 , \2057 );
and \U$2016 ( \2201 , \2197 , \2200 );
and \U$2017 ( \2202 , \2187 , \2200 );
or \U$2018 ( \2203 , \2198 , \2201 , \2202 );
xor \U$2019 ( \2204 , \2050 , \2060 );
xor \U$2020 ( \2205 , \2204 , \2063 );
and \U$2021 ( \2206 , \2203 , \2205 );
xor \U$2022 ( \2207 , \2068 , \2070 );
and \U$2023 ( \2208 , \2205 , \2207 );
and \U$2024 ( \2209 , \2203 , \2207 );
or \U$2025 ( \2210 , \2206 , \2208 , \2209 );
xor \U$2026 ( \2211 , \2066 , \2071 );
xor \U$2027 ( \2212 , \2211 , \2074 );
and \U$2028 ( \2213 , \2210 , \2212 );
xor \U$2029 ( \2214 , \1918 , \1928 );
xor \U$2030 ( \2215 , \2214 , \1931 );
and \U$2031 ( \2216 , \2212 , \2215 );
and \U$2032 ( \2217 , \2210 , \2215 );
or \U$2033 ( \2218 , \2213 , \2216 , \2217 );
and \U$2034 ( \2219 , \2083 , \2218 );
xor \U$2035 ( \2220 , \2083 , \2218 );
xor \U$2036 ( \2221 , \2210 , \2212 );
xor \U$2037 ( \2222 , \2221 , \2215 );
and \U$2038 ( \2223 , \701 , \911 );
and \U$2039 ( \2224 , \620 , \909 );
nor \U$2040 ( \2225 , \2223 , \2224 );
xnor \U$2041 ( \2226 , \2225 , \815 );
and \U$2042 ( \2227 , \839 , \738 );
and \U$2043 ( \2228 , \776 , \736 );
nor \U$2044 ( \2229 , \2227 , \2228 );
xnor \U$2045 ( \2230 , \2229 , \665 );
and \U$2046 ( \2231 , \2226 , \2230 );
and \U$2047 ( \2232 , \1102 , \602 );
and \U$2048 ( \2233 , \903 , \600 );
nor \U$2049 ( \2234 , \2232 , \2233 );
xnor \U$2050 ( \2235 , \2234 , \558 );
and \U$2051 ( \2236 , \2230 , \2235 );
and \U$2052 ( \2237 , \2226 , \2235 );
or \U$2053 ( \2238 , \2231 , \2236 , \2237 );
and \U$2054 ( \2239 , \342 , \1474 );
and \U$2055 ( \2240 , \351 , \1472 );
nor \U$2056 ( \2241 , \2239 , \2240 );
xnor \U$2057 ( \2242 , \2241 , \1360 );
and \U$2058 ( \2243 , \444 , \1277 );
and \U$2059 ( \2244 , \359 , \1275 );
nor \U$2060 ( \2245 , \2243 , \2244 );
xnor \U$2061 ( \2246 , \2245 , \1173 );
and \U$2062 ( \2247 , \2242 , \2246 );
and \U$2063 ( \2248 , \591 , \1059 );
and \U$2064 ( \2249 , \494 , \1057 );
nor \U$2065 ( \2250 , \2248 , \2249 );
xnor \U$2066 ( \2251 , \2250 , \981 );
and \U$2067 ( \2252 , \2246 , \2251 );
and \U$2068 ( \2253 , \2242 , \2251 );
or \U$2069 ( \2254 , \2247 , \2252 , \2253 );
and \U$2070 ( \2255 , \2238 , \2254 );
xor \U$2071 ( \2256 , \1829 , \2117 );
xor \U$2072 ( \2257 , \2117 , \2118 );
not \U$2073 ( \2258 , \2257 );
and \U$2074 ( \2259 , \2256 , \2258 );
and \U$2075 ( \2260 , \289 , \2259 );
not \U$2076 ( \2261 , \2260 );
xnor \U$2077 ( \2262 , \2261 , \2121 );
and \U$2078 ( \2263 , \304 , \1952 );
and \U$2079 ( \2264 , \313 , \1950 );
nor \U$2080 ( \2265 , \2263 , \2264 );
xnor \U$2081 ( \2266 , \2265 , \1832 );
and \U$2082 ( \2267 , \2262 , \2266 );
and \U$2083 ( \2268 , \322 , \1739 );
and \U$2084 ( \2269 , \331 , \1737 );
nor \U$2085 ( \2270 , \2268 , \2269 );
xnor \U$2086 ( \2271 , \2270 , \1607 );
and \U$2087 ( \2272 , \2266 , \2271 );
and \U$2088 ( \2273 , \2262 , \2271 );
or \U$2089 ( \2274 , \2267 , \2272 , \2273 );
and \U$2090 ( \2275 , \2254 , \2274 );
and \U$2091 ( \2276 , \2238 , \2274 );
or \U$2092 ( \2277 , \2255 , \2275 , \2276 );
and \U$2093 ( \2278 , \1297 , \502 );
and \U$2094 ( \2279 , \1191 , \500 );
nor \U$2095 ( \2280 , \2278 , \2279 );
xnor \U$2096 ( \2281 , \2280 , \453 );
and \U$2097 ( \2282 , \1420 , \296 );
and \U$2098 ( \2283 , \1303 , \294 );
nor \U$2099 ( \2284 , \2282 , \2283 );
xnor \U$2100 ( \2285 , \2284 , \301 );
and \U$2101 ( \2286 , \2281 , \2285 );
and \U$2102 ( \2287 , \1768 , \310 );
and \U$2103 ( \2288 , \1536 , \308 );
nor \U$2104 ( \2289 , \2287 , \2288 );
xnor \U$2105 ( \2290 , \2289 , \318 );
and \U$2106 ( \2291 , \2285 , \2290 );
and \U$2107 ( \2292 , \2281 , \2290 );
or \U$2108 ( \2293 , \2286 , \2291 , \2292 );
and \U$2109 ( \2294 , \2021 , \328 );
and \U$2110 ( \2295 , \1777 , \326 );
nor \U$2111 ( \2296 , \2294 , \2295 );
xnor \U$2112 ( \2297 , \2296 , \336 );
and \U$2113 ( \2298 , \2159 , \348 );
and \U$2114 ( \2299 , \2027 , \346 );
nor \U$2115 ( \2300 , \2298 , \2299 );
xnor \U$2116 ( \2301 , \2300 , \356 );
and \U$2117 ( \2302 , \2297 , \2301 );
_DC g128 ( \2303_nG128 , RIb4c2c60_60 , \287 );
buf \U$2118 ( \2304 , \2303_nG128 );
and \U$2119 ( \2305 , \2304 , \343 );
and \U$2120 ( \2306 , \2301 , \2305 );
and \U$2121 ( \2307 , \2297 , \2305 );
or \U$2122 ( \2308 , \2302 , \2306 , \2307 );
and \U$2123 ( \2309 , \2293 , \2308 );
xor \U$2124 ( \2310 , \2152 , \2156 );
xor \U$2125 ( \2311 , \2310 , \2160 );
and \U$2126 ( \2312 , \2308 , \2311 );
and \U$2127 ( \2313 , \2293 , \2311 );
or \U$2128 ( \2314 , \2309 , \2312 , \2313 );
and \U$2129 ( \2315 , \2277 , \2314 );
xor \U$2130 ( \2316 , \2087 , \2091 );
xor \U$2131 ( \2317 , \2316 , \2096 );
xor \U$2132 ( \2318 , \2103 , \2107 );
xor \U$2133 ( \2319 , \2318 , \2112 );
and \U$2134 ( \2320 , \2317 , \2319 );
xor \U$2135 ( \2321 , \2167 , \2171 );
xor \U$2136 ( \2322 , \2321 , \2176 );
and \U$2137 ( \2323 , \2319 , \2322 );
and \U$2138 ( \2324 , \2317 , \2322 );
or \U$2139 ( \2325 , \2320 , \2323 , \2324 );
and \U$2140 ( \2326 , \2314 , \2325 );
and \U$2141 ( \2327 , \2277 , \2325 );
or \U$2142 ( \2328 , \2315 , \2326 , \2327 );
xor \U$2143 ( \2329 , \1955 , \1959 );
xor \U$2144 ( \2330 , \2329 , \1964 );
xor \U$2145 ( \2331 , \2139 , \2141 );
xor \U$2146 ( \2332 , \2331 , \2144 );
and \U$2147 ( \2333 , \2330 , \2332 );
xor \U$2148 ( \2334 , \2163 , \2179 );
xor \U$2149 ( \2335 , \2334 , \2181 );
and \U$2150 ( \2336 , \2332 , \2335 );
and \U$2151 ( \2337 , \2330 , \2335 );
or \U$2152 ( \2338 , \2333 , \2336 , \2337 );
and \U$2153 ( \2339 , \2328 , \2338 );
xor \U$2154 ( \2340 , \2019 , \2029 );
xor \U$2155 ( \2341 , \2340 , \2034 );
and \U$2156 ( \2342 , \2338 , \2341 );
and \U$2157 ( \2343 , \2328 , \2341 );
or \U$2158 ( \2344 , \2339 , \2342 , \2343 );
xor \U$2159 ( \2345 , \1967 , \1983 );
xor \U$2160 ( \2346 , \2345 , \2000 );
xor \U$2161 ( \2347 , \2137 , \2147 );
xor \U$2162 ( \2348 , \2347 , \2184 );
and \U$2163 ( \2349 , \2346 , \2348 );
xor \U$2164 ( \2350 , \2189 , \2191 );
xor \U$2165 ( \2351 , \2350 , \2194 );
and \U$2166 ( \2352 , \2348 , \2351 );
and \U$2167 ( \2353 , \2346 , \2351 );
or \U$2168 ( \2354 , \2349 , \2352 , \2353 );
and \U$2169 ( \2355 , \2344 , \2354 );
xor \U$2170 ( \2356 , \2003 , \2037 );
xor \U$2171 ( \2357 , \2356 , \2047 );
and \U$2172 ( \2358 , \2354 , \2357 );
and \U$2173 ( \2359 , \2344 , \2357 );
or \U$2174 ( \2360 , \2355 , \2358 , \2359 );
xor \U$2175 ( \2361 , \2203 , \2205 );
xor \U$2176 ( \2362 , \2361 , \2207 );
and \U$2177 ( \2363 , \2360 , \2362 );
and \U$2178 ( \2364 , \2222 , \2363 );
xor \U$2179 ( \2365 , \2222 , \2363 );
xor \U$2180 ( \2366 , \2360 , \2362 );
buf \U$2181 ( \2367 , RIa166c70_30);
buf \U$2182 ( \2368 , RIb4ca4d8_31);
and \U$2183 ( \2369 , \2367 , \2368 );
not \U$2184 ( \2370 , \2369 );
and \U$2185 ( \2371 , \2118 , \2370 );
not \U$2186 ( \2372 , \2371 );
and \U$2187 ( \2373 , \313 , \2259 );
and \U$2188 ( \2374 , \289 , \2257 );
nor \U$2189 ( \2375 , \2373 , \2374 );
xnor \U$2190 ( \2376 , \2375 , \2121 );
and \U$2191 ( \2377 , \2372 , \2376 );
and \U$2192 ( \2378 , \331 , \1952 );
and \U$2193 ( \2379 , \304 , \1950 );
nor \U$2194 ( \2380 , \2378 , \2379 );
xnor \U$2195 ( \2381 , \2380 , \1832 );
and \U$2196 ( \2382 , \2376 , \2381 );
and \U$2197 ( \2383 , \2372 , \2381 );
or \U$2198 ( \2384 , \2377 , \2382 , \2383 );
and \U$2199 ( \2385 , \351 , \1739 );
and \U$2200 ( \2386 , \322 , \1737 );
nor \U$2201 ( \2387 , \2385 , \2386 );
xnor \U$2202 ( \2388 , \2387 , \1607 );
and \U$2203 ( \2389 , \359 , \1474 );
and \U$2204 ( \2390 , \342 , \1472 );
nor \U$2205 ( \2391 , \2389 , \2390 );
xnor \U$2206 ( \2392 , \2391 , \1360 );
and \U$2207 ( \2393 , \2388 , \2392 );
and \U$2208 ( \2394 , \494 , \1277 );
and \U$2209 ( \2395 , \444 , \1275 );
nor \U$2210 ( \2396 , \2394 , \2395 );
xnor \U$2211 ( \2397 , \2396 , \1173 );
and \U$2212 ( \2398 , \2392 , \2397 );
and \U$2213 ( \2399 , \2388 , \2397 );
or \U$2214 ( \2400 , \2393 , \2398 , \2399 );
and \U$2215 ( \2401 , \2384 , \2400 );
and \U$2216 ( \2402 , \620 , \1059 );
and \U$2217 ( \2403 , \591 , \1057 );
nor \U$2218 ( \2404 , \2402 , \2403 );
xnor \U$2219 ( \2405 , \2404 , \981 );
and \U$2220 ( \2406 , \776 , \911 );
and \U$2221 ( \2407 , \701 , \909 );
nor \U$2222 ( \2408 , \2406 , \2407 );
xnor \U$2223 ( \2409 , \2408 , \815 );
and \U$2224 ( \2410 , \2405 , \2409 );
and \U$2225 ( \2411 , \903 , \738 );
and \U$2226 ( \2412 , \839 , \736 );
nor \U$2227 ( \2413 , \2411 , \2412 );
xnor \U$2228 ( \2414 , \2413 , \665 );
and \U$2229 ( \2415 , \2409 , \2414 );
and \U$2230 ( \2416 , \2405 , \2414 );
or \U$2231 ( \2417 , \2410 , \2415 , \2416 );
and \U$2232 ( \2418 , \2400 , \2417 );
and \U$2233 ( \2419 , \2384 , \2417 );
or \U$2234 ( \2420 , \2401 , \2418 , \2419 );
xor \U$2235 ( \2421 , \2226 , \2230 );
xor \U$2236 ( \2422 , \2421 , \2235 );
xor \U$2237 ( \2423 , \2281 , \2285 );
xor \U$2238 ( \2424 , \2423 , \2290 );
and \U$2239 ( \2425 , \2422 , \2424 );
xor \U$2240 ( \2426 , \2297 , \2301 );
xor \U$2241 ( \2427 , \2426 , \2305 );
and \U$2242 ( \2428 , \2424 , \2427 );
and \U$2243 ( \2429 , \2422 , \2427 );
or \U$2244 ( \2430 , \2425 , \2428 , \2429 );
and \U$2245 ( \2431 , \2420 , \2430 );
and \U$2246 ( \2432 , \1777 , \310 );
and \U$2247 ( \2433 , \1768 , \308 );
nor \U$2248 ( \2434 , \2432 , \2433 );
xnor \U$2249 ( \2435 , \2434 , \318 );
and \U$2250 ( \2436 , \2027 , \328 );
and \U$2251 ( \2437 , \2021 , \326 );
nor \U$2252 ( \2438 , \2436 , \2437 );
xnor \U$2253 ( \2439 , \2438 , \336 );
and \U$2254 ( \2440 , \2435 , \2439 );
and \U$2255 ( \2441 , \2304 , \348 );
and \U$2256 ( \2442 , \2159 , \346 );
nor \U$2257 ( \2443 , \2441 , \2442 );
xnor \U$2258 ( \2444 , \2443 , \356 );
and \U$2259 ( \2445 , \2439 , \2444 );
and \U$2260 ( \2446 , \2435 , \2444 );
or \U$2261 ( \2447 , \2440 , \2445 , \2446 );
and \U$2262 ( \2448 , \1191 , \602 );
and \U$2263 ( \2449 , \1102 , \600 );
nor \U$2264 ( \2450 , \2448 , \2449 );
xnor \U$2265 ( \2451 , \2450 , \558 );
and \U$2266 ( \2452 , \1303 , \502 );
and \U$2267 ( \2453 , \1297 , \500 );
nor \U$2268 ( \2454 , \2452 , \2453 );
xnor \U$2269 ( \2455 , \2454 , \453 );
and \U$2270 ( \2456 , \2451 , \2455 );
and \U$2271 ( \2457 , \1536 , \296 );
and \U$2272 ( \2458 , \1420 , \294 );
nor \U$2273 ( \2459 , \2457 , \2458 );
xnor \U$2274 ( \2460 , \2459 , \301 );
and \U$2275 ( \2461 , \2455 , \2460 );
and \U$2276 ( \2462 , \2451 , \2460 );
or \U$2277 ( \2463 , \2456 , \2461 , \2462 );
or \U$2278 ( \2464 , \2447 , \2463 );
and \U$2279 ( \2465 , \2430 , \2464 );
and \U$2280 ( \2466 , \2420 , \2464 );
or \U$2281 ( \2467 , \2431 , \2465 , \2466 );
xor \U$2282 ( \2468 , \2122 , \2126 );
xor \U$2283 ( \2469 , \2468 , \2131 );
xor \U$2284 ( \2470 , \2293 , \2308 );
xor \U$2285 ( \2471 , \2470 , \2311 );
and \U$2286 ( \2472 , \2469 , \2471 );
xor \U$2287 ( \2473 , \2317 , \2319 );
xor \U$2288 ( \2474 , \2473 , \2322 );
and \U$2289 ( \2475 , \2471 , \2474 );
and \U$2290 ( \2476 , \2469 , \2474 );
or \U$2291 ( \2477 , \2472 , \2475 , \2476 );
and \U$2292 ( \2478 , \2467 , \2477 );
xor \U$2293 ( \2479 , \2099 , \2115 );
xor \U$2294 ( \2480 , \2479 , \2134 );
and \U$2295 ( \2481 , \2477 , \2480 );
and \U$2296 ( \2482 , \2467 , \2480 );
or \U$2297 ( \2483 , \2478 , \2481 , \2482 );
xor \U$2298 ( \2484 , \2328 , \2338 );
xor \U$2299 ( \2485 , \2484 , \2341 );
and \U$2300 ( \2486 , \2483 , \2485 );
xor \U$2301 ( \2487 , \2346 , \2348 );
xor \U$2302 ( \2488 , \2487 , \2351 );
and \U$2303 ( \2489 , \2485 , \2488 );
and \U$2304 ( \2490 , \2483 , \2488 );
or \U$2305 ( \2491 , \2486 , \2489 , \2490 );
xor \U$2306 ( \2492 , \2344 , \2354 );
xor \U$2307 ( \2493 , \2492 , \2357 );
and \U$2308 ( \2494 , \2491 , \2493 );
xor \U$2309 ( \2495 , \2187 , \2197 );
xor \U$2310 ( \2496 , \2495 , \2200 );
and \U$2311 ( \2497 , \2493 , \2496 );
and \U$2312 ( \2498 , \2491 , \2496 );
or \U$2313 ( \2499 , \2494 , \2497 , \2498 );
and \U$2314 ( \2500 , \2366 , \2499 );
xor \U$2315 ( \2501 , \2366 , \2499 );
xor \U$2316 ( \2502 , \2491 , \2493 );
xor \U$2317 ( \2503 , \2502 , \2496 );
and \U$2318 ( \2504 , \1297 , \602 );
and \U$2319 ( \2505 , \1191 , \600 );
nor \U$2320 ( \2506 , \2504 , \2505 );
xnor \U$2321 ( \2507 , \2506 , \558 );
and \U$2322 ( \2508 , \1420 , \502 );
and \U$2323 ( \2509 , \1303 , \500 );
nor \U$2324 ( \2510 , \2508 , \2509 );
xnor \U$2325 ( \2511 , \2510 , \453 );
and \U$2326 ( \2512 , \2507 , \2511 );
and \U$2327 ( \2513 , \1768 , \296 );
and \U$2328 ( \2514 , \1536 , \294 );
nor \U$2329 ( \2515 , \2513 , \2514 );
xnor \U$2330 ( \2516 , \2515 , \301 );
and \U$2331 ( \2517 , \2511 , \2516 );
and \U$2332 ( \2518 , \2507 , \2516 );
or \U$2333 ( \2519 , \2512 , \2517 , \2518 );
and \U$2334 ( \2520 , \2021 , \310 );
and \U$2335 ( \2521 , \1777 , \308 );
nor \U$2336 ( \2522 , \2520 , \2521 );
xnor \U$2337 ( \2523 , \2522 , \318 );
and \U$2338 ( \2524 , \2159 , \328 );
and \U$2339 ( \2525 , \2027 , \326 );
nor \U$2340 ( \2526 , \2524 , \2525 );
xnor \U$2341 ( \2527 , \2526 , \336 );
and \U$2342 ( \2528 , \2523 , \2527 );
_DC g127 ( \2529_nG127 , RIb4c2be8_61 , \287 );
buf \U$2343 ( \2530 , \2529_nG127 );
and \U$2344 ( \2531 , \2530 , \348 );
and \U$2345 ( \2532 , \2304 , \346 );
nor \U$2346 ( \2533 , \2531 , \2532 );
xnor \U$2347 ( \2534 , \2533 , \356 );
and \U$2348 ( \2535 , \2527 , \2534 );
and \U$2349 ( \2536 , \2523 , \2534 );
or \U$2350 ( \2537 , \2528 , \2535 , \2536 );
and \U$2351 ( \2538 , \2519 , \2537 );
_DC g126 ( \2539_nG126 , RIb4c2b70_62 , \287 );
buf \U$2352 ( \2540 , \2539_nG126 );
and \U$2353 ( \2541 , \2540 , \343 );
buf \U$2354 ( \2542 , \2541 );
and \U$2355 ( \2543 , \2537 , \2542 );
and \U$2356 ( \2544 , \2519 , \2542 );
or \U$2357 ( \2545 , \2538 , \2543 , \2544 );
xor \U$2358 ( \2546 , \2118 , \2367 );
xor \U$2359 ( \2547 , \2367 , \2368 );
not \U$2360 ( \2548 , \2547 );
and \U$2361 ( \2549 , \2546 , \2548 );
and \U$2362 ( \2550 , \289 , \2549 );
not \U$2363 ( \2551 , \2550 );
xnor \U$2364 ( \2552 , \2551 , \2371 );
and \U$2365 ( \2553 , \304 , \2259 );
and \U$2366 ( \2554 , \313 , \2257 );
nor \U$2367 ( \2555 , \2553 , \2554 );
xnor \U$2368 ( \2556 , \2555 , \2121 );
and \U$2369 ( \2557 , \2552 , \2556 );
and \U$2370 ( \2558 , \322 , \1952 );
and \U$2371 ( \2559 , \331 , \1950 );
nor \U$2372 ( \2560 , \2558 , \2559 );
xnor \U$2373 ( \2561 , \2560 , \1832 );
and \U$2374 ( \2562 , \2556 , \2561 );
and \U$2375 ( \2563 , \2552 , \2561 );
or \U$2376 ( \2564 , \2557 , \2562 , \2563 );
and \U$2377 ( \2565 , \342 , \1739 );
and \U$2378 ( \2566 , \351 , \1737 );
nor \U$2379 ( \2567 , \2565 , \2566 );
xnor \U$2380 ( \2568 , \2567 , \1607 );
and \U$2381 ( \2569 , \444 , \1474 );
and \U$2382 ( \2570 , \359 , \1472 );
nor \U$2383 ( \2571 , \2569 , \2570 );
xnor \U$2384 ( \2572 , \2571 , \1360 );
and \U$2385 ( \2573 , \2568 , \2572 );
and \U$2386 ( \2574 , \591 , \1277 );
and \U$2387 ( \2575 , \494 , \1275 );
nor \U$2388 ( \2576 , \2574 , \2575 );
xnor \U$2389 ( \2577 , \2576 , \1173 );
and \U$2390 ( \2578 , \2572 , \2577 );
and \U$2391 ( \2579 , \2568 , \2577 );
or \U$2392 ( \2580 , \2573 , \2578 , \2579 );
and \U$2393 ( \2581 , \2564 , \2580 );
and \U$2394 ( \2582 , \701 , \1059 );
and \U$2395 ( \2583 , \620 , \1057 );
nor \U$2396 ( \2584 , \2582 , \2583 );
xnor \U$2397 ( \2585 , \2584 , \981 );
and \U$2398 ( \2586 , \839 , \911 );
and \U$2399 ( \2587 , \776 , \909 );
nor \U$2400 ( \2588 , \2586 , \2587 );
xnor \U$2401 ( \2589 , \2588 , \815 );
and \U$2402 ( \2590 , \2585 , \2589 );
and \U$2403 ( \2591 , \1102 , \738 );
and \U$2404 ( \2592 , \903 , \736 );
nor \U$2405 ( \2593 , \2591 , \2592 );
xnor \U$2406 ( \2594 , \2593 , \665 );
and \U$2407 ( \2595 , \2589 , \2594 );
and \U$2408 ( \2596 , \2585 , \2594 );
or \U$2409 ( \2597 , \2590 , \2595 , \2596 );
and \U$2410 ( \2598 , \2580 , \2597 );
and \U$2411 ( \2599 , \2564 , \2597 );
or \U$2412 ( \2600 , \2581 , \2598 , \2599 );
and \U$2413 ( \2601 , \2545 , \2600 );
and \U$2414 ( \2602 , \2530 , \343 );
xor \U$2415 ( \2603 , \2435 , \2439 );
xor \U$2416 ( \2604 , \2603 , \2444 );
and \U$2417 ( \2605 , \2602 , \2604 );
xor \U$2418 ( \2606 , \2451 , \2455 );
xor \U$2419 ( \2607 , \2606 , \2460 );
and \U$2420 ( \2608 , \2604 , \2607 );
and \U$2421 ( \2609 , \2602 , \2607 );
or \U$2422 ( \2610 , \2605 , \2608 , \2609 );
and \U$2423 ( \2611 , \2600 , \2610 );
and \U$2424 ( \2612 , \2545 , \2610 );
or \U$2425 ( \2613 , \2601 , \2611 , \2612 );
xor \U$2426 ( \2614 , \2372 , \2376 );
xor \U$2427 ( \2615 , \2614 , \2381 );
xor \U$2428 ( \2616 , \2388 , \2392 );
xor \U$2429 ( \2617 , \2616 , \2397 );
and \U$2430 ( \2618 , \2615 , \2617 );
xor \U$2431 ( \2619 , \2405 , \2409 );
xor \U$2432 ( \2620 , \2619 , \2414 );
and \U$2433 ( \2621 , \2617 , \2620 );
and \U$2434 ( \2622 , \2615 , \2620 );
or \U$2435 ( \2623 , \2618 , \2621 , \2622 );
xor \U$2436 ( \2624 , \2242 , \2246 );
xor \U$2437 ( \2625 , \2624 , \2251 );
and \U$2438 ( \2626 , \2623 , \2625 );
xor \U$2439 ( \2627 , \2262 , \2266 );
xor \U$2440 ( \2628 , \2627 , \2271 );
and \U$2441 ( \2629 , \2625 , \2628 );
and \U$2442 ( \2630 , \2623 , \2628 );
or \U$2443 ( \2631 , \2626 , \2629 , \2630 );
and \U$2444 ( \2632 , \2613 , \2631 );
xor \U$2445 ( \2633 , \2384 , \2400 );
xor \U$2446 ( \2634 , \2633 , \2417 );
xor \U$2447 ( \2635 , \2422 , \2424 );
xor \U$2448 ( \2636 , \2635 , \2427 );
and \U$2449 ( \2637 , \2634 , \2636 );
xnor \U$2450 ( \2638 , \2447 , \2463 );
and \U$2451 ( \2639 , \2636 , \2638 );
and \U$2452 ( \2640 , \2634 , \2638 );
or \U$2453 ( \2641 , \2637 , \2639 , \2640 );
and \U$2454 ( \2642 , \2631 , \2641 );
and \U$2455 ( \2643 , \2613 , \2641 );
or \U$2456 ( \2644 , \2632 , \2642 , \2643 );
xor \U$2457 ( \2645 , \2238 , \2254 );
xor \U$2458 ( \2646 , \2645 , \2274 );
xor \U$2459 ( \2647 , \2420 , \2430 );
xor \U$2460 ( \2648 , \2647 , \2464 );
and \U$2461 ( \2649 , \2646 , \2648 );
xor \U$2462 ( \2650 , \2469 , \2471 );
xor \U$2463 ( \2651 , \2650 , \2474 );
and \U$2464 ( \2652 , \2648 , \2651 );
and \U$2465 ( \2653 , \2646 , \2651 );
or \U$2466 ( \2654 , \2649 , \2652 , \2653 );
and \U$2467 ( \2655 , \2644 , \2654 );
xor \U$2468 ( \2656 , \2330 , \2332 );
xor \U$2469 ( \2657 , \2656 , \2335 );
and \U$2470 ( \2658 , \2654 , \2657 );
and \U$2471 ( \2659 , \2644 , \2657 );
or \U$2472 ( \2660 , \2655 , \2658 , \2659 );
xor \U$2473 ( \2661 , \2277 , \2314 );
xor \U$2474 ( \2662 , \2661 , \2325 );
xor \U$2475 ( \2663 , \2467 , \2477 );
xor \U$2476 ( \2664 , \2663 , \2480 );
and \U$2477 ( \2665 , \2662 , \2664 );
and \U$2478 ( \2666 , \2660 , \2665 );
xor \U$2479 ( \2667 , \2483 , \2485 );
xor \U$2480 ( \2668 , \2667 , \2488 );
and \U$2481 ( \2669 , \2665 , \2668 );
and \U$2482 ( \2670 , \2660 , \2668 );
or \U$2483 ( \2671 , \2666 , \2669 , \2670 );
and \U$2484 ( \2672 , \2503 , \2671 );
xor \U$2485 ( \2673 , \2503 , \2671 );
xor \U$2486 ( \2674 , \2660 , \2665 );
xor \U$2487 ( \2675 , \2674 , \2668 );
and \U$2488 ( \2676 , \620 , \1277 );
and \U$2489 ( \2677 , \591 , \1275 );
nor \U$2490 ( \2678 , \2676 , \2677 );
xnor \U$2491 ( \2679 , \2678 , \1173 );
and \U$2492 ( \2680 , \776 , \1059 );
and \U$2493 ( \2681 , \701 , \1057 );
nor \U$2494 ( \2682 , \2680 , \2681 );
xnor \U$2495 ( \2683 , \2682 , \981 );
and \U$2496 ( \2684 , \2679 , \2683 );
and \U$2497 ( \2685 , \903 , \911 );
and \U$2498 ( \2686 , \839 , \909 );
nor \U$2499 ( \2687 , \2685 , \2686 );
xnor \U$2500 ( \2688 , \2687 , \815 );
and \U$2501 ( \2689 , \2683 , \2688 );
and \U$2502 ( \2690 , \2679 , \2688 );
or \U$2503 ( \2691 , \2684 , \2689 , \2690 );
not \U$2504 ( \2692 , \2368 );
and \U$2505 ( \2693 , \313 , \2549 );
and \U$2506 ( \2694 , \289 , \2547 );
nor \U$2507 ( \2695 , \2693 , \2694 );
xnor \U$2508 ( \2696 , \2695 , \2371 );
and \U$2509 ( \2697 , \2692 , \2696 );
and \U$2510 ( \2698 , \331 , \2259 );
and \U$2511 ( \2699 , \304 , \2257 );
nor \U$2512 ( \2700 , \2698 , \2699 );
xnor \U$2513 ( \2701 , \2700 , \2121 );
and \U$2514 ( \2702 , \2696 , \2701 );
and \U$2515 ( \2703 , \2692 , \2701 );
or \U$2516 ( \2704 , \2697 , \2702 , \2703 );
and \U$2517 ( \2705 , \2691 , \2704 );
and \U$2518 ( \2706 , \351 , \1952 );
and \U$2519 ( \2707 , \322 , \1950 );
nor \U$2520 ( \2708 , \2706 , \2707 );
xnor \U$2521 ( \2709 , \2708 , \1832 );
and \U$2522 ( \2710 , \359 , \1739 );
and \U$2523 ( \2711 , \342 , \1737 );
nor \U$2524 ( \2712 , \2710 , \2711 );
xnor \U$2525 ( \2713 , \2712 , \1607 );
and \U$2526 ( \2714 , \2709 , \2713 );
and \U$2527 ( \2715 , \494 , \1474 );
and \U$2528 ( \2716 , \444 , \1472 );
nor \U$2529 ( \2717 , \2715 , \2716 );
xnor \U$2530 ( \2718 , \2717 , \1360 );
and \U$2531 ( \2719 , \2713 , \2718 );
and \U$2532 ( \2720 , \2709 , \2718 );
or \U$2533 ( \2721 , \2714 , \2719 , \2720 );
and \U$2534 ( \2722 , \2704 , \2721 );
and \U$2535 ( \2723 , \2691 , \2721 );
or \U$2536 ( \2724 , \2705 , \2722 , \2723 );
and \U$2537 ( \2725 , \1777 , \296 );
and \U$2538 ( \2726 , \1768 , \294 );
nor \U$2539 ( \2727 , \2725 , \2726 );
xnor \U$2540 ( \2728 , \2727 , \301 );
and \U$2541 ( \2729 , \2027 , \310 );
and \U$2542 ( \2730 , \2021 , \308 );
nor \U$2543 ( \2731 , \2729 , \2730 );
xnor \U$2544 ( \2732 , \2731 , \318 );
and \U$2545 ( \2733 , \2728 , \2732 );
and \U$2546 ( \2734 , \2304 , \328 );
and \U$2547 ( \2735 , \2159 , \326 );
nor \U$2548 ( \2736 , \2734 , \2735 );
xnor \U$2549 ( \2737 , \2736 , \336 );
and \U$2550 ( \2738 , \2732 , \2737 );
and \U$2551 ( \2739 , \2728 , \2737 );
or \U$2552 ( \2740 , \2733 , \2738 , \2739 );
and \U$2553 ( \2741 , \1191 , \738 );
and \U$2554 ( \2742 , \1102 , \736 );
nor \U$2555 ( \2743 , \2741 , \2742 );
xnor \U$2556 ( \2744 , \2743 , \665 );
and \U$2557 ( \2745 , \1303 , \602 );
and \U$2558 ( \2746 , \1297 , \600 );
nor \U$2559 ( \2747 , \2745 , \2746 );
xnor \U$2560 ( \2748 , \2747 , \558 );
and \U$2561 ( \2749 , \2744 , \2748 );
and \U$2562 ( \2750 , \1536 , \502 );
and \U$2563 ( \2751 , \1420 , \500 );
nor \U$2564 ( \2752 , \2750 , \2751 );
xnor \U$2565 ( \2753 , \2752 , \453 );
and \U$2566 ( \2754 , \2748 , \2753 );
and \U$2567 ( \2755 , \2744 , \2753 );
or \U$2568 ( \2756 , \2749 , \2754 , \2755 );
and \U$2569 ( \2757 , \2740 , \2756 );
and \U$2570 ( \2758 , \2540 , \348 );
and \U$2571 ( \2759 , \2530 , \346 );
nor \U$2572 ( \2760 , \2758 , \2759 );
xnor \U$2573 ( \2761 , \2760 , \356 );
_DC g125 ( \2762_nG125 , RIb4c2af8_63 , \287 );
buf \U$2574 ( \2763 , \2762_nG125 );
and \U$2575 ( \2764 , \2763 , \343 );
or \U$2576 ( \2765 , \2761 , \2764 );
and \U$2577 ( \2766 , \2756 , \2765 );
and \U$2578 ( \2767 , \2740 , \2765 );
or \U$2579 ( \2768 , \2757 , \2766 , \2767 );
and \U$2580 ( \2769 , \2724 , \2768 );
xor \U$2581 ( \2770 , \2507 , \2511 );
xor \U$2582 ( \2771 , \2770 , \2516 );
xor \U$2583 ( \2772 , \2523 , \2527 );
xor \U$2584 ( \2773 , \2772 , \2534 );
and \U$2585 ( \2774 , \2771 , \2773 );
not \U$2586 ( \2775 , \2541 );
and \U$2587 ( \2776 , \2773 , \2775 );
and \U$2588 ( \2777 , \2771 , \2775 );
or \U$2589 ( \2778 , \2774 , \2776 , \2777 );
and \U$2590 ( \2779 , \2768 , \2778 );
and \U$2591 ( \2780 , \2724 , \2778 );
or \U$2592 ( \2781 , \2769 , \2779 , \2780 );
xor \U$2593 ( \2782 , \2552 , \2556 );
xor \U$2594 ( \2783 , \2782 , \2561 );
xor \U$2595 ( \2784 , \2568 , \2572 );
xor \U$2596 ( \2785 , \2784 , \2577 );
and \U$2597 ( \2786 , \2783 , \2785 );
xor \U$2598 ( \2787 , \2585 , \2589 );
xor \U$2599 ( \2788 , \2787 , \2594 );
and \U$2600 ( \2789 , \2785 , \2788 );
and \U$2601 ( \2790 , \2783 , \2788 );
or \U$2602 ( \2791 , \2786 , \2789 , \2790 );
xor \U$2603 ( \2792 , \2602 , \2604 );
xor \U$2604 ( \2793 , \2792 , \2607 );
and \U$2605 ( \2794 , \2791 , \2793 );
xor \U$2606 ( \2795 , \2615 , \2617 );
xor \U$2607 ( \2796 , \2795 , \2620 );
and \U$2608 ( \2797 , \2793 , \2796 );
and \U$2609 ( \2798 , \2791 , \2796 );
or \U$2610 ( \2799 , \2794 , \2797 , \2798 );
and \U$2611 ( \2800 , \2781 , \2799 );
xor \U$2612 ( \2801 , \2634 , \2636 );
xor \U$2613 ( \2802 , \2801 , \2638 );
and \U$2614 ( \2803 , \2799 , \2802 );
and \U$2615 ( \2804 , \2781 , \2802 );
or \U$2616 ( \2805 , \2800 , \2803 , \2804 );
xor \U$2617 ( \2806 , \2613 , \2631 );
xor \U$2618 ( \2807 , \2806 , \2641 );
and \U$2619 ( \2808 , \2805 , \2807 );
xor \U$2620 ( \2809 , \2646 , \2648 );
xor \U$2621 ( \2810 , \2809 , \2651 );
and \U$2622 ( \2811 , \2807 , \2810 );
and \U$2623 ( \2812 , \2805 , \2810 );
or \U$2624 ( \2813 , \2808 , \2811 , \2812 );
xor \U$2625 ( \2814 , \2644 , \2654 );
xor \U$2626 ( \2815 , \2814 , \2657 );
and \U$2627 ( \2816 , \2813 , \2815 );
xor \U$2628 ( \2817 , \2662 , \2664 );
and \U$2629 ( \2818 , \2815 , \2817 );
and \U$2630 ( \2819 , \2813 , \2817 );
or \U$2631 ( \2820 , \2816 , \2818 , \2819 );
and \U$2632 ( \2821 , \2675 , \2820 );
xor \U$2633 ( \2822 , \2675 , \2820 );
xor \U$2634 ( \2823 , \2813 , \2815 );
xor \U$2635 ( \2824 , \2823 , \2817 );
and \U$2636 ( \2825 , \1768 , \502 );
and \U$2637 ( \2826 , \1536 , \500 );
nor \U$2638 ( \2827 , \2825 , \2826 );
xnor \U$2639 ( \2828 , \2827 , \453 );
and \U$2640 ( \2829 , \2021 , \296 );
and \U$2641 ( \2830 , \1777 , \294 );
nor \U$2642 ( \2831 , \2829 , \2830 );
xnor \U$2643 ( \2832 , \2831 , \301 );
and \U$2644 ( \2833 , \2828 , \2832 );
and \U$2645 ( \2834 , \2159 , \310 );
and \U$2646 ( \2835 , \2027 , \308 );
nor \U$2647 ( \2836 , \2834 , \2835 );
xnor \U$2648 ( \2837 , \2836 , \318 );
and \U$2649 ( \2838 , \2832 , \2837 );
and \U$2650 ( \2839 , \2828 , \2837 );
or \U$2651 ( \2840 , \2833 , \2838 , \2839 );
and \U$2652 ( \2841 , \2530 , \328 );
and \U$2653 ( \2842 , \2304 , \326 );
nor \U$2654 ( \2843 , \2841 , \2842 );
xnor \U$2655 ( \2844 , \2843 , \336 );
and \U$2656 ( \2845 , \2763 , \348 );
and \U$2657 ( \2846 , \2540 , \346 );
nor \U$2658 ( \2847 , \2845 , \2846 );
xnor \U$2659 ( \2848 , \2847 , \356 );
and \U$2660 ( \2849 , \2844 , \2848 );
_HMUX g124_GF_PartitionCandidate ( \2850_nG124 , RIb4bfab0_64 , 1'b1 , \287 );
buf \U$2662 ( \2851 , \2850_nG124 );
nand \U$2663 ( \2852 , \2851 , \343 );
not \U$2664 ( \2853 , \2852 );
and \U$2665 ( \2854 , \2848 , \2853 );
and \U$2666 ( \2855 , \2844 , \2853 );
or \U$2667 ( \2856 , \2849 , \2854 , \2855 );
and \U$2668 ( \2857 , \2840 , \2856 );
and \U$2669 ( \2858 , \1102 , \911 );
and \U$2670 ( \2859 , \903 , \909 );
nor \U$2671 ( \2860 , \2858 , \2859 );
xnor \U$2672 ( \2861 , \2860 , \815 );
and \U$2673 ( \2862 , \1297 , \738 );
and \U$2674 ( \2863 , \1191 , \736 );
nor \U$2675 ( \2864 , \2862 , \2863 );
xnor \U$2676 ( \2865 , \2864 , \665 );
and \U$2677 ( \2866 , \2861 , \2865 );
and \U$2678 ( \2867 , \1420 , \602 );
and \U$2679 ( \2868 , \1303 , \600 );
nor \U$2680 ( \2869 , \2867 , \2868 );
xnor \U$2681 ( \2870 , \2869 , \558 );
and \U$2682 ( \2871 , \2865 , \2870 );
and \U$2683 ( \2872 , \2861 , \2870 );
or \U$2684 ( \2873 , \2866 , \2871 , \2872 );
and \U$2685 ( \2874 , \2856 , \2873 );
and \U$2686 ( \2875 , \2840 , \2873 );
or \U$2687 ( \2876 , \2857 , \2874 , \2875 );
and \U$2688 ( \2877 , \591 , \1474 );
and \U$2689 ( \2878 , \494 , \1472 );
nor \U$2690 ( \2879 , \2877 , \2878 );
xnor \U$2691 ( \2880 , \2879 , \1360 );
and \U$2692 ( \2881 , \701 , \1277 );
and \U$2693 ( \2882 , \620 , \1275 );
nor \U$2694 ( \2883 , \2881 , \2882 );
xnor \U$2695 ( \2884 , \2883 , \1173 );
and \U$2696 ( \2885 , \2880 , \2884 );
and \U$2697 ( \2886 , \839 , \1059 );
and \U$2698 ( \2887 , \776 , \1057 );
nor \U$2699 ( \2888 , \2886 , \2887 );
xnor \U$2700 ( \2889 , \2888 , \981 );
and \U$2701 ( \2890 , \2884 , \2889 );
and \U$2702 ( \2891 , \2880 , \2889 );
or \U$2703 ( \2892 , \2885 , \2890 , \2891 );
and \U$2704 ( \2893 , \322 , \2259 );
and \U$2705 ( \2894 , \331 , \2257 );
nor \U$2706 ( \2895 , \2893 , \2894 );
xnor \U$2707 ( \2896 , \2895 , \2121 );
and \U$2708 ( \2897 , \342 , \1952 );
and \U$2709 ( \2898 , \351 , \1950 );
nor \U$2710 ( \2899 , \2897 , \2898 );
xnor \U$2711 ( \2900 , \2899 , \1832 );
and \U$2712 ( \2901 , \2896 , \2900 );
and \U$2713 ( \2902 , \444 , \1739 );
and \U$2714 ( \2903 , \359 , \1737 );
nor \U$2715 ( \2904 , \2902 , \2903 );
xnor \U$2716 ( \2905 , \2904 , \1607 );
and \U$2717 ( \2906 , \2900 , \2905 );
and \U$2718 ( \2907 , \2896 , \2905 );
or \U$2719 ( \2908 , \2901 , \2906 , \2907 );
and \U$2720 ( \2909 , \2892 , \2908 );
buf \U$2721 ( \2910 , RIb4ca460_32);
xor \U$2722 ( \2911 , \2368 , \2910 );
not \U$2723 ( \2912 , \2910 );
and \U$2724 ( \2913 , \2911 , \2912 );
and \U$2725 ( \2914 , \289 , \2913 );
not \U$2726 ( \2915 , \2914 );
xnor \U$2727 ( \2916 , \2915 , \2368 );
and \U$2728 ( \2917 , \304 , \2549 );
and \U$2729 ( \2918 , \313 , \2547 );
nor \U$2730 ( \2919 , \2917 , \2918 );
xnor \U$2731 ( \2920 , \2919 , \2371 );
and \U$2732 ( \2921 , \2916 , \2920 );
and \U$2733 ( \2922 , \2908 , \2921 );
and \U$2734 ( \2923 , \2892 , \2921 );
or \U$2735 ( \2924 , \2909 , \2922 , \2923 );
and \U$2736 ( \2925 , \2876 , \2924 );
xor \U$2737 ( \2926 , \2728 , \2732 );
xor \U$2738 ( \2927 , \2926 , \2737 );
xor \U$2739 ( \2928 , \2744 , \2748 );
xor \U$2740 ( \2929 , \2928 , \2753 );
and \U$2741 ( \2930 , \2927 , \2929 );
xnor \U$2742 ( \2931 , \2761 , \2764 );
and \U$2743 ( \2932 , \2929 , \2931 );
and \U$2744 ( \2933 , \2927 , \2931 );
or \U$2745 ( \2934 , \2930 , \2932 , \2933 );
and \U$2746 ( \2935 , \2924 , \2934 );
and \U$2747 ( \2936 , \2876 , \2934 );
or \U$2748 ( \2937 , \2925 , \2935 , \2936 );
xor \U$2749 ( \2938 , \2679 , \2683 );
xor \U$2750 ( \2939 , \2938 , \2688 );
xor \U$2751 ( \2940 , \2692 , \2696 );
xor \U$2752 ( \2941 , \2940 , \2701 );
and \U$2753 ( \2942 , \2939 , \2941 );
xor \U$2754 ( \2943 , \2709 , \2713 );
xor \U$2755 ( \2944 , \2943 , \2718 );
and \U$2756 ( \2945 , \2941 , \2944 );
and \U$2757 ( \2946 , \2939 , \2944 );
or \U$2758 ( \2947 , \2942 , \2945 , \2946 );
xor \U$2759 ( \2948 , \2783 , \2785 );
xor \U$2760 ( \2949 , \2948 , \2788 );
and \U$2761 ( \2950 , \2947 , \2949 );
xor \U$2762 ( \2951 , \2771 , \2773 );
xor \U$2763 ( \2952 , \2951 , \2775 );
and \U$2764 ( \2953 , \2949 , \2952 );
and \U$2765 ( \2954 , \2947 , \2952 );
or \U$2766 ( \2955 , \2950 , \2953 , \2954 );
and \U$2767 ( \2956 , \2937 , \2955 );
xor \U$2768 ( \2957 , \2519 , \2537 );
xor \U$2769 ( \2958 , \2957 , \2542 );
and \U$2770 ( \2959 , \2955 , \2958 );
and \U$2771 ( \2960 , \2937 , \2958 );
or \U$2772 ( \2961 , \2956 , \2959 , \2960 );
xor \U$2773 ( \2962 , \2564 , \2580 );
xor \U$2774 ( \2963 , \2962 , \2597 );
xor \U$2775 ( \2964 , \2724 , \2768 );
xor \U$2776 ( \2965 , \2964 , \2778 );
and \U$2777 ( \2966 , \2963 , \2965 );
xor \U$2778 ( \2967 , \2791 , \2793 );
xor \U$2779 ( \2968 , \2967 , \2796 );
and \U$2780 ( \2969 , \2965 , \2968 );
and \U$2781 ( \2970 , \2963 , \2968 );
or \U$2782 ( \2971 , \2966 , \2969 , \2970 );
and \U$2783 ( \2972 , \2961 , \2971 );
xor \U$2784 ( \2973 , \2623 , \2625 );
xor \U$2785 ( \2974 , \2973 , \2628 );
and \U$2786 ( \2975 , \2971 , \2974 );
and \U$2787 ( \2976 , \2961 , \2974 );
or \U$2788 ( \2977 , \2972 , \2975 , \2976 );
xor \U$2789 ( \2978 , \2545 , \2600 );
xor \U$2790 ( \2979 , \2978 , \2610 );
xor \U$2791 ( \2980 , \2781 , \2799 );
xor \U$2792 ( \2981 , \2980 , \2802 );
and \U$2793 ( \2982 , \2979 , \2981 );
and \U$2794 ( \2983 , \2977 , \2982 );
xor \U$2795 ( \2984 , \2805 , \2807 );
xor \U$2796 ( \2985 , \2984 , \2810 );
and \U$2797 ( \2986 , \2982 , \2985 );
and \U$2798 ( \2987 , \2977 , \2985 );
or \U$2799 ( \2988 , \2983 , \2986 , \2987 );
and \U$2800 ( \2989 , \2824 , \2988 );
xor \U$2801 ( \2990 , \2824 , \2988 );
xor \U$2802 ( \2991 , \2977 , \2982 );
xor \U$2803 ( \2992 , \2991 , \2985 );
and \U$2804 ( \2993 , \359 , \1952 );
and \U$2805 ( \2994 , \342 , \1950 );
nor \U$2806 ( \2995 , \2993 , \2994 );
xnor \U$2807 ( \2996 , \2995 , \1832 );
and \U$2808 ( \2997 , \494 , \1739 );
and \U$2809 ( \2998 , \444 , \1737 );
nor \U$2810 ( \2999 , \2997 , \2998 );
xnor \U$2811 ( \3000 , \2999 , \1607 );
and \U$2812 ( \3001 , \2996 , \3000 );
and \U$2813 ( \3002 , \620 , \1474 );
and \U$2814 ( \3003 , \591 , \1472 );
nor \U$2815 ( \3004 , \3002 , \3003 );
xnor \U$2816 ( \3005 , \3004 , \1360 );
and \U$2817 ( \3006 , \3000 , \3005 );
and \U$2818 ( \3007 , \2996 , \3005 );
or \U$2819 ( \3008 , \3001 , \3006 , \3007 );
and \U$2820 ( \3009 , \313 , \2913 );
and \U$2821 ( \3010 , \289 , \2910 );
nor \U$2822 ( \3011 , \3009 , \3010 );
xnor \U$2823 ( \3012 , \3011 , \2368 );
and \U$2824 ( \3013 , \331 , \2549 );
and \U$2825 ( \3014 , \304 , \2547 );
nor \U$2826 ( \3015 , \3013 , \3014 );
xnor \U$2827 ( \3016 , \3015 , \2371 );
and \U$2828 ( \3017 , \3012 , \3016 );
and \U$2829 ( \3018 , \351 , \2259 );
and \U$2830 ( \3019 , \322 , \2257 );
nor \U$2831 ( \3020 , \3018 , \3019 );
xnor \U$2832 ( \3021 , \3020 , \2121 );
and \U$2833 ( \3022 , \3016 , \3021 );
and \U$2834 ( \3023 , \3012 , \3021 );
or \U$2835 ( \3024 , \3017 , \3022 , \3023 );
and \U$2836 ( \3025 , \3008 , \3024 );
and \U$2837 ( \3026 , \776 , \1277 );
and \U$2838 ( \3027 , \701 , \1275 );
nor \U$2839 ( \3028 , \3026 , \3027 );
xnor \U$2840 ( \3029 , \3028 , \1173 );
and \U$2841 ( \3030 , \903 , \1059 );
and \U$2842 ( \3031 , \839 , \1057 );
nor \U$2843 ( \3032 , \3030 , \3031 );
xnor \U$2844 ( \3033 , \3032 , \981 );
and \U$2845 ( \3034 , \3029 , \3033 );
and \U$2846 ( \3035 , \1191 , \911 );
and \U$2847 ( \3036 , \1102 , \909 );
nor \U$2848 ( \3037 , \3035 , \3036 );
xnor \U$2849 ( \3038 , \3037 , \815 );
and \U$2850 ( \3039 , \3033 , \3038 );
and \U$2851 ( \3040 , \3029 , \3038 );
or \U$2852 ( \3041 , \3034 , \3039 , \3040 );
and \U$2853 ( \3042 , \3024 , \3041 );
and \U$2854 ( \3043 , \3008 , \3041 );
or \U$2855 ( \3044 , \3025 , \3042 , \3043 );
xor \U$2856 ( \3045 , \2828 , \2832 );
xor \U$2857 ( \3046 , \3045 , \2837 );
xor \U$2858 ( \3047 , \2880 , \2884 );
xor \U$2859 ( \3048 , \3047 , \2889 );
and \U$2860 ( \3049 , \3046 , \3048 );
xor \U$2861 ( \3050 , \2861 , \2865 );
xor \U$2862 ( \3051 , \3050 , \2870 );
and \U$2863 ( \3052 , \3048 , \3051 );
and \U$2864 ( \3053 , \3046 , \3051 );
or \U$2865 ( \3054 , \3049 , \3052 , \3053 );
and \U$2866 ( \3055 , \3044 , \3054 );
and \U$2867 ( \3056 , \1303 , \738 );
and \U$2868 ( \3057 , \1297 , \736 );
nor \U$2869 ( \3058 , \3056 , \3057 );
xnor \U$2870 ( \3059 , \3058 , \665 );
and \U$2871 ( \3060 , \1536 , \602 );
and \U$2872 ( \3061 , \1420 , \600 );
nor \U$2873 ( \3062 , \3060 , \3061 );
xnor \U$2874 ( \3063 , \3062 , \558 );
and \U$2875 ( \3064 , \3059 , \3063 );
and \U$2876 ( \3065 , \1777 , \502 );
and \U$2877 ( \3066 , \1768 , \500 );
nor \U$2878 ( \3067 , \3065 , \3066 );
xnor \U$2879 ( \3068 , \3067 , \453 );
and \U$2880 ( \3069 , \3063 , \3068 );
and \U$2881 ( \3070 , \3059 , \3068 );
or \U$2882 ( \3071 , \3064 , \3069 , \3070 );
and \U$2883 ( \3072 , \2027 , \296 );
and \U$2884 ( \3073 , \2021 , \294 );
nor \U$2885 ( \3074 , \3072 , \3073 );
xnor \U$2886 ( \3075 , \3074 , \301 );
and \U$2887 ( \3076 , \2304 , \310 );
and \U$2888 ( \3077 , \2159 , \308 );
nor \U$2889 ( \3078 , \3076 , \3077 );
xnor \U$2890 ( \3079 , \3078 , \318 );
and \U$2891 ( \3080 , \3075 , \3079 );
and \U$2892 ( \3081 , \2540 , \328 );
and \U$2893 ( \3082 , \2530 , \326 );
nor \U$2894 ( \3083 , \3081 , \3082 );
xnor \U$2895 ( \3084 , \3083 , \336 );
and \U$2896 ( \3085 , \3079 , \3084 );
and \U$2897 ( \3086 , \3075 , \3084 );
or \U$2898 ( \3087 , \3080 , \3085 , \3086 );
and \U$2899 ( \3088 , \3071 , \3087 );
xor \U$2900 ( \3089 , \2844 , \2848 );
xor \U$2901 ( \3090 , \3089 , \2853 );
and \U$2902 ( \3091 , \3087 , \3090 );
and \U$2903 ( \3092 , \3071 , \3090 );
or \U$2904 ( \3093 , \3088 , \3091 , \3092 );
and \U$2905 ( \3094 , \3054 , \3093 );
and \U$2906 ( \3095 , \3044 , \3093 );
or \U$2907 ( \3096 , \3055 , \3094 , \3095 );
xor \U$2908 ( \3097 , \2840 , \2856 );
xor \U$2909 ( \3098 , \3097 , \2873 );
xor \U$2910 ( \3099 , \2939 , \2941 );
xor \U$2911 ( \3100 , \3099 , \2944 );
and \U$2912 ( \3101 , \3098 , \3100 );
xor \U$2913 ( \3102 , \2927 , \2929 );
xor \U$2914 ( \3103 , \3102 , \2931 );
and \U$2915 ( \3104 , \3100 , \3103 );
and \U$2916 ( \3105 , \3098 , \3103 );
or \U$2917 ( \3106 , \3101 , \3104 , \3105 );
and \U$2918 ( \3107 , \3096 , \3106 );
xor \U$2919 ( \3108 , \2740 , \2756 );
xor \U$2920 ( \3109 , \3108 , \2765 );
and \U$2921 ( \3110 , \3106 , \3109 );
and \U$2922 ( \3111 , \3096 , \3109 );
or \U$2923 ( \3112 , \3107 , \3110 , \3111 );
xor \U$2924 ( \3113 , \2691 , \2704 );
xor \U$2925 ( \3114 , \3113 , \2721 );
xor \U$2926 ( \3115 , \2876 , \2924 );
xor \U$2927 ( \3116 , \3115 , \2934 );
and \U$2928 ( \3117 , \3114 , \3116 );
xor \U$2929 ( \3118 , \2947 , \2949 );
xor \U$2930 ( \3119 , \3118 , \2952 );
and \U$2931 ( \3120 , \3116 , \3119 );
and \U$2932 ( \3121 , \3114 , \3119 );
or \U$2933 ( \3122 , \3117 , \3120 , \3121 );
and \U$2934 ( \3123 , \3112 , \3122 );
xor \U$2935 ( \3124 , \2963 , \2965 );
xor \U$2936 ( \3125 , \3124 , \2968 );
and \U$2937 ( \3126 , \3122 , \3125 );
and \U$2938 ( \3127 , \3112 , \3125 );
or \U$2939 ( \3128 , \3123 , \3126 , \3127 );
xor \U$2940 ( \3129 , \2961 , \2971 );
xor \U$2941 ( \3130 , \3129 , \2974 );
and \U$2942 ( \3131 , \3128 , \3130 );
xor \U$2943 ( \3132 , \2979 , \2981 );
and \U$2944 ( \3133 , \3130 , \3132 );
and \U$2945 ( \3134 , \3128 , \3132 );
or \U$2946 ( \3135 , \3131 , \3133 , \3134 );
and \U$2947 ( \3136 , \2992 , \3135 );
xor \U$2948 ( \3137 , \2992 , \3135 );
xor \U$2949 ( \3138 , \3128 , \3130 );
xor \U$2950 ( \3139 , \3138 , \3132 );
and \U$2951 ( \3140 , \342 , \2259 );
and \U$2952 ( \3141 , \351 , \2257 );
nor \U$2953 ( \3142 , \3140 , \3141 );
xnor \U$2954 ( \3143 , \3142 , \2121 );
and \U$2955 ( \3144 , \444 , \1952 );
and \U$2956 ( \3145 , \359 , \1950 );
nor \U$2957 ( \3146 , \3144 , \3145 );
xnor \U$2958 ( \3147 , \3146 , \1832 );
and \U$2959 ( \3148 , \3143 , \3147 );
and \U$2960 ( \3149 , \591 , \1739 );
and \U$2961 ( \3150 , \494 , \1737 );
nor \U$2962 ( \3151 , \3149 , \3150 );
xnor \U$2963 ( \3152 , \3151 , \1607 );
and \U$2964 ( \3153 , \3147 , \3152 );
and \U$2965 ( \3154 , \3143 , \3152 );
or \U$2966 ( \3155 , \3148 , \3153 , \3154 );
and \U$2967 ( \3156 , \701 , \1474 );
and \U$2968 ( \3157 , \620 , \1472 );
nor \U$2969 ( \3158 , \3156 , \3157 );
xnor \U$2970 ( \3159 , \3158 , \1360 );
and \U$2971 ( \3160 , \839 , \1277 );
and \U$2972 ( \3161 , \776 , \1275 );
nor \U$2973 ( \3162 , \3160 , \3161 );
xnor \U$2974 ( \3163 , \3162 , \1173 );
and \U$2975 ( \3164 , \3159 , \3163 );
and \U$2976 ( \3165 , \1102 , \1059 );
and \U$2977 ( \3166 , \903 , \1057 );
nor \U$2978 ( \3167 , \3165 , \3166 );
xnor \U$2979 ( \3168 , \3167 , \981 );
and \U$2980 ( \3169 , \3163 , \3168 );
and \U$2981 ( \3170 , \3159 , \3168 );
or \U$2982 ( \3171 , \3164 , \3169 , \3170 );
and \U$2983 ( \3172 , \3155 , \3171 );
and \U$2984 ( \3173 , \304 , \2913 );
and \U$2985 ( \3174 , \313 , \2910 );
nor \U$2986 ( \3175 , \3173 , \3174 );
xnor \U$2987 ( \3176 , \3175 , \2368 );
and \U$2988 ( \3177 , \322 , \2549 );
and \U$2989 ( \3178 , \331 , \2547 );
nor \U$2990 ( \3179 , \3177 , \3178 );
xnor \U$2991 ( \3180 , \3179 , \2371 );
and \U$2992 ( \3181 , \3176 , \3180 );
and \U$2993 ( \3182 , \3180 , \356 );
and \U$2994 ( \3183 , \3176 , \356 );
or \U$2995 ( \3184 , \3181 , \3182 , \3183 );
and \U$2996 ( \3185 , \3171 , \3184 );
and \U$2997 ( \3186 , \3155 , \3184 );
or \U$2998 ( \3187 , \3172 , \3185 , \3186 );
and \U$2999 ( \3188 , \2021 , \502 );
and \U$3000 ( \3189 , \1777 , \500 );
nor \U$3001 ( \3190 , \3188 , \3189 );
xnor \U$3002 ( \3191 , \3190 , \453 );
and \U$3003 ( \3192 , \2159 , \296 );
and \U$3004 ( \3193 , \2027 , \294 );
nor \U$3005 ( \3194 , \3192 , \3193 );
xnor \U$3006 ( \3195 , \3194 , \301 );
and \U$3007 ( \3196 , \3191 , \3195 );
and \U$3008 ( \3197 , \2530 , \310 );
and \U$3009 ( \3198 , \2304 , \308 );
nor \U$3010 ( \3199 , \3197 , \3198 );
xnor \U$3011 ( \3200 , \3199 , \318 );
and \U$3012 ( \3201 , \3195 , \3200 );
and \U$3013 ( \3202 , \3191 , \3200 );
or \U$3014 ( \3203 , \3196 , \3201 , \3202 );
and \U$3015 ( \3204 , \1297 , \911 );
and \U$3016 ( \3205 , \1191 , \909 );
nor \U$3017 ( \3206 , \3204 , \3205 );
xnor \U$3018 ( \3207 , \3206 , \815 );
and \U$3019 ( \3208 , \1420 , \738 );
and \U$3020 ( \3209 , \1303 , \736 );
nor \U$3021 ( \3210 , \3208 , \3209 );
xnor \U$3022 ( \3211 , \3210 , \665 );
and \U$3023 ( \3212 , \3207 , \3211 );
and \U$3024 ( \3213 , \1768 , \602 );
and \U$3025 ( \3214 , \1536 , \600 );
nor \U$3026 ( \3215 , \3213 , \3214 );
xnor \U$3027 ( \3216 , \3215 , \558 );
and \U$3028 ( \3217 , \3211 , \3216 );
and \U$3029 ( \3218 , \3207 , \3216 );
or \U$3030 ( \3219 , \3212 , \3217 , \3218 );
and \U$3031 ( \3220 , \3203 , \3219 );
and \U$3032 ( \3221 , \2851 , \348 );
and \U$3033 ( \3222 , \2763 , \346 );
nor \U$3034 ( \3223 , \3221 , \3222 );
xnor \U$3035 ( \3224 , \3223 , \356 );
and \U$3036 ( \3225 , \3219 , \3224 );
and \U$3037 ( \3226 , \3203 , \3224 );
or \U$3038 ( \3227 , \3220 , \3225 , \3226 );
and \U$3039 ( \3228 , \3187 , \3227 );
xor \U$3040 ( \3229 , \3059 , \3063 );
xor \U$3041 ( \3230 , \3229 , \3068 );
xor \U$3042 ( \3231 , \3075 , \3079 );
xor \U$3043 ( \3232 , \3231 , \3084 );
and \U$3044 ( \3233 , \3230 , \3232 );
xor \U$3045 ( \3234 , \3029 , \3033 );
xor \U$3046 ( \3235 , \3234 , \3038 );
and \U$3047 ( \3236 , \3232 , \3235 );
and \U$3048 ( \3237 , \3230 , \3235 );
or \U$3049 ( \3238 , \3233 , \3236 , \3237 );
and \U$3050 ( \3239 , \3227 , \3238 );
and \U$3051 ( \3240 , \3187 , \3238 );
or \U$3052 ( \3241 , \3228 , \3239 , \3240 );
xor \U$3053 ( \3242 , \2896 , \2900 );
xor \U$3054 ( \3243 , \3242 , \2905 );
xor \U$3055 ( \3244 , \3046 , \3048 );
xor \U$3056 ( \3245 , \3244 , \3051 );
and \U$3057 ( \3246 , \3243 , \3245 );
xor \U$3058 ( \3247 , \2916 , \2920 );
and \U$3059 ( \3248 , \3245 , \3247 );
and \U$3060 ( \3249 , \3243 , \3247 );
or \U$3061 ( \3250 , \3246 , \3248 , \3249 );
and \U$3062 ( \3251 , \3241 , \3250 );
xor \U$3063 ( \3252 , \3008 , \3024 );
xor \U$3064 ( \3253 , \3252 , \3041 );
xor \U$3065 ( \3254 , \3071 , \3087 );
xor \U$3066 ( \3255 , \3254 , \3090 );
and \U$3067 ( \3256 , \3253 , \3255 );
and \U$3068 ( \3257 , \3250 , \3256 );
and \U$3069 ( \3258 , \3241 , \3256 );
or \U$3070 ( \3259 , \3251 , \3257 , \3258 );
xor \U$3071 ( \3260 , \2892 , \2908 );
xor \U$3072 ( \3261 , \3260 , \2921 );
xor \U$3073 ( \3262 , \3044 , \3054 );
xor \U$3074 ( \3263 , \3262 , \3093 );
and \U$3075 ( \3264 , \3261 , \3263 );
xor \U$3076 ( \3265 , \3098 , \3100 );
xor \U$3077 ( \3266 , \3265 , \3103 );
and \U$3078 ( \3267 , \3263 , \3266 );
and \U$3079 ( \3268 , \3261 , \3266 );
or \U$3080 ( \3269 , \3264 , \3267 , \3268 );
and \U$3081 ( \3270 , \3259 , \3269 );
xor \U$3082 ( \3271 , \3114 , \3116 );
xor \U$3083 ( \3272 , \3271 , \3119 );
and \U$3084 ( \3273 , \3269 , \3272 );
and \U$3085 ( \3274 , \3259 , \3272 );
or \U$3086 ( \3275 , \3270 , \3273 , \3274 );
xor \U$3087 ( \3276 , \2937 , \2955 );
xor \U$3088 ( \3277 , \3276 , \2958 );
and \U$3089 ( \3278 , \3275 , \3277 );
xor \U$3090 ( \3279 , \3112 , \3122 );
xor \U$3091 ( \3280 , \3279 , \3125 );
and \U$3092 ( \3281 , \3277 , \3280 );
and \U$3093 ( \3282 , \3275 , \3280 );
or \U$3094 ( \3283 , \3278 , \3281 , \3282 );
and \U$3095 ( \3284 , \3139 , \3283 );
xor \U$3096 ( \3285 , \3139 , \3283 );
xor \U$3097 ( \3286 , \3275 , \3277 );
xor \U$3098 ( \3287 , \3286 , \3280 );
and \U$3099 ( \3288 , \903 , \1277 );
and \U$3100 ( \3289 , \839 , \1275 );
nor \U$3101 ( \3290 , \3288 , \3289 );
xnor \U$3102 ( \3291 , \3290 , \1173 );
and \U$3103 ( \3292 , \1191 , \1059 );
and \U$3104 ( \3293 , \1102 , \1057 );
nor \U$3105 ( \3294 , \3292 , \3293 );
xnor \U$3106 ( \3295 , \3294 , \981 );
and \U$3107 ( \3296 , \3291 , \3295 );
and \U$3108 ( \3297 , \1303 , \911 );
and \U$3109 ( \3298 , \1297 , \909 );
nor \U$3110 ( \3299 , \3297 , \3298 );
xnor \U$3111 ( \3300 , \3299 , \815 );
and \U$3112 ( \3301 , \3295 , \3300 );
and \U$3113 ( \3302 , \3291 , \3300 );
or \U$3114 ( \3303 , \3296 , \3301 , \3302 );
and \U$3115 ( \3304 , \494 , \1952 );
and \U$3116 ( \3305 , \444 , \1950 );
nor \U$3117 ( \3306 , \3304 , \3305 );
xnor \U$3118 ( \3307 , \3306 , \1832 );
and \U$3119 ( \3308 , \620 , \1739 );
and \U$3120 ( \3309 , \591 , \1737 );
nor \U$3121 ( \3310 , \3308 , \3309 );
xnor \U$3122 ( \3311 , \3310 , \1607 );
and \U$3123 ( \3312 , \3307 , \3311 );
and \U$3124 ( \3313 , \776 , \1474 );
and \U$3125 ( \3314 , \701 , \1472 );
nor \U$3126 ( \3315 , \3313 , \3314 );
xnor \U$3127 ( \3316 , \3315 , \1360 );
and \U$3128 ( \3317 , \3311 , \3316 );
and \U$3129 ( \3318 , \3307 , \3316 );
or \U$3130 ( \3319 , \3312 , \3317 , \3318 );
and \U$3131 ( \3320 , \3303 , \3319 );
and \U$3132 ( \3321 , \331 , \2913 );
and \U$3133 ( \3322 , \304 , \2910 );
nor \U$3134 ( \3323 , \3321 , \3322 );
xnor \U$3135 ( \3324 , \3323 , \2368 );
and \U$3136 ( \3325 , \351 , \2549 );
and \U$3137 ( \3326 , \322 , \2547 );
nor \U$3138 ( \3327 , \3325 , \3326 );
xnor \U$3139 ( \3328 , \3327 , \2371 );
and \U$3140 ( \3329 , \3324 , \3328 );
and \U$3141 ( \3330 , \359 , \2259 );
and \U$3142 ( \3331 , \342 , \2257 );
nor \U$3143 ( \3332 , \3330 , \3331 );
xnor \U$3144 ( \3333 , \3332 , \2121 );
and \U$3145 ( \3334 , \3328 , \3333 );
and \U$3146 ( \3335 , \3324 , \3333 );
or \U$3147 ( \3336 , \3329 , \3334 , \3335 );
and \U$3148 ( \3337 , \3319 , \3336 );
and \U$3149 ( \3338 , \3303 , \3336 );
or \U$3150 ( \3339 , \3320 , \3337 , \3338 );
and \U$3151 ( \3340 , \2304 , \296 );
and \U$3152 ( \3341 , \2159 , \294 );
nor \U$3153 ( \3342 , \3340 , \3341 );
xnor \U$3154 ( \3343 , \3342 , \301 );
and \U$3155 ( \3344 , \2540 , \310 );
and \U$3156 ( \3345 , \2530 , \308 );
nor \U$3157 ( \3346 , \3344 , \3345 );
xnor \U$3158 ( \3347 , \3346 , \318 );
and \U$3159 ( \3348 , \3343 , \3347 );
and \U$3160 ( \3349 , \2851 , \328 );
and \U$3161 ( \3350 , \2763 , \326 );
nor \U$3162 ( \3351 , \3349 , \3350 );
xnor \U$3163 ( \3352 , \3351 , \336 );
and \U$3164 ( \3353 , \3347 , \3352 );
and \U$3165 ( \3354 , \3343 , \3352 );
or \U$3166 ( \3355 , \3348 , \3353 , \3354 );
and \U$3167 ( \3356 , \1536 , \738 );
and \U$3168 ( \3357 , \1420 , \736 );
nor \U$3169 ( \3358 , \3356 , \3357 );
xnor \U$3170 ( \3359 , \3358 , \665 );
and \U$3171 ( \3360 , \1777 , \602 );
and \U$3172 ( \3361 , \1768 , \600 );
nor \U$3173 ( \3362 , \3360 , \3361 );
xnor \U$3174 ( \3363 , \3362 , \558 );
and \U$3175 ( \3364 , \3359 , \3363 );
and \U$3176 ( \3365 , \2027 , \502 );
and \U$3177 ( \3366 , \2021 , \500 );
nor \U$3178 ( \3367 , \3365 , \3366 );
xnor \U$3179 ( \3368 , \3367 , \453 );
and \U$3180 ( \3369 , \3363 , \3368 );
and \U$3181 ( \3370 , \3359 , \3368 );
or \U$3182 ( \3371 , \3364 , \3369 , \3370 );
and \U$3183 ( \3372 , \3355 , \3371 );
and \U$3184 ( \3373 , \2763 , \328 );
and \U$3185 ( \3374 , \2540 , \326 );
nor \U$3186 ( \3375 , \3373 , \3374 );
xnor \U$3187 ( \3376 , \3375 , \336 );
and \U$3188 ( \3377 , \3371 , \3376 );
and \U$3189 ( \3378 , \3355 , \3376 );
or \U$3190 ( \3379 , \3372 , \3377 , \3378 );
and \U$3191 ( \3380 , \3339 , \3379 );
nand \U$3192 ( \3381 , \2851 , \346 );
xnor \U$3193 ( \3382 , \3381 , \356 );
xor \U$3194 ( \3383 , \3191 , \3195 );
xor \U$3195 ( \3384 , \3383 , \3200 );
and \U$3196 ( \3385 , \3382 , \3384 );
xor \U$3197 ( \3386 , \3207 , \3211 );
xor \U$3198 ( \3387 , \3386 , \3216 );
and \U$3199 ( \3388 , \3384 , \3387 );
and \U$3200 ( \3389 , \3382 , \3387 );
or \U$3201 ( \3390 , \3385 , \3388 , \3389 );
and \U$3202 ( \3391 , \3379 , \3390 );
and \U$3203 ( \3392 , \3339 , \3390 );
or \U$3204 ( \3393 , \3380 , \3391 , \3392 );
xor \U$3205 ( \3394 , \3143 , \3147 );
xor \U$3206 ( \3395 , \3394 , \3152 );
xor \U$3207 ( \3396 , \3159 , \3163 );
xor \U$3208 ( \3397 , \3396 , \3168 );
and \U$3209 ( \3398 , \3395 , \3397 );
xor \U$3210 ( \3399 , \3176 , \3180 );
xor \U$3211 ( \3400 , \3399 , \356 );
and \U$3212 ( \3401 , \3397 , \3400 );
and \U$3213 ( \3402 , \3395 , \3400 );
or \U$3214 ( \3403 , \3398 , \3401 , \3402 );
xor \U$3215 ( \3404 , \2996 , \3000 );
xor \U$3216 ( \3405 , \3404 , \3005 );
and \U$3217 ( \3406 , \3403 , \3405 );
xor \U$3218 ( \3407 , \3012 , \3016 );
xor \U$3219 ( \3408 , \3407 , \3021 );
and \U$3220 ( \3409 , \3405 , \3408 );
and \U$3221 ( \3410 , \3403 , \3408 );
or \U$3222 ( \3411 , \3406 , \3409 , \3410 );
and \U$3223 ( \3412 , \3393 , \3411 );
xor \U$3224 ( \3413 , \3155 , \3171 );
xor \U$3225 ( \3414 , \3413 , \3184 );
xor \U$3226 ( \3415 , \3203 , \3219 );
xor \U$3227 ( \3416 , \3415 , \3224 );
and \U$3228 ( \3417 , \3414 , \3416 );
xor \U$3229 ( \3418 , \3230 , \3232 );
xor \U$3230 ( \3419 , \3418 , \3235 );
and \U$3231 ( \3420 , \3416 , \3419 );
and \U$3232 ( \3421 , \3414 , \3419 );
or \U$3233 ( \3422 , \3417 , \3420 , \3421 );
and \U$3234 ( \3423 , \3411 , \3422 );
and \U$3235 ( \3424 , \3393 , \3422 );
or \U$3236 ( \3425 , \3412 , \3423 , \3424 );
xor \U$3237 ( \3426 , \3187 , \3227 );
xor \U$3238 ( \3427 , \3426 , \3238 );
xor \U$3239 ( \3428 , \3243 , \3245 );
xor \U$3240 ( \3429 , \3428 , \3247 );
and \U$3241 ( \3430 , \3427 , \3429 );
xor \U$3242 ( \3431 , \3253 , \3255 );
and \U$3243 ( \3432 , \3429 , \3431 );
and \U$3244 ( \3433 , \3427 , \3431 );
or \U$3245 ( \3434 , \3430 , \3432 , \3433 );
and \U$3246 ( \3435 , \3425 , \3434 );
xor \U$3247 ( \3436 , \3261 , \3263 );
xor \U$3248 ( \3437 , \3436 , \3266 );
and \U$3249 ( \3438 , \3434 , \3437 );
and \U$3250 ( \3439 , \3425 , \3437 );
or \U$3251 ( \3440 , \3435 , \3438 , \3439 );
xor \U$3252 ( \3441 , \3096 , \3106 );
xor \U$3253 ( \3442 , \3441 , \3109 );
and \U$3254 ( \3443 , \3440 , \3442 );
xor \U$3255 ( \3444 , \3259 , \3269 );
xor \U$3256 ( \3445 , \3444 , \3272 );
and \U$3257 ( \3446 , \3442 , \3445 );
and \U$3258 ( \3447 , \3440 , \3445 );
or \U$3259 ( \3448 , \3443 , \3446 , \3447 );
and \U$3260 ( \3449 , \3287 , \3448 );
xor \U$3261 ( \3450 , \3287 , \3448 );
xor \U$3262 ( \3451 , \3440 , \3442 );
xor \U$3263 ( \3452 , \3451 , \3445 );
and \U$3264 ( \3453 , \839 , \1474 );
and \U$3265 ( \3454 , \776 , \1472 );
nor \U$3266 ( \3455 , \3453 , \3454 );
xnor \U$3267 ( \3456 , \3455 , \1360 );
and \U$3268 ( \3457 , \1102 , \1277 );
and \U$3269 ( \3458 , \903 , \1275 );
nor \U$3270 ( \3459 , \3457 , \3458 );
xnor \U$3271 ( \3460 , \3459 , \1173 );
and \U$3272 ( \3461 , \3456 , \3460 );
and \U$3273 ( \3462 , \1297 , \1059 );
and \U$3274 ( \3463 , \1191 , \1057 );
nor \U$3275 ( \3464 , \3462 , \3463 );
xnor \U$3276 ( \3465 , \3464 , \981 );
and \U$3277 ( \3466 , \3460 , \3465 );
and \U$3278 ( \3467 , \3456 , \3465 );
or \U$3279 ( \3468 , \3461 , \3466 , \3467 );
and \U$3280 ( \3469 , \444 , \2259 );
and \U$3281 ( \3470 , \359 , \2257 );
nor \U$3282 ( \3471 , \3469 , \3470 );
xnor \U$3283 ( \3472 , \3471 , \2121 );
and \U$3284 ( \3473 , \591 , \1952 );
and \U$3285 ( \3474 , \494 , \1950 );
nor \U$3286 ( \3475 , \3473 , \3474 );
xnor \U$3287 ( \3476 , \3475 , \1832 );
and \U$3288 ( \3477 , \3472 , \3476 );
and \U$3289 ( \3478 , \701 , \1739 );
and \U$3290 ( \3479 , \620 , \1737 );
nor \U$3291 ( \3480 , \3478 , \3479 );
xnor \U$3292 ( \3481 , \3480 , \1607 );
and \U$3293 ( \3482 , \3476 , \3481 );
and \U$3294 ( \3483 , \3472 , \3481 );
or \U$3295 ( \3484 , \3477 , \3482 , \3483 );
and \U$3296 ( \3485 , \3468 , \3484 );
and \U$3297 ( \3486 , \322 , \2913 );
and \U$3298 ( \3487 , \331 , \2910 );
nor \U$3299 ( \3488 , \3486 , \3487 );
xnor \U$3300 ( \3489 , \3488 , \2368 );
and \U$3301 ( \3490 , \342 , \2549 );
and \U$3302 ( \3491 , \351 , \2547 );
nor \U$3303 ( \3492 , \3490 , \3491 );
xnor \U$3304 ( \3493 , \3492 , \2371 );
and \U$3305 ( \3494 , \3489 , \3493 );
and \U$3306 ( \3495 , \3493 , \336 );
and \U$3307 ( \3496 , \3489 , \336 );
or \U$3308 ( \3497 , \3494 , \3495 , \3496 );
and \U$3309 ( \3498 , \3484 , \3497 );
and \U$3310 ( \3499 , \3468 , \3497 );
or \U$3311 ( \3500 , \3485 , \3498 , \3499 );
and \U$3312 ( \3501 , \1420 , \911 );
and \U$3313 ( \3502 , \1303 , \909 );
nor \U$3314 ( \3503 , \3501 , \3502 );
xnor \U$3315 ( \3504 , \3503 , \815 );
and \U$3316 ( \3505 , \1768 , \738 );
and \U$3317 ( \3506 , \1536 , \736 );
nor \U$3318 ( \3507 , \3505 , \3506 );
xnor \U$3319 ( \3508 , \3507 , \665 );
and \U$3320 ( \3509 , \3504 , \3508 );
and \U$3321 ( \3510 , \2021 , \602 );
and \U$3322 ( \3511 , \1777 , \600 );
nor \U$3323 ( \3512 , \3510 , \3511 );
xnor \U$3324 ( \3513 , \3512 , \558 );
and \U$3325 ( \3514 , \3508 , \3513 );
and \U$3326 ( \3515 , \3504 , \3513 );
or \U$3327 ( \3516 , \3509 , \3514 , \3515 );
and \U$3328 ( \3517 , \2159 , \502 );
and \U$3329 ( \3518 , \2027 , \500 );
nor \U$3330 ( \3519 , \3517 , \3518 );
xnor \U$3331 ( \3520 , \3519 , \453 );
and \U$3332 ( \3521 , \2530 , \296 );
and \U$3333 ( \3522 , \2304 , \294 );
nor \U$3334 ( \3523 , \3521 , \3522 );
xnor \U$3335 ( \3524 , \3523 , \301 );
and \U$3336 ( \3525 , \3520 , \3524 );
and \U$3337 ( \3526 , \2763 , \310 );
and \U$3338 ( \3527 , \2540 , \308 );
nor \U$3339 ( \3528 , \3526 , \3527 );
xnor \U$3340 ( \3529 , \3528 , \318 );
and \U$3341 ( \3530 , \3524 , \3529 );
and \U$3342 ( \3531 , \3520 , \3529 );
or \U$3343 ( \3532 , \3525 , \3530 , \3531 );
and \U$3344 ( \3533 , \3516 , \3532 );
xor \U$3345 ( \3534 , \3343 , \3347 );
xor \U$3346 ( \3535 , \3534 , \3352 );
and \U$3347 ( \3536 , \3532 , \3535 );
and \U$3348 ( \3537 , \3516 , \3535 );
or \U$3349 ( \3538 , \3533 , \3536 , \3537 );
and \U$3350 ( \3539 , \3500 , \3538 );
xor \U$3351 ( \3540 , \3291 , \3295 );
xor \U$3352 ( \3541 , \3540 , \3300 );
xor \U$3353 ( \3542 , \3307 , \3311 );
xor \U$3354 ( \3543 , \3542 , \3316 );
and \U$3355 ( \3544 , \3541 , \3543 );
xor \U$3356 ( \3545 , \3359 , \3363 );
xor \U$3357 ( \3546 , \3545 , \3368 );
and \U$3358 ( \3547 , \3543 , \3546 );
and \U$3359 ( \3548 , \3541 , \3546 );
or \U$3360 ( \3549 , \3544 , \3547 , \3548 );
and \U$3361 ( \3550 , \3538 , \3549 );
and \U$3362 ( \3551 , \3500 , \3549 );
or \U$3363 ( \3552 , \3539 , \3550 , \3551 );
xor \U$3364 ( \3553 , \3355 , \3371 );
xor \U$3365 ( \3554 , \3553 , \3376 );
xor \U$3366 ( \3555 , \3395 , \3397 );
xor \U$3367 ( \3556 , \3555 , \3400 );
and \U$3368 ( \3557 , \3554 , \3556 );
xor \U$3369 ( \3558 , \3382 , \3384 );
xor \U$3370 ( \3559 , \3558 , \3387 );
and \U$3371 ( \3560 , \3556 , \3559 );
and \U$3372 ( \3561 , \3554 , \3559 );
or \U$3373 ( \3562 , \3557 , \3560 , \3561 );
and \U$3374 ( \3563 , \3552 , \3562 );
xor \U$3375 ( \3564 , \3414 , \3416 );
xor \U$3376 ( \3565 , \3564 , \3419 );
and \U$3377 ( \3566 , \3562 , \3565 );
and \U$3378 ( \3567 , \3552 , \3565 );
or \U$3379 ( \3568 , \3563 , \3566 , \3567 );
xor \U$3380 ( \3569 , \3339 , \3379 );
xor \U$3381 ( \3570 , \3569 , \3390 );
xor \U$3382 ( \3571 , \3403 , \3405 );
xor \U$3383 ( \3572 , \3571 , \3408 );
and \U$3384 ( \3573 , \3570 , \3572 );
and \U$3385 ( \3574 , \3568 , \3573 );
xor \U$3386 ( \3575 , \3427 , \3429 );
xor \U$3387 ( \3576 , \3575 , \3431 );
and \U$3388 ( \3577 , \3573 , \3576 );
and \U$3389 ( \3578 , \3568 , \3576 );
or \U$3390 ( \3579 , \3574 , \3577 , \3578 );
xor \U$3391 ( \3580 , \3241 , \3250 );
xor \U$3392 ( \3581 , \3580 , \3256 );
and \U$3393 ( \3582 , \3579 , \3581 );
xor \U$3394 ( \3583 , \3425 , \3434 );
xor \U$3395 ( \3584 , \3583 , \3437 );
and \U$3396 ( \3585 , \3581 , \3584 );
and \U$3397 ( \3586 , \3579 , \3584 );
or \U$3398 ( \3587 , \3582 , \3585 , \3586 );
and \U$3399 ( \3588 , \3452 , \3587 );
xor \U$3400 ( \3589 , \3452 , \3587 );
xor \U$3401 ( \3590 , \3579 , \3581 );
xor \U$3402 ( \3591 , \3590 , \3584 );
and \U$3403 ( \3592 , \351 , \2913 );
and \U$3404 ( \3593 , \322 , \2910 );
nor \U$3405 ( \3594 , \3592 , \3593 );
xnor \U$3406 ( \3595 , \3594 , \2368 );
and \U$3407 ( \3596 , \359 , \2549 );
and \U$3408 ( \3597 , \342 , \2547 );
nor \U$3409 ( \3598 , \3596 , \3597 );
xnor \U$3410 ( \3599 , \3598 , \2371 );
and \U$3411 ( \3600 , \3595 , \3599 );
and \U$3412 ( \3601 , \494 , \2259 );
and \U$3413 ( \3602 , \444 , \2257 );
nor \U$3414 ( \3603 , \3601 , \3602 );
xnor \U$3415 ( \3604 , \3603 , \2121 );
and \U$3416 ( \3605 , \3599 , \3604 );
and \U$3417 ( \3606 , \3595 , \3604 );
or \U$3418 ( \3607 , \3600 , \3605 , \3606 );
and \U$3419 ( \3608 , \1191 , \1277 );
and \U$3420 ( \3609 , \1102 , \1275 );
nor \U$3421 ( \3610 , \3608 , \3609 );
xnor \U$3422 ( \3611 , \3610 , \1173 );
and \U$3423 ( \3612 , \1303 , \1059 );
and \U$3424 ( \3613 , \1297 , \1057 );
nor \U$3425 ( \3614 , \3612 , \3613 );
xnor \U$3426 ( \3615 , \3614 , \981 );
and \U$3427 ( \3616 , \3611 , \3615 );
and \U$3428 ( \3617 , \1536 , \911 );
and \U$3429 ( \3618 , \1420 , \909 );
nor \U$3430 ( \3619 , \3617 , \3618 );
xnor \U$3431 ( \3620 , \3619 , \815 );
and \U$3432 ( \3621 , \3615 , \3620 );
and \U$3433 ( \3622 , \3611 , \3620 );
or \U$3434 ( \3623 , \3616 , \3621 , \3622 );
and \U$3435 ( \3624 , \3607 , \3623 );
and \U$3436 ( \3625 , \620 , \1952 );
and \U$3437 ( \3626 , \591 , \1950 );
nor \U$3438 ( \3627 , \3625 , \3626 );
xnor \U$3439 ( \3628 , \3627 , \1832 );
and \U$3440 ( \3629 , \776 , \1739 );
and \U$3441 ( \3630 , \701 , \1737 );
nor \U$3442 ( \3631 , \3629 , \3630 );
xnor \U$3443 ( \3632 , \3631 , \1607 );
and \U$3444 ( \3633 , \3628 , \3632 );
and \U$3445 ( \3634 , \903 , \1474 );
and \U$3446 ( \3635 , \839 , \1472 );
nor \U$3447 ( \3636 , \3634 , \3635 );
xnor \U$3448 ( \3637 , \3636 , \1360 );
and \U$3449 ( \3638 , \3632 , \3637 );
and \U$3450 ( \3639 , \3628 , \3637 );
or \U$3451 ( \3640 , \3633 , \3638 , \3639 );
and \U$3452 ( \3641 , \3623 , \3640 );
and \U$3453 ( \3642 , \3607 , \3640 );
or \U$3454 ( \3643 , \3624 , \3641 , \3642 );
xor \U$3455 ( \3644 , \3456 , \3460 );
xor \U$3456 ( \3645 , \3644 , \3465 );
xor \U$3457 ( \3646 , \3472 , \3476 );
xor \U$3458 ( \3647 , \3646 , \3481 );
and \U$3459 ( \3648 , \3645 , \3647 );
xor \U$3460 ( \3649 , \3504 , \3508 );
xor \U$3461 ( \3650 , \3649 , \3513 );
and \U$3462 ( \3651 , \3647 , \3650 );
and \U$3463 ( \3652 , \3645 , \3650 );
or \U$3464 ( \3653 , \3648 , \3651 , \3652 );
and \U$3465 ( \3654 , \3643 , \3653 );
and \U$3466 ( \3655 , \1777 , \738 );
and \U$3467 ( \3656 , \1768 , \736 );
nor \U$3468 ( \3657 , \3655 , \3656 );
xnor \U$3469 ( \3658 , \3657 , \665 );
and \U$3470 ( \3659 , \2027 , \602 );
and \U$3471 ( \3660 , \2021 , \600 );
nor \U$3472 ( \3661 , \3659 , \3660 );
xnor \U$3473 ( \3662 , \3661 , \558 );
and \U$3474 ( \3663 , \3658 , \3662 );
and \U$3475 ( \3664 , \2304 , \502 );
and \U$3476 ( \3665 , \2159 , \500 );
nor \U$3477 ( \3666 , \3664 , \3665 );
xnor \U$3478 ( \3667 , \3666 , \453 );
and \U$3479 ( \3668 , \3662 , \3667 );
and \U$3480 ( \3669 , \3658 , \3667 );
or \U$3481 ( \3670 , \3663 , \3668 , \3669 );
nand \U$3482 ( \3671 , \2851 , \326 );
xnor \U$3483 ( \3672 , \3671 , \336 );
and \U$3484 ( \3673 , \3670 , \3672 );
xor \U$3485 ( \3674 , \3520 , \3524 );
xor \U$3486 ( \3675 , \3674 , \3529 );
and \U$3487 ( \3676 , \3672 , \3675 );
and \U$3488 ( \3677 , \3670 , \3675 );
or \U$3489 ( \3678 , \3673 , \3676 , \3677 );
and \U$3490 ( \3679 , \3653 , \3678 );
and \U$3491 ( \3680 , \3643 , \3678 );
or \U$3492 ( \3681 , \3654 , \3679 , \3680 );
xor \U$3493 ( \3682 , \3324 , \3328 );
xor \U$3494 ( \3683 , \3682 , \3333 );
xor \U$3495 ( \3684 , \3516 , \3532 );
xor \U$3496 ( \3685 , \3684 , \3535 );
and \U$3497 ( \3686 , \3683 , \3685 );
xor \U$3498 ( \3687 , \3541 , \3543 );
xor \U$3499 ( \3688 , \3687 , \3546 );
and \U$3500 ( \3689 , \3685 , \3688 );
and \U$3501 ( \3690 , \3683 , \3688 );
or \U$3502 ( \3691 , \3686 , \3689 , \3690 );
and \U$3503 ( \3692 , \3681 , \3691 );
xor \U$3504 ( \3693 , \3303 , \3319 );
xor \U$3505 ( \3694 , \3693 , \3336 );
and \U$3506 ( \3695 , \3691 , \3694 );
and \U$3507 ( \3696 , \3681 , \3694 );
or \U$3508 ( \3697 , \3692 , \3695 , \3696 );
xor \U$3509 ( \3698 , \3552 , \3562 );
xor \U$3510 ( \3699 , \3698 , \3565 );
and \U$3511 ( \3700 , \3697 , \3699 );
xor \U$3512 ( \3701 , \3570 , \3572 );
and \U$3513 ( \3702 , \3699 , \3701 );
and \U$3514 ( \3703 , \3697 , \3701 );
or \U$3515 ( \3704 , \3700 , \3702 , \3703 );
xor \U$3516 ( \3705 , \3393 , \3411 );
xor \U$3517 ( \3706 , \3705 , \3422 );
and \U$3518 ( \3707 , \3704 , \3706 );
xor \U$3519 ( \3708 , \3568 , \3573 );
xor \U$3520 ( \3709 , \3708 , \3576 );
and \U$3521 ( \3710 , \3706 , \3709 );
and \U$3522 ( \3711 , \3704 , \3709 );
or \U$3523 ( \3712 , \3707 , \3710 , \3711 );
and \U$3524 ( \3713 , \3591 , \3712 );
xor \U$3525 ( \3714 , \3591 , \3712 );
xor \U$3526 ( \3715 , \3704 , \3706 );
xor \U$3527 ( \3716 , \3715 , \3709 );
and \U$3528 ( \3717 , \1768 , \911 );
and \U$3529 ( \3718 , \1536 , \909 );
nor \U$3530 ( \3719 , \3717 , \3718 );
xnor \U$3531 ( \3720 , \3719 , \815 );
and \U$3532 ( \3721 , \2021 , \738 );
and \U$3533 ( \3722 , \1777 , \736 );
nor \U$3534 ( \3723 , \3721 , \3722 );
xnor \U$3535 ( \3724 , \3723 , \665 );
and \U$3536 ( \3725 , \3720 , \3724 );
and \U$3537 ( \3726 , \2159 , \602 );
and \U$3538 ( \3727 , \2027 , \600 );
nor \U$3539 ( \3728 , \3726 , \3727 );
xnor \U$3540 ( \3729 , \3728 , \558 );
and \U$3541 ( \3730 , \3724 , \3729 );
and \U$3542 ( \3731 , \3720 , \3729 );
or \U$3543 ( \3732 , \3725 , \3730 , \3731 );
and \U$3544 ( \3733 , \2530 , \502 );
and \U$3545 ( \3734 , \2304 , \500 );
nor \U$3546 ( \3735 , \3733 , \3734 );
xnor \U$3547 ( \3736 , \3735 , \453 );
and \U$3548 ( \3737 , \2763 , \296 );
and \U$3549 ( \3738 , \2540 , \294 );
nor \U$3550 ( \3739 , \3737 , \3738 );
xnor \U$3551 ( \3740 , \3739 , \301 );
and \U$3552 ( \3741 , \3736 , \3740 );
nand \U$3553 ( \3742 , \2851 , \308 );
xnor \U$3554 ( \3743 , \3742 , \318 );
and \U$3555 ( \3744 , \3740 , \3743 );
and \U$3556 ( \3745 , \3736 , \3743 );
or \U$3557 ( \3746 , \3741 , \3744 , \3745 );
and \U$3558 ( \3747 , \3732 , \3746 );
and \U$3559 ( \3748 , \2540 , \296 );
and \U$3560 ( \3749 , \2530 , \294 );
nor \U$3561 ( \3750 , \3748 , \3749 );
xnor \U$3562 ( \3751 , \3750 , \301 );
and \U$3563 ( \3752 , \3746 , \3751 );
and \U$3564 ( \3753 , \3732 , \3751 );
or \U$3565 ( \3754 , \3747 , \3752 , \3753 );
and \U$3566 ( \3755 , \1102 , \1474 );
and \U$3567 ( \3756 , \903 , \1472 );
nor \U$3568 ( \3757 , \3755 , \3756 );
xnor \U$3569 ( \3758 , \3757 , \1360 );
and \U$3570 ( \3759 , \1297 , \1277 );
and \U$3571 ( \3760 , \1191 , \1275 );
nor \U$3572 ( \3761 , \3759 , \3760 );
xnor \U$3573 ( \3762 , \3761 , \1173 );
and \U$3574 ( \3763 , \3758 , \3762 );
and \U$3575 ( \3764 , \1420 , \1059 );
and \U$3576 ( \3765 , \1303 , \1057 );
nor \U$3577 ( \3766 , \3764 , \3765 );
xnor \U$3578 ( \3767 , \3766 , \981 );
and \U$3579 ( \3768 , \3762 , \3767 );
and \U$3580 ( \3769 , \3758 , \3767 );
or \U$3581 ( \3770 , \3763 , \3768 , \3769 );
and \U$3582 ( \3771 , \342 , \2913 );
and \U$3583 ( \3772 , \351 , \2910 );
nor \U$3584 ( \3773 , \3771 , \3772 );
xnor \U$3585 ( \3774 , \3773 , \2368 );
and \U$3586 ( \3775 , \444 , \2549 );
and \U$3587 ( \3776 , \359 , \2547 );
nor \U$3588 ( \3777 , \3775 , \3776 );
xnor \U$3589 ( \3778 , \3777 , \2371 );
and \U$3590 ( \3779 , \3774 , \3778 );
and \U$3591 ( \3780 , \3778 , \318 );
and \U$3592 ( \3781 , \3774 , \318 );
or \U$3593 ( \3782 , \3779 , \3780 , \3781 );
and \U$3594 ( \3783 , \3770 , \3782 );
and \U$3595 ( \3784 , \591 , \2259 );
and \U$3596 ( \3785 , \494 , \2257 );
nor \U$3597 ( \3786 , \3784 , \3785 );
xnor \U$3598 ( \3787 , \3786 , \2121 );
and \U$3599 ( \3788 , \701 , \1952 );
and \U$3600 ( \3789 , \620 , \1950 );
nor \U$3601 ( \3790 , \3788 , \3789 );
xnor \U$3602 ( \3791 , \3790 , \1832 );
and \U$3603 ( \3792 , \3787 , \3791 );
and \U$3604 ( \3793 , \839 , \1739 );
and \U$3605 ( \3794 , \776 , \1737 );
nor \U$3606 ( \3795 , \3793 , \3794 );
xnor \U$3607 ( \3796 , \3795 , \1607 );
and \U$3608 ( \3797 , \3791 , \3796 );
and \U$3609 ( \3798 , \3787 , \3796 );
or \U$3610 ( \3799 , \3792 , \3797 , \3798 );
and \U$3611 ( \3800 , \3782 , \3799 );
and \U$3612 ( \3801 , \3770 , \3799 );
or \U$3613 ( \3802 , \3783 , \3800 , \3801 );
and \U$3614 ( \3803 , \3754 , \3802 );
and \U$3615 ( \3804 , \2851 , \310 );
and \U$3616 ( \3805 , \2763 , \308 );
nor \U$3617 ( \3806 , \3804 , \3805 );
xnor \U$3618 ( \3807 , \3806 , \318 );
xor \U$3619 ( \3808 , \3658 , \3662 );
xor \U$3620 ( \3809 , \3808 , \3667 );
and \U$3621 ( \3810 , \3807 , \3809 );
xor \U$3622 ( \3811 , \3611 , \3615 );
xor \U$3623 ( \3812 , \3811 , \3620 );
and \U$3624 ( \3813 , \3809 , \3812 );
and \U$3625 ( \3814 , \3807 , \3812 );
or \U$3626 ( \3815 , \3810 , \3813 , \3814 );
and \U$3627 ( \3816 , \3802 , \3815 );
and \U$3628 ( \3817 , \3754 , \3815 );
or \U$3629 ( \3818 , \3803 , \3816 , \3817 );
xor \U$3630 ( \3819 , \3489 , \3493 );
xor \U$3631 ( \3820 , \3819 , \336 );
xor \U$3632 ( \3821 , \3645 , \3647 );
xor \U$3633 ( \3822 , \3821 , \3650 );
and \U$3634 ( \3823 , \3820 , \3822 );
xor \U$3635 ( \3824 , \3670 , \3672 );
xor \U$3636 ( \3825 , \3824 , \3675 );
and \U$3637 ( \3826 , \3822 , \3825 );
and \U$3638 ( \3827 , \3820 , \3825 );
or \U$3639 ( \3828 , \3823 , \3826 , \3827 );
and \U$3640 ( \3829 , \3818 , \3828 );
xor \U$3641 ( \3830 , \3468 , \3484 );
xor \U$3642 ( \3831 , \3830 , \3497 );
and \U$3643 ( \3832 , \3828 , \3831 );
and \U$3644 ( \3833 , \3818 , \3831 );
or \U$3645 ( \3834 , \3829 , \3832 , \3833 );
xor \U$3646 ( \3835 , \3643 , \3653 );
xor \U$3647 ( \3836 , \3835 , \3678 );
xor \U$3648 ( \3837 , \3683 , \3685 );
xor \U$3649 ( \3838 , \3837 , \3688 );
and \U$3650 ( \3839 , \3836 , \3838 );
and \U$3651 ( \3840 , \3834 , \3839 );
xor \U$3652 ( \3841 , \3554 , \3556 );
xor \U$3653 ( \3842 , \3841 , \3559 );
and \U$3654 ( \3843 , \3839 , \3842 );
and \U$3655 ( \3844 , \3834 , \3842 );
or \U$3656 ( \3845 , \3840 , \3843 , \3844 );
xor \U$3657 ( \3846 , \3500 , \3538 );
xor \U$3658 ( \3847 , \3846 , \3549 );
xor \U$3659 ( \3848 , \3681 , \3691 );
xor \U$3660 ( \3849 , \3848 , \3694 );
and \U$3661 ( \3850 , \3847 , \3849 );
and \U$3662 ( \3851 , \3845 , \3850 );
xor \U$3663 ( \3852 , \3697 , \3699 );
xor \U$3664 ( \3853 , \3852 , \3701 );
and \U$3665 ( \3854 , \3850 , \3853 );
and \U$3666 ( \3855 , \3845 , \3853 );
or \U$3667 ( \3856 , \3851 , \3854 , \3855 );
and \U$3668 ( \3857 , \3716 , \3856 );
xor \U$3669 ( \3858 , \3716 , \3856 );
xor \U$3670 ( \3859 , \3845 , \3850 );
xor \U$3671 ( \3860 , \3859 , \3853 );
and \U$3672 ( \3861 , \776 , \1952 );
and \U$3673 ( \3862 , \701 , \1950 );
nor \U$3674 ( \3863 , \3861 , \3862 );
xnor \U$3675 ( \3864 , \3863 , \1832 );
and \U$3676 ( \3865 , \903 , \1739 );
and \U$3677 ( \3866 , \839 , \1737 );
nor \U$3678 ( \3867 , \3865 , \3866 );
xnor \U$3679 ( \3868 , \3867 , \1607 );
and \U$3680 ( \3869 , \3864 , \3868 );
and \U$3681 ( \3870 , \1191 , \1474 );
and \U$3682 ( \3871 , \1102 , \1472 );
nor \U$3683 ( \3872 , \3870 , \3871 );
xnor \U$3684 ( \3873 , \3872 , \1360 );
and \U$3685 ( \3874 , \3868 , \3873 );
and \U$3686 ( \3875 , \3864 , \3873 );
or \U$3687 ( \3876 , \3869 , \3874 , \3875 );
and \U$3688 ( \3877 , \359 , \2913 );
and \U$3689 ( \3878 , \342 , \2910 );
nor \U$3690 ( \3879 , \3877 , \3878 );
xnor \U$3691 ( \3880 , \3879 , \2368 );
and \U$3692 ( \3881 , \494 , \2549 );
and \U$3693 ( \3882 , \444 , \2547 );
nor \U$3694 ( \3883 , \3881 , \3882 );
xnor \U$3695 ( \3884 , \3883 , \2371 );
and \U$3696 ( \3885 , \3880 , \3884 );
and \U$3697 ( \3886 , \620 , \2259 );
and \U$3698 ( \3887 , \591 , \2257 );
nor \U$3699 ( \3888 , \3886 , \3887 );
xnor \U$3700 ( \3889 , \3888 , \2121 );
and \U$3701 ( \3890 , \3884 , \3889 );
and \U$3702 ( \3891 , \3880 , \3889 );
or \U$3703 ( \3892 , \3885 , \3890 , \3891 );
and \U$3704 ( \3893 , \3876 , \3892 );
and \U$3705 ( \3894 , \1303 , \1277 );
and \U$3706 ( \3895 , \1297 , \1275 );
nor \U$3707 ( \3896 , \3894 , \3895 );
xnor \U$3708 ( \3897 , \3896 , \1173 );
and \U$3709 ( \3898 , \1536 , \1059 );
and \U$3710 ( \3899 , \1420 , \1057 );
nor \U$3711 ( \3900 , \3898 , \3899 );
xnor \U$3712 ( \3901 , \3900 , \981 );
and \U$3713 ( \3902 , \3897 , \3901 );
and \U$3714 ( \3903 , \1777 , \911 );
and \U$3715 ( \3904 , \1768 , \909 );
nor \U$3716 ( \3905 , \3903 , \3904 );
xnor \U$3717 ( \3906 , \3905 , \815 );
and \U$3718 ( \3907 , \3901 , \3906 );
and \U$3719 ( \3908 , \3897 , \3906 );
or \U$3720 ( \3909 , \3902 , \3907 , \3908 );
and \U$3721 ( \3910 , \3892 , \3909 );
and \U$3722 ( \3911 , \3876 , \3909 );
or \U$3723 ( \3912 , \3893 , \3910 , \3911 );
xor \U$3724 ( \3913 , \3758 , \3762 );
xor \U$3725 ( \3914 , \3913 , \3767 );
xor \U$3726 ( \3915 , \3774 , \3778 );
xor \U$3727 ( \3916 , \3915 , \318 );
and \U$3728 ( \3917 , \3914 , \3916 );
xor \U$3729 ( \3918 , \3787 , \3791 );
xor \U$3730 ( \3919 , \3918 , \3796 );
and \U$3731 ( \3920 , \3916 , \3919 );
and \U$3732 ( \3921 , \3914 , \3919 );
or \U$3733 ( \3922 , \3917 , \3920 , \3921 );
and \U$3734 ( \3923 , \3912 , \3922 );
and \U$3735 ( \3924 , \2027 , \738 );
and \U$3736 ( \3925 , \2021 , \736 );
nor \U$3737 ( \3926 , \3924 , \3925 );
xnor \U$3738 ( \3927 , \3926 , \665 );
and \U$3739 ( \3928 , \2304 , \602 );
and \U$3740 ( \3929 , \2159 , \600 );
nor \U$3741 ( \3930 , \3928 , \3929 );
xnor \U$3742 ( \3931 , \3930 , \558 );
and \U$3743 ( \3932 , \3927 , \3931 );
and \U$3744 ( \3933 , \2540 , \502 );
and \U$3745 ( \3934 , \2530 , \500 );
nor \U$3746 ( \3935 , \3933 , \3934 );
xnor \U$3747 ( \3936 , \3935 , \453 );
and \U$3748 ( \3937 , \3931 , \3936 );
and \U$3749 ( \3938 , \3927 , \3936 );
or \U$3750 ( \3939 , \3932 , \3937 , \3938 );
xor \U$3751 ( \3940 , \3720 , \3724 );
xor \U$3752 ( \3941 , \3940 , \3729 );
and \U$3753 ( \3942 , \3939 , \3941 );
xor \U$3754 ( \3943 , \3736 , \3740 );
xor \U$3755 ( \3944 , \3943 , \3743 );
and \U$3756 ( \3945 , \3941 , \3944 );
and \U$3757 ( \3946 , \3939 , \3944 );
or \U$3758 ( \3947 , \3942 , \3945 , \3946 );
and \U$3759 ( \3948 , \3922 , \3947 );
and \U$3760 ( \3949 , \3912 , \3947 );
or \U$3761 ( \3950 , \3923 , \3948 , \3949 );
xor \U$3762 ( \3951 , \3595 , \3599 );
xor \U$3763 ( \3952 , \3951 , \3604 );
xor \U$3764 ( \3953 , \3628 , \3632 );
xor \U$3765 ( \3954 , \3953 , \3637 );
and \U$3766 ( \3955 , \3952 , \3954 );
xor \U$3767 ( \3956 , \3807 , \3809 );
xor \U$3768 ( \3957 , \3956 , \3812 );
and \U$3769 ( \3958 , \3954 , \3957 );
and \U$3770 ( \3959 , \3952 , \3957 );
or \U$3771 ( \3960 , \3955 , \3958 , \3959 );
and \U$3772 ( \3961 , \3950 , \3960 );
xor \U$3773 ( \3962 , \3607 , \3623 );
xor \U$3774 ( \3963 , \3962 , \3640 );
and \U$3775 ( \3964 , \3960 , \3963 );
and \U$3776 ( \3965 , \3950 , \3963 );
or \U$3777 ( \3966 , \3961 , \3964 , \3965 );
xor \U$3778 ( \3967 , \3818 , \3828 );
xor \U$3779 ( \3968 , \3967 , \3831 );
and \U$3780 ( \3969 , \3966 , \3968 );
xor \U$3781 ( \3970 , \3836 , \3838 );
and \U$3782 ( \3971 , \3968 , \3970 );
and \U$3783 ( \3972 , \3966 , \3970 );
or \U$3784 ( \3973 , \3969 , \3971 , \3972 );
xor \U$3785 ( \3974 , \3834 , \3839 );
xor \U$3786 ( \3975 , \3974 , \3842 );
and \U$3787 ( \3976 , \3973 , \3975 );
xor \U$3788 ( \3977 , \3847 , \3849 );
and \U$3789 ( \3978 , \3975 , \3977 );
and \U$3790 ( \3979 , \3973 , \3977 );
or \U$3791 ( \3980 , \3976 , \3978 , \3979 );
and \U$3792 ( \3981 , \3860 , \3980 );
xor \U$3793 ( \3982 , \3860 , \3980 );
xor \U$3794 ( \3983 , \3973 , \3975 );
xor \U$3795 ( \3984 , \3983 , \3977 );
and \U$3796 ( \3985 , \701 , \2259 );
and \U$3797 ( \3986 , \620 , \2257 );
nor \U$3798 ( \3987 , \3985 , \3986 );
xnor \U$3799 ( \3988 , \3987 , \2121 );
and \U$3800 ( \3989 , \839 , \1952 );
and \U$3801 ( \3990 , \776 , \1950 );
nor \U$3802 ( \3991 , \3989 , \3990 );
xnor \U$3803 ( \3992 , \3991 , \1832 );
and \U$3804 ( \3993 , \3988 , \3992 );
and \U$3805 ( \3994 , \1102 , \1739 );
and \U$3806 ( \3995 , \903 , \1737 );
nor \U$3807 ( \3996 , \3994 , \3995 );
xnor \U$3808 ( \3997 , \3996 , \1607 );
and \U$3809 ( \3998 , \3992 , \3997 );
and \U$3810 ( \3999 , \3988 , \3997 );
or \U$3811 ( \4000 , \3993 , \3998 , \3999 );
and \U$3812 ( \4001 , \444 , \2913 );
and \U$3813 ( \4002 , \359 , \2910 );
nor \U$3814 ( \4003 , \4001 , \4002 );
xnor \U$3815 ( \4004 , \4003 , \2368 );
and \U$3816 ( \4005 , \591 , \2549 );
and \U$3817 ( \4006 , \494 , \2547 );
nor \U$3818 ( \4007 , \4005 , \4006 );
xnor \U$3819 ( \4008 , \4007 , \2371 );
and \U$3820 ( \4009 , \4004 , \4008 );
and \U$3821 ( \4010 , \4008 , \301 );
and \U$3822 ( \4011 , \4004 , \301 );
or \U$3823 ( \4012 , \4009 , \4010 , \4011 );
and \U$3824 ( \4013 , \4000 , \4012 );
and \U$3825 ( \4014 , \1297 , \1474 );
and \U$3826 ( \4015 , \1191 , \1472 );
nor \U$3827 ( \4016 , \4014 , \4015 );
xnor \U$3828 ( \4017 , \4016 , \1360 );
and \U$3829 ( \4018 , \1420 , \1277 );
and \U$3830 ( \4019 , \1303 , \1275 );
nor \U$3831 ( \4020 , \4018 , \4019 );
xnor \U$3832 ( \4021 , \4020 , \1173 );
and \U$3833 ( \4022 , \4017 , \4021 );
and \U$3834 ( \4023 , \1768 , \1059 );
and \U$3835 ( \4024 , \1536 , \1057 );
nor \U$3836 ( \4025 , \4023 , \4024 );
xnor \U$3837 ( \4026 , \4025 , \981 );
and \U$3838 ( \4027 , \4021 , \4026 );
and \U$3839 ( \4028 , \4017 , \4026 );
or \U$3840 ( \4029 , \4022 , \4027 , \4028 );
and \U$3841 ( \4030 , \4012 , \4029 );
and \U$3842 ( \4031 , \4000 , \4029 );
or \U$3843 ( \4032 , \4013 , \4030 , \4031 );
and \U$3844 ( \4033 , \2021 , \911 );
and \U$3845 ( \4034 , \1777 , \909 );
nor \U$3846 ( \4035 , \4033 , \4034 );
xnor \U$3847 ( \4036 , \4035 , \815 );
and \U$3848 ( \4037 , \2159 , \738 );
and \U$3849 ( \4038 , \2027 , \736 );
nor \U$3850 ( \4039 , \4037 , \4038 );
xnor \U$3851 ( \4040 , \4039 , \665 );
and \U$3852 ( \4041 , \4036 , \4040 );
and \U$3853 ( \4042 , \2530 , \602 );
and \U$3854 ( \4043 , \2304 , \600 );
nor \U$3855 ( \4044 , \4042 , \4043 );
xnor \U$3856 ( \4045 , \4044 , \558 );
and \U$3857 ( \4046 , \4040 , \4045 );
and \U$3858 ( \4047 , \4036 , \4045 );
or \U$3859 ( \4048 , \4041 , \4046 , \4047 );
and \U$3860 ( \4049 , \2763 , \502 );
and \U$3861 ( \4050 , \2540 , \500 );
nor \U$3862 ( \4051 , \4049 , \4050 );
xnor \U$3863 ( \4052 , \4051 , \453 );
nand \U$3864 ( \4053 , \2851 , \294 );
xnor \U$3865 ( \4054 , \4053 , \301 );
and \U$3866 ( \4055 , \4052 , \4054 );
and \U$3867 ( \4056 , \4048 , \4055 );
and \U$3868 ( \4057 , \2851 , \296 );
and \U$3869 ( \4058 , \2763 , \294 );
nor \U$3870 ( \4059 , \4057 , \4058 );
xnor \U$3871 ( \4060 , \4059 , \301 );
and \U$3872 ( \4061 , \4055 , \4060 );
and \U$3873 ( \4062 , \4048 , \4060 );
or \U$3874 ( \4063 , \4056 , \4061 , \4062 );
and \U$3875 ( \4064 , \4032 , \4063 );
xor \U$3876 ( \4065 , \3864 , \3868 );
xor \U$3877 ( \4066 , \4065 , \3873 );
xor \U$3878 ( \4067 , \3927 , \3931 );
xor \U$3879 ( \4068 , \4067 , \3936 );
and \U$3880 ( \4069 , \4066 , \4068 );
xor \U$3881 ( \4070 , \3897 , \3901 );
xor \U$3882 ( \4071 , \4070 , \3906 );
and \U$3883 ( \4072 , \4068 , \4071 );
and \U$3884 ( \4073 , \4066 , \4071 );
or \U$3885 ( \4074 , \4069 , \4072 , \4073 );
and \U$3886 ( \4075 , \4063 , \4074 );
and \U$3887 ( \4076 , \4032 , \4074 );
or \U$3888 ( \4077 , \4064 , \4075 , \4076 );
xor \U$3889 ( \4078 , \3876 , \3892 );
xor \U$3890 ( \4079 , \4078 , \3909 );
xor \U$3891 ( \4080 , \3914 , \3916 );
xor \U$3892 ( \4081 , \4080 , \3919 );
and \U$3893 ( \4082 , \4079 , \4081 );
xor \U$3894 ( \4083 , \3939 , \3941 );
xor \U$3895 ( \4084 , \4083 , \3944 );
and \U$3896 ( \4085 , \4081 , \4084 );
and \U$3897 ( \4086 , \4079 , \4084 );
or \U$3898 ( \4087 , \4082 , \4085 , \4086 );
and \U$3899 ( \4088 , \4077 , \4087 );
xor \U$3900 ( \4089 , \3732 , \3746 );
xor \U$3901 ( \4090 , \4089 , \3751 );
and \U$3902 ( \4091 , \4087 , \4090 );
and \U$3903 ( \4092 , \4077 , \4090 );
or \U$3904 ( \4093 , \4088 , \4091 , \4092 );
xor \U$3905 ( \4094 , \3770 , \3782 );
xor \U$3906 ( \4095 , \4094 , \3799 );
xor \U$3907 ( \4096 , \3912 , \3922 );
xor \U$3908 ( \4097 , \4096 , \3947 );
and \U$3909 ( \4098 , \4095 , \4097 );
xor \U$3910 ( \4099 , \3952 , \3954 );
xor \U$3911 ( \4100 , \4099 , \3957 );
and \U$3912 ( \4101 , \4097 , \4100 );
and \U$3913 ( \4102 , \4095 , \4100 );
or \U$3914 ( \4103 , \4098 , \4101 , \4102 );
and \U$3915 ( \4104 , \4093 , \4103 );
xor \U$3916 ( \4105 , \3820 , \3822 );
xor \U$3917 ( \4106 , \4105 , \3825 );
and \U$3918 ( \4107 , \4103 , \4106 );
and \U$3919 ( \4108 , \4093 , \4106 );
or \U$3920 ( \4109 , \4104 , \4107 , \4108 );
xor \U$3921 ( \4110 , \3754 , \3802 );
xor \U$3922 ( \4111 , \4110 , \3815 );
xor \U$3923 ( \4112 , \3950 , \3960 );
xor \U$3924 ( \4113 , \4112 , \3963 );
and \U$3925 ( \4114 , \4111 , \4113 );
and \U$3926 ( \4115 , \4109 , \4114 );
xor \U$3927 ( \4116 , \3966 , \3968 );
xor \U$3928 ( \4117 , \4116 , \3970 );
and \U$3929 ( \4118 , \4114 , \4117 );
and \U$3930 ( \4119 , \4109 , \4117 );
or \U$3931 ( \4120 , \4115 , \4118 , \4119 );
and \U$3932 ( \4121 , \3984 , \4120 );
xor \U$3933 ( \4122 , \3984 , \4120 );
xor \U$3934 ( \4123 , \4109 , \4114 );
xor \U$3935 ( \4124 , \4123 , \4117 );
and \U$3936 ( \4125 , \903 , \1952 );
and \U$3937 ( \4126 , \839 , \1950 );
nor \U$3938 ( \4127 , \4125 , \4126 );
xnor \U$3939 ( \4128 , \4127 , \1832 );
and \U$3940 ( \4129 , \1191 , \1739 );
and \U$3941 ( \4130 , \1102 , \1737 );
nor \U$3942 ( \4131 , \4129 , \4130 );
xnor \U$3943 ( \4132 , \4131 , \1607 );
and \U$3944 ( \4133 , \4128 , \4132 );
and \U$3945 ( \4134 , \1303 , \1474 );
and \U$3946 ( \4135 , \1297 , \1472 );
nor \U$3947 ( \4136 , \4134 , \4135 );
xnor \U$3948 ( \4137 , \4136 , \1360 );
and \U$3949 ( \4138 , \4132 , \4137 );
and \U$3950 ( \4139 , \4128 , \4137 );
or \U$3951 ( \4140 , \4133 , \4138 , \4139 );
and \U$3952 ( \4141 , \1536 , \1277 );
and \U$3953 ( \4142 , \1420 , \1275 );
nor \U$3954 ( \4143 , \4141 , \4142 );
xnor \U$3955 ( \4144 , \4143 , \1173 );
and \U$3956 ( \4145 , \1777 , \1059 );
and \U$3957 ( \4146 , \1768 , \1057 );
nor \U$3958 ( \4147 , \4145 , \4146 );
xnor \U$3959 ( \4148 , \4147 , \981 );
and \U$3960 ( \4149 , \4144 , \4148 );
and \U$3961 ( \4150 , \2027 , \911 );
and \U$3962 ( \4151 , \2021 , \909 );
nor \U$3963 ( \4152 , \4150 , \4151 );
xnor \U$3964 ( \4153 , \4152 , \815 );
and \U$3965 ( \4154 , \4148 , \4153 );
and \U$3966 ( \4155 , \4144 , \4153 );
or \U$3967 ( \4156 , \4149 , \4154 , \4155 );
and \U$3968 ( \4157 , \4140 , \4156 );
and \U$3969 ( \4158 , \494 , \2913 );
and \U$3970 ( \4159 , \444 , \2910 );
nor \U$3971 ( \4160 , \4158 , \4159 );
xnor \U$3972 ( \4161 , \4160 , \2368 );
and \U$3973 ( \4162 , \620 , \2549 );
and \U$3974 ( \4163 , \591 , \2547 );
nor \U$3975 ( \4164 , \4162 , \4163 );
xnor \U$3976 ( \4165 , \4164 , \2371 );
and \U$3977 ( \4166 , \4161 , \4165 );
and \U$3978 ( \4167 , \776 , \2259 );
and \U$3979 ( \4168 , \701 , \2257 );
nor \U$3980 ( \4169 , \4167 , \4168 );
xnor \U$3981 ( \4170 , \4169 , \2121 );
and \U$3982 ( \4171 , \4165 , \4170 );
and \U$3983 ( \4172 , \4161 , \4170 );
or \U$3984 ( \4173 , \4166 , \4171 , \4172 );
and \U$3985 ( \4174 , \4156 , \4173 );
and \U$3986 ( \4175 , \4140 , \4173 );
or \U$3987 ( \4176 , \4157 , \4174 , \4175 );
xor \U$3988 ( \4177 , \3988 , \3992 );
xor \U$3989 ( \4178 , \4177 , \3997 );
xor \U$3990 ( \4179 , \4004 , \4008 );
xor \U$3991 ( \4180 , \4179 , \301 );
and \U$3992 ( \4181 , \4178 , \4180 );
xor \U$3993 ( \4182 , \4017 , \4021 );
xor \U$3994 ( \4183 , \4182 , \4026 );
and \U$3995 ( \4184 , \4180 , \4183 );
and \U$3996 ( \4185 , \4178 , \4183 );
or \U$3997 ( \4186 , \4181 , \4184 , \4185 );
and \U$3998 ( \4187 , \4176 , \4186 );
and \U$3999 ( \4188 , \2304 , \738 );
and \U$4000 ( \4189 , \2159 , \736 );
nor \U$4001 ( \4190 , \4188 , \4189 );
xnor \U$4002 ( \4191 , \4190 , \665 );
and \U$4003 ( \4192 , \2540 , \602 );
and \U$4004 ( \4193 , \2530 , \600 );
nor \U$4005 ( \4194 , \4192 , \4193 );
xnor \U$4006 ( \4195 , \4194 , \558 );
and \U$4007 ( \4196 , \4191 , \4195 );
and \U$4008 ( \4197 , \2851 , \502 );
and \U$4009 ( \4198 , \2763 , \500 );
nor \U$4010 ( \4199 , \4197 , \4198 );
xnor \U$4011 ( \4200 , \4199 , \453 );
and \U$4012 ( \4201 , \4195 , \4200 );
and \U$4013 ( \4202 , \4191 , \4200 );
or \U$4014 ( \4203 , \4196 , \4201 , \4202 );
xor \U$4015 ( \4204 , \4036 , \4040 );
xor \U$4016 ( \4205 , \4204 , \4045 );
and \U$4017 ( \4206 , \4203 , \4205 );
xor \U$4018 ( \4207 , \4052 , \4054 );
and \U$4019 ( \4208 , \4205 , \4207 );
and \U$4020 ( \4209 , \4203 , \4207 );
or \U$4021 ( \4210 , \4206 , \4208 , \4209 );
and \U$4022 ( \4211 , \4186 , \4210 );
and \U$4023 ( \4212 , \4176 , \4210 );
or \U$4024 ( \4213 , \4187 , \4211 , \4212 );
xor \U$4025 ( \4214 , \3880 , \3884 );
xor \U$4026 ( \4215 , \4214 , \3889 );
xor \U$4027 ( \4216 , \4048 , \4055 );
xor \U$4028 ( \4217 , \4216 , \4060 );
and \U$4029 ( \4218 , \4215 , \4217 );
xor \U$4030 ( \4219 , \4066 , \4068 );
xor \U$4031 ( \4220 , \4219 , \4071 );
and \U$4032 ( \4221 , \4217 , \4220 );
and \U$4033 ( \4222 , \4215 , \4220 );
or \U$4034 ( \4223 , \4218 , \4221 , \4222 );
and \U$4035 ( \4224 , \4213 , \4223 );
xor \U$4036 ( \4225 , \4079 , \4081 );
xor \U$4037 ( \4226 , \4225 , \4084 );
and \U$4038 ( \4227 , \4223 , \4226 );
and \U$4039 ( \4228 , \4213 , \4226 );
or \U$4040 ( \4229 , \4224 , \4227 , \4228 );
xor \U$4041 ( \4230 , \4077 , \4087 );
xor \U$4042 ( \4231 , \4230 , \4090 );
and \U$4043 ( \4232 , \4229 , \4231 );
xor \U$4044 ( \4233 , \4095 , \4097 );
xor \U$4045 ( \4234 , \4233 , \4100 );
and \U$4046 ( \4235 , \4231 , \4234 );
and \U$4047 ( \4236 , \4229 , \4234 );
or \U$4048 ( \4237 , \4232 , \4235 , \4236 );
xor \U$4049 ( \4238 , \4093 , \4103 );
xor \U$4050 ( \4239 , \4238 , \4106 );
and \U$4051 ( \4240 , \4237 , \4239 );
xor \U$4052 ( \4241 , \4111 , \4113 );
and \U$4053 ( \4242 , \4239 , \4241 );
and \U$4054 ( \4243 , \4237 , \4241 );
or \U$4055 ( \4244 , \4240 , \4242 , \4243 );
and \U$4056 ( \4245 , \4124 , \4244 );
xor \U$4057 ( \4246 , \4124 , \4244 );
xor \U$4058 ( \4247 , \4237 , \4239 );
xor \U$4059 ( \4248 , \4247 , \4241 );
and \U$4060 ( \4249 , \839 , \2259 );
and \U$4061 ( \4250 , \776 , \2257 );
nor \U$4062 ( \4251 , \4249 , \4250 );
xnor \U$4063 ( \4252 , \4251 , \2121 );
and \U$4064 ( \4253 , \1102 , \1952 );
and \U$4065 ( \4254 , \903 , \1950 );
nor \U$4066 ( \4255 , \4253 , \4254 );
xnor \U$4067 ( \4256 , \4255 , \1832 );
and \U$4068 ( \4257 , \4252 , \4256 );
and \U$4069 ( \4258 , \1297 , \1739 );
and \U$4070 ( \4259 , \1191 , \1737 );
nor \U$4071 ( \4260 , \4258 , \4259 );
xnor \U$4072 ( \4261 , \4260 , \1607 );
and \U$4073 ( \4262 , \4256 , \4261 );
and \U$4074 ( \4263 , \4252 , \4261 );
or \U$4075 ( \4264 , \4257 , \4262 , \4263 );
and \U$4076 ( \4265 , \1420 , \1474 );
and \U$4077 ( \4266 , \1303 , \1472 );
nor \U$4078 ( \4267 , \4265 , \4266 );
xnor \U$4079 ( \4268 , \4267 , \1360 );
and \U$4080 ( \4269 , \1768 , \1277 );
and \U$4081 ( \4270 , \1536 , \1275 );
nor \U$4082 ( \4271 , \4269 , \4270 );
xnor \U$4083 ( \4272 , \4271 , \1173 );
and \U$4084 ( \4273 , \4268 , \4272 );
and \U$4085 ( \4274 , \2021 , \1059 );
and \U$4086 ( \4275 , \1777 , \1057 );
nor \U$4087 ( \4276 , \4274 , \4275 );
xnor \U$4088 ( \4277 , \4276 , \981 );
and \U$4089 ( \4278 , \4272 , \4277 );
and \U$4090 ( \4279 , \4268 , \4277 );
or \U$4091 ( \4280 , \4273 , \4278 , \4279 );
and \U$4092 ( \4281 , \4264 , \4280 );
and \U$4093 ( \4282 , \591 , \2913 );
and \U$4094 ( \4283 , \494 , \2910 );
nor \U$4095 ( \4284 , \4282 , \4283 );
xnor \U$4096 ( \4285 , \4284 , \2368 );
and \U$4097 ( \4286 , \701 , \2549 );
and \U$4098 ( \4287 , \620 , \2547 );
nor \U$4099 ( \4288 , \4286 , \4287 );
xnor \U$4100 ( \4289 , \4288 , \2371 );
and \U$4101 ( \4290 , \4285 , \4289 );
and \U$4102 ( \4291 , \4289 , \453 );
and \U$4103 ( \4292 , \4285 , \453 );
or \U$4104 ( \4293 , \4290 , \4291 , \4292 );
and \U$4105 ( \4294 , \4280 , \4293 );
and \U$4106 ( \4295 , \4264 , \4293 );
or \U$4107 ( \4296 , \4281 , \4294 , \4295 );
and \U$4108 ( \4297 , \2159 , \911 );
and \U$4109 ( \4298 , \2027 , \909 );
nor \U$4110 ( \4299 , \4297 , \4298 );
xnor \U$4111 ( \4300 , \4299 , \815 );
and \U$4112 ( \4301 , \2530 , \738 );
and \U$4113 ( \4302 , \2304 , \736 );
nor \U$4114 ( \4303 , \4301 , \4302 );
xnor \U$4115 ( \4304 , \4303 , \665 );
and \U$4116 ( \4305 , \4300 , \4304 );
and \U$4117 ( \4306 , \2763 , \602 );
and \U$4118 ( \4307 , \2540 , \600 );
nor \U$4119 ( \4308 , \4306 , \4307 );
xnor \U$4120 ( \4309 , \4308 , \558 );
and \U$4121 ( \4310 , \4304 , \4309 );
and \U$4122 ( \4311 , \4300 , \4309 );
or \U$4123 ( \4312 , \4305 , \4310 , \4311 );
xor \U$4124 ( \4313 , \4144 , \4148 );
xor \U$4125 ( \4314 , \4313 , \4153 );
and \U$4126 ( \4315 , \4312 , \4314 );
xor \U$4127 ( \4316 , \4191 , \4195 );
xor \U$4128 ( \4317 , \4316 , \4200 );
and \U$4129 ( \4318 , \4314 , \4317 );
and \U$4130 ( \4319 , \4312 , \4317 );
or \U$4131 ( \4320 , \4315 , \4318 , \4319 );
and \U$4132 ( \4321 , \4296 , \4320 );
xor \U$4133 ( \4322 , \4128 , \4132 );
xor \U$4134 ( \4323 , \4322 , \4137 );
xor \U$4135 ( \4324 , \4161 , \4165 );
xor \U$4136 ( \4325 , \4324 , \4170 );
and \U$4137 ( \4326 , \4323 , \4325 );
and \U$4138 ( \4327 , \4320 , \4326 );
and \U$4139 ( \4328 , \4296 , \4326 );
or \U$4140 ( \4329 , \4321 , \4327 , \4328 );
xor \U$4141 ( \4330 , \4140 , \4156 );
xor \U$4142 ( \4331 , \4330 , \4173 );
xor \U$4143 ( \4332 , \4178 , \4180 );
xor \U$4144 ( \4333 , \4332 , \4183 );
and \U$4145 ( \4334 , \4331 , \4333 );
xor \U$4146 ( \4335 , \4203 , \4205 );
xor \U$4147 ( \4336 , \4335 , \4207 );
and \U$4148 ( \4337 , \4333 , \4336 );
and \U$4149 ( \4338 , \4331 , \4336 );
or \U$4150 ( \4339 , \4334 , \4337 , \4338 );
and \U$4151 ( \4340 , \4329 , \4339 );
xor \U$4152 ( \4341 , \4000 , \4012 );
xor \U$4153 ( \4342 , \4341 , \4029 );
and \U$4154 ( \4343 , \4339 , \4342 );
and \U$4155 ( \4344 , \4329 , \4342 );
or \U$4156 ( \4345 , \4340 , \4343 , \4344 );
xor \U$4157 ( \4346 , \4176 , \4186 );
xor \U$4158 ( \4347 , \4346 , \4210 );
xor \U$4159 ( \4348 , \4215 , \4217 );
xor \U$4160 ( \4349 , \4348 , \4220 );
and \U$4161 ( \4350 , \4347 , \4349 );
and \U$4162 ( \4351 , \4345 , \4350 );
xor \U$4163 ( \4352 , \4032 , \4063 );
xor \U$4164 ( \4353 , \4352 , \4074 );
and \U$4165 ( \4354 , \4350 , \4353 );
and \U$4166 ( \4355 , \4345 , \4353 );
or \U$4167 ( \4356 , \4351 , \4354 , \4355 );
xor \U$4168 ( \4357 , \4229 , \4231 );
xor \U$4169 ( \4358 , \4357 , \4234 );
and \U$4170 ( \4359 , \4356 , \4358 );
and \U$4171 ( \4360 , \4248 , \4359 );
xor \U$4172 ( \4361 , \4248 , \4359 );
xor \U$4173 ( \4362 , \4356 , \4358 );
xor \U$4174 ( \4363 , \4345 , \4350 );
xor \U$4175 ( \4364 , \4363 , \4353 );
xor \U$4176 ( \4365 , \4213 , \4223 );
xor \U$4177 ( \4366 , \4365 , \4226 );
and \U$4178 ( \4367 , \4364 , \4366 );
and \U$4179 ( \4368 , \4362 , \4367 );
xor \U$4180 ( \4369 , \4362 , \4367 );
xor \U$4181 ( \4370 , \4364 , \4366 );
and \U$4182 ( \4371 , \620 , \2913 );
and \U$4183 ( \4372 , \591 , \2910 );
nor \U$4184 ( \4373 , \4371 , \4372 );
xnor \U$4185 ( \4374 , \4373 , \2368 );
and \U$4186 ( \4375 , \776 , \2549 );
and \U$4187 ( \4376 , \701 , \2547 );
nor \U$4188 ( \4377 , \4375 , \4376 );
xnor \U$4189 ( \4378 , \4377 , \2371 );
and \U$4190 ( \4379 , \4374 , \4378 );
and \U$4191 ( \4380 , \903 , \2259 );
and \U$4192 ( \4381 , \839 , \2257 );
nor \U$4193 ( \4382 , \4380 , \4381 );
xnor \U$4194 ( \4383 , \4382 , \2121 );
and \U$4195 ( \4384 , \4378 , \4383 );
and \U$4196 ( \4385 , \4374 , \4383 );
or \U$4197 ( \4386 , \4379 , \4384 , \4385 );
and \U$4198 ( \4387 , \1777 , \1277 );
and \U$4199 ( \4388 , \1768 , \1275 );
nor \U$4200 ( \4389 , \4387 , \4388 );
xnor \U$4201 ( \4390 , \4389 , \1173 );
and \U$4202 ( \4391 , \2027 , \1059 );
and \U$4203 ( \4392 , \2021 , \1057 );
nor \U$4204 ( \4393 , \4391 , \4392 );
xnor \U$4205 ( \4394 , \4393 , \981 );
and \U$4206 ( \4395 , \4390 , \4394 );
and \U$4207 ( \4396 , \2304 , \911 );
and \U$4208 ( \4397 , \2159 , \909 );
nor \U$4209 ( \4398 , \4396 , \4397 );
xnor \U$4210 ( \4399 , \4398 , \815 );
and \U$4211 ( \4400 , \4394 , \4399 );
and \U$4212 ( \4401 , \4390 , \4399 );
or \U$4213 ( \4402 , \4395 , \4400 , \4401 );
and \U$4214 ( \4403 , \4386 , \4402 );
and \U$4215 ( \4404 , \1191 , \1952 );
and \U$4216 ( \4405 , \1102 , \1950 );
nor \U$4217 ( \4406 , \4404 , \4405 );
xnor \U$4218 ( \4407 , \4406 , \1832 );
and \U$4219 ( \4408 , \1303 , \1739 );
and \U$4220 ( \4409 , \1297 , \1737 );
nor \U$4221 ( \4410 , \4408 , \4409 );
xnor \U$4222 ( \4411 , \4410 , \1607 );
and \U$4223 ( \4412 , \4407 , \4411 );
and \U$4224 ( \4413 , \1536 , \1474 );
and \U$4225 ( \4414 , \1420 , \1472 );
nor \U$4226 ( \4415 , \4413 , \4414 );
xnor \U$4227 ( \4416 , \4415 , \1360 );
and \U$4228 ( \4417 , \4411 , \4416 );
and \U$4229 ( \4418 , \4407 , \4416 );
or \U$4230 ( \4419 , \4412 , \4417 , \4418 );
and \U$4231 ( \4420 , \4402 , \4419 );
and \U$4232 ( \4421 , \4386 , \4419 );
or \U$4233 ( \4422 , \4403 , \4420 , \4421 );
nand \U$4234 ( \4423 , \2851 , \500 );
xnor \U$4235 ( \4424 , \4423 , \453 );
xor \U$4236 ( \4425 , \4268 , \4272 );
xor \U$4237 ( \4426 , \4425 , \4277 );
and \U$4238 ( \4427 , \4424 , \4426 );
xor \U$4239 ( \4428 , \4300 , \4304 );
xor \U$4240 ( \4429 , \4428 , \4309 );
and \U$4241 ( \4430 , \4426 , \4429 );
and \U$4242 ( \4431 , \4424 , \4429 );
or \U$4243 ( \4432 , \4427 , \4430 , \4431 );
and \U$4244 ( \4433 , \4422 , \4432 );
xor \U$4245 ( \4434 , \4252 , \4256 );
xor \U$4246 ( \4435 , \4434 , \4261 );
xor \U$4247 ( \4436 , \4285 , \4289 );
xor \U$4248 ( \4437 , \4436 , \453 );
and \U$4249 ( \4438 , \4435 , \4437 );
and \U$4250 ( \4439 , \4432 , \4438 );
and \U$4251 ( \4440 , \4422 , \4438 );
or \U$4252 ( \4441 , \4433 , \4439 , \4440 );
xor \U$4253 ( \4442 , \4264 , \4280 );
xor \U$4254 ( \4443 , \4442 , \4293 );
xor \U$4255 ( \4444 , \4312 , \4314 );
xor \U$4256 ( \4445 , \4444 , \4317 );
and \U$4257 ( \4446 , \4443 , \4445 );
xor \U$4258 ( \4447 , \4323 , \4325 );
and \U$4259 ( \4448 , \4445 , \4447 );
and \U$4260 ( \4449 , \4443 , \4447 );
or \U$4261 ( \4450 , \4446 , \4448 , \4449 );
and \U$4262 ( \4451 , \4441 , \4450 );
xor \U$4263 ( \4452 , \4331 , \4333 );
xor \U$4264 ( \4453 , \4452 , \4336 );
and \U$4265 ( \4454 , \4450 , \4453 );
and \U$4266 ( \4455 , \4441 , \4453 );
or \U$4267 ( \4456 , \4451 , \4454 , \4455 );
xor \U$4268 ( \4457 , \4329 , \4339 );
xor \U$4269 ( \4458 , \4457 , \4342 );
and \U$4270 ( \4459 , \4456 , \4458 );
xor \U$4271 ( \4460 , \4347 , \4349 );
and \U$4272 ( \4461 , \4458 , \4460 );
and \U$4273 ( \4462 , \4456 , \4460 );
or \U$4274 ( \4463 , \4459 , \4461 , \4462 );
and \U$4275 ( \4464 , \4370 , \4463 );
xor \U$4276 ( \4465 , \4370 , \4463 );
xor \U$4277 ( \4466 , \4456 , \4458 );
xor \U$4278 ( \4467 , \4466 , \4460 );
and \U$4279 ( \4468 , \2530 , \911 );
and \U$4280 ( \4469 , \2304 , \909 );
nor \U$4281 ( \4470 , \4468 , \4469 );
xnor \U$4282 ( \4471 , \4470 , \815 );
and \U$4283 ( \4472 , \2763 , \738 );
and \U$4284 ( \4473 , \2540 , \736 );
nor \U$4285 ( \4474 , \4472 , \4473 );
xnor \U$4286 ( \4475 , \4474 , \665 );
and \U$4287 ( \4476 , \4471 , \4475 );
nand \U$4288 ( \4477 , \2851 , \600 );
xnor \U$4289 ( \4478 , \4477 , \558 );
and \U$4290 ( \4479 , \4475 , \4478 );
and \U$4291 ( \4480 , \4471 , \4478 );
or \U$4292 ( \4481 , \4476 , \4479 , \4480 );
and \U$4293 ( \4482 , \2540 , \738 );
and \U$4294 ( \4483 , \2530 , \736 );
nor \U$4295 ( \4484 , \4482 , \4483 );
xnor \U$4296 ( \4485 , \4484 , \665 );
and \U$4297 ( \4486 , \4481 , \4485 );
and \U$4298 ( \4487 , \2851 , \602 );
and \U$4299 ( \4488 , \2763 , \600 );
nor \U$4300 ( \4489 , \4487 , \4488 );
xnor \U$4301 ( \4490 , \4489 , \558 );
and \U$4302 ( \4491 , \4485 , \4490 );
and \U$4303 ( \4492 , \4481 , \4490 );
or \U$4304 ( \4493 , \4486 , \4491 , \4492 );
and \U$4305 ( \4494 , \701 , \2913 );
and \U$4306 ( \4495 , \620 , \2910 );
nor \U$4307 ( \4496 , \4494 , \4495 );
xnor \U$4308 ( \4497 , \4496 , \2368 );
and \U$4309 ( \4498 , \839 , \2549 );
and \U$4310 ( \4499 , \776 , \2547 );
nor \U$4311 ( \4500 , \4498 , \4499 );
xnor \U$4312 ( \4501 , \4500 , \2371 );
and \U$4313 ( \4502 , \4497 , \4501 );
and \U$4314 ( \4503 , \4501 , \558 );
and \U$4315 ( \4504 , \4497 , \558 );
or \U$4316 ( \4505 , \4502 , \4503 , \4504 );
and \U$4317 ( \4506 , \1102 , \2259 );
and \U$4318 ( \4507 , \903 , \2257 );
nor \U$4319 ( \4508 , \4506 , \4507 );
xnor \U$4320 ( \4509 , \4508 , \2121 );
and \U$4321 ( \4510 , \1297 , \1952 );
and \U$4322 ( \4511 , \1191 , \1950 );
nor \U$4323 ( \4512 , \4510 , \4511 );
xnor \U$4324 ( \4513 , \4512 , \1832 );
and \U$4325 ( \4514 , \4509 , \4513 );
and \U$4326 ( \4515 , \1420 , \1739 );
and \U$4327 ( \4516 , \1303 , \1737 );
nor \U$4328 ( \4517 , \4515 , \4516 );
xnor \U$4329 ( \4518 , \4517 , \1607 );
and \U$4330 ( \4519 , \4513 , \4518 );
and \U$4331 ( \4520 , \4509 , \4518 );
or \U$4332 ( \4521 , \4514 , \4519 , \4520 );
and \U$4333 ( \4522 , \4505 , \4521 );
and \U$4334 ( \4523 , \1768 , \1474 );
and \U$4335 ( \4524 , \1536 , \1472 );
nor \U$4336 ( \4525 , \4523 , \4524 );
xnor \U$4337 ( \4526 , \4525 , \1360 );
and \U$4338 ( \4527 , \2021 , \1277 );
and \U$4339 ( \4528 , \1777 , \1275 );
nor \U$4340 ( \4529 , \4527 , \4528 );
xnor \U$4341 ( \4530 , \4529 , \1173 );
and \U$4342 ( \4531 , \4526 , \4530 );
and \U$4343 ( \4532 , \2159 , \1059 );
and \U$4344 ( \4533 , \2027 , \1057 );
nor \U$4345 ( \4534 , \4532 , \4533 );
xnor \U$4346 ( \4535 , \4534 , \981 );
and \U$4347 ( \4536 , \4530 , \4535 );
and \U$4348 ( \4537 , \4526 , \4535 );
or \U$4349 ( \4538 , \4531 , \4536 , \4537 );
and \U$4350 ( \4539 , \4521 , \4538 );
and \U$4351 ( \4540 , \4505 , \4538 );
or \U$4352 ( \4541 , \4522 , \4539 , \4540 );
and \U$4353 ( \4542 , \4493 , \4541 );
xor \U$4354 ( \4543 , \4374 , \4378 );
xor \U$4355 ( \4544 , \4543 , \4383 );
xor \U$4356 ( \4545 , \4390 , \4394 );
xor \U$4357 ( \4546 , \4545 , \4399 );
and \U$4358 ( \4547 , \4544 , \4546 );
xor \U$4359 ( \4548 , \4407 , \4411 );
xor \U$4360 ( \4549 , \4548 , \4416 );
and \U$4361 ( \4550 , \4546 , \4549 );
and \U$4362 ( \4551 , \4544 , \4549 );
or \U$4363 ( \4552 , \4547 , \4550 , \4551 );
and \U$4364 ( \4553 , \4541 , \4552 );
and \U$4365 ( \4554 , \4493 , \4552 );
or \U$4366 ( \4555 , \4542 , \4553 , \4554 );
xor \U$4367 ( \4556 , \4386 , \4402 );
xor \U$4368 ( \4557 , \4556 , \4419 );
xor \U$4369 ( \4558 , \4424 , \4426 );
xor \U$4370 ( \4559 , \4558 , \4429 );
and \U$4371 ( \4560 , \4557 , \4559 );
xor \U$4372 ( \4561 , \4435 , \4437 );
and \U$4373 ( \4562 , \4559 , \4561 );
and \U$4374 ( \4563 , \4557 , \4561 );
or \U$4375 ( \4564 , \4560 , \4562 , \4563 );
and \U$4376 ( \4565 , \4555 , \4564 );
xor \U$4377 ( \4566 , \4443 , \4445 );
xor \U$4378 ( \4567 , \4566 , \4447 );
and \U$4379 ( \4568 , \4564 , \4567 );
and \U$4380 ( \4569 , \4555 , \4567 );
or \U$4381 ( \4570 , \4565 , \4568 , \4569 );
xor \U$4382 ( \4571 , \4296 , \4320 );
xor \U$4383 ( \4572 , \4571 , \4326 );
and \U$4384 ( \4573 , \4570 , \4572 );
xor \U$4385 ( \4574 , \4441 , \4450 );
xor \U$4386 ( \4575 , \4574 , \4453 );
and \U$4387 ( \4576 , \4572 , \4575 );
and \U$4388 ( \4577 , \4570 , \4575 );
or \U$4389 ( \4578 , \4573 , \4576 , \4577 );
and \U$4390 ( \4579 , \4467 , \4578 );
xor \U$4391 ( \4580 , \4467 , \4578 );
xor \U$4392 ( \4581 , \4570 , \4572 );
xor \U$4393 ( \4582 , \4581 , \4575 );
and \U$4394 ( \4583 , \2027 , \1277 );
and \U$4395 ( \4584 , \2021 , \1275 );
nor \U$4396 ( \4585 , \4583 , \4584 );
xnor \U$4397 ( \4586 , \4585 , \1173 );
and \U$4398 ( \4587 , \2304 , \1059 );
and \U$4399 ( \4588 , \2159 , \1057 );
nor \U$4400 ( \4589 , \4587 , \4588 );
xnor \U$4401 ( \4590 , \4589 , \981 );
and \U$4402 ( \4591 , \4586 , \4590 );
and \U$4403 ( \4592 , \2540 , \911 );
and \U$4404 ( \4593 , \2530 , \909 );
nor \U$4405 ( \4594 , \4592 , \4593 );
xnor \U$4406 ( \4595 , \4594 , \815 );
and \U$4407 ( \4596 , \4590 , \4595 );
and \U$4408 ( \4597 , \4586 , \4595 );
or \U$4409 ( \4598 , \4591 , \4596 , \4597 );
and \U$4410 ( \4599 , \776 , \2913 );
and \U$4411 ( \4600 , \701 , \2910 );
nor \U$4412 ( \4601 , \4599 , \4600 );
xnor \U$4413 ( \4602 , \4601 , \2368 );
and \U$4414 ( \4603 , \903 , \2549 );
and \U$4415 ( \4604 , \839 , \2547 );
nor \U$4416 ( \4605 , \4603 , \4604 );
xnor \U$4417 ( \4606 , \4605 , \2371 );
and \U$4418 ( \4607 , \4602 , \4606 );
and \U$4419 ( \4608 , \1191 , \2259 );
and \U$4420 ( \4609 , \1102 , \2257 );
nor \U$4421 ( \4610 , \4608 , \4609 );
xnor \U$4422 ( \4611 , \4610 , \2121 );
and \U$4423 ( \4612 , \4606 , \4611 );
and \U$4424 ( \4613 , \4602 , \4611 );
or \U$4425 ( \4614 , \4607 , \4612 , \4613 );
and \U$4426 ( \4615 , \4598 , \4614 );
and \U$4427 ( \4616 , \1303 , \1952 );
and \U$4428 ( \4617 , \1297 , \1950 );
nor \U$4429 ( \4618 , \4616 , \4617 );
xnor \U$4430 ( \4619 , \4618 , \1832 );
and \U$4431 ( \4620 , \1536 , \1739 );
and \U$4432 ( \4621 , \1420 , \1737 );
nor \U$4433 ( \4622 , \4620 , \4621 );
xnor \U$4434 ( \4623 , \4622 , \1607 );
and \U$4435 ( \4624 , \4619 , \4623 );
and \U$4436 ( \4625 , \1777 , \1474 );
and \U$4437 ( \4626 , \1768 , \1472 );
nor \U$4438 ( \4627 , \4625 , \4626 );
xnor \U$4439 ( \4628 , \4627 , \1360 );
and \U$4440 ( \4629 , \4623 , \4628 );
and \U$4441 ( \4630 , \4619 , \4628 );
or \U$4442 ( \4631 , \4624 , \4629 , \4630 );
and \U$4443 ( \4632 , \4614 , \4631 );
and \U$4444 ( \4633 , \4598 , \4631 );
or \U$4445 ( \4634 , \4615 , \4632 , \4633 );
xor \U$4446 ( \4635 , \4509 , \4513 );
xor \U$4447 ( \4636 , \4635 , \4518 );
xor \U$4448 ( \4637 , \4471 , \4475 );
xor \U$4449 ( \4638 , \4637 , \4478 );
and \U$4450 ( \4639 , \4636 , \4638 );
xor \U$4451 ( \4640 , \4526 , \4530 );
xor \U$4452 ( \4641 , \4640 , \4535 );
and \U$4453 ( \4642 , \4638 , \4641 );
and \U$4454 ( \4643 , \4636 , \4641 );
or \U$4455 ( \4644 , \4639 , \4642 , \4643 );
and \U$4456 ( \4645 , \4634 , \4644 );
xor \U$4457 ( \4646 , \4544 , \4546 );
xor \U$4458 ( \4647 , \4646 , \4549 );
and \U$4459 ( \4648 , \4644 , \4647 );
and \U$4460 ( \4649 , \4634 , \4647 );
or \U$4461 ( \4650 , \4645 , \4648 , \4649 );
xor \U$4462 ( \4651 , \4493 , \4541 );
xor \U$4463 ( \4652 , \4651 , \4552 );
and \U$4464 ( \4653 , \4650 , \4652 );
xor \U$4465 ( \4654 , \4557 , \4559 );
xor \U$4466 ( \4655 , \4654 , \4561 );
and \U$4467 ( \4656 , \4652 , \4655 );
and \U$4468 ( \4657 , \4650 , \4655 );
or \U$4469 ( \4658 , \4653 , \4656 , \4657 );
xor \U$4470 ( \4659 , \4422 , \4432 );
xor \U$4471 ( \4660 , \4659 , \4438 );
and \U$4472 ( \4661 , \4658 , \4660 );
xor \U$4473 ( \4662 , \4555 , \4564 );
xor \U$4474 ( \4663 , \4662 , \4567 );
and \U$4475 ( \4664 , \4660 , \4663 );
and \U$4476 ( \4665 , \4658 , \4663 );
or \U$4477 ( \4666 , \4661 , \4664 , \4665 );
and \U$4478 ( \4667 , \4582 , \4666 );
xor \U$4479 ( \4668 , \4582 , \4666 );
xor \U$4480 ( \4669 , \4658 , \4660 );
xor \U$4481 ( \4670 , \4669 , \4663 );
and \U$4482 ( \4671 , \839 , \2913 );
and \U$4483 ( \4672 , \776 , \2910 );
nor \U$4484 ( \4673 , \4671 , \4672 );
xnor \U$4485 ( \4674 , \4673 , \2368 );
and \U$4486 ( \4675 , \1102 , \2549 );
and \U$4487 ( \4676 , \903 , \2547 );
nor \U$4488 ( \4677 , \4675 , \4676 );
xnor \U$4489 ( \4678 , \4677 , \2371 );
and \U$4490 ( \4679 , \4674 , \4678 );
and \U$4491 ( \4680 , \4678 , \665 );
and \U$4492 ( \4681 , \4674 , \665 );
or \U$4493 ( \4682 , \4679 , \4680 , \4681 );
and \U$4494 ( \4683 , \2021 , \1474 );
and \U$4495 ( \4684 , \1777 , \1472 );
nor \U$4496 ( \4685 , \4683 , \4684 );
xnor \U$4497 ( \4686 , \4685 , \1360 );
and \U$4498 ( \4687 , \2159 , \1277 );
and \U$4499 ( \4688 , \2027 , \1275 );
nor \U$4500 ( \4689 , \4687 , \4688 );
xnor \U$4501 ( \4690 , \4689 , \1173 );
and \U$4502 ( \4691 , \4686 , \4690 );
and \U$4503 ( \4692 , \2530 , \1059 );
and \U$4504 ( \4693 , \2304 , \1057 );
nor \U$4505 ( \4694 , \4692 , \4693 );
xnor \U$4506 ( \4695 , \4694 , \981 );
and \U$4507 ( \4696 , \4690 , \4695 );
and \U$4508 ( \4697 , \4686 , \4695 );
or \U$4509 ( \4698 , \4691 , \4696 , \4697 );
and \U$4510 ( \4699 , \4682 , \4698 );
and \U$4511 ( \4700 , \1297 , \2259 );
and \U$4512 ( \4701 , \1191 , \2257 );
nor \U$4513 ( \4702 , \4700 , \4701 );
xnor \U$4514 ( \4703 , \4702 , \2121 );
and \U$4515 ( \4704 , \1420 , \1952 );
and \U$4516 ( \4705 , \1303 , \1950 );
nor \U$4517 ( \4706 , \4704 , \4705 );
xnor \U$4518 ( \4707 , \4706 , \1832 );
and \U$4519 ( \4708 , \4703 , \4707 );
and \U$4520 ( \4709 , \1768 , \1739 );
and \U$4521 ( \4710 , \1536 , \1737 );
nor \U$4522 ( \4711 , \4709 , \4710 );
xnor \U$4523 ( \4712 , \4711 , \1607 );
and \U$4524 ( \4713 , \4707 , \4712 );
and \U$4525 ( \4714 , \4703 , \4712 );
or \U$4526 ( \4715 , \4708 , \4713 , \4714 );
and \U$4527 ( \4716 , \4698 , \4715 );
and \U$4528 ( \4717 , \4682 , \4715 );
or \U$4529 ( \4718 , \4699 , \4716 , \4717 );
and \U$4530 ( \4719 , \2851 , \738 );
and \U$4531 ( \4720 , \2763 , \736 );
nor \U$4532 ( \4721 , \4719 , \4720 );
xnor \U$4533 ( \4722 , \4721 , \665 );
xor \U$4534 ( \4723 , \4586 , \4590 );
xor \U$4535 ( \4724 , \4723 , \4595 );
and \U$4536 ( \4725 , \4722 , \4724 );
xor \U$4537 ( \4726 , \4619 , \4623 );
xor \U$4538 ( \4727 , \4726 , \4628 );
and \U$4539 ( \4728 , \4724 , \4727 );
and \U$4540 ( \4729 , \4722 , \4727 );
or \U$4541 ( \4730 , \4725 , \4728 , \4729 );
and \U$4542 ( \4731 , \4718 , \4730 );
xor \U$4543 ( \4732 , \4497 , \4501 );
xor \U$4544 ( \4733 , \4732 , \558 );
and \U$4545 ( \4734 , \4730 , \4733 );
and \U$4546 ( \4735 , \4718 , \4733 );
or \U$4547 ( \4736 , \4731 , \4734 , \4735 );
xor \U$4548 ( \4737 , \4598 , \4614 );
xor \U$4549 ( \4738 , \4737 , \4631 );
xor \U$4550 ( \4739 , \4636 , \4638 );
xor \U$4551 ( \4740 , \4739 , \4641 );
and \U$4552 ( \4741 , \4738 , \4740 );
and \U$4553 ( \4742 , \4736 , \4741 );
xor \U$4554 ( \4743 , \4481 , \4485 );
xor \U$4555 ( \4744 , \4743 , \4490 );
and \U$4556 ( \4745 , \4741 , \4744 );
and \U$4557 ( \4746 , \4736 , \4744 );
or \U$4558 ( \4747 , \4742 , \4745 , \4746 );
xor \U$4559 ( \4748 , \4505 , \4521 );
xor \U$4560 ( \4749 , \4748 , \4538 );
xor \U$4561 ( \4750 , \4634 , \4644 );
xor \U$4562 ( \4751 , \4750 , \4647 );
and \U$4563 ( \4752 , \4749 , \4751 );
and \U$4564 ( \4753 , \4747 , \4752 );
xor \U$4565 ( \4754 , \4650 , \4652 );
xor \U$4566 ( \4755 , \4754 , \4655 );
and \U$4567 ( \4756 , \4752 , \4755 );
and \U$4568 ( \4757 , \4747 , \4755 );
or \U$4569 ( \4758 , \4753 , \4756 , \4757 );
and \U$4570 ( \4759 , \4670 , \4758 );
xor \U$4571 ( \4760 , \4670 , \4758 );
xor \U$4572 ( \4761 , \4747 , \4752 );
xor \U$4573 ( \4762 , \4761 , \4755 );
and \U$4574 ( \4763 , \1536 , \1952 );
and \U$4575 ( \4764 , \1420 , \1950 );
nor \U$4576 ( \4765 , \4763 , \4764 );
xnor \U$4577 ( \4766 , \4765 , \1832 );
and \U$4578 ( \4767 , \1777 , \1739 );
and \U$4579 ( \4768 , \1768 , \1737 );
nor \U$4580 ( \4769 , \4767 , \4768 );
xnor \U$4581 ( \4770 , \4769 , \1607 );
and \U$4582 ( \4771 , \4766 , \4770 );
and \U$4583 ( \4772 , \2027 , \1474 );
and \U$4584 ( \4773 , \2021 , \1472 );
nor \U$4585 ( \4774 , \4772 , \4773 );
xnor \U$4586 ( \4775 , \4774 , \1360 );
and \U$4587 ( \4776 , \4770 , \4775 );
and \U$4588 ( \4777 , \4766 , \4775 );
or \U$4589 ( \4778 , \4771 , \4776 , \4777 );
and \U$4590 ( \4779 , \903 , \2913 );
and \U$4591 ( \4780 , \839 , \2910 );
nor \U$4592 ( \4781 , \4779 , \4780 );
xnor \U$4593 ( \4782 , \4781 , \2368 );
and \U$4594 ( \4783 , \1191 , \2549 );
and \U$4595 ( \4784 , \1102 , \2547 );
nor \U$4596 ( \4785 , \4783 , \4784 );
xnor \U$4597 ( \4786 , \4785 , \2371 );
and \U$4598 ( \4787 , \4782 , \4786 );
and \U$4599 ( \4788 , \1303 , \2259 );
and \U$4600 ( \4789 , \1297 , \2257 );
nor \U$4601 ( \4790 , \4788 , \4789 );
xnor \U$4602 ( \4791 , \4790 , \2121 );
and \U$4603 ( \4792 , \4786 , \4791 );
and \U$4604 ( \4793 , \4782 , \4791 );
or \U$4605 ( \4794 , \4787 , \4792 , \4793 );
and \U$4606 ( \4795 , \4778 , \4794 );
and \U$4607 ( \4796 , \2304 , \1277 );
and \U$4608 ( \4797 , \2159 , \1275 );
nor \U$4609 ( \4798 , \4796 , \4797 );
xnor \U$4610 ( \4799 , \4798 , \1173 );
and \U$4611 ( \4800 , \2540 , \1059 );
and \U$4612 ( \4801 , \2530 , \1057 );
nor \U$4613 ( \4802 , \4800 , \4801 );
xnor \U$4614 ( \4803 , \4802 , \981 );
and \U$4615 ( \4804 , \4799 , \4803 );
and \U$4616 ( \4805 , \2851 , \911 );
and \U$4617 ( \4806 , \2763 , \909 );
nor \U$4618 ( \4807 , \4805 , \4806 );
xnor \U$4619 ( \4808 , \4807 , \815 );
and \U$4620 ( \4809 , \4803 , \4808 );
and \U$4621 ( \4810 , \4799 , \4808 );
or \U$4622 ( \4811 , \4804 , \4809 , \4810 );
and \U$4623 ( \4812 , \4794 , \4811 );
and \U$4624 ( \4813 , \4778 , \4811 );
or \U$4625 ( \4814 , \4795 , \4812 , \4813 );
and \U$4626 ( \4815 , \2763 , \911 );
and \U$4627 ( \4816 , \2540 , \909 );
nor \U$4628 ( \4817 , \4815 , \4816 );
xnor \U$4629 ( \4818 , \4817 , \815 );
nand \U$4630 ( \4819 , \2851 , \736 );
xnor \U$4631 ( \4820 , \4819 , \665 );
and \U$4632 ( \4821 , \4818 , \4820 );
xor \U$4633 ( \4822 , \4686 , \4690 );
xor \U$4634 ( \4823 , \4822 , \4695 );
and \U$4635 ( \4824 , \4820 , \4823 );
and \U$4636 ( \4825 , \4818 , \4823 );
or \U$4637 ( \4826 , \4821 , \4824 , \4825 );
and \U$4638 ( \4827 , \4814 , \4826 );
xor \U$4639 ( \4828 , \4602 , \4606 );
xor \U$4640 ( \4829 , \4828 , \4611 );
and \U$4641 ( \4830 , \4826 , \4829 );
and \U$4642 ( \4831 , \4814 , \4829 );
or \U$4643 ( \4832 , \4827 , \4830 , \4831 );
xor \U$4644 ( \4833 , \4718 , \4730 );
xor \U$4645 ( \4834 , \4833 , \4733 );
and \U$4646 ( \4835 , \4832 , \4834 );
xor \U$4647 ( \4836 , \4738 , \4740 );
and \U$4648 ( \4837 , \4834 , \4836 );
and \U$4649 ( \4838 , \4832 , \4836 );
or \U$4650 ( \4839 , \4835 , \4837 , \4838 );
xor \U$4651 ( \4840 , \4736 , \4741 );
xor \U$4652 ( \4841 , \4840 , \4744 );
and \U$4653 ( \4842 , \4839 , \4841 );
xor \U$4654 ( \4843 , \4749 , \4751 );
and \U$4655 ( \4844 , \4841 , \4843 );
and \U$4656 ( \4845 , \4839 , \4843 );
or \U$4657 ( \4846 , \4842 , \4844 , \4845 );
and \U$4658 ( \4847 , \4762 , \4846 );
xor \U$4659 ( \4848 , \4762 , \4846 );
xor \U$4660 ( \4849 , \4839 , \4841 );
xor \U$4661 ( \4850 , \4849 , \4843 );
and \U$4662 ( \4851 , \1420 , \2259 );
and \U$4663 ( \4852 , \1303 , \2257 );
nor \U$4664 ( \4853 , \4851 , \4852 );
xnor \U$4665 ( \4854 , \4853 , \2121 );
and \U$4666 ( \4855 , \1768 , \1952 );
and \U$4667 ( \4856 , \1536 , \1950 );
nor \U$4668 ( \4857 , \4855 , \4856 );
xnor \U$4669 ( \4858 , \4857 , \1832 );
and \U$4670 ( \4859 , \4854 , \4858 );
and \U$4671 ( \4860 , \2021 , \1739 );
and \U$4672 ( \4861 , \1777 , \1737 );
nor \U$4673 ( \4862 , \4860 , \4861 );
xnor \U$4674 ( \4863 , \4862 , \1607 );
and \U$4675 ( \4864 , \4858 , \4863 );
and \U$4676 ( \4865 , \4854 , \4863 );
or \U$4677 ( \4866 , \4859 , \4864 , \4865 );
and \U$4678 ( \4867 , \1102 , \2913 );
and \U$4679 ( \4868 , \903 , \2910 );
nor \U$4680 ( \4869 , \4867 , \4868 );
xnor \U$4681 ( \4870 , \4869 , \2368 );
and \U$4682 ( \4871 , \1297 , \2549 );
and \U$4683 ( \4872 , \1191 , \2547 );
nor \U$4684 ( \4873 , \4871 , \4872 );
xnor \U$4685 ( \4874 , \4873 , \2371 );
and \U$4686 ( \4875 , \4870 , \4874 );
and \U$4687 ( \4876 , \4874 , \815 );
and \U$4688 ( \4877 , \4870 , \815 );
or \U$4689 ( \4878 , \4875 , \4876 , \4877 );
and \U$4690 ( \4879 , \4866 , \4878 );
and \U$4691 ( \4880 , \2159 , \1474 );
and \U$4692 ( \4881 , \2027 , \1472 );
nor \U$4693 ( \4882 , \4880 , \4881 );
xnor \U$4694 ( \4883 , \4882 , \1360 );
and \U$4695 ( \4884 , \2530 , \1277 );
and \U$4696 ( \4885 , \2304 , \1275 );
nor \U$4697 ( \4886 , \4884 , \4885 );
xnor \U$4698 ( \4887 , \4886 , \1173 );
and \U$4699 ( \4888 , \4883 , \4887 );
and \U$4700 ( \4889 , \2763 , \1059 );
and \U$4701 ( \4890 , \2540 , \1057 );
nor \U$4702 ( \4891 , \4889 , \4890 );
xnor \U$4703 ( \4892 , \4891 , \981 );
and \U$4704 ( \4893 , \4887 , \4892 );
and \U$4705 ( \4894 , \4883 , \4892 );
or \U$4706 ( \4895 , \4888 , \4893 , \4894 );
and \U$4707 ( \4896 , \4878 , \4895 );
and \U$4708 ( \4897 , \4866 , \4895 );
or \U$4709 ( \4898 , \4879 , \4896 , \4897 );
xor \U$4710 ( \4899 , \4766 , \4770 );
xor \U$4711 ( \4900 , \4899 , \4775 );
xor \U$4712 ( \4901 , \4782 , \4786 );
xor \U$4713 ( \4902 , \4901 , \4791 );
and \U$4714 ( \4903 , \4900 , \4902 );
xor \U$4715 ( \4904 , \4799 , \4803 );
xor \U$4716 ( \4905 , \4904 , \4808 );
and \U$4717 ( \4906 , \4902 , \4905 );
and \U$4718 ( \4907 , \4900 , \4905 );
or \U$4719 ( \4908 , \4903 , \4906 , \4907 );
and \U$4720 ( \4909 , \4898 , \4908 );
xor \U$4721 ( \4910 , \4703 , \4707 );
xor \U$4722 ( \4911 , \4910 , \4712 );
and \U$4723 ( \4912 , \4908 , \4911 );
and \U$4724 ( \4913 , \4898 , \4911 );
or \U$4725 ( \4914 , \4909 , \4912 , \4913 );
xor \U$4726 ( \4915 , \4674 , \4678 );
xor \U$4727 ( \4916 , \4915 , \665 );
xor \U$4728 ( \4917 , \4778 , \4794 );
xor \U$4729 ( \4918 , \4917 , \4811 );
and \U$4730 ( \4919 , \4916 , \4918 );
xor \U$4731 ( \4920 , \4818 , \4820 );
xor \U$4732 ( \4921 , \4920 , \4823 );
and \U$4733 ( \4922 , \4918 , \4921 );
and \U$4734 ( \4923 , \4916 , \4921 );
or \U$4735 ( \4924 , \4919 , \4922 , \4923 );
and \U$4736 ( \4925 , \4914 , \4924 );
xor \U$4737 ( \4926 , \4722 , \4724 );
xor \U$4738 ( \4927 , \4926 , \4727 );
and \U$4739 ( \4928 , \4924 , \4927 );
and \U$4740 ( \4929 , \4914 , \4927 );
or \U$4741 ( \4930 , \4925 , \4928 , \4929 );
xor \U$4742 ( \4931 , \4682 , \4698 );
xor \U$4743 ( \4932 , \4931 , \4715 );
xor \U$4744 ( \4933 , \4814 , \4826 );
xor \U$4745 ( \4934 , \4933 , \4829 );
and \U$4746 ( \4935 , \4932 , \4934 );
and \U$4747 ( \4936 , \4930 , \4935 );
xor \U$4748 ( \4937 , \4832 , \4834 );
xor \U$4749 ( \4938 , \4937 , \4836 );
and \U$4750 ( \4939 , \4935 , \4938 );
and \U$4751 ( \4940 , \4930 , \4938 );
or \U$4752 ( \4941 , \4936 , \4939 , \4940 );
and \U$4753 ( \4942 , \4850 , \4941 );
xor \U$4754 ( \4943 , \4850 , \4941 );
xor \U$4755 ( \4944 , \4930 , \4935 );
xor \U$4756 ( \4945 , \4944 , \4938 );
and \U$4757 ( \4946 , \1191 , \2913 );
and \U$4758 ( \4947 , \1102 , \2910 );
nor \U$4759 ( \4948 , \4946 , \4947 );
xnor \U$4760 ( \4949 , \4948 , \2368 );
and \U$4761 ( \4950 , \1303 , \2549 );
and \U$4762 ( \4951 , \1297 , \2547 );
nor \U$4763 ( \4952 , \4950 , \4951 );
xnor \U$4764 ( \4953 , \4952 , \2371 );
and \U$4765 ( \4954 , \4949 , \4953 );
and \U$4766 ( \4955 , \1536 , \2259 );
and \U$4767 ( \4956 , \1420 , \2257 );
nor \U$4768 ( \4957 , \4955 , \4956 );
xnor \U$4769 ( \4958 , \4957 , \2121 );
and \U$4770 ( \4959 , \4953 , \4958 );
and \U$4771 ( \4960 , \4949 , \4958 );
or \U$4772 ( \4961 , \4954 , \4959 , \4960 );
and \U$4773 ( \4962 , \1777 , \1952 );
and \U$4774 ( \4963 , \1768 , \1950 );
nor \U$4775 ( \4964 , \4962 , \4963 );
xnor \U$4776 ( \4965 , \4964 , \1832 );
and \U$4777 ( \4966 , \2027 , \1739 );
and \U$4778 ( \4967 , \2021 , \1737 );
nor \U$4779 ( \4968 , \4966 , \4967 );
xnor \U$4780 ( \4969 , \4968 , \1607 );
and \U$4781 ( \4970 , \4965 , \4969 );
and \U$4782 ( \4971 , \2304 , \1474 );
and \U$4783 ( \4972 , \2159 , \1472 );
nor \U$4784 ( \4973 , \4971 , \4972 );
xnor \U$4785 ( \4974 , \4973 , \1360 );
and \U$4786 ( \4975 , \4969 , \4974 );
and \U$4787 ( \4976 , \4965 , \4974 );
or \U$4788 ( \4977 , \4970 , \4975 , \4976 );
and \U$4789 ( \4978 , \4961 , \4977 );
and \U$4790 ( \4979 , \2540 , \1277 );
and \U$4791 ( \4980 , \2530 , \1275 );
nor \U$4792 ( \4981 , \4979 , \4980 );
xnor \U$4793 ( \4982 , \4981 , \1173 );
and \U$4794 ( \4983 , \2851 , \1059 );
and \U$4795 ( \4984 , \2763 , \1057 );
nor \U$4796 ( \4985 , \4983 , \4984 );
xnor \U$4797 ( \4986 , \4985 , \981 );
and \U$4798 ( \4987 , \4982 , \4986 );
and \U$4799 ( \4988 , \4977 , \4987 );
and \U$4800 ( \4989 , \4961 , \4987 );
or \U$4801 ( \4990 , \4978 , \4988 , \4989 );
nand \U$4802 ( \4991 , \2851 , \909 );
xnor \U$4803 ( \4992 , \4991 , \815 );
xor \U$4804 ( \4993 , \4854 , \4858 );
xor \U$4805 ( \4994 , \4993 , \4863 );
and \U$4806 ( \4995 , \4992 , \4994 );
xor \U$4807 ( \4996 , \4883 , \4887 );
xor \U$4808 ( \4997 , \4996 , \4892 );
and \U$4809 ( \4998 , \4994 , \4997 );
and \U$4810 ( \4999 , \4992 , \4997 );
or \U$4811 ( \5000 , \4995 , \4998 , \4999 );
and \U$4812 ( \5001 , \4990 , \5000 );
xor \U$4813 ( \5002 , \4900 , \4902 );
xor \U$4814 ( \5003 , \5002 , \4905 );
and \U$4815 ( \5004 , \5000 , \5003 );
and \U$4816 ( \5005 , \4990 , \5003 );
or \U$4817 ( \5006 , \5001 , \5004 , \5005 );
xor \U$4818 ( \5007 , \4898 , \4908 );
xor \U$4819 ( \5008 , \5007 , \4911 );
and \U$4820 ( \5009 , \5006 , \5008 );
xor \U$4821 ( \5010 , \4916 , \4918 );
xor \U$4822 ( \5011 , \5010 , \4921 );
and \U$4823 ( \5012 , \5008 , \5011 );
and \U$4824 ( \5013 , \5006 , \5011 );
or \U$4825 ( \5014 , \5009 , \5012 , \5013 );
xor \U$4826 ( \5015 , \4914 , \4924 );
xor \U$4827 ( \5016 , \5015 , \4927 );
and \U$4828 ( \5017 , \5014 , \5016 );
xor \U$4829 ( \5018 , \4932 , \4934 );
and \U$4830 ( \5019 , \5016 , \5018 );
and \U$4831 ( \5020 , \5014 , \5018 );
or \U$4832 ( \5021 , \5017 , \5019 , \5020 );
and \U$4833 ( \5022 , \4945 , \5021 );
xor \U$4834 ( \5023 , \4945 , \5021 );
xor \U$4835 ( \5024 , \5014 , \5016 );
xor \U$4836 ( \5025 , \5024 , \5018 );
and \U$4837 ( \5026 , \2530 , \1474 );
and \U$4838 ( \5027 , \2304 , \1472 );
nor \U$4839 ( \5028 , \5026 , \5027 );
xnor \U$4840 ( \5029 , \5028 , \1360 );
and \U$4841 ( \5030 , \2763 , \1277 );
and \U$4842 ( \5031 , \2540 , \1275 );
nor \U$4843 ( \5032 , \5030 , \5031 );
xnor \U$4844 ( \5033 , \5032 , \1173 );
and \U$4845 ( \5034 , \5029 , \5033 );
nand \U$4846 ( \5035 , \2851 , \1057 );
xnor \U$4847 ( \5036 , \5035 , \981 );
and \U$4848 ( \5037 , \5033 , \5036 );
and \U$4849 ( \5038 , \5029 , \5036 );
or \U$4850 ( \5039 , \5034 , \5037 , \5038 );
and \U$4851 ( \5040 , \1297 , \2913 );
and \U$4852 ( \5041 , \1191 , \2910 );
nor \U$4853 ( \5042 , \5040 , \5041 );
xnor \U$4854 ( \5043 , \5042 , \2368 );
and \U$4855 ( \5044 , \1420 , \2549 );
and \U$4856 ( \5045 , \1303 , \2547 );
nor \U$4857 ( \5046 , \5044 , \5045 );
xnor \U$4858 ( \5047 , \5046 , \2371 );
and \U$4859 ( \5048 , \5043 , \5047 );
and \U$4860 ( \5049 , \5047 , \981 );
and \U$4861 ( \5050 , \5043 , \981 );
or \U$4862 ( \5051 , \5048 , \5049 , \5050 );
and \U$4863 ( \5052 , \5039 , \5051 );
and \U$4864 ( \5053 , \1768 , \2259 );
and \U$4865 ( \5054 , \1536 , \2257 );
nor \U$4866 ( \5055 , \5053 , \5054 );
xnor \U$4867 ( \5056 , \5055 , \2121 );
and \U$4868 ( \5057 , \2021 , \1952 );
and \U$4869 ( \5058 , \1777 , \1950 );
nor \U$4870 ( \5059 , \5057 , \5058 );
xnor \U$4871 ( \5060 , \5059 , \1832 );
and \U$4872 ( \5061 , \5056 , \5060 );
and \U$4873 ( \5062 , \2159 , \1739 );
and \U$4874 ( \5063 , \2027 , \1737 );
nor \U$4875 ( \5064 , \5062 , \5063 );
xnor \U$4876 ( \5065 , \5064 , \1607 );
and \U$4877 ( \5066 , \5060 , \5065 );
and \U$4878 ( \5067 , \5056 , \5065 );
or \U$4879 ( \5068 , \5061 , \5066 , \5067 );
and \U$4880 ( \5069 , \5051 , \5068 );
and \U$4881 ( \5070 , \5039 , \5068 );
or \U$4882 ( \5071 , \5052 , \5069 , \5070 );
xor \U$4883 ( \5072 , \4949 , \4953 );
xor \U$4884 ( \5073 , \5072 , \4958 );
xor \U$4885 ( \5074 , \4965 , \4969 );
xor \U$4886 ( \5075 , \5074 , \4974 );
and \U$4887 ( \5076 , \5073 , \5075 );
xor \U$4888 ( \5077 , \4982 , \4986 );
and \U$4889 ( \5078 , \5075 , \5077 );
and \U$4890 ( \5079 , \5073 , \5077 );
or \U$4891 ( \5080 , \5076 , \5078 , \5079 );
and \U$4892 ( \5081 , \5071 , \5080 );
xor \U$4893 ( \5082 , \4870 , \4874 );
xor \U$4894 ( \5083 , \5082 , \815 );
and \U$4895 ( \5084 , \5080 , \5083 );
and \U$4896 ( \5085 , \5071 , \5083 );
or \U$4897 ( \5086 , \5081 , \5084 , \5085 );
xor \U$4898 ( \5087 , \4961 , \4977 );
xor \U$4899 ( \5088 , \5087 , \4987 );
xor \U$4900 ( \5089 , \4992 , \4994 );
xor \U$4901 ( \5090 , \5089 , \4997 );
and \U$4902 ( \5091 , \5088 , \5090 );
and \U$4903 ( \5092 , \5086 , \5091 );
xor \U$4904 ( \5093 , \4866 , \4878 );
xor \U$4905 ( \5094 , \5093 , \4895 );
and \U$4906 ( \5095 , \5091 , \5094 );
and \U$4907 ( \5096 , \5086 , \5094 );
or \U$4908 ( \5097 , \5092 , \5095 , \5096 );
xor \U$4909 ( \5098 , \5006 , \5008 );
xor \U$4910 ( \5099 , \5098 , \5011 );
and \U$4911 ( \5100 , \5097 , \5099 );
and \U$4912 ( \5101 , \5025 , \5100 );
xor \U$4913 ( \5102 , \5025 , \5100 );
xor \U$4914 ( \5103 , \5097 , \5099 );
xor \U$4915 ( \5104 , \5086 , \5091 );
xor \U$4916 ( \5105 , \5104 , \5094 );
xor \U$4917 ( \5106 , \4990 , \5000 );
xor \U$4918 ( \5107 , \5106 , \5003 );
and \U$4919 ( \5108 , \5105 , \5107 );
and \U$4920 ( \5109 , \5103 , \5108 );
xor \U$4921 ( \5110 , \5103 , \5108 );
xor \U$4922 ( \5111 , \5105 , \5107 );
and \U$4923 ( \5112 , \1303 , \2913 );
and \U$4924 ( \5113 , \1297 , \2910 );
nor \U$4925 ( \5114 , \5112 , \5113 );
xnor \U$4926 ( \5115 , \5114 , \2368 );
and \U$4927 ( \5116 , \1536 , \2549 );
and \U$4928 ( \5117 , \1420 , \2547 );
nor \U$4929 ( \5118 , \5116 , \5117 );
xnor \U$4930 ( \5119 , \5118 , \2371 );
and \U$4931 ( \5120 , \5115 , \5119 );
and \U$4932 ( \5121 , \1777 , \2259 );
and \U$4933 ( \5122 , \1768 , \2257 );
nor \U$4934 ( \5123 , \5121 , \5122 );
xnor \U$4935 ( \5124 , \5123 , \2121 );
and \U$4936 ( \5125 , \5119 , \5124 );
and \U$4937 ( \5126 , \5115 , \5124 );
or \U$4938 ( \5127 , \5120 , \5125 , \5126 );
and \U$4939 ( \5128 , \2027 , \1952 );
and \U$4940 ( \5129 , \2021 , \1950 );
nor \U$4941 ( \5130 , \5128 , \5129 );
xnor \U$4942 ( \5131 , \5130 , \1832 );
and \U$4943 ( \5132 , \2304 , \1739 );
and \U$4944 ( \5133 , \2159 , \1737 );
nor \U$4945 ( \5134 , \5132 , \5133 );
xnor \U$4946 ( \5135 , \5134 , \1607 );
and \U$4947 ( \5136 , \5131 , \5135 );
and \U$4948 ( \5137 , \2540 , \1474 );
and \U$4949 ( \5138 , \2530 , \1472 );
nor \U$4950 ( \5139 , \5137 , \5138 );
xnor \U$4951 ( \5140 , \5139 , \1360 );
and \U$4952 ( \5141 , \5135 , \5140 );
and \U$4953 ( \5142 , \5131 , \5140 );
or \U$4954 ( \5143 , \5136 , \5141 , \5142 );
and \U$4955 ( \5144 , \5127 , \5143 );
xor \U$4956 ( \5145 , \5029 , \5033 );
xor \U$4957 ( \5146 , \5145 , \5036 );
and \U$4958 ( \5147 , \5143 , \5146 );
and \U$4959 ( \5148 , \5127 , \5146 );
or \U$4960 ( \5149 , \5144 , \5147 , \5148 );
xor \U$4961 ( \5150 , \5043 , \5047 );
xor \U$4962 ( \5151 , \5150 , \981 );
xor \U$4963 ( \5152 , \5056 , \5060 );
xor \U$4964 ( \5153 , \5152 , \5065 );
and \U$4965 ( \5154 , \5151 , \5153 );
and \U$4966 ( \5155 , \5149 , \5154 );
xor \U$4967 ( \5156 , \5073 , \5075 );
xor \U$4968 ( \5157 , \5156 , \5077 );
and \U$4969 ( \5158 , \5154 , \5157 );
and \U$4970 ( \5159 , \5149 , \5157 );
or \U$4971 ( \5160 , \5155 , \5158 , \5159 );
xor \U$4972 ( \5161 , \5071 , \5080 );
xor \U$4973 ( \5162 , \5161 , \5083 );
and \U$4974 ( \5163 , \5160 , \5162 );
xor \U$4975 ( \5164 , \5088 , \5090 );
and \U$4976 ( \5165 , \5162 , \5164 );
and \U$4977 ( \5166 , \5160 , \5164 );
or \U$4978 ( \5167 , \5163 , \5165 , \5166 );
and \U$4979 ( \5168 , \5111 , \5167 );
xor \U$4980 ( \5169 , \5111 , \5167 );
xor \U$4981 ( \5170 , \5160 , \5162 );
xor \U$4982 ( \5171 , \5170 , \5164 );
and \U$4983 ( \5172 , \1420 , \2913 );
and \U$4984 ( \5173 , \1303 , \2910 );
nor \U$4985 ( \5174 , \5172 , \5173 );
xnor \U$4986 ( \5175 , \5174 , \2368 );
and \U$4987 ( \5176 , \1768 , \2549 );
and \U$4988 ( \5177 , \1536 , \2547 );
nor \U$4989 ( \5178 , \5176 , \5177 );
xnor \U$4990 ( \5179 , \5178 , \2371 );
and \U$4991 ( \5180 , \5175 , \5179 );
and \U$4992 ( \5181 , \5179 , \1173 );
and \U$4993 ( \5182 , \5175 , \1173 );
or \U$4994 ( \5183 , \5180 , \5181 , \5182 );
and \U$4995 ( \5184 , \2021 , \2259 );
and \U$4996 ( \5185 , \1777 , \2257 );
nor \U$4997 ( \5186 , \5184 , \5185 );
xnor \U$4998 ( \5187 , \5186 , \2121 );
and \U$4999 ( \5188 , \2159 , \1952 );
and \U$5000 ( \5189 , \2027 , \1950 );
nor \U$5001 ( \5190 , \5188 , \5189 );
xnor \U$5002 ( \5191 , \5190 , \1832 );
and \U$5003 ( \5192 , \5187 , \5191 );
and \U$5004 ( \5193 , \2530 , \1739 );
and \U$5005 ( \5194 , \2304 , \1737 );
nor \U$5006 ( \5195 , \5193 , \5194 );
xnor \U$5007 ( \5196 , \5195 , \1607 );
and \U$5008 ( \5197 , \5191 , \5196 );
and \U$5009 ( \5198 , \5187 , \5196 );
or \U$5010 ( \5199 , \5192 , \5197 , \5198 );
and \U$5011 ( \5200 , \5183 , \5199 );
and \U$5012 ( \5201 , \2851 , \1277 );
and \U$5013 ( \5202 , \2763 , \1275 );
nor \U$5014 ( \5203 , \5201 , \5202 );
xnor \U$5015 ( \5204 , \5203 , \1173 );
and \U$5016 ( \5205 , \5199 , \5204 );
and \U$5017 ( \5206 , \5183 , \5204 );
or \U$5018 ( \5207 , \5200 , \5205 , \5206 );
xor \U$5019 ( \5208 , \5127 , \5143 );
xor \U$5020 ( \5209 , \5208 , \5146 );
and \U$5021 ( \5210 , \5207 , \5209 );
xor \U$5022 ( \5211 , \5151 , \5153 );
and \U$5023 ( \5212 , \5209 , \5211 );
and \U$5024 ( \5213 , \5207 , \5211 );
or \U$5025 ( \5214 , \5210 , \5212 , \5213 );
xor \U$5026 ( \5215 , \5039 , \5051 );
xor \U$5027 ( \5216 , \5215 , \5068 );
and \U$5028 ( \5217 , \5214 , \5216 );
xor \U$5029 ( \5218 , \5149 , \5154 );
xor \U$5030 ( \5219 , \5218 , \5157 );
and \U$5031 ( \5220 , \5216 , \5219 );
and \U$5032 ( \5221 , \5214 , \5219 );
or \U$5033 ( \5222 , \5217 , \5220 , \5221 );
and \U$5034 ( \5223 , \5171 , \5222 );
xor \U$5035 ( \5224 , \5171 , \5222 );
xor \U$5036 ( \5225 , \5214 , \5216 );
xor \U$5037 ( \5226 , \5225 , \5219 );
and \U$5038 ( \5227 , \2304 , \1952 );
and \U$5039 ( \5228 , \2159 , \1950 );
nor \U$5040 ( \5229 , \5227 , \5228 );
xnor \U$5041 ( \5230 , \5229 , \1832 );
and \U$5042 ( \5231 , \2540 , \1739 );
and \U$5043 ( \5232 , \2530 , \1737 );
nor \U$5044 ( \5233 , \5231 , \5232 );
xnor \U$5045 ( \5234 , \5233 , \1607 );
and \U$5046 ( \5235 , \5230 , \5234 );
and \U$5047 ( \5236 , \2851 , \1474 );
and \U$5048 ( \5237 , \2763 , \1472 );
nor \U$5049 ( \5238 , \5236 , \5237 );
xnor \U$5050 ( \5239 , \5238 , \1360 );
and \U$5051 ( \5240 , \5234 , \5239 );
and \U$5052 ( \5241 , \5230 , \5239 );
or \U$5053 ( \5242 , \5235 , \5240 , \5241 );
and \U$5054 ( \5243 , \1536 , \2913 );
and \U$5055 ( \5244 , \1420 , \2910 );
nor \U$5056 ( \5245 , \5243 , \5244 );
xnor \U$5057 ( \5246 , \5245 , \2368 );
and \U$5058 ( \5247 , \1777 , \2549 );
and \U$5059 ( \5248 , \1768 , \2547 );
nor \U$5060 ( \5249 , \5247 , \5248 );
xnor \U$5061 ( \5250 , \5249 , \2371 );
and \U$5062 ( \5251 , \5246 , \5250 );
and \U$5063 ( \5252 , \2027 , \2259 );
and \U$5064 ( \5253 , \2021 , \2257 );
nor \U$5065 ( \5254 , \5252 , \5253 );
xnor \U$5066 ( \5255 , \5254 , \2121 );
and \U$5067 ( \5256 , \5250 , \5255 );
and \U$5068 ( \5257 , \5246 , \5255 );
or \U$5069 ( \5258 , \5251 , \5256 , \5257 );
and \U$5070 ( \5259 , \5242 , \5258 );
and \U$5071 ( \5260 , \2763 , \1474 );
and \U$5072 ( \5261 , \2540 , \1472 );
nor \U$5073 ( \5262 , \5260 , \5261 );
xnor \U$5074 ( \5263 , \5262 , \1360 );
and \U$5075 ( \5264 , \5258 , \5263 );
and \U$5076 ( \5265 , \5242 , \5263 );
or \U$5077 ( \5266 , \5259 , \5264 , \5265 );
nand \U$5078 ( \5267 , \2851 , \1275 );
xnor \U$5079 ( \5268 , \5267 , \1173 );
xor \U$5080 ( \5269 , \5175 , \5179 );
xor \U$5081 ( \5270 , \5269 , \1173 );
and \U$5082 ( \5271 , \5268 , \5270 );
xor \U$5083 ( \5272 , \5187 , \5191 );
xor \U$5084 ( \5273 , \5272 , \5196 );
and \U$5085 ( \5274 , \5270 , \5273 );
and \U$5086 ( \5275 , \5268 , \5273 );
or \U$5087 ( \5276 , \5271 , \5274 , \5275 );
and \U$5088 ( \5277 , \5266 , \5276 );
xor \U$5089 ( \5278 , \5131 , \5135 );
xor \U$5090 ( \5279 , \5278 , \5140 );
and \U$5091 ( \5280 , \5276 , \5279 );
and \U$5092 ( \5281 , \5266 , \5279 );
or \U$5093 ( \5282 , \5277 , \5280 , \5281 );
xor \U$5094 ( \5283 , \5115 , \5119 );
xor \U$5095 ( \5284 , \5283 , \5124 );
xor \U$5096 ( \5285 , \5183 , \5199 );
xor \U$5097 ( \5286 , \5285 , \5204 );
and \U$5098 ( \5287 , \5284 , \5286 );
and \U$5099 ( \5288 , \5282 , \5287 );
xor \U$5100 ( \5289 , \5207 , \5209 );
xor \U$5101 ( \5290 , \5289 , \5211 );
and \U$5102 ( \5291 , \5287 , \5290 );
and \U$5103 ( \5292 , \5282 , \5290 );
or \U$5104 ( \5293 , \5288 , \5291 , \5292 );
and \U$5105 ( \5294 , \5226 , \5293 );
xor \U$5106 ( \5295 , \5226 , \5293 );
xor \U$5107 ( \5296 , \5282 , \5287 );
xor \U$5108 ( \5297 , \5296 , \5290 );
and \U$5109 ( \5298 , \2159 , \2259 );
and \U$5110 ( \5299 , \2027 , \2257 );
nor \U$5111 ( \5300 , \5298 , \5299 );
xnor \U$5112 ( \5301 , \5300 , \2121 );
and \U$5113 ( \5302 , \2530 , \1952 );
and \U$5114 ( \5303 , \2304 , \1950 );
nor \U$5115 ( \5304 , \5302 , \5303 );
xnor \U$5116 ( \5305 , \5304 , \1832 );
and \U$5117 ( \5306 , \5301 , \5305 );
and \U$5118 ( \5307 , \2763 , \1739 );
and \U$5119 ( \5308 , \2540 , \1737 );
nor \U$5120 ( \5309 , \5307 , \5308 );
xnor \U$5121 ( \5310 , \5309 , \1607 );
and \U$5122 ( \5311 , \5305 , \5310 );
and \U$5123 ( \5312 , \5301 , \5310 );
or \U$5124 ( \5313 , \5306 , \5311 , \5312 );
and \U$5125 ( \5314 , \1768 , \2913 );
and \U$5126 ( \5315 , \1536 , \2910 );
nor \U$5127 ( \5316 , \5314 , \5315 );
xnor \U$5128 ( \5317 , \5316 , \2368 );
and \U$5129 ( \5318 , \2021 , \2549 );
and \U$5130 ( \5319 , \1777 , \2547 );
nor \U$5131 ( \5320 , \5318 , \5319 );
xnor \U$5132 ( \5321 , \5320 , \2371 );
and \U$5133 ( \5322 , \5317 , \5321 );
and \U$5134 ( \5323 , \5321 , \1360 );
and \U$5135 ( \5324 , \5317 , \1360 );
or \U$5136 ( \5325 , \5322 , \5323 , \5324 );
and \U$5137 ( \5326 , \5313 , \5325 );
xor \U$5138 ( \5327 , \5230 , \5234 );
xor \U$5139 ( \5328 , \5327 , \5239 );
and \U$5140 ( \5329 , \5325 , \5328 );
and \U$5141 ( \5330 , \5313 , \5328 );
or \U$5142 ( \5331 , \5326 , \5329 , \5330 );
xor \U$5143 ( \5332 , \5242 , \5258 );
xor \U$5144 ( \5333 , \5332 , \5263 );
and \U$5145 ( \5334 , \5331 , \5333 );
xor \U$5146 ( \5335 , \5268 , \5270 );
xor \U$5147 ( \5336 , \5335 , \5273 );
and \U$5148 ( \5337 , \5333 , \5336 );
and \U$5149 ( \5338 , \5331 , \5336 );
or \U$5150 ( \5339 , \5334 , \5337 , \5338 );
xor \U$5151 ( \5340 , \5266 , \5276 );
xor \U$5152 ( \5341 , \5340 , \5279 );
and \U$5153 ( \5342 , \5339 , \5341 );
xor \U$5154 ( \5343 , \5284 , \5286 );
and \U$5155 ( \5344 , \5341 , \5343 );
and \U$5156 ( \5345 , \5339 , \5343 );
or \U$5157 ( \5346 , \5342 , \5344 , \5345 );
and \U$5158 ( \5347 , \5297 , \5346 );
xor \U$5159 ( \5348 , \5297 , \5346 );
xor \U$5160 ( \5349 , \5339 , \5341 );
xor \U$5161 ( \5350 , \5349 , \5343 );
and \U$5162 ( \5351 , \1777 , \2913 );
and \U$5163 ( \5352 , \1768 , \2910 );
nor \U$5164 ( \5353 , \5351 , \5352 );
xnor \U$5165 ( \5354 , \5353 , \2368 );
and \U$5166 ( \5355 , \2027 , \2549 );
and \U$5167 ( \5356 , \2021 , \2547 );
nor \U$5168 ( \5357 , \5355 , \5356 );
xnor \U$5169 ( \5358 , \5357 , \2371 );
and \U$5170 ( \5359 , \5354 , \5358 );
and \U$5171 ( \5360 , \2304 , \2259 );
and \U$5172 ( \5361 , \2159 , \2257 );
nor \U$5173 ( \5362 , \5360 , \5361 );
xnor \U$5174 ( \5363 , \5362 , \2121 );
and \U$5175 ( \5364 , \5358 , \5363 );
and \U$5176 ( \5365 , \5354 , \5363 );
or \U$5177 ( \5366 , \5359 , \5364 , \5365 );
nand \U$5178 ( \5367 , \2851 , \1472 );
xnor \U$5179 ( \5368 , \5367 , \1360 );
and \U$5180 ( \5369 , \5366 , \5368 );
xor \U$5181 ( \5370 , \5301 , \5305 );
xor \U$5182 ( \5371 , \5370 , \5310 );
and \U$5183 ( \5372 , \5368 , \5371 );
and \U$5184 ( \5373 , \5366 , \5371 );
or \U$5185 ( \5374 , \5369 , \5372 , \5373 );
xor \U$5186 ( \5375 , \5246 , \5250 );
xor \U$5187 ( \5376 , \5375 , \5255 );
and \U$5188 ( \5377 , \5374 , \5376 );
xor \U$5189 ( \5378 , \5313 , \5325 );
xor \U$5190 ( \5379 , \5378 , \5328 );
and \U$5191 ( \5380 , \5376 , \5379 );
and \U$5192 ( \5381 , \5374 , \5379 );
or \U$5193 ( \5382 , \5377 , \5380 , \5381 );
xor \U$5194 ( \5383 , \5331 , \5333 );
xor \U$5195 ( \5384 , \5383 , \5336 );
and \U$5196 ( \5385 , \5382 , \5384 );
and \U$5197 ( \5386 , \5350 , \5385 );
xor \U$5198 ( \5387 , \5350 , \5385 );
xor \U$5199 ( \5388 , \5382 , \5384 );
and \U$5200 ( \5389 , \2530 , \2259 );
and \U$5201 ( \5390 , \2304 , \2257 );
nor \U$5202 ( \5391 , \5389 , \5390 );
xnor \U$5203 ( \5392 , \5391 , \2121 );
and \U$5204 ( \5393 , \2763 , \1952 );
and \U$5205 ( \5394 , \2540 , \1950 );
nor \U$5206 ( \5395 , \5393 , \5394 );
xnor \U$5207 ( \5396 , \5395 , \1832 );
and \U$5208 ( \5397 , \5392 , \5396 );
nand \U$5209 ( \5398 , \2851 , \1737 );
xnor \U$5210 ( \5399 , \5398 , \1607 );
and \U$5211 ( \5400 , \5396 , \5399 );
and \U$5212 ( \5401 , \5392 , \5399 );
or \U$5213 ( \5402 , \5397 , \5400 , \5401 );
and \U$5214 ( \5403 , \2021 , \2913 );
and \U$5215 ( \5404 , \1777 , \2910 );
nor \U$5216 ( \5405 , \5403 , \5404 );
xnor \U$5217 ( \5406 , \5405 , \2368 );
and \U$5218 ( \5407 , \2159 , \2549 );
and \U$5219 ( \5408 , \2027 , \2547 );
nor \U$5220 ( \5409 , \5407 , \5408 );
xnor \U$5221 ( \5410 , \5409 , \2371 );
and \U$5222 ( \5411 , \5406 , \5410 );
and \U$5223 ( \5412 , \5410 , \1607 );
and \U$5224 ( \5413 , \5406 , \1607 );
or \U$5225 ( \5414 , \5411 , \5412 , \5413 );
and \U$5226 ( \5415 , \5402 , \5414 );
and \U$5227 ( \5416 , \2540 , \1952 );
and \U$5228 ( \5417 , \2530 , \1950 );
nor \U$5229 ( \5418 , \5416 , \5417 );
xnor \U$5230 ( \5419 , \5418 , \1832 );
and \U$5231 ( \5420 , \5414 , \5419 );
and \U$5232 ( \5421 , \5402 , \5419 );
or \U$5233 ( \5422 , \5415 , \5420 , \5421 );
and \U$5234 ( \5423 , \2851 , \1739 );
and \U$5235 ( \5424 , \2763 , \1737 );
nor \U$5236 ( \5425 , \5423 , \5424 );
xnor \U$5237 ( \5426 , \5425 , \1607 );
xor \U$5238 ( \5427 , \5354 , \5358 );
xor \U$5239 ( \5428 , \5427 , \5363 );
and \U$5240 ( \5429 , \5426 , \5428 );
and \U$5241 ( \5430 , \5422 , \5429 );
xor \U$5242 ( \5431 , \5317 , \5321 );
xor \U$5243 ( \5432 , \5431 , \1360 );
and \U$5244 ( \5433 , \5429 , \5432 );
and \U$5245 ( \5434 , \5422 , \5432 );
or \U$5246 ( \5435 , \5430 , \5433 , \5434 );
xor \U$5247 ( \5436 , \5374 , \5376 );
xor \U$5248 ( \5437 , \5436 , \5379 );
and \U$5249 ( \5438 , \5435 , \5437 );
and \U$5250 ( \5439 , \5388 , \5438 );
xor \U$5251 ( \5440 , \5388 , \5438 );
xor \U$5252 ( \5441 , \5435 , \5437 );
xor \U$5253 ( \5442 , \5366 , \5368 );
xor \U$5254 ( \5443 , \5442 , \5371 );
xor \U$5255 ( \5444 , \5422 , \5429 );
xor \U$5256 ( \5445 , \5444 , \5432 );
and \U$5257 ( \5446 , \5443 , \5445 );
and \U$5258 ( \5447 , \5441 , \5446 );
xor \U$5259 ( \5448 , \5441 , \5446 );
xor \U$5260 ( \5449 , \5443 , \5445 );
and \U$5261 ( \5450 , \2027 , \2913 );
and \U$5262 ( \5451 , \2021 , \2910 );
nor \U$5263 ( \5452 , \5450 , \5451 );
xnor \U$5264 ( \5453 , \5452 , \2368 );
and \U$5265 ( \5454 , \2304 , \2549 );
and \U$5266 ( \5455 , \2159 , \2547 );
nor \U$5267 ( \5456 , \5454 , \5455 );
xnor \U$5268 ( \5457 , \5456 , \2371 );
and \U$5269 ( \5458 , \5453 , \5457 );
and \U$5270 ( \5459 , \2540 , \2259 );
and \U$5271 ( \5460 , \2530 , \2257 );
nor \U$5272 ( \5461 , \5459 , \5460 );
xnor \U$5273 ( \5462 , \5461 , \2121 );
and \U$5274 ( \5463 , \5457 , \5462 );
and \U$5275 ( \5464 , \5453 , \5462 );
or \U$5276 ( \5465 , \5458 , \5463 , \5464 );
xor \U$5277 ( \5466 , \5392 , \5396 );
xor \U$5278 ( \5467 , \5466 , \5399 );
and \U$5279 ( \5468 , \5465 , \5467 );
xor \U$5280 ( \5469 , \5406 , \5410 );
xor \U$5281 ( \5470 , \5469 , \1607 );
and \U$5282 ( \5471 , \5467 , \5470 );
and \U$5283 ( \5472 , \5465 , \5470 );
or \U$5284 ( \5473 , \5468 , \5471 , \5472 );
xor \U$5285 ( \5474 , \5402 , \5414 );
xor \U$5286 ( \5475 , \5474 , \5419 );
and \U$5287 ( \5476 , \5473 , \5475 );
xor \U$5288 ( \5477 , \5426 , \5428 );
and \U$5289 ( \5478 , \5475 , \5477 );
and \U$5290 ( \5479 , \5473 , \5477 );
or \U$5291 ( \5480 , \5476 , \5478 , \5479 );
and \U$5292 ( \5481 , \5449 , \5480 );
xor \U$5293 ( \5482 , \5449 , \5480 );
xor \U$5294 ( \5483 , \5473 , \5475 );
xor \U$5295 ( \5484 , \5483 , \5477 );
and \U$5296 ( \5485 , \2159 , \2913 );
and \U$5297 ( \5486 , \2027 , \2910 );
nor \U$5298 ( \5487 , \5485 , \5486 );
xnor \U$5299 ( \5488 , \5487 , \2368 );
and \U$5300 ( \5489 , \2530 , \2549 );
and \U$5301 ( \5490 , \2304 , \2547 );
nor \U$5302 ( \5491 , \5489 , \5490 );
xnor \U$5303 ( \5492 , \5491 , \2371 );
and \U$5304 ( \5493 , \5488 , \5492 );
and \U$5305 ( \5494 , \5492 , \1832 );
and \U$5306 ( \5495 , \5488 , \1832 );
or \U$5307 ( \5496 , \5493 , \5494 , \5495 );
and \U$5308 ( \5497 , \2763 , \2259 );
and \U$5309 ( \5498 , \2540 , \2257 );
nor \U$5310 ( \5499 , \5497 , \5498 );
xnor \U$5311 ( \5500 , \5499 , \2121 );
nand \U$5312 ( \5501 , \2851 , \1950 );
xnor \U$5313 ( \5502 , \5501 , \1832 );
and \U$5314 ( \5503 , \5500 , \5502 );
and \U$5315 ( \5504 , \5496 , \5503 );
and \U$5316 ( \5505 , \2851 , \1952 );
and \U$5317 ( \5506 , \2763 , \1950 );
nor \U$5318 ( \5507 , \5505 , \5506 );
xnor \U$5319 ( \5508 , \5507 , \1832 );
and \U$5320 ( \5509 , \5503 , \5508 );
and \U$5321 ( \5510 , \5496 , \5508 );
or \U$5322 ( \5511 , \5504 , \5509 , \5510 );
xor \U$5323 ( \5512 , \5465 , \5467 );
xor \U$5324 ( \5513 , \5512 , \5470 );
and \U$5325 ( \5514 , \5511 , \5513 );
and \U$5326 ( \5515 , \5484 , \5514 );
xor \U$5327 ( \5516 , \5484 , \5514 );
xor \U$5328 ( \5517 , \5511 , \5513 );
xor \U$5329 ( \5518 , \5453 , \5457 );
xor \U$5330 ( \5519 , \5518 , \5462 );
xor \U$5331 ( \5520 , \5496 , \5503 );
xor \U$5332 ( \5521 , \5520 , \5508 );
and \U$5333 ( \5522 , \5519 , \5521 );
and \U$5334 ( \5523 , \5517 , \5522 );
xor \U$5335 ( \5524 , \5517 , \5522 );
xor \U$5336 ( \5525 , \5519 , \5521 );
and \U$5337 ( \5526 , \2304 , \2913 );
and \U$5338 ( \5527 , \2159 , \2910 );
nor \U$5339 ( \5528 , \5526 , \5527 );
xnor \U$5340 ( \5529 , \5528 , \2368 );
and \U$5341 ( \5530 , \2540 , \2549 );
and \U$5342 ( \5531 , \2530 , \2547 );
nor \U$5343 ( \5532 , \5530 , \5531 );
xnor \U$5344 ( \5533 , \5532 , \2371 );
and \U$5345 ( \5534 , \5529 , \5533 );
and \U$5346 ( \5535 , \2851 , \2259 );
and \U$5347 ( \5536 , \2763 , \2257 );
nor \U$5348 ( \5537 , \5535 , \5536 );
xnor \U$5349 ( \5538 , \5537 , \2121 );
and \U$5350 ( \5539 , \5533 , \5538 );
and \U$5351 ( \5540 , \5529 , \5538 );
or \U$5352 ( \5541 , \5534 , \5539 , \5540 );
xor \U$5353 ( \5542 , \5488 , \5492 );
xor \U$5354 ( \5543 , \5542 , \1832 );
and \U$5355 ( \5544 , \5541 , \5543 );
xor \U$5356 ( \5545 , \5500 , \5502 );
and \U$5357 ( \5546 , \5543 , \5545 );
and \U$5358 ( \5547 , \5541 , \5545 );
or \U$5359 ( \5548 , \5544 , \5546 , \5547 );
and \U$5360 ( \5549 , \5525 , \5548 );
xor \U$5361 ( \5550 , \5525 , \5548 );
xor \U$5362 ( \5551 , \5541 , \5543 );
xor \U$5363 ( \5552 , \5551 , \5545 );
and \U$5364 ( \5553 , \2530 , \2913 );
and \U$5365 ( \5554 , \2304 , \2910 );
nor \U$5366 ( \5555 , \5553 , \5554 );
xnor \U$5367 ( \5556 , \5555 , \2368 );
and \U$5368 ( \5557 , \2763 , \2549 );
and \U$5369 ( \5558 , \2540 , \2547 );
nor \U$5370 ( \5559 , \5557 , \5558 );
xnor \U$5371 ( \5560 , \5559 , \2371 );
and \U$5372 ( \5561 , \5556 , \5560 );
and \U$5373 ( \5562 , \5560 , \2121 );
and \U$5374 ( \5563 , \5556 , \2121 );
or \U$5375 ( \5564 , \5561 , \5562 , \5563 );
xor \U$5376 ( \5565 , \5529 , \5533 );
xor \U$5377 ( \5566 , \5565 , \5538 );
and \U$5378 ( \5567 , \5564 , \5566 );
and \U$5379 ( \5568 , \5552 , \5567 );
xor \U$5380 ( \5569 , \5552 , \5567 );
xor \U$5381 ( \5570 , \5564 , \5566 );
nand \U$5382 ( \5571 , \2851 , \2257 );
xnor \U$5383 ( \5572 , \5571 , \2121 );
xor \U$5384 ( \5573 , \5556 , \5560 );
xor \U$5385 ( \5574 , \5573 , \2121 );
and \U$5386 ( \5575 , \5572 , \5574 );
and \U$5387 ( \5576 , \5570 , \5575 );
xor \U$5388 ( \5577 , \5570 , \5575 );
xor \U$5389 ( \5578 , \5572 , \5574 );
and \U$5390 ( \5579 , \2540 , \2913 );
and \U$5391 ( \5580 , \2530 , \2910 );
nor \U$5392 ( \5581 , \5579 , \5580 );
xnor \U$5393 ( \5582 , \5581 , \2368 );
and \U$5394 ( \5583 , \2851 , \2549 );
and \U$5395 ( \5584 , \2763 , \2547 );
nor \U$5396 ( \5585 , \5583 , \5584 );
xnor \U$5397 ( \5586 , \5585 , \2371 );
and \U$5398 ( \5587 , \5582 , \5586 );
and \U$5399 ( \5588 , \5578 , \5587 );
xor \U$5400 ( \5589 , \5578 , \5587 );
xor \U$5401 ( \5590 , \5582 , \5586 );
and \U$5402 ( \5591 , \2763 , \2913 );
and \U$5403 ( \5592 , \2540 , \2910 );
nor \U$5404 ( \5593 , \5591 , \5592 );
xnor \U$5405 ( \5594 , \5593 , \2368 );
and \U$5406 ( \5595 , \5594 , \2371 );
and \U$5407 ( \5596 , \5590 , \5595 );
xor \U$5408 ( \5597 , \5590 , \5595 );
nand \U$5409 ( \5598 , \2851 , \2547 );
xnor \U$5410 ( \5599 , \5598 , \2371 );
xor \U$5411 ( \5600 , \5594 , \2371 );
and \U$5412 ( \5601 , \5599 , \5600 );
xor \U$5413 ( \5602 , \5599 , \5600 );
and \U$5414 ( \5603 , \2851 , \2913 );
and \U$5415 ( \5604 , \2763 , \2910 );
nor \U$5416 ( \5605 , \5603 , \5604 );
xnor \U$5417 ( \5606 , \5605 , \2368 );
nand \U$5418 ( \5607 , \2851 , \2910 );
xnor \U$5419 ( \5608 , \5607 , \2368 );
and \U$5420 ( \5609 , \5608 , \2368 );
and \U$5421 ( \5610 , \5606 , \5609 );
and \U$5422 ( \5611 , \5602 , \5610 );
or \U$5423 ( \5612 , \5601 , \5611 );
and \U$5424 ( \5613 , \5597 , \5612 );
or \U$5425 ( \5614 , \5596 , \5613 );
and \U$5426 ( \5615 , \5589 , \5614 );
or \U$5427 ( \5616 , \5588 , \5615 );
and \U$5428 ( \5617 , \5577 , \5616 );
or \U$5429 ( \5618 , \5576 , \5617 );
and \U$5430 ( \5619 , \5569 , \5618 );
or \U$5431 ( \5620 , \5568 , \5619 );
and \U$5432 ( \5621 , \5550 , \5620 );
or \U$5433 ( \5622 , \5549 , \5621 );
and \U$5434 ( \5623 , \5524 , \5622 );
or \U$5435 ( \5624 , \5523 , \5623 );
and \U$5436 ( \5625 , \5516 , \5624 );
or \U$5437 ( \5626 , \5515 , \5625 );
and \U$5438 ( \5627 , \5482 , \5626 );
or \U$5439 ( \5628 , \5481 , \5627 );
and \U$5440 ( \5629 , \5448 , \5628 );
or \U$5441 ( \5630 , \5447 , \5629 );
and \U$5442 ( \5631 , \5440 , \5630 );
or \U$5443 ( \5632 , \5439 , \5631 );
and \U$5444 ( \5633 , \5387 , \5632 );
or \U$5445 ( \5634 , \5386 , \5633 );
and \U$5446 ( \5635 , \5348 , \5634 );
or \U$5447 ( \5636 , \5347 , \5635 );
and \U$5448 ( \5637 , \5295 , \5636 );
or \U$5449 ( \5638 , \5294 , \5637 );
and \U$5450 ( \5639 , \5224 , \5638 );
or \U$5451 ( \5640 , \5223 , \5639 );
and \U$5452 ( \5641 , \5169 , \5640 );
or \U$5453 ( \5642 , \5168 , \5641 );
and \U$5454 ( \5643 , \5110 , \5642 );
or \U$5455 ( \5644 , \5109 , \5643 );
and \U$5456 ( \5645 , \5102 , \5644 );
or \U$5457 ( \5646 , \5101 , \5645 );
and \U$5458 ( \5647 , \5023 , \5646 );
or \U$5459 ( \5648 , \5022 , \5647 );
and \U$5460 ( \5649 , \4943 , \5648 );
or \U$5461 ( \5650 , \4942 , \5649 );
and \U$5462 ( \5651 , \4848 , \5650 );
or \U$5463 ( \5652 , \4847 , \5651 );
and \U$5464 ( \5653 , \4760 , \5652 );
or \U$5465 ( \5654 , \4759 , \5653 );
and \U$5466 ( \5655 , \4668 , \5654 );
or \U$5467 ( \5656 , \4667 , \5655 );
and \U$5468 ( \5657 , \4580 , \5656 );
or \U$5469 ( \5658 , \4579 , \5657 );
and \U$5470 ( \5659 , \4465 , \5658 );
or \U$5471 ( \5660 , \4464 , \5659 );
and \U$5472 ( \5661 , \4369 , \5660 );
or \U$5473 ( \5662 , \4368 , \5661 );
and \U$5474 ( \5663 , \4361 , \5662 );
or \U$5475 ( \5664 , \4360 , \5663 );
and \U$5476 ( \5665 , \4246 , \5664 );
or \U$5477 ( \5666 , \4245 , \5665 );
and \U$5478 ( \5667 , \4122 , \5666 );
or \U$5479 ( \5668 , \4121 , \5667 );
and \U$5480 ( \5669 , \3982 , \5668 );
or \U$5481 ( \5670 , \3981 , \5669 );
and \U$5482 ( \5671 , \3858 , \5670 );
or \U$5483 ( \5672 , \3857 , \5671 );
and \U$5484 ( \5673 , \3714 , \5672 );
or \U$5485 ( \5674 , \3713 , \5673 );
and \U$5486 ( \5675 , \3589 , \5674 );
or \U$5487 ( \5676 , \3588 , \5675 );
and \U$5488 ( \5677 , \3450 , \5676 );
or \U$5489 ( \5678 , \3449 , \5677 );
and \U$5490 ( \5679 , \3285 , \5678 );
or \U$5491 ( \5680 , \3284 , \5679 );
and \U$5492 ( \5681 , \3137 , \5680 );
or \U$5493 ( \5682 , \3136 , \5681 );
and \U$5494 ( \5683 , \2990 , \5682 );
or \U$5495 ( \5684 , \2989 , \5683 );
and \U$5496 ( \5685 , \2822 , \5684 );
or \U$5497 ( \5686 , \2821 , \5685 );
and \U$5498 ( \5687 , \2673 , \5686 );
or \U$5499 ( \5688 , \2672 , \5687 );
and \U$5500 ( \5689 , \2501 , \5688 );
or \U$5501 ( \5690 , \2500 , \5689 );
and \U$5502 ( \5691 , \2365 , \5690 );
or \U$5503 ( \5692 , \2364 , \5691 );
and \U$5504 ( \5693 , \2220 , \5692 );
or \U$5505 ( \5694 , \2219 , \5693 );
and \U$5506 ( \5695 , \2082 , \5694 );
or \U$5507 ( \5696 , \2081 , \5695 );
and \U$5508 ( \5697 , \1947 , \5696 );
or \U$5509 ( \5698 , \1946 , \5697 );
and \U$5510 ( \5699 , \1826 , \5698 );
or \U$5511 ( \5700 , \1825 , \5699 );
and \U$5512 ( \5701 , \1701 , \5700 );
or \U$5513 ( \5702 , \1700 , \5701 );
and \U$5514 ( \5703 , \1585 , \5702 );
or \U$5515 ( \5704 , \1584 , \5703 );
and \U$5516 ( \5705 , \1469 , \5704 );
or \U$5517 ( \5706 , \1468 , \5705 );
and \U$5518 ( \5707 , \1354 , \5706 );
or \U$5519 ( \5708 , \1353 , \5707 );
and \U$5520 ( \5709 , \1238 , \5708 );
or \U$5521 ( \5710 , \1237 , \5709 );
and \U$5522 ( \5711 , \1054 , \5710 );
or \U$5523 ( \5712 , \1053 , \5711 );
and \U$5524 ( \5713 , \975 , \5712 );
or \U$5525 ( \5714 , \974 , \5713 );
and \U$5526 ( \5715 , \891 , \5714 );
or \U$5527 ( \5716 , \890 , \5715 );
and \U$5528 ( \5717 , \809 , \5716 );
or \U$5529 ( \5718 , \808 , \5717 );
and \U$5530 ( \5719 , \733 , \5718 );
or \U$5531 ( \5720 , \732 , \5719 );
and \U$5532 ( \5721 , \658 , \5720 );
or \U$5533 ( \5722 , \657 , \5721 );
and \U$5534 ( \5723 , \536 , \5722 );
or \U$5535 ( \5724 , \535 , \5723 );
xor \U$5536 ( \5725 , \482 , \5724 );
buf g16bf_GF_PartitionCandidate( \5726_nG16bf , \5725 );
buf \U$5537 ( \5727 , \5726_nG16bf );
xor \U$5538 ( \5728 , \536 , \5722 );
buf g16c2_GF_PartitionCandidate( \5729_nG16c2 , \5728 );
buf \U$5539 ( \5730 , \5729_nG16c2 );
xor \U$5540 ( \5731 , \658 , \5720 );
buf g16c5_GF_PartitionCandidate( \5732_nG16c5 , \5731 );
buf \U$5541 ( \5733 , \5732_nG16c5 );
and \U$5542 ( \5734 , \5730 , \5733 );
not \U$5543 ( \5735 , \5734 );
and \U$5544 ( \5736 , \5727 , \5735 );
buf \U$5545 ( \5737 , RIb4bfa38_65);
xor \U$5546 ( \5738 , \4369 , \5660 );
buf g171f_GF_PartitionCandidate( \5739_nG171f , \5738 );
buf \U$5547 ( \5740 , \5739_nG171f );
xor \U$5548 ( \5741 , \4465 , \5658 );
buf g1722_GF_PartitionCandidate( \5742_nG1722 , \5741 );
buf \U$5549 ( \5743 , \5742_nG1722 );
xor \U$5550 ( \5744 , \5740 , \5743 );
xor \U$5551 ( \5745 , \4580 , \5656 );
buf g1725_GF_PartitionCandidate( \5746_nG1725 , \5745 );
buf \U$5552 ( \5747 , \5746_nG1725 );
xor \U$5553 ( \5748 , \5743 , \5747 );
not \U$5554 ( \5749 , \5748 );
and \U$5555 ( \5750 , \5744 , \5749 );
and \U$5556 ( \5751 , \5737 , \5750 );
not \U$5557 ( \5752 , \5751 );
and \U$5558 ( \5753 , \5743 , \5747 );
not \U$5559 ( \5754 , \5753 );
and \U$5560 ( \5755 , \5740 , \5754 );
xnor \U$5561 ( \5756 , \5752 , \5755 );
and \U$5562 ( \5757 , \5736 , \5756 );
buf \U$5563 ( \5758 , RIb4bf948_67);
xor \U$5564 ( \5759 , \4246 , \5664 );
buf g1719_GF_PartitionCandidate( \5760_nG1719 , \5759 );
buf \U$5565 ( \5761 , \5760_nG1719 );
xor \U$5566 ( \5762 , \4361 , \5662 );
buf g171c_GF_PartitionCandidate( \5763_nG171c , \5762 );
buf \U$5567 ( \5764 , \5763_nG171c );
xor \U$5568 ( \5765 , \5761 , \5764 );
xor \U$5569 ( \5766 , \5764 , \5740 );
not \U$5570 ( \5767 , \5766 );
and \U$5571 ( \5768 , \5765 , \5767 );
and \U$5572 ( \5769 , \5758 , \5768 );
buf \U$5573 ( \5770 , RIb4bf9c0_66);
and \U$5574 ( \5771 , \5770 , \5766 );
nor \U$5575 ( \5772 , \5769 , \5771 );
and \U$5576 ( \5773 , \5764 , \5740 );
not \U$5577 ( \5774 , \5773 );
and \U$5578 ( \5775 , \5761 , \5774 );
xnor \U$5579 ( \5776 , \5772 , \5775 );
and \U$5580 ( \5777 , \5756 , \5776 );
and \U$5581 ( \5778 , \5736 , \5776 );
or \U$5582 ( \5779 , \5757 , \5777 , \5778 );
buf \U$5583 ( \5780 , RIb4bf858_69);
xor \U$5584 ( \5781 , \3982 , \5668 );
buf g1713_GF_PartitionCandidate( \5782_nG1713 , \5781 );
buf \U$5585 ( \5783 , \5782_nG1713 );
xor \U$5586 ( \5784 , \4122 , \5666 );
buf g1716_GF_PartitionCandidate( \5785_nG1716 , \5784 );
buf \U$5587 ( \5786 , \5785_nG1716 );
xor \U$5588 ( \5787 , \5783 , \5786 );
xor \U$5589 ( \5788 , \5786 , \5761 );
not \U$5590 ( \5789 , \5788 );
and \U$5591 ( \5790 , \5787 , \5789 );
and \U$5592 ( \5791 , \5780 , \5790 );
buf \U$5593 ( \5792 , RIb4bf8d0_68);
and \U$5594 ( \5793 , \5792 , \5788 );
nor \U$5595 ( \5794 , \5791 , \5793 );
and \U$5596 ( \5795 , \5786 , \5761 );
not \U$5597 ( \5796 , \5795 );
and \U$5598 ( \5797 , \5783 , \5796 );
xnor \U$5599 ( \5798 , \5794 , \5797 );
buf \U$5600 ( \5799 , RIb4bf768_71);
xor \U$5601 ( \5800 , \3714 , \5672 );
buf g170d_GF_PartitionCandidate( \5801_nG170d , \5800 );
buf \U$5602 ( \5802 , \5801_nG170d );
xor \U$5603 ( \5803 , \3858 , \5670 );
buf g1710_GF_PartitionCandidate( \5804_nG1710 , \5803 );
buf \U$5604 ( \5805 , \5804_nG1710 );
xor \U$5605 ( \5806 , \5802 , \5805 );
xor \U$5606 ( \5807 , \5805 , \5783 );
not \U$5607 ( \5808 , \5807 );
and \U$5608 ( \5809 , \5806 , \5808 );
and \U$5609 ( \5810 , \5799 , \5809 );
buf \U$5610 ( \5811 , RIb4bf7e0_70);
and \U$5611 ( \5812 , \5811 , \5807 );
nor \U$5612 ( \5813 , \5810 , \5812 );
and \U$5613 ( \5814 , \5805 , \5783 );
not \U$5614 ( \5815 , \5814 );
and \U$5615 ( \5816 , \5802 , \5815 );
xnor \U$5616 ( \5817 , \5813 , \5816 );
and \U$5617 ( \5818 , \5798 , \5817 );
buf \U$5618 ( \5819 , RIb4bf678_73);
xor \U$5619 ( \5820 , \3450 , \5676 );
buf g1707_GF_PartitionCandidate( \5821_nG1707 , \5820 );
buf \U$5620 ( \5822 , \5821_nG1707 );
xor \U$5621 ( \5823 , \3589 , \5674 );
buf g170a_GF_PartitionCandidate( \5824_nG170a , \5823 );
buf \U$5622 ( \5825 , \5824_nG170a );
xor \U$5623 ( \5826 , \5822 , \5825 );
xor \U$5624 ( \5827 , \5825 , \5802 );
not \U$5625 ( \5828 , \5827 );
and \U$5626 ( \5829 , \5826 , \5828 );
and \U$5627 ( \5830 , \5819 , \5829 );
buf \U$5628 ( \5831 , RIb4bf6f0_72);
and \U$5629 ( \5832 , \5831 , \5827 );
nor \U$5630 ( \5833 , \5830 , \5832 );
and \U$5631 ( \5834 , \5825 , \5802 );
not \U$5632 ( \5835 , \5834 );
and \U$5633 ( \5836 , \5822 , \5835 );
xnor \U$5634 ( \5837 , \5833 , \5836 );
and \U$5635 ( \5838 , \5817 , \5837 );
and \U$5636 ( \5839 , \5798 , \5837 );
or \U$5637 ( \5840 , \5818 , \5838 , \5839 );
and \U$5638 ( \5841 , \5779 , \5840 );
buf \U$5639 ( \5842 , RIb4bf588_75);
xor \U$5640 ( \5843 , \3137 , \5680 );
buf g1701_GF_PartitionCandidate( \5844_nG1701 , \5843 );
buf \U$5641 ( \5845 , \5844_nG1701 );
xor \U$5642 ( \5846 , \3285 , \5678 );
buf g1704_GF_PartitionCandidate( \5847_nG1704 , \5846 );
buf \U$5643 ( \5848 , \5847_nG1704 );
xor \U$5644 ( \5849 , \5845 , \5848 );
xor \U$5645 ( \5850 , \5848 , \5822 );
not \U$5646 ( \5851 , \5850 );
and \U$5647 ( \5852 , \5849 , \5851 );
and \U$5648 ( \5853 , \5842 , \5852 );
buf \U$5649 ( \5854 , RIb4bf600_74);
and \U$5650 ( \5855 , \5854 , \5850 );
nor \U$5651 ( \5856 , \5853 , \5855 );
and \U$5652 ( \5857 , \5848 , \5822 );
not \U$5653 ( \5858 , \5857 );
and \U$5654 ( \5859 , \5845 , \5858 );
xnor \U$5655 ( \5860 , \5856 , \5859 );
buf \U$5656 ( \5861 , RIb4bf498_77);
xor \U$5657 ( \5862 , \2822 , \5684 );
buf g16fb_GF_PartitionCandidate( \5863_nG16fb , \5862 );
buf \U$5658 ( \5864 , \5863_nG16fb );
xor \U$5659 ( \5865 , \2990 , \5682 );
buf g16fe_GF_PartitionCandidate( \5866_nG16fe , \5865 );
buf \U$5660 ( \5867 , \5866_nG16fe );
xor \U$5661 ( \5868 , \5864 , \5867 );
xor \U$5662 ( \5869 , \5867 , \5845 );
not \U$5663 ( \5870 , \5869 );
and \U$5664 ( \5871 , \5868 , \5870 );
and \U$5665 ( \5872 , \5861 , \5871 );
buf \U$5666 ( \5873 , RIb4bf510_76);
and \U$5667 ( \5874 , \5873 , \5869 );
nor \U$5668 ( \5875 , \5872 , \5874 );
and \U$5669 ( \5876 , \5867 , \5845 );
not \U$5670 ( \5877 , \5876 );
and \U$5671 ( \5878 , \5864 , \5877 );
xnor \U$5672 ( \5879 , \5875 , \5878 );
and \U$5673 ( \5880 , \5860 , \5879 );
buf \U$5674 ( \5881 , RIb4bf3a8_79);
xor \U$5675 ( \5882 , \2501 , \5688 );
buf g16f5_GF_PartitionCandidate( \5883_nG16f5 , \5882 );
buf \U$5676 ( \5884 , \5883_nG16f5 );
xor \U$5677 ( \5885 , \2673 , \5686 );
buf g16f8_GF_PartitionCandidate( \5886_nG16f8 , \5885 );
buf \U$5678 ( \5887 , \5886_nG16f8 );
xor \U$5679 ( \5888 , \5884 , \5887 );
xor \U$5680 ( \5889 , \5887 , \5864 );
not \U$5681 ( \5890 , \5889 );
and \U$5682 ( \5891 , \5888 , \5890 );
and \U$5683 ( \5892 , \5881 , \5891 );
buf \U$5684 ( \5893 , RIb4bf420_78);
and \U$5685 ( \5894 , \5893 , \5889 );
nor \U$5686 ( \5895 , \5892 , \5894 );
and \U$5687 ( \5896 , \5887 , \5864 );
not \U$5688 ( \5897 , \5896 );
and \U$5689 ( \5898 , \5884 , \5897 );
xnor \U$5690 ( \5899 , \5895 , \5898 );
and \U$5691 ( \5900 , \5879 , \5899 );
and \U$5692 ( \5901 , \5860 , \5899 );
or \U$5693 ( \5902 , \5880 , \5900 , \5901 );
and \U$5694 ( \5903 , \5840 , \5902 );
and \U$5695 ( \5904 , \5779 , \5902 );
or \U$5696 ( \5905 , \5841 , \5903 , \5904 );
buf \U$5697 ( \5906 , RIb4bf2b8_81);
xor \U$5698 ( \5907 , \2220 , \5692 );
buf g16ef_GF_PartitionCandidate( \5908_nG16ef , \5907 );
buf \U$5699 ( \5909 , \5908_nG16ef );
xor \U$5700 ( \5910 , \2365 , \5690 );
buf g16f2_GF_PartitionCandidate( \5911_nG16f2 , \5910 );
buf \U$5701 ( \5912 , \5911_nG16f2 );
xor \U$5702 ( \5913 , \5909 , \5912 );
xor \U$5703 ( \5914 , \5912 , \5884 );
not \U$5704 ( \5915 , \5914 );
and \U$5705 ( \5916 , \5913 , \5915 );
and \U$5706 ( \5917 , \5906 , \5916 );
buf \U$5707 ( \5918 , RIb4bf330_80);
and \U$5708 ( \5919 , \5918 , \5914 );
nor \U$5709 ( \5920 , \5917 , \5919 );
and \U$5710 ( \5921 , \5912 , \5884 );
not \U$5711 ( \5922 , \5921 );
and \U$5712 ( \5923 , \5909 , \5922 );
xnor \U$5713 ( \5924 , \5920 , \5923 );
buf \U$5714 ( \5925 , RIb4bf1c8_83);
xor \U$5715 ( \5926 , \1947 , \5696 );
buf g16e9_GF_PartitionCandidate( \5927_nG16e9 , \5926 );
buf \U$5716 ( \5928 , \5927_nG16e9 );
xor \U$5717 ( \5929 , \2082 , \5694 );
buf g16ec_GF_PartitionCandidate( \5930_nG16ec , \5929 );
buf \U$5718 ( \5931 , \5930_nG16ec );
xor \U$5719 ( \5932 , \5928 , \5931 );
xor \U$5720 ( \5933 , \5931 , \5909 );
not \U$5721 ( \5934 , \5933 );
and \U$5722 ( \5935 , \5932 , \5934 );
and \U$5723 ( \5936 , \5925 , \5935 );
buf \U$5724 ( \5937 , RIb4bf240_82);
and \U$5725 ( \5938 , \5937 , \5933 );
nor \U$5726 ( \5939 , \5936 , \5938 );
and \U$5727 ( \5940 , \5931 , \5909 );
not \U$5728 ( \5941 , \5940 );
and \U$5729 ( \5942 , \5928 , \5941 );
xnor \U$5730 ( \5943 , \5939 , \5942 );
and \U$5731 ( \5944 , \5924 , \5943 );
buf \U$5732 ( \5945 , RIb4bf0d8_85);
xor \U$5733 ( \5946 , \1701 , \5700 );
buf g16e3_GF_PartitionCandidate( \5947_nG16e3 , \5946 );
buf \U$5734 ( \5948 , \5947_nG16e3 );
xor \U$5735 ( \5949 , \1826 , \5698 );
buf g16e6_GF_PartitionCandidate( \5950_nG16e6 , \5949 );
buf \U$5736 ( \5951 , \5950_nG16e6 );
xor \U$5737 ( \5952 , \5948 , \5951 );
xor \U$5738 ( \5953 , \5951 , \5928 );
not \U$5739 ( \5954 , \5953 );
and \U$5740 ( \5955 , \5952 , \5954 );
and \U$5741 ( \5956 , \5945 , \5955 );
buf \U$5742 ( \5957 , RIb4bf150_84);
and \U$5743 ( \5958 , \5957 , \5953 );
nor \U$5744 ( \5959 , \5956 , \5958 );
and \U$5745 ( \5960 , \5951 , \5928 );
not \U$5746 ( \5961 , \5960 );
and \U$5747 ( \5962 , \5948 , \5961 );
xnor \U$5748 ( \5963 , \5959 , \5962 );
and \U$5749 ( \5964 , \5943 , \5963 );
and \U$5750 ( \5965 , \5924 , \5963 );
or \U$5751 ( \5966 , \5944 , \5964 , \5965 );
buf \U$5752 ( \5967 , RIb4befe8_87);
xor \U$5753 ( \5968 , \1469 , \5704 );
buf g16dd_GF_PartitionCandidate( \5969_nG16dd , \5968 );
buf \U$5754 ( \5970 , \5969_nG16dd );
xor \U$5755 ( \5971 , \1585 , \5702 );
buf g16e0_GF_PartitionCandidate( \5972_nG16e0 , \5971 );
buf \U$5756 ( \5973 , \5972_nG16e0 );
xor \U$5757 ( \5974 , \5970 , \5973 );
xor \U$5758 ( \5975 , \5973 , \5948 );
not \U$5759 ( \5976 , \5975 );
and \U$5760 ( \5977 , \5974 , \5976 );
and \U$5761 ( \5978 , \5967 , \5977 );
buf \U$5762 ( \5979 , RIb4bf060_86);
and \U$5763 ( \5980 , \5979 , \5975 );
nor \U$5764 ( \5981 , \5978 , \5980 );
and \U$5765 ( \5982 , \5973 , \5948 );
not \U$5766 ( \5983 , \5982 );
and \U$5767 ( \5984 , \5970 , \5983 );
xnor \U$5768 ( \5985 , \5981 , \5984 );
buf \U$5769 ( \5986 , RIb4beef8_89);
xor \U$5770 ( \5987 , \1238 , \5708 );
buf g16d7_GF_PartitionCandidate( \5988_nG16d7 , \5987 );
buf \U$5771 ( \5989 , \5988_nG16d7 );
xor \U$5772 ( \5990 , \1354 , \5706 );
buf g16da_GF_PartitionCandidate( \5991_nG16da , \5990 );
buf \U$5773 ( \5992 , \5991_nG16da );
xor \U$5774 ( \5993 , \5989 , \5992 );
xor \U$5775 ( \5994 , \5992 , \5970 );
not \U$5776 ( \5995 , \5994 );
and \U$5777 ( \5996 , \5993 , \5995 );
and \U$5778 ( \5997 , \5986 , \5996 );
buf \U$5779 ( \5998 , RIb4bef70_88);
and \U$5780 ( \5999 , \5998 , \5994 );
nor \U$5781 ( \6000 , \5997 , \5999 );
and \U$5782 ( \6001 , \5992 , \5970 );
not \U$5783 ( \6002 , \6001 );
and \U$5784 ( \6003 , \5989 , \6002 );
xnor \U$5785 ( \6004 , \6000 , \6003 );
and \U$5786 ( \6005 , \5985 , \6004 );
buf \U$5787 ( \6006 , RIb4bc1f8_91);
xor \U$5788 ( \6007 , \975 , \5712 );
buf g16d1_GF_PartitionCandidate( \6008_nG16d1 , \6007 );
buf \U$5789 ( \6009 , \6008_nG16d1 );
xor \U$5790 ( \6010 , \1054 , \5710 );
buf g16d4_GF_PartitionCandidate( \6011_nG16d4 , \6010 );
buf \U$5791 ( \6012 , \6011_nG16d4 );
xor \U$5792 ( \6013 , \6009 , \6012 );
xor \U$5793 ( \6014 , \6012 , \5989 );
not \U$5794 ( \6015 , \6014 );
and \U$5795 ( \6016 , \6013 , \6015 );
and \U$5796 ( \6017 , \6006 , \6016 );
buf \U$5797 ( \6018 , RIb4bee80_90);
and \U$5798 ( \6019 , \6018 , \6014 );
nor \U$5799 ( \6020 , \6017 , \6019 );
and \U$5800 ( \6021 , \6012 , \5989 );
not \U$5801 ( \6022 , \6021 );
and \U$5802 ( \6023 , \6009 , \6022 );
xnor \U$5803 ( \6024 , \6020 , \6023 );
and \U$5804 ( \6025 , \6004 , \6024 );
and \U$5805 ( \6026 , \5985 , \6024 );
or \U$5806 ( \6027 , \6005 , \6025 , \6026 );
and \U$5807 ( \6028 , \5966 , \6027 );
buf \U$5808 ( \6029 , RIb4bc108_93);
xor \U$5809 ( \6030 , \809 , \5716 );
buf g16cb_GF_PartitionCandidate( \6031_nG16cb , \6030 );
buf \U$5810 ( \6032 , \6031_nG16cb );
xor \U$5811 ( \6033 , \891 , \5714 );
buf g16ce_GF_PartitionCandidate( \6034_nG16ce , \6033 );
buf \U$5812 ( \6035 , \6034_nG16ce );
xor \U$5813 ( \6036 , \6032 , \6035 );
xor \U$5814 ( \6037 , \6035 , \6009 );
not \U$5815 ( \6038 , \6037 );
and \U$5816 ( \6039 , \6036 , \6038 );
and \U$5817 ( \6040 , \6029 , \6039 );
buf \U$5818 ( \6041 , RIb4bc180_92);
and \U$5819 ( \6042 , \6041 , \6037 );
nor \U$5820 ( \6043 , \6040 , \6042 );
and \U$5821 ( \6044 , \6035 , \6009 );
not \U$5822 ( \6045 , \6044 );
and \U$5823 ( \6046 , \6032 , \6045 );
xnor \U$5824 ( \6047 , \6043 , \6046 );
buf \U$5825 ( \6048 , RIb4bc018_95);
xor \U$5826 ( \6049 , \733 , \5718 );
buf g16c8_GF_PartitionCandidate( \6050_nG16c8 , \6049 );
buf \U$5827 ( \6051 , \6050_nG16c8 );
xor \U$5828 ( \6052 , \5733 , \6051 );
xor \U$5829 ( \6053 , \6051 , \6032 );
not \U$5830 ( \6054 , \6053 );
and \U$5831 ( \6055 , \6052 , \6054 );
and \U$5832 ( \6056 , \6048 , \6055 );
buf \U$5833 ( \6057 , RIb4bc090_94);
and \U$5834 ( \6058 , \6057 , \6053 );
nor \U$5835 ( \6059 , \6056 , \6058 );
and \U$5836 ( \6060 , \6051 , \6032 );
not \U$5837 ( \6061 , \6060 );
and \U$5838 ( \6062 , \5733 , \6061 );
xnor \U$5839 ( \6063 , \6059 , \6062 );
and \U$5840 ( \6064 , \6047 , \6063 );
buf \U$5841 ( \6065 , RIb4bbfa0_96);
xor \U$5842 ( \6066 , \5730 , \5733 );
nand \U$5843 ( \6067 , \6065 , \6066 );
xnor \U$5844 ( \6068 , \6067 , \5736 );
and \U$5845 ( \6069 , \6063 , \6068 );
and \U$5846 ( \6070 , \6047 , \6068 );
or \U$5847 ( \6071 , \6064 , \6069 , \6070 );
and \U$5848 ( \6072 , \6027 , \6071 );
and \U$5849 ( \6073 , \5966 , \6071 );
or \U$5850 ( \6074 , \6028 , \6072 , \6073 );
and \U$5851 ( \6075 , \5905 , \6074 );
and \U$5852 ( \6076 , \6057 , \6055 );
and \U$5853 ( \6077 , \6029 , \6053 );
nor \U$5854 ( \6078 , \6076 , \6077 );
xnor \U$5855 ( \6079 , \6078 , \6062 );
xor \U$5856 ( \6080 , \5727 , \5730 );
not \U$5857 ( \6081 , \6066 );
and \U$5858 ( \6082 , \6080 , \6081 );
and \U$5859 ( \6083 , \6065 , \6082 );
and \U$5860 ( \6084 , \6048 , \6066 );
nor \U$5861 ( \6085 , \6083 , \6084 );
xnor \U$5862 ( \6086 , \6085 , \5736 );
xor \U$5863 ( \6087 , \6079 , \6086 );
and \U$5864 ( \6088 , \5998 , \5996 );
and \U$5865 ( \6089 , \5967 , \5994 );
nor \U$5866 ( \6090 , \6088 , \6089 );
xnor \U$5867 ( \6091 , \6090 , \6003 );
and \U$5868 ( \6092 , \6018 , \6016 );
and \U$5869 ( \6093 , \5986 , \6014 );
nor \U$5870 ( \6094 , \6092 , \6093 );
xnor \U$5871 ( \6095 , \6094 , \6023 );
xor \U$5872 ( \6096 , \6091 , \6095 );
and \U$5873 ( \6097 , \6041 , \6039 );
and \U$5874 ( \6098 , \6006 , \6037 );
nor \U$5875 ( \6099 , \6097 , \6098 );
xnor \U$5876 ( \6100 , \6099 , \6046 );
xor \U$5877 ( \6101 , \6096 , \6100 );
and \U$5878 ( \6102 , \6087 , \6101 );
and \U$5879 ( \6103 , \5937 , \5935 );
and \U$5880 ( \6104 , \5906 , \5933 );
nor \U$5881 ( \6105 , \6103 , \6104 );
xnor \U$5882 ( \6106 , \6105 , \5942 );
and \U$5883 ( \6107 , \5957 , \5955 );
and \U$5884 ( \6108 , \5925 , \5953 );
nor \U$5885 ( \6109 , \6107 , \6108 );
xnor \U$5886 ( \6110 , \6109 , \5962 );
xor \U$5887 ( \6111 , \6106 , \6110 );
and \U$5888 ( \6112 , \5979 , \5977 );
and \U$5889 ( \6113 , \5945 , \5975 );
nor \U$5890 ( \6114 , \6112 , \6113 );
xnor \U$5891 ( \6115 , \6114 , \5984 );
xor \U$5892 ( \6116 , \6111 , \6115 );
and \U$5893 ( \6117 , \6101 , \6116 );
and \U$5894 ( \6118 , \6087 , \6116 );
or \U$5895 ( \6119 , \6102 , \6117 , \6118 );
and \U$5896 ( \6120 , \6074 , \6119 );
and \U$5897 ( \6121 , \5905 , \6119 );
or \U$5898 ( \6122 , \6075 , \6120 , \6121 );
and \U$5899 ( \6123 , \5873 , \5871 );
and \U$5900 ( \6124 , \5842 , \5869 );
nor \U$5901 ( \6125 , \6123 , \6124 );
xnor \U$5902 ( \6126 , \6125 , \5878 );
and \U$5903 ( \6127 , \5893 , \5891 );
and \U$5904 ( \6128 , \5861 , \5889 );
nor \U$5905 ( \6129 , \6127 , \6128 );
xnor \U$5906 ( \6130 , \6129 , \5898 );
xor \U$5907 ( \6131 , \6126 , \6130 );
and \U$5908 ( \6132 , \5918 , \5916 );
and \U$5909 ( \6133 , \5881 , \5914 );
nor \U$5910 ( \6134 , \6132 , \6133 );
xnor \U$5911 ( \6135 , \6134 , \5923 );
xor \U$5912 ( \6136 , \6131 , \6135 );
and \U$5913 ( \6137 , \5811 , \5809 );
and \U$5914 ( \6138 , \5780 , \5807 );
nor \U$5915 ( \6139 , \6137 , \6138 );
xnor \U$5916 ( \6140 , \6139 , \5816 );
and \U$5917 ( \6141 , \5831 , \5829 );
and \U$5918 ( \6142 , \5799 , \5827 );
nor \U$5919 ( \6143 , \6141 , \6142 );
xnor \U$5920 ( \6144 , \6143 , \5836 );
xor \U$5921 ( \6145 , \6140 , \6144 );
and \U$5922 ( \6146 , \5854 , \5852 );
and \U$5923 ( \6147 , \5819 , \5850 );
nor \U$5924 ( \6148 , \6146 , \6147 );
xnor \U$5925 ( \6149 , \6148 , \5859 );
xor \U$5926 ( \6150 , \6145 , \6149 );
and \U$5927 ( \6151 , \6136 , \6150 );
not \U$5928 ( \6152 , \5755 );
and \U$5929 ( \6153 , \5770 , \5768 );
and \U$5930 ( \6154 , \5737 , \5766 );
nor \U$5931 ( \6155 , \6153 , \6154 );
xnor \U$5932 ( \6156 , \6155 , \5775 );
xor \U$5933 ( \6157 , \6152 , \6156 );
and \U$5934 ( \6158 , \5792 , \5790 );
and \U$5935 ( \6159 , \5758 , \5788 );
nor \U$5936 ( \6160 , \6158 , \6159 );
xnor \U$5937 ( \6161 , \6160 , \5797 );
xor \U$5938 ( \6162 , \6157 , \6161 );
and \U$5939 ( \6163 , \6150 , \6162 );
and \U$5940 ( \6164 , \6136 , \6162 );
or \U$5941 ( \6165 , \6151 , \6163 , \6164 );
and \U$5942 ( \6166 , \289 , \328 );
not \U$5943 ( \6167 , \6166 );
xnor \U$5944 ( \6168 , \6167 , \336 );
and \U$5945 ( \6169 , \304 , \348 );
and \U$5946 ( \6170 , \313 , \346 );
nor \U$5947 ( \6171 , \6169 , \6170 );
xnor \U$5948 ( \6172 , \6171 , \356 );
and \U$5949 ( \6173 , \6168 , \6172 );
and \U$5950 ( \6174 , \331 , \343 );
and \U$5951 ( \6175 , \6172 , \6174 );
and \U$5952 ( \6176 , \6168 , \6174 );
or \U$5953 ( \6177 , \6173 , \6175 , \6176 );
and \U$5954 ( \6178 , \412 , \416 );
and \U$5955 ( \6179 , \416 , \421 );
and \U$5956 ( \6180 , \412 , \421 );
or \U$5957 ( \6181 , \6178 , \6179 , \6180 );
xor \U$5958 ( \6182 , \6168 , \6172 );
xor \U$5959 ( \6183 , \6182 , \6174 );
or \U$5960 ( \6184 , \6181 , \6183 );
xor \U$5961 ( \6185 , \6177 , \6184 );
not \U$5962 ( \6186 , \336 );
and \U$5963 ( \6187 , \313 , \348 );
and \U$5964 ( \6188 , \289 , \346 );
nor \U$5965 ( \6189 , \6187 , \6188 );
xnor \U$5966 ( \6190 , \6189 , \356 );
xor \U$5967 ( \6191 , \6186 , \6190 );
and \U$5968 ( \6192 , \304 , \343 );
xor \U$5969 ( \6193 , \6191 , \6192 );
xor \U$5970 ( \6194 , \6185 , \6193 );
and \U$5971 ( \6195 , \427 , \428 );
and \U$5972 ( \6196 , \428 , \430 );
and \U$5973 ( \6197 , \427 , \430 );
or \U$5974 ( \6198 , \6195 , \6196 , \6197 );
and \U$5975 ( \6199 , \411 , \422 );
and \U$5976 ( \6200 , \422 , \431 );
and \U$5977 ( \6201 , \411 , \431 );
or \U$5978 ( \6202 , \6199 , \6200 , \6201 );
and \U$5979 ( \6203 , \6198 , \6202 );
xnor \U$5980 ( \6204 , \6181 , \6183 );
and \U$5981 ( \6205 , \6202 , \6204 );
and \U$5982 ( \6206 , \6198 , \6204 );
or \U$5983 ( \6207 , \6203 , \6205 , \6206 );
xor \U$5984 ( \6208 , \6194 , \6207 );
xor \U$5985 ( \6209 , \6198 , \6202 );
xor \U$5986 ( \6210 , \6209 , \6204 );
and \U$5987 ( \6211 , \407 , \432 );
and \U$5988 ( \6212 , \6210 , \6211 );
xor \U$5989 ( \6213 , \6210 , \6211 );
and \U$5990 ( \6214 , \433 , \481 );
and \U$5991 ( \6215 , \482 , \5724 );
or \U$5992 ( \6216 , \6214 , \6215 );
and \U$5993 ( \6217 , \6213 , \6216 );
or \U$5994 ( \6218 , \6212 , \6217 );
xor \U$5995 ( \6219 , \6208 , \6218 );
buf g16b9_GF_PartitionCandidate( \6220_nG16b9 , \6219 );
buf \U$5996 ( \6221 , \6220_nG16b9 );
xor \U$5997 ( \6222 , \6213 , \6216 );
buf g16bc_GF_PartitionCandidate( \6223_nG16bc , \6222 );
buf \U$5998 ( \6224 , \6223_nG16bc );
and \U$5999 ( \6225 , \6224 , \5727 );
not \U$6000 ( \6226 , \6225 );
and \U$6001 ( \6227 , \6221 , \6226 );
and \U$6002 ( \6228 , \5737 , \5768 );
not \U$6003 ( \6229 , \6228 );
xnor \U$6004 ( \6230 , \6229 , \5775 );
xor \U$6005 ( \6231 , \6227 , \6230 );
and \U$6006 ( \6232 , \5758 , \5790 );
and \U$6007 ( \6233 , \5770 , \5788 );
nor \U$6008 ( \6234 , \6232 , \6233 );
xnor \U$6009 ( \6235 , \6234 , \5797 );
xor \U$6010 ( \6236 , \6231 , \6235 );
and \U$6011 ( \6237 , \6165 , \6236 );
and \U$6012 ( \6238 , \5906 , \5935 );
and \U$6013 ( \6239 , \5918 , \5933 );
nor \U$6014 ( \6240 , \6238 , \6239 );
xnor \U$6015 ( \6241 , \6240 , \5942 );
and \U$6016 ( \6242 , \5925 , \5955 );
and \U$6017 ( \6243 , \5937 , \5953 );
nor \U$6018 ( \6244 , \6242 , \6243 );
xnor \U$6019 ( \6245 , \6244 , \5962 );
xor \U$6020 ( \6246 , \6241 , \6245 );
and \U$6021 ( \6247 , \5945 , \5977 );
and \U$6022 ( \6248 , \5957 , \5975 );
nor \U$6023 ( \6249 , \6247 , \6248 );
xnor \U$6024 ( \6250 , \6249 , \5984 );
xor \U$6025 ( \6251 , \6246 , \6250 );
and \U$6026 ( \6252 , \5842 , \5871 );
and \U$6027 ( \6253 , \5854 , \5869 );
nor \U$6028 ( \6254 , \6252 , \6253 );
xnor \U$6029 ( \6255 , \6254 , \5878 );
and \U$6030 ( \6256 , \5861 , \5891 );
and \U$6031 ( \6257 , \5873 , \5889 );
nor \U$6032 ( \6258 , \6256 , \6257 );
xnor \U$6033 ( \6259 , \6258 , \5898 );
xor \U$6034 ( \6260 , \6255 , \6259 );
and \U$6035 ( \6261 , \5881 , \5916 );
and \U$6036 ( \6262 , \5893 , \5914 );
nor \U$6037 ( \6263 , \6261 , \6262 );
xnor \U$6038 ( \6264 , \6263 , \5923 );
xor \U$6039 ( \6265 , \6260 , \6264 );
xor \U$6040 ( \6266 , \6251 , \6265 );
and \U$6041 ( \6267 , \5780 , \5809 );
and \U$6042 ( \6268 , \5792 , \5807 );
nor \U$6043 ( \6269 , \6267 , \6268 );
xnor \U$6044 ( \6270 , \6269 , \5816 );
and \U$6045 ( \6271 , \5799 , \5829 );
and \U$6046 ( \6272 , \5811 , \5827 );
nor \U$6047 ( \6273 , \6271 , \6272 );
xnor \U$6048 ( \6274 , \6273 , \5836 );
xor \U$6049 ( \6275 , \6270 , \6274 );
and \U$6050 ( \6276 , \5819 , \5852 );
and \U$6051 ( \6277 , \5831 , \5850 );
nor \U$6052 ( \6278 , \6276 , \6277 );
xnor \U$6053 ( \6279 , \6278 , \5859 );
xor \U$6054 ( \6280 , \6275 , \6279 );
xor \U$6055 ( \6281 , \6266 , \6280 );
and \U$6056 ( \6282 , \6236 , \6281 );
and \U$6057 ( \6283 , \6165 , \6281 );
or \U$6058 ( \6284 , \6237 , \6282 , \6283 );
and \U$6059 ( \6285 , \6122 , \6284 );
and \U$6060 ( \6286 , \6029 , \6055 );
and \U$6061 ( \6287 , \6041 , \6053 );
nor \U$6062 ( \6288 , \6286 , \6287 );
xnor \U$6063 ( \6289 , \6288 , \6062 );
and \U$6064 ( \6290 , \6048 , \6082 );
and \U$6065 ( \6291 , \6057 , \6066 );
nor \U$6066 ( \6292 , \6290 , \6291 );
xnor \U$6067 ( \6293 , \6292 , \5736 );
xor \U$6068 ( \6294 , \6289 , \6293 );
xor \U$6069 ( \6295 , \6224 , \5727 );
nand \U$6070 ( \6296 , \6065 , \6295 );
xnor \U$6071 ( \6297 , \6296 , \6227 );
xor \U$6072 ( \6298 , \6294 , \6297 );
and \U$6073 ( \6299 , \5967 , \5996 );
and \U$6074 ( \6300 , \5979 , \5994 );
nor \U$6075 ( \6301 , \6299 , \6300 );
xnor \U$6076 ( \6302 , \6301 , \6003 );
and \U$6077 ( \6303 , \5986 , \6016 );
and \U$6078 ( \6304 , \5998 , \6014 );
nor \U$6079 ( \6305 , \6303 , \6304 );
xnor \U$6080 ( \6306 , \6305 , \6023 );
xor \U$6081 ( \6307 , \6302 , \6306 );
and \U$6082 ( \6308 , \6006 , \6039 );
and \U$6083 ( \6309 , \6018 , \6037 );
nor \U$6084 ( \6310 , \6308 , \6309 );
xnor \U$6085 ( \6311 , \6310 , \6046 );
xor \U$6086 ( \6312 , \6307 , \6311 );
xnor \U$6087 ( \6313 , \6298 , \6312 );
and \U$6088 ( \6314 , \6106 , \6110 );
and \U$6089 ( \6315 , \6110 , \6115 );
and \U$6090 ( \6316 , \6106 , \6115 );
or \U$6091 ( \6317 , \6314 , \6315 , \6316 );
and \U$6092 ( \6318 , \6091 , \6095 );
and \U$6093 ( \6319 , \6095 , \6100 );
and \U$6094 ( \6320 , \6091 , \6100 );
or \U$6095 ( \6321 , \6318 , \6319 , \6320 );
xor \U$6096 ( \6322 , \6317 , \6321 );
and \U$6097 ( \6323 , \6079 , \6086 );
xor \U$6098 ( \6324 , \6322 , \6323 );
and \U$6099 ( \6325 , \6313 , \6324 );
and \U$6100 ( \6326 , \6152 , \6156 );
and \U$6101 ( \6327 , \6156 , \6161 );
and \U$6102 ( \6328 , \6152 , \6161 );
or \U$6103 ( \6329 , \6326 , \6327 , \6328 );
and \U$6104 ( \6330 , \6140 , \6144 );
and \U$6105 ( \6331 , \6144 , \6149 );
and \U$6106 ( \6332 , \6140 , \6149 );
or \U$6107 ( \6333 , \6330 , \6331 , \6332 );
xor \U$6108 ( \6334 , \6329 , \6333 );
and \U$6109 ( \6335 , \6126 , \6130 );
and \U$6110 ( \6336 , \6130 , \6135 );
and \U$6111 ( \6337 , \6126 , \6135 );
or \U$6112 ( \6338 , \6335 , \6336 , \6337 );
xor \U$6113 ( \6339 , \6334 , \6338 );
and \U$6114 ( \6340 , \6324 , \6339 );
and \U$6115 ( \6341 , \6313 , \6339 );
or \U$6116 ( \6342 , \6325 , \6340 , \6341 );
and \U$6117 ( \6343 , \6284 , \6342 );
and \U$6118 ( \6344 , \6122 , \6342 );
or \U$6119 ( \6345 , \6285 , \6343 , \6344 );
and \U$6120 ( \6346 , \6241 , \6245 );
and \U$6121 ( \6347 , \6245 , \6250 );
and \U$6122 ( \6348 , \6241 , \6250 );
or \U$6123 ( \6349 , \6346 , \6347 , \6348 );
and \U$6124 ( \6350 , \6302 , \6306 );
and \U$6125 ( \6351 , \6306 , \6311 );
and \U$6126 ( \6352 , \6302 , \6311 );
or \U$6127 ( \6353 , \6350 , \6351 , \6352 );
xor \U$6128 ( \6354 , \6349 , \6353 );
and \U$6129 ( \6355 , \6289 , \6293 );
and \U$6130 ( \6356 , \6293 , \6297 );
and \U$6131 ( \6357 , \6289 , \6297 );
or \U$6132 ( \6358 , \6355 , \6356 , \6357 );
xor \U$6133 ( \6359 , \6354 , \6358 );
and \U$6134 ( \6360 , \6227 , \6230 );
and \U$6135 ( \6361 , \6230 , \6235 );
and \U$6136 ( \6362 , \6227 , \6235 );
or \U$6137 ( \6363 , \6360 , \6361 , \6362 );
and \U$6138 ( \6364 , \6270 , \6274 );
and \U$6139 ( \6365 , \6274 , \6279 );
and \U$6140 ( \6366 , \6270 , \6279 );
or \U$6141 ( \6367 , \6364 , \6365 , \6366 );
xor \U$6142 ( \6368 , \6363 , \6367 );
and \U$6143 ( \6369 , \6255 , \6259 );
and \U$6144 ( \6370 , \6259 , \6264 );
and \U$6145 ( \6371 , \6255 , \6264 );
or \U$6146 ( \6372 , \6369 , \6370 , \6371 );
xor \U$6147 ( \6373 , \6368 , \6372 );
xor \U$6148 ( \6374 , \6359 , \6373 );
and \U$6149 ( \6375 , \6251 , \6265 );
and \U$6150 ( \6376 , \6265 , \6280 );
and \U$6151 ( \6377 , \6251 , \6280 );
or \U$6152 ( \6378 , \6375 , \6376 , \6377 );
and \U$6153 ( \6379 , \5873 , \5891 );
and \U$6154 ( \6380 , \5842 , \5889 );
nor \U$6155 ( \6381 , \6379 , \6380 );
xnor \U$6156 ( \6382 , \6381 , \5898 );
and \U$6157 ( \6383 , \5893 , \5916 );
and \U$6158 ( \6384 , \5861 , \5914 );
nor \U$6159 ( \6385 , \6383 , \6384 );
xnor \U$6160 ( \6386 , \6385 , \5923 );
xor \U$6161 ( \6387 , \6382 , \6386 );
and \U$6162 ( \6388 , \5918 , \5935 );
and \U$6163 ( \6389 , \5881 , \5933 );
nor \U$6164 ( \6390 , \6388 , \6389 );
xnor \U$6165 ( \6391 , \6390 , \5942 );
xor \U$6166 ( \6392 , \6387 , \6391 );
and \U$6167 ( \6393 , \5811 , \5829 );
and \U$6168 ( \6394 , \5780 , \5827 );
nor \U$6169 ( \6395 , \6393 , \6394 );
xnor \U$6170 ( \6396 , \6395 , \5836 );
and \U$6171 ( \6397 , \5831 , \5852 );
and \U$6172 ( \6398 , \5799 , \5850 );
nor \U$6173 ( \6399 , \6397 , \6398 );
xnor \U$6174 ( \6400 , \6399 , \5859 );
xor \U$6175 ( \6401 , \6396 , \6400 );
and \U$6176 ( \6402 , \5854 , \5871 );
and \U$6177 ( \6403 , \5819 , \5869 );
nor \U$6178 ( \6404 , \6402 , \6403 );
xnor \U$6179 ( \6405 , \6404 , \5878 );
xor \U$6180 ( \6406 , \6401 , \6405 );
xor \U$6181 ( \6407 , \6392 , \6406 );
not \U$6182 ( \6408 , \5775 );
and \U$6183 ( \6409 , \5770 , \5790 );
and \U$6184 ( \6410 , \5737 , \5788 );
nor \U$6185 ( \6411 , \6409 , \6410 );
xnor \U$6186 ( \6412 , \6411 , \5797 );
xor \U$6187 ( \6413 , \6408 , \6412 );
and \U$6188 ( \6414 , \5792 , \5809 );
and \U$6189 ( \6415 , \5758 , \5807 );
nor \U$6190 ( \6416 , \6414 , \6415 );
xnor \U$6191 ( \6417 , \6416 , \5816 );
xor \U$6192 ( \6418 , \6413 , \6417 );
xor \U$6193 ( \6419 , \6407 , \6418 );
xor \U$6194 ( \6420 , \6378 , \6419 );
and \U$6195 ( \6421 , \6057 , \6082 );
and \U$6196 ( \6422 , \6029 , \6066 );
nor \U$6197 ( \6423 , \6421 , \6422 );
xnor \U$6198 ( \6424 , \6423 , \5736 );
xor \U$6199 ( \6425 , \6221 , \6224 );
not \U$6200 ( \6426 , \6295 );
and \U$6201 ( \6427 , \6425 , \6426 );
and \U$6202 ( \6428 , \6065 , \6427 );
and \U$6203 ( \6429 , \6048 , \6295 );
nor \U$6204 ( \6430 , \6428 , \6429 );
xnor \U$6205 ( \6431 , \6430 , \6227 );
xor \U$6206 ( \6432 , \6424 , \6431 );
and \U$6207 ( \6433 , \5998 , \6016 );
and \U$6208 ( \6434 , \5967 , \6014 );
nor \U$6209 ( \6435 , \6433 , \6434 );
xnor \U$6210 ( \6436 , \6435 , \6023 );
and \U$6211 ( \6437 , \6018 , \6039 );
and \U$6212 ( \6438 , \5986 , \6037 );
nor \U$6213 ( \6439 , \6437 , \6438 );
xnor \U$6214 ( \6440 , \6439 , \6046 );
xor \U$6215 ( \6441 , \6436 , \6440 );
and \U$6216 ( \6442 , \6041 , \6055 );
and \U$6217 ( \6443 , \6006 , \6053 );
nor \U$6218 ( \6444 , \6442 , \6443 );
xnor \U$6219 ( \6445 , \6444 , \6062 );
xor \U$6220 ( \6446 , \6441 , \6445 );
xor \U$6221 ( \6447 , \6432 , \6446 );
and \U$6222 ( \6448 , \5937 , \5955 );
and \U$6223 ( \6449 , \5906 , \5953 );
nor \U$6224 ( \6450 , \6448 , \6449 );
xnor \U$6225 ( \6451 , \6450 , \5962 );
and \U$6226 ( \6452 , \5957 , \5977 );
and \U$6227 ( \6453 , \5925 , \5975 );
nor \U$6228 ( \6454 , \6452 , \6453 );
xnor \U$6229 ( \6455 , \6454 , \5984 );
xor \U$6230 ( \6456 , \6451 , \6455 );
and \U$6231 ( \6457 , \5979 , \5996 );
and \U$6232 ( \6458 , \5945 , \5994 );
nor \U$6233 ( \6459 , \6457 , \6458 );
xnor \U$6234 ( \6460 , \6459 , \6003 );
xor \U$6235 ( \6461 , \6456 , \6460 );
xor \U$6236 ( \6462 , \6447 , \6461 );
xor \U$6237 ( \6463 , \6420 , \6462 );
and \U$6238 ( \6464 , \6374 , \6463 );
and \U$6239 ( \6465 , \6329 , \6333 );
and \U$6240 ( \6466 , \6333 , \6338 );
and \U$6241 ( \6467 , \6329 , \6338 );
or \U$6242 ( \6468 , \6465 , \6466 , \6467 );
and \U$6243 ( \6469 , \6317 , \6321 );
and \U$6244 ( \6470 , \6321 , \6323 );
and \U$6245 ( \6471 , \6317 , \6323 );
or \U$6246 ( \6472 , \6469 , \6470 , \6471 );
xor \U$6247 ( \6473 , \6468 , \6472 );
or \U$6248 ( \6474 , \6298 , \6312 );
xor \U$6249 ( \6475 , \6473 , \6474 );
and \U$6250 ( \6476 , \6463 , \6475 );
and \U$6251 ( \6477 , \6374 , \6475 );
or \U$6252 ( \6478 , \6464 , \6476 , \6477 );
and \U$6253 ( \6479 , \6345 , \6478 );
and \U$6254 ( \6480 , \6029 , \6082 );
and \U$6255 ( \6481 , \6041 , \6066 );
nor \U$6256 ( \6482 , \6480 , \6481 );
xnor \U$6257 ( \6483 , \6482 , \5736 );
and \U$6258 ( \6484 , \6048 , \6427 );
and \U$6259 ( \6485 , \6057 , \6295 );
nor \U$6260 ( \6486 , \6484 , \6485 );
xnor \U$6261 ( \6487 , \6486 , \6227 );
xor \U$6262 ( \6488 , \6483 , \6487 );
and \U$6263 ( \6489 , \6186 , \6190 );
and \U$6264 ( \6490 , \6190 , \6192 );
and \U$6265 ( \6491 , \6186 , \6192 );
or \U$6266 ( \6492 , \6489 , \6490 , \6491 );
and \U$6267 ( \6493 , \289 , \348 );
not \U$6268 ( \6494 , \6493 );
xnor \U$6269 ( \6495 , \6494 , \356 );
and \U$6270 ( \6496 , \313 , \343 );
xnor \U$6271 ( \6497 , \6495 , \6496 );
xor \U$6272 ( \6498 , \6492 , \6497 );
and \U$6273 ( \6499 , \6177 , \6184 );
and \U$6274 ( \6500 , \6184 , \6193 );
and \U$6275 ( \6501 , \6177 , \6193 );
or \U$6276 ( \6502 , \6499 , \6500 , \6501 );
xor \U$6277 ( \6503 , \6498 , \6502 );
and \U$6278 ( \6504 , \6194 , \6207 );
and \U$6279 ( \6505 , \6208 , \6218 );
or \U$6280 ( \6506 , \6504 , \6505 );
xor \U$6281 ( \6507 , \6503 , \6506 );
buf g16b6_GF_PartitionCandidate( \6508_nG16b6 , \6507 );
buf \U$6282 ( \6509 , \6508_nG16b6 );
xor \U$6283 ( \6510 , \6509 , \6221 );
nand \U$6284 ( \6511 , \6065 , \6510 );
or \U$6285 ( \6512 , \6495 , \6496 );
not \U$6286 ( \6513 , \356 );
xor \U$6287 ( \6514 , \6512 , \6513 );
and \U$6288 ( \6515 , \289 , \343 );
xor \U$6289 ( \6516 , \6514 , \6515 );
and \U$6290 ( \6517 , \6492 , \6497 );
xor \U$6291 ( \6518 , \6516 , \6517 );
and \U$6292 ( \6519 , \6498 , \6502 );
and \U$6293 ( \6520 , \6503 , \6506 );
or \U$6294 ( \6521 , \6519 , \6520 );
xor \U$6295 ( \6522 , \6518 , \6521 );
buf g16b3_GF_PartitionCandidate( \6523_nG16b3 , \6522 );
buf \U$6296 ( \6524 , \6523_nG16b3 );
and \U$6297 ( \6525 , \6509 , \6221 );
not \U$6298 ( \6526 , \6525 );
and \U$6299 ( \6527 , \6524 , \6526 );
xnor \U$6300 ( \6528 , \6511 , \6527 );
xor \U$6301 ( \6529 , \6488 , \6528 );
and \U$6302 ( \6530 , \5967 , \6016 );
and \U$6303 ( \6531 , \5979 , \6014 );
nor \U$6304 ( \6532 , \6530 , \6531 );
xnor \U$6305 ( \6533 , \6532 , \6023 );
and \U$6306 ( \6534 , \5986 , \6039 );
and \U$6307 ( \6535 , \5998 , \6037 );
nor \U$6308 ( \6536 , \6534 , \6535 );
xnor \U$6309 ( \6537 , \6536 , \6046 );
xor \U$6310 ( \6538 , \6533 , \6537 );
and \U$6311 ( \6539 , \6006 , \6055 );
and \U$6312 ( \6540 , \6018 , \6053 );
nor \U$6313 ( \6541 , \6539 , \6540 );
xnor \U$6314 ( \6542 , \6541 , \6062 );
xor \U$6315 ( \6543 , \6538 , \6542 );
xnor \U$6316 ( \6544 , \6529 , \6543 );
and \U$6317 ( \6545 , \6451 , \6455 );
and \U$6318 ( \6546 , \6455 , \6460 );
and \U$6319 ( \6547 , \6451 , \6460 );
or \U$6320 ( \6548 , \6545 , \6546 , \6547 );
and \U$6321 ( \6549 , \6436 , \6440 );
and \U$6322 ( \6550 , \6440 , \6445 );
and \U$6323 ( \6551 , \6436 , \6445 );
or \U$6324 ( \6552 , \6549 , \6550 , \6551 );
xor \U$6325 ( \6553 , \6548 , \6552 );
and \U$6326 ( \6554 , \6424 , \6431 );
xor \U$6327 ( \6555 , \6553 , \6554 );
xor \U$6328 ( \6556 , \6544 , \6555 );
and \U$6329 ( \6557 , \6408 , \6412 );
and \U$6330 ( \6558 , \6412 , \6417 );
and \U$6331 ( \6559 , \6408 , \6417 );
or \U$6332 ( \6560 , \6557 , \6558 , \6559 );
and \U$6333 ( \6561 , \6396 , \6400 );
and \U$6334 ( \6562 , \6400 , \6405 );
and \U$6335 ( \6563 , \6396 , \6405 );
or \U$6336 ( \6564 , \6561 , \6562 , \6563 );
xor \U$6337 ( \6565 , \6560 , \6564 );
and \U$6338 ( \6566 , \6382 , \6386 );
and \U$6339 ( \6567 , \6386 , \6391 );
and \U$6340 ( \6568 , \6382 , \6391 );
or \U$6341 ( \6569 , \6566 , \6567 , \6568 );
xor \U$6342 ( \6570 , \6565 , \6569 );
xor \U$6343 ( \6571 , \6556 , \6570 );
and \U$6344 ( \6572 , \6392 , \6406 );
and \U$6345 ( \6573 , \6406 , \6418 );
and \U$6346 ( \6574 , \6392 , \6418 );
or \U$6347 ( \6575 , \6572 , \6573 , \6574 );
and \U$6348 ( \6576 , \5737 , \5790 );
not \U$6349 ( \6577 , \6576 );
xnor \U$6350 ( \6578 , \6577 , \5797 );
xor \U$6351 ( \6579 , \6527 , \6578 );
and \U$6352 ( \6580 , \5758 , \5809 );
and \U$6353 ( \6581 , \5770 , \5807 );
nor \U$6354 ( \6582 , \6580 , \6581 );
xnor \U$6355 ( \6583 , \6582 , \5816 );
xor \U$6356 ( \6584 , \6579 , \6583 );
xor \U$6357 ( \6585 , \6575 , \6584 );
and \U$6358 ( \6586 , \5906 , \5955 );
and \U$6359 ( \6587 , \5918 , \5953 );
nor \U$6360 ( \6588 , \6586 , \6587 );
xnor \U$6361 ( \6589 , \6588 , \5962 );
and \U$6362 ( \6590 , \5925 , \5977 );
and \U$6363 ( \6591 , \5937 , \5975 );
nor \U$6364 ( \6592 , \6590 , \6591 );
xnor \U$6365 ( \6593 , \6592 , \5984 );
xor \U$6366 ( \6594 , \6589 , \6593 );
and \U$6367 ( \6595 , \5945 , \5996 );
and \U$6368 ( \6596 , \5957 , \5994 );
nor \U$6369 ( \6597 , \6595 , \6596 );
xnor \U$6370 ( \6598 , \6597 , \6003 );
xor \U$6371 ( \6599 , \6594 , \6598 );
and \U$6372 ( \6600 , \5842 , \5891 );
and \U$6373 ( \6601 , \5854 , \5889 );
nor \U$6374 ( \6602 , \6600 , \6601 );
xnor \U$6375 ( \6603 , \6602 , \5898 );
and \U$6376 ( \6604 , \5861 , \5916 );
and \U$6377 ( \6605 , \5873 , \5914 );
nor \U$6378 ( \6606 , \6604 , \6605 );
xnor \U$6379 ( \6607 , \6606 , \5923 );
xor \U$6380 ( \6608 , \6603 , \6607 );
and \U$6381 ( \6609 , \5881 , \5935 );
and \U$6382 ( \6610 , \5893 , \5933 );
nor \U$6383 ( \6611 , \6609 , \6610 );
xnor \U$6384 ( \6612 , \6611 , \5942 );
xor \U$6385 ( \6613 , \6608 , \6612 );
xor \U$6386 ( \6614 , \6599 , \6613 );
and \U$6387 ( \6615 , \5780 , \5829 );
and \U$6388 ( \6616 , \5792 , \5827 );
nor \U$6389 ( \6617 , \6615 , \6616 );
xnor \U$6390 ( \6618 , \6617 , \5836 );
and \U$6391 ( \6619 , \5799 , \5852 );
and \U$6392 ( \6620 , \5811 , \5850 );
nor \U$6393 ( \6621 , \6619 , \6620 );
xnor \U$6394 ( \6622 , \6621 , \5859 );
xor \U$6395 ( \6623 , \6618 , \6622 );
and \U$6396 ( \6624 , \5819 , \5871 );
and \U$6397 ( \6625 , \5831 , \5869 );
nor \U$6398 ( \6626 , \6624 , \6625 );
xnor \U$6399 ( \6627 , \6626 , \5878 );
xor \U$6400 ( \6628 , \6623 , \6627 );
xor \U$6401 ( \6629 , \6614 , \6628 );
xor \U$6402 ( \6630 , \6585 , \6629 );
xor \U$6403 ( \6631 , \6571 , \6630 );
and \U$6404 ( \6632 , \6363 , \6367 );
and \U$6405 ( \6633 , \6367 , \6372 );
and \U$6406 ( \6634 , \6363 , \6372 );
or \U$6407 ( \6635 , \6632 , \6633 , \6634 );
and \U$6408 ( \6636 , \6349 , \6353 );
and \U$6409 ( \6637 , \6353 , \6358 );
and \U$6410 ( \6638 , \6349 , \6358 );
or \U$6411 ( \6639 , \6636 , \6637 , \6638 );
xor \U$6412 ( \6640 , \6635 , \6639 );
and \U$6413 ( \6641 , \6432 , \6446 );
and \U$6414 ( \6642 , \6446 , \6461 );
and \U$6415 ( \6643 , \6432 , \6461 );
or \U$6416 ( \6644 , \6641 , \6642 , \6643 );
xor \U$6417 ( \6645 , \6640 , \6644 );
xor \U$6418 ( \6646 , \6631 , \6645 );
and \U$6419 ( \6647 , \6478 , \6646 );
and \U$6420 ( \6648 , \6345 , \6646 );
or \U$6421 ( \6649 , \6479 , \6647 , \6648 );
and \U$6422 ( \6650 , \6635 , \6639 );
and \U$6423 ( \6651 , \6639 , \6644 );
and \U$6424 ( \6652 , \6635 , \6644 );
or \U$6425 ( \6653 , \6650 , \6651 , \6652 );
and \U$6426 ( \6654 , \6575 , \6584 );
and \U$6427 ( \6655 , \6584 , \6629 );
and \U$6428 ( \6656 , \6575 , \6629 );
or \U$6429 ( \6657 , \6654 , \6655 , \6656 );
xor \U$6430 ( \6658 , \6653 , \6657 );
and \U$6431 ( \6659 , \6544 , \6555 );
and \U$6432 ( \6660 , \6555 , \6570 );
and \U$6433 ( \6661 , \6544 , \6570 );
or \U$6434 ( \6662 , \6659 , \6660 , \6661 );
xor \U$6435 ( \6663 , \6658 , \6662 );
xor \U$6436 ( \6664 , \6649 , \6663 );
and \U$6437 ( \6665 , \6468 , \6472 );
and \U$6438 ( \6666 , \6472 , \6474 );
and \U$6439 ( \6667 , \6468 , \6474 );
or \U$6440 ( \6668 , \6665 , \6666 , \6667 );
and \U$6441 ( \6669 , \6378 , \6419 );
and \U$6442 ( \6670 , \6419 , \6462 );
and \U$6443 ( \6671 , \6378 , \6462 );
or \U$6444 ( \6672 , \6669 , \6670 , \6671 );
and \U$6445 ( \6673 , \6668 , \6672 );
and \U$6446 ( \6674 , \6359 , \6373 );
and \U$6447 ( \6675 , \6672 , \6674 );
and \U$6448 ( \6676 , \6668 , \6674 );
or \U$6449 ( \6677 , \6673 , \6675 , \6676 );
and \U$6450 ( \6678 , \6571 , \6630 );
and \U$6451 ( \6679 , \6630 , \6645 );
and \U$6452 ( \6680 , \6571 , \6645 );
or \U$6453 ( \6681 , \6678 , \6679 , \6680 );
xor \U$6454 ( \6682 , \6677 , \6681 );
and \U$6455 ( \6683 , \6589 , \6593 );
and \U$6456 ( \6684 , \6593 , \6598 );
and \U$6457 ( \6685 , \6589 , \6598 );
or \U$6458 ( \6686 , \6683 , \6684 , \6685 );
and \U$6459 ( \6687 , \6533 , \6537 );
and \U$6460 ( \6688 , \6537 , \6542 );
and \U$6461 ( \6689 , \6533 , \6542 );
or \U$6462 ( \6690 , \6687 , \6688 , \6689 );
xor \U$6463 ( \6691 , \6686 , \6690 );
and \U$6464 ( \6692 , \6483 , \6487 );
and \U$6465 ( \6693 , \6487 , \6528 );
and \U$6466 ( \6694 , \6483 , \6528 );
or \U$6467 ( \6695 , \6692 , \6693 , \6694 );
xor \U$6468 ( \6696 , \6691 , \6695 );
and \U$6469 ( \6697 , \6527 , \6578 );
and \U$6470 ( \6698 , \6578 , \6583 );
and \U$6471 ( \6699 , \6527 , \6583 );
or \U$6472 ( \6700 , \6697 , \6698 , \6699 );
and \U$6473 ( \6701 , \6618 , \6622 );
and \U$6474 ( \6702 , \6622 , \6627 );
and \U$6475 ( \6703 , \6618 , \6627 );
or \U$6476 ( \6704 , \6701 , \6702 , \6703 );
xor \U$6477 ( \6705 , \6700 , \6704 );
and \U$6478 ( \6706 , \6603 , \6607 );
and \U$6479 ( \6707 , \6607 , \6612 );
and \U$6480 ( \6708 , \6603 , \6612 );
or \U$6481 ( \6709 , \6706 , \6707 , \6708 );
xor \U$6482 ( \6710 , \6705 , \6709 );
xor \U$6483 ( \6711 , \6696 , \6710 );
and \U$6484 ( \6712 , \6599 , \6613 );
and \U$6485 ( \6713 , \6613 , \6628 );
and \U$6486 ( \6714 , \6599 , \6628 );
or \U$6487 ( \6715 , \6712 , \6713 , \6714 );
and \U$6488 ( \6716 , \5873 , \5916 );
and \U$6489 ( \6717 , \5842 , \5914 );
nor \U$6490 ( \6718 , \6716 , \6717 );
xnor \U$6491 ( \6719 , \6718 , \5923 );
and \U$6492 ( \6720 , \5893 , \5935 );
and \U$6493 ( \6721 , \5861 , \5933 );
nor \U$6494 ( \6722 , \6720 , \6721 );
xnor \U$6495 ( \6723 , \6722 , \5942 );
xor \U$6496 ( \6724 , \6719 , \6723 );
and \U$6497 ( \6725 , \5918 , \5955 );
and \U$6498 ( \6726 , \5881 , \5953 );
nor \U$6499 ( \6727 , \6725 , \6726 );
xnor \U$6500 ( \6728 , \6727 , \5962 );
xor \U$6501 ( \6729 , \6724 , \6728 );
and \U$6502 ( \6730 , \5811 , \5852 );
and \U$6503 ( \6731 , \5780 , \5850 );
nor \U$6504 ( \6732 , \6730 , \6731 );
xnor \U$6505 ( \6733 , \6732 , \5859 );
and \U$6506 ( \6734 , \5831 , \5871 );
and \U$6507 ( \6735 , \5799 , \5869 );
nor \U$6508 ( \6736 , \6734 , \6735 );
xnor \U$6509 ( \6737 , \6736 , \5878 );
xor \U$6510 ( \6738 , \6733 , \6737 );
and \U$6511 ( \6739 , \5854 , \5891 );
and \U$6512 ( \6740 , \5819 , \5889 );
nor \U$6513 ( \6741 , \6739 , \6740 );
xnor \U$6514 ( \6742 , \6741 , \5898 );
xor \U$6515 ( \6743 , \6738 , \6742 );
xor \U$6516 ( \6744 , \6729 , \6743 );
not \U$6517 ( \6745 , \5797 );
and \U$6518 ( \6746 , \5770 , \5809 );
and \U$6519 ( \6747 , \5737 , \5807 );
nor \U$6520 ( \6748 , \6746 , \6747 );
xnor \U$6521 ( \6749 , \6748 , \5816 );
xor \U$6522 ( \6750 , \6745 , \6749 );
and \U$6523 ( \6751 , \5792 , \5829 );
and \U$6524 ( \6752 , \5758 , \5827 );
nor \U$6525 ( \6753 , \6751 , \6752 );
xnor \U$6526 ( \6754 , \6753 , \5836 );
xor \U$6527 ( \6755 , \6750 , \6754 );
xor \U$6528 ( \6756 , \6744 , \6755 );
xor \U$6529 ( \6757 , \6715 , \6756 );
and \U$6530 ( \6758 , \6057 , \6427 );
and \U$6531 ( \6759 , \6029 , \6295 );
nor \U$6532 ( \6760 , \6758 , \6759 );
xnor \U$6533 ( \6761 , \6760 , \6227 );
xor \U$6534 ( \6762 , \6524 , \6509 );
not \U$6535 ( \6763 , \6510 );
and \U$6536 ( \6764 , \6762 , \6763 );
and \U$6537 ( \6765 , \6065 , \6764 );
and \U$6538 ( \6766 , \6048 , \6510 );
nor \U$6539 ( \6767 , \6765 , \6766 );
xnor \U$6540 ( \6768 , \6767 , \6527 );
xor \U$6541 ( \6769 , \6761 , \6768 );
and \U$6542 ( \6770 , \5998 , \6039 );
and \U$6543 ( \6771 , \5967 , \6037 );
nor \U$6544 ( \6772 , \6770 , \6771 );
xnor \U$6545 ( \6773 , \6772 , \6046 );
and \U$6546 ( \6774 , \6018 , \6055 );
and \U$6547 ( \6775 , \5986 , \6053 );
nor \U$6548 ( \6776 , \6774 , \6775 );
xnor \U$6549 ( \6777 , \6776 , \6062 );
xor \U$6550 ( \6778 , \6773 , \6777 );
and \U$6551 ( \6779 , \6041 , \6082 );
and \U$6552 ( \6780 , \6006 , \6066 );
nor \U$6553 ( \6781 , \6779 , \6780 );
xnor \U$6554 ( \6782 , \6781 , \5736 );
xor \U$6555 ( \6783 , \6778 , \6782 );
xor \U$6556 ( \6784 , \6769 , \6783 );
and \U$6557 ( \6785 , \5937 , \5977 );
and \U$6558 ( \6786 , \5906 , \5975 );
nor \U$6559 ( \6787 , \6785 , \6786 );
xnor \U$6560 ( \6788 , \6787 , \5984 );
and \U$6561 ( \6789 , \5957 , \5996 );
and \U$6562 ( \6790 , \5925 , \5994 );
nor \U$6563 ( \6791 , \6789 , \6790 );
xnor \U$6564 ( \6792 , \6791 , \6003 );
xor \U$6565 ( \6793 , \6788 , \6792 );
and \U$6566 ( \6794 , \5979 , \6016 );
and \U$6567 ( \6795 , \5945 , \6014 );
nor \U$6568 ( \6796 , \6794 , \6795 );
xnor \U$6569 ( \6797 , \6796 , \6023 );
xor \U$6570 ( \6798 , \6793 , \6797 );
xor \U$6571 ( \6799 , \6784 , \6798 );
xor \U$6572 ( \6800 , \6757 , \6799 );
xor \U$6573 ( \6801 , \6711 , \6800 );
and \U$6574 ( \6802 , \6560 , \6564 );
and \U$6575 ( \6803 , \6564 , \6569 );
and \U$6576 ( \6804 , \6560 , \6569 );
or \U$6577 ( \6805 , \6802 , \6803 , \6804 );
and \U$6578 ( \6806 , \6548 , \6552 );
and \U$6579 ( \6807 , \6552 , \6554 );
and \U$6580 ( \6808 , \6548 , \6554 );
or \U$6581 ( \6809 , \6806 , \6807 , \6808 );
xor \U$6582 ( \6810 , \6805 , \6809 );
or \U$6583 ( \6811 , \6529 , \6543 );
xor \U$6584 ( \6812 , \6810 , \6811 );
xor \U$6585 ( \6813 , \6801 , \6812 );
xor \U$6586 ( \6814 , \6682 , \6813 );
xor \U$6587 ( \6815 , \6664 , \6814 );
xor \U$6588 ( \6816 , \4668 , \5654 );
buf g1728_GF_PartitionCandidate( \6817_nG1728 , \6816 );
buf \U$6589 ( \6818 , \6817_nG1728 );
xor \U$6590 ( \6819 , \4760 , \5652 );
buf g172b_GF_PartitionCandidate( \6820_nG172b , \6819 );
buf \U$6591 ( \6821 , \6820_nG172b );
and \U$6592 ( \6822 , \6818 , \6821 );
not \U$6593 ( \6823 , \6822 );
and \U$6594 ( \6824 , \5747 , \6823 );
not \U$6595 ( \6825 , \6824 );
and \U$6596 ( \6826 , \5770 , \5750 );
and \U$6597 ( \6827 , \5737 , \5748 );
nor \U$6598 ( \6828 , \6826 , \6827 );
xnor \U$6599 ( \6829 , \6828 , \5755 );
and \U$6600 ( \6830 , \6825 , \6829 );
and \U$6601 ( \6831 , \5792 , \5768 );
and \U$6602 ( \6832 , \5758 , \5766 );
nor \U$6603 ( \6833 , \6831 , \6832 );
xnor \U$6604 ( \6834 , \6833 , \5775 );
and \U$6605 ( \6835 , \6829 , \6834 );
and \U$6606 ( \6836 , \6825 , \6834 );
or \U$6607 ( \6837 , \6830 , \6835 , \6836 );
and \U$6608 ( \6838 , \5811 , \5790 );
and \U$6609 ( \6839 , \5780 , \5788 );
nor \U$6610 ( \6840 , \6838 , \6839 );
xnor \U$6611 ( \6841 , \6840 , \5797 );
and \U$6612 ( \6842 , \5831 , \5809 );
and \U$6613 ( \6843 , \5799 , \5807 );
nor \U$6614 ( \6844 , \6842 , \6843 );
xnor \U$6615 ( \6845 , \6844 , \5816 );
and \U$6616 ( \6846 , \6841 , \6845 );
and \U$6617 ( \6847 , \5854 , \5829 );
and \U$6618 ( \6848 , \5819 , \5827 );
nor \U$6619 ( \6849 , \6847 , \6848 );
xnor \U$6620 ( \6850 , \6849 , \5836 );
and \U$6621 ( \6851 , \6845 , \6850 );
and \U$6622 ( \6852 , \6841 , \6850 );
or \U$6623 ( \6853 , \6846 , \6851 , \6852 );
and \U$6624 ( \6854 , \6837 , \6853 );
and \U$6625 ( \6855 , \5873 , \5852 );
and \U$6626 ( \6856 , \5842 , \5850 );
nor \U$6627 ( \6857 , \6855 , \6856 );
xnor \U$6628 ( \6858 , \6857 , \5859 );
and \U$6629 ( \6859 , \5893 , \5871 );
and \U$6630 ( \6860 , \5861 , \5869 );
nor \U$6631 ( \6861 , \6859 , \6860 );
xnor \U$6632 ( \6862 , \6861 , \5878 );
and \U$6633 ( \6863 , \6858 , \6862 );
and \U$6634 ( \6864 , \5918 , \5891 );
and \U$6635 ( \6865 , \5881 , \5889 );
nor \U$6636 ( \6866 , \6864 , \6865 );
xnor \U$6637 ( \6867 , \6866 , \5898 );
and \U$6638 ( \6868 , \6862 , \6867 );
and \U$6639 ( \6869 , \6858 , \6867 );
or \U$6640 ( \6870 , \6863 , \6868 , \6869 );
and \U$6641 ( \6871 , \6853 , \6870 );
and \U$6642 ( \6872 , \6837 , \6870 );
or \U$6643 ( \6873 , \6854 , \6871 , \6872 );
and \U$6644 ( \6874 , \5937 , \5916 );
and \U$6645 ( \6875 , \5906 , \5914 );
nor \U$6646 ( \6876 , \6874 , \6875 );
xnor \U$6647 ( \6877 , \6876 , \5923 );
and \U$6648 ( \6878 , \5957 , \5935 );
and \U$6649 ( \6879 , \5925 , \5933 );
nor \U$6650 ( \6880 , \6878 , \6879 );
xnor \U$6651 ( \6881 , \6880 , \5942 );
and \U$6652 ( \6882 , \6877 , \6881 );
and \U$6653 ( \6883 , \5979 , \5955 );
and \U$6654 ( \6884 , \5945 , \5953 );
nor \U$6655 ( \6885 , \6883 , \6884 );
xnor \U$6656 ( \6886 , \6885 , \5962 );
and \U$6657 ( \6887 , \6881 , \6886 );
and \U$6658 ( \6888 , \6877 , \6886 );
or \U$6659 ( \6889 , \6882 , \6887 , \6888 );
and \U$6660 ( \6890 , \5998 , \5977 );
and \U$6661 ( \6891 , \5967 , \5975 );
nor \U$6662 ( \6892 , \6890 , \6891 );
xnor \U$6663 ( \6893 , \6892 , \5984 );
and \U$6664 ( \6894 , \6018 , \5996 );
and \U$6665 ( \6895 , \5986 , \5994 );
nor \U$6666 ( \6896 , \6894 , \6895 );
xnor \U$6667 ( \6897 , \6896 , \6003 );
and \U$6668 ( \6898 , \6893 , \6897 );
and \U$6669 ( \6899 , \6041 , \6016 );
and \U$6670 ( \6900 , \6006 , \6014 );
nor \U$6671 ( \6901 , \6899 , \6900 );
xnor \U$6672 ( \6902 , \6901 , \6023 );
and \U$6673 ( \6903 , \6897 , \6902 );
and \U$6674 ( \6904 , \6893 , \6902 );
or \U$6675 ( \6905 , \6898 , \6903 , \6904 );
and \U$6676 ( \6906 , \6889 , \6905 );
and \U$6677 ( \6907 , \6057 , \6039 );
and \U$6678 ( \6908 , \6029 , \6037 );
nor \U$6679 ( \6909 , \6907 , \6908 );
xnor \U$6680 ( \6910 , \6909 , \6046 );
and \U$6681 ( \6911 , \6065 , \6055 );
and \U$6682 ( \6912 , \6048 , \6053 );
nor \U$6683 ( \6913 , \6911 , \6912 );
xnor \U$6684 ( \6914 , \6913 , \6062 );
and \U$6685 ( \6915 , \6910 , \6914 );
and \U$6686 ( \6916 , \6905 , \6915 );
and \U$6687 ( \6917 , \6889 , \6915 );
or \U$6688 ( \6918 , \6906 , \6916 , \6917 );
and \U$6689 ( \6919 , \6873 , \6918 );
xor \U$6690 ( \6920 , \6047 , \6063 );
xor \U$6691 ( \6921 , \6920 , \6068 );
xor \U$6692 ( \6922 , \5985 , \6004 );
xor \U$6693 ( \6923 , \6922 , \6024 );
or \U$6694 ( \6924 , \6921 , \6923 );
and \U$6695 ( \6925 , \6918 , \6924 );
and \U$6696 ( \6926 , \6873 , \6924 );
or \U$6697 ( \6927 , \6919 , \6925 , \6926 );
xor \U$6698 ( \6928 , \5924 , \5943 );
xor \U$6699 ( \6929 , \6928 , \5963 );
xor \U$6700 ( \6930 , \5860 , \5879 );
xor \U$6701 ( \6931 , \6930 , \5899 );
and \U$6702 ( \6932 , \6929 , \6931 );
xor \U$6703 ( \6933 , \5798 , \5817 );
xor \U$6704 ( \6934 , \6933 , \5837 );
and \U$6705 ( \6935 , \6931 , \6934 );
and \U$6706 ( \6936 , \6929 , \6934 );
or \U$6707 ( \6937 , \6932 , \6935 , \6936 );
xor \U$6708 ( \6938 , \6136 , \6150 );
xor \U$6709 ( \6939 , \6938 , \6162 );
and \U$6710 ( \6940 , \6937 , \6939 );
xor \U$6711 ( \6941 , \6087 , \6101 );
xor \U$6712 ( \6942 , \6941 , \6116 );
and \U$6713 ( \6943 , \6939 , \6942 );
and \U$6714 ( \6944 , \6937 , \6942 );
or \U$6715 ( \6945 , \6940 , \6943 , \6944 );
and \U$6716 ( \6946 , \6927 , \6945 );
xor \U$6717 ( \6947 , \5966 , \6027 );
xor \U$6718 ( \6948 , \6947 , \6071 );
xor \U$6719 ( \6949 , \5779 , \5840 );
xor \U$6720 ( \6950 , \6949 , \5902 );
and \U$6721 ( \6951 , \6948 , \6950 );
and \U$6722 ( \6952 , \6945 , \6951 );
and \U$6723 ( \6953 , \6927 , \6951 );
or \U$6724 ( \6954 , \6946 , \6952 , \6953 );
xor \U$6725 ( \6955 , \6313 , \6324 );
xor \U$6726 ( \6956 , \6955 , \6339 );
xor \U$6727 ( \6957 , \6165 , \6236 );
xor \U$6728 ( \6958 , \6957 , \6281 );
and \U$6729 ( \6959 , \6956 , \6958 );
xor \U$6730 ( \6960 , \5905 , \6074 );
xor \U$6731 ( \6961 , \6960 , \6119 );
and \U$6732 ( \6962 , \6958 , \6961 );
and \U$6733 ( \6963 , \6956 , \6961 );
or \U$6734 ( \6964 , \6959 , \6962 , \6963 );
and \U$6735 ( \6965 , \6954 , \6964 );
xor \U$6736 ( \6966 , \6374 , \6463 );
xor \U$6737 ( \6967 , \6966 , \6475 );
and \U$6738 ( \6968 , \6964 , \6967 );
and \U$6739 ( \6969 , \6954 , \6967 );
or \U$6740 ( \6970 , \6965 , \6968 , \6969 );
xor \U$6741 ( \6971 , \6668 , \6672 );
xor \U$6742 ( \6972 , \6971 , \6674 );
and \U$6743 ( \6973 , \6970 , \6972 );
xor \U$6744 ( \6974 , \6345 , \6478 );
xor \U$6745 ( \6975 , \6974 , \6646 );
and \U$6746 ( \6976 , \6972 , \6975 );
and \U$6747 ( \6977 , \6970 , \6975 );
or \U$6748 ( \6978 , \6973 , \6976 , \6977 );
nand \U$6749 ( \6979 , \6815 , \6978 );
nor \U$6750 ( \6980 , \6815 , \6978 );
not \U$6751 ( \6981 , \6980 );
nand \U$6752 ( \6982 , \6979 , \6981 );
xor \U$6753 ( \6983 , \5606 , \5609 );
buf g176d_GF_PartitionCandidate( \6984_nG176d , \6983 );
buf \U$6754 ( \6985 , \6984_nG176d );
xor \U$6755 ( \6986 , \5608 , \2368 );
buf g1770_GF_PartitionCandidate( \6987_nG1770 , \6986 );
buf \U$6756 ( \6988 , \6987_nG1770 );
xor \U$6757 ( \6989 , \6985 , \6988 );
not \U$6758 ( \6990 , \6988 );
and \U$6759 ( \6991 , \6989 , \6990 );
and \U$6760 ( \6992 , \5799 , \6991 );
and \U$6761 ( \6993 , \5811 , \6988 );
nor \U$6762 ( \6994 , \6992 , \6993 );
xnor \U$6763 ( \6995 , \6994 , \6985 );
and \U$6764 ( \6996 , \5755 , \6995 );
xor \U$6765 ( \6997 , \5597 , \5612 );
buf g1767_GF_PartitionCandidate( \6998_nG1767 , \6997 );
buf \U$6766 ( \6999 , \6998_nG1767 );
xor \U$6767 ( \7000 , \5602 , \5610 );
buf g176a_GF_PartitionCandidate( \7001_nG176a , \7000 );
buf \U$6768 ( \7002 , \7001_nG176a );
xor \U$6769 ( \7003 , \6999 , \7002 );
xor \U$6770 ( \7004 , \7002 , \6985 );
not \U$6771 ( \7005 , \7004 );
and \U$6772 ( \7006 , \7003 , \7005 );
and \U$6773 ( \7007 , \5819 , \7006 );
and \U$6774 ( \7008 , \5831 , \7004 );
nor \U$6775 ( \7009 , \7007 , \7008 );
and \U$6776 ( \7010 , \7002 , \6985 );
not \U$6777 ( \7011 , \7010 );
and \U$6778 ( \7012 , \6999 , \7011 );
xnor \U$6779 ( \7013 , \7009 , \7012 );
and \U$6780 ( \7014 , \6995 , \7013 );
and \U$6781 ( \7015 , \5755 , \7013 );
or \U$6782 ( \7016 , \6996 , \7014 , \7015 );
xor \U$6783 ( \7017 , \5577 , \5616 );
buf g1761_GF_PartitionCandidate( \7018_nG1761 , \7017 );
buf \U$6784 ( \7019 , \7018_nG1761 );
xor \U$6785 ( \7020 , \5589 , \5614 );
buf g1764_GF_PartitionCandidate( \7021_nG1764 , \7020 );
buf \U$6786 ( \7022 , \7021_nG1764 );
xor \U$6787 ( \7023 , \7019 , \7022 );
xor \U$6788 ( \7024 , \7022 , \6999 );
not \U$6789 ( \7025 , \7024 );
and \U$6790 ( \7026 , \7023 , \7025 );
and \U$6791 ( \7027 , \5842 , \7026 );
and \U$6792 ( \7028 , \5854 , \7024 );
nor \U$6793 ( \7029 , \7027 , \7028 );
and \U$6794 ( \7030 , \7022 , \6999 );
not \U$6795 ( \7031 , \7030 );
and \U$6796 ( \7032 , \7019 , \7031 );
xnor \U$6797 ( \7033 , \7029 , \7032 );
xor \U$6798 ( \7034 , \5550 , \5620 );
buf g175b_GF_PartitionCandidate( \7035_nG175b , \7034 );
buf \U$6799 ( \7036 , \7035_nG175b );
xor \U$6800 ( \7037 , \5569 , \5618 );
buf g175e_GF_PartitionCandidate( \7038_nG175e , \7037 );
buf \U$6801 ( \7039 , \7038_nG175e );
xor \U$6802 ( \7040 , \7036 , \7039 );
xor \U$6803 ( \7041 , \7039 , \7019 );
not \U$6804 ( \7042 , \7041 );
and \U$6805 ( \7043 , \7040 , \7042 );
and \U$6806 ( \7044 , \5861 , \7043 );
and \U$6807 ( \7045 , \5873 , \7041 );
nor \U$6808 ( \7046 , \7044 , \7045 );
and \U$6809 ( \7047 , \7039 , \7019 );
not \U$6810 ( \7048 , \7047 );
and \U$6811 ( \7049 , \7036 , \7048 );
xnor \U$6812 ( \7050 , \7046 , \7049 );
and \U$6813 ( \7051 , \7033 , \7050 );
xor \U$6814 ( \7052 , \5516 , \5624 );
buf g1755_GF_PartitionCandidate( \7053_nG1755 , \7052 );
buf \U$6815 ( \7054 , \7053_nG1755 );
xor \U$6816 ( \7055 , \5524 , \5622 );
buf g1758_GF_PartitionCandidate( \7056_nG1758 , \7055 );
buf \U$6817 ( \7057 , \7056_nG1758 );
xor \U$6818 ( \7058 , \7054 , \7057 );
xor \U$6819 ( \7059 , \7057 , \7036 );
not \U$6820 ( \7060 , \7059 );
and \U$6821 ( \7061 , \7058 , \7060 );
and \U$6822 ( \7062 , \5881 , \7061 );
and \U$6823 ( \7063 , \5893 , \7059 );
nor \U$6824 ( \7064 , \7062 , \7063 );
and \U$6825 ( \7065 , \7057 , \7036 );
not \U$6826 ( \7066 , \7065 );
and \U$6827 ( \7067 , \7054 , \7066 );
xnor \U$6828 ( \7068 , \7064 , \7067 );
and \U$6829 ( \7069 , \7050 , \7068 );
and \U$6830 ( \7070 , \7033 , \7068 );
or \U$6831 ( \7071 , \7051 , \7069 , \7070 );
and \U$6832 ( \7072 , \7016 , \7071 );
xor \U$6833 ( \7073 , \5448 , \5628 );
buf g174f_GF_PartitionCandidate( \7074_nG174f , \7073 );
buf \U$6834 ( \7075 , \7074_nG174f );
xor \U$6835 ( \7076 , \5482 , \5626 );
buf g1752_GF_PartitionCandidate( \7077_nG1752 , \7076 );
buf \U$6836 ( \7078 , \7077_nG1752 );
xor \U$6837 ( \7079 , \7075 , \7078 );
xor \U$6838 ( \7080 , \7078 , \7054 );
not \U$6839 ( \7081 , \7080 );
and \U$6840 ( \7082 , \7079 , \7081 );
and \U$6841 ( \7083 , \5906 , \7082 );
and \U$6842 ( \7084 , \5918 , \7080 );
nor \U$6843 ( \7085 , \7083 , \7084 );
and \U$6844 ( \7086 , \7078 , \7054 );
not \U$6845 ( \7087 , \7086 );
and \U$6846 ( \7088 , \7075 , \7087 );
xnor \U$6847 ( \7089 , \7085 , \7088 );
xor \U$6848 ( \7090 , \5387 , \5632 );
buf g1749_GF_PartitionCandidate( \7091_nG1749 , \7090 );
buf \U$6849 ( \7092 , \7091_nG1749 );
xor \U$6850 ( \7093 , \5440 , \5630 );
buf g174c_GF_PartitionCandidate( \7094_nG174c , \7093 );
buf \U$6851 ( \7095 , \7094_nG174c );
xor \U$6852 ( \7096 , \7092 , \7095 );
xor \U$6853 ( \7097 , \7095 , \7075 );
not \U$6854 ( \7098 , \7097 );
and \U$6855 ( \7099 , \7096 , \7098 );
and \U$6856 ( \7100 , \5925 , \7099 );
and \U$6857 ( \7101 , \5937 , \7097 );
nor \U$6858 ( \7102 , \7100 , \7101 );
and \U$6859 ( \7103 , \7095 , \7075 );
not \U$6860 ( \7104 , \7103 );
and \U$6861 ( \7105 , \7092 , \7104 );
xnor \U$6862 ( \7106 , \7102 , \7105 );
and \U$6863 ( \7107 , \7089 , \7106 );
xor \U$6864 ( \7108 , \5295 , \5636 );
buf g1743_GF_PartitionCandidate( \7109_nG1743 , \7108 );
buf \U$6865 ( \7110 , \7109_nG1743 );
xor \U$6866 ( \7111 , \5348 , \5634 );
buf g1746_GF_PartitionCandidate( \7112_nG1746 , \7111 );
buf \U$6867 ( \7113 , \7112_nG1746 );
xor \U$6868 ( \7114 , \7110 , \7113 );
xor \U$6869 ( \7115 , \7113 , \7092 );
not \U$6870 ( \7116 , \7115 );
and \U$6871 ( \7117 , \7114 , \7116 );
and \U$6872 ( \7118 , \5945 , \7117 );
and \U$6873 ( \7119 , \5957 , \7115 );
nor \U$6874 ( \7120 , \7118 , \7119 );
and \U$6875 ( \7121 , \7113 , \7092 );
not \U$6876 ( \7122 , \7121 );
and \U$6877 ( \7123 , \7110 , \7122 );
xnor \U$6878 ( \7124 , \7120 , \7123 );
and \U$6879 ( \7125 , \7106 , \7124 );
and \U$6880 ( \7126 , \7089 , \7124 );
or \U$6881 ( \7127 , \7107 , \7125 , \7126 );
and \U$6882 ( \7128 , \7071 , \7127 );
and \U$6883 ( \7129 , \7016 , \7127 );
or \U$6884 ( \7130 , \7072 , \7128 , \7129 );
xor \U$6885 ( \7131 , \5169 , \5640 );
buf g173d_GF_PartitionCandidate( \7132_nG173d , \7131 );
buf \U$6886 ( \7133 , \7132_nG173d );
xor \U$6887 ( \7134 , \5224 , \5638 );
buf g1740_GF_PartitionCandidate( \7135_nG1740 , \7134 );
buf \U$6888 ( \7136 , \7135_nG1740 );
xor \U$6889 ( \7137 , \7133 , \7136 );
xor \U$6890 ( \7138 , \7136 , \7110 );
not \U$6891 ( \7139 , \7138 );
and \U$6892 ( \7140 , \7137 , \7139 );
and \U$6893 ( \7141 , \5967 , \7140 );
and \U$6894 ( \7142 , \5979 , \7138 );
nor \U$6895 ( \7143 , \7141 , \7142 );
and \U$6896 ( \7144 , \7136 , \7110 );
not \U$6897 ( \7145 , \7144 );
and \U$6898 ( \7146 , \7133 , \7145 );
xnor \U$6899 ( \7147 , \7143 , \7146 );
xor \U$6900 ( \7148 , \5102 , \5644 );
buf g1737_GF_PartitionCandidate( \7149_nG1737 , \7148 );
buf \U$6901 ( \7150 , \7149_nG1737 );
xor \U$6902 ( \7151 , \5110 , \5642 );
buf g173a_GF_PartitionCandidate( \7152_nG173a , \7151 );
buf \U$6903 ( \7153 , \7152_nG173a );
xor \U$6904 ( \7154 , \7150 , \7153 );
xor \U$6905 ( \7155 , \7153 , \7133 );
not \U$6906 ( \7156 , \7155 );
and \U$6907 ( \7157 , \7154 , \7156 );
and \U$6908 ( \7158 , \5986 , \7157 );
and \U$6909 ( \7159 , \5998 , \7155 );
nor \U$6910 ( \7160 , \7158 , \7159 );
and \U$6911 ( \7161 , \7153 , \7133 );
not \U$6912 ( \7162 , \7161 );
and \U$6913 ( \7163 , \7150 , \7162 );
xnor \U$6914 ( \7164 , \7160 , \7163 );
and \U$6915 ( \7165 , \7147 , \7164 );
xor \U$6916 ( \7166 , \4943 , \5648 );
buf g1731_GF_PartitionCandidate( \7167_nG1731 , \7166 );
buf \U$6917 ( \7168 , \7167_nG1731 );
xor \U$6918 ( \7169 , \5023 , \5646 );
buf g1734_GF_PartitionCandidate( \7170_nG1734 , \7169 );
buf \U$6919 ( \7171 , \7170_nG1734 );
xor \U$6920 ( \7172 , \7168 , \7171 );
xor \U$6921 ( \7173 , \7171 , \7150 );
not \U$6922 ( \7174 , \7173 );
and \U$6923 ( \7175 , \7172 , \7174 );
and \U$6924 ( \7176 , \6006 , \7175 );
and \U$6925 ( \7177 , \6018 , \7173 );
nor \U$6926 ( \7178 , \7176 , \7177 );
and \U$6927 ( \7179 , \7171 , \7150 );
not \U$6928 ( \7180 , \7179 );
and \U$6929 ( \7181 , \7168 , \7180 );
xnor \U$6930 ( \7182 , \7178 , \7181 );
and \U$6931 ( \7183 , \7164 , \7182 );
and \U$6932 ( \7184 , \7147 , \7182 );
or \U$6933 ( \7185 , \7165 , \7183 , \7184 );
xor \U$6934 ( \7186 , \4848 , \5650 );
buf g172e_GF_PartitionCandidate( \7187_nG172e , \7186 );
buf \U$6935 ( \7188 , \7187_nG172e );
xor \U$6936 ( \7189 , \6821 , \7188 );
xor \U$6937 ( \7190 , \7188 , \7168 );
not \U$6938 ( \7191 , \7190 );
and \U$6939 ( \7192 , \7189 , \7191 );
and \U$6940 ( \7193 , \6029 , \7192 );
and \U$6941 ( \7194 , \6041 , \7190 );
nor \U$6942 ( \7195 , \7193 , \7194 );
and \U$6943 ( \7196 , \7188 , \7168 );
not \U$6944 ( \7197 , \7196 );
and \U$6945 ( \7198 , \6821 , \7197 );
xnor \U$6946 ( \7199 , \7195 , \7198 );
xor \U$6947 ( \7200 , \5747 , \6818 );
xor \U$6948 ( \7201 , \6818 , \6821 );
not \U$6949 ( \7202 , \7201 );
and \U$6950 ( \7203 , \7200 , \7202 );
and \U$6951 ( \7204 , \6048 , \7203 );
and \U$6952 ( \7205 , \6057 , \7201 );
nor \U$6953 ( \7206 , \7204 , \7205 );
xnor \U$6954 ( \7207 , \7206 , \6824 );
and \U$6955 ( \7208 , \7199 , \7207 );
nand \U$6956 ( \7209 , \6065 , \5748 );
xnor \U$6957 ( \7210 , \7209 , \5755 );
and \U$6958 ( \7211 , \7207 , \7210 );
and \U$6959 ( \7212 , \7199 , \7210 );
or \U$6960 ( \7213 , \7208 , \7211 , \7212 );
and \U$6961 ( \7214 , \7185 , \7213 );
and \U$6962 ( \7215 , \6057 , \7203 );
and \U$6963 ( \7216 , \6029 , \7201 );
nor \U$6964 ( \7217 , \7215 , \7216 );
xnor \U$6965 ( \7218 , \7217 , \6824 );
and \U$6966 ( \7219 , \7213 , \7218 );
and \U$6967 ( \7220 , \7185 , \7218 );
or \U$6968 ( \7221 , \7214 , \7219 , \7220 );
and \U$6969 ( \7222 , \7130 , \7221 );
and \U$6970 ( \7223 , \6065 , \5750 );
and \U$6971 ( \7224 , \6048 , \5748 );
nor \U$6972 ( \7225 , \7223 , \7224 );
xnor \U$6973 ( \7226 , \7225 , \5755 );
and \U$6974 ( \7227 , \5998 , \7157 );
and \U$6975 ( \7228 , \5967 , \7155 );
nor \U$6976 ( \7229 , \7227 , \7228 );
xnor \U$6977 ( \7230 , \7229 , \7163 );
and \U$6978 ( \7231 , \6018 , \7175 );
and \U$6979 ( \7232 , \5986 , \7173 );
nor \U$6980 ( \7233 , \7231 , \7232 );
xnor \U$6981 ( \7234 , \7233 , \7181 );
xor \U$6982 ( \7235 , \7230 , \7234 );
and \U$6983 ( \7236 , \6041 , \7192 );
and \U$6984 ( \7237 , \6006 , \7190 );
nor \U$6985 ( \7238 , \7236 , \7237 );
xnor \U$6986 ( \7239 , \7238 , \7198 );
xor \U$6987 ( \7240 , \7235 , \7239 );
and \U$6988 ( \7241 , \7226 , \7240 );
and \U$6989 ( \7242 , \5937 , \7099 );
and \U$6990 ( \7243 , \5906 , \7097 );
nor \U$6991 ( \7244 , \7242 , \7243 );
xnor \U$6992 ( \7245 , \7244 , \7105 );
and \U$6993 ( \7246 , \5957 , \7117 );
and \U$6994 ( \7247 , \5925 , \7115 );
nor \U$6995 ( \7248 , \7246 , \7247 );
xnor \U$6996 ( \7249 , \7248 , \7123 );
xor \U$6997 ( \7250 , \7245 , \7249 );
and \U$6998 ( \7251 , \5979 , \7140 );
and \U$6999 ( \7252 , \5945 , \7138 );
nor \U$7000 ( \7253 , \7251 , \7252 );
xnor \U$7001 ( \7254 , \7253 , \7146 );
xor \U$7002 ( \7255 , \7250 , \7254 );
and \U$7003 ( \7256 , \7240 , \7255 );
and \U$7004 ( \7257 , \7226 , \7255 );
or \U$7005 ( \7258 , \7241 , \7256 , \7257 );
and \U$7006 ( \7259 , \7221 , \7258 );
and \U$7007 ( \7260 , \7130 , \7258 );
or \U$7008 ( \7261 , \7222 , \7259 , \7260 );
and \U$7009 ( \7262 , \5780 , \6991 );
and \U$7010 ( \7263 , \5792 , \6988 );
nor \U$7011 ( \7264 , \7262 , \7263 );
xnor \U$7012 ( \7265 , \7264 , \6985 );
xor \U$7013 ( \7266 , \5775 , \7265 );
and \U$7014 ( \7267 , \5799 , \7006 );
and \U$7015 ( \7268 , \5811 , \7004 );
nor \U$7016 ( \7269 , \7267 , \7268 );
xnor \U$7017 ( \7270 , \7269 , \7012 );
xor \U$7018 ( \7271 , \7266 , \7270 );
and \U$7019 ( \7272 , \5945 , \7140 );
and \U$7020 ( \7273 , \5957 , \7138 );
nor \U$7021 ( \7274 , \7272 , \7273 );
xnor \U$7022 ( \7275 , \7274 , \7146 );
and \U$7023 ( \7276 , \5967 , \7157 );
and \U$7024 ( \7277 , \5979 , \7155 );
nor \U$7025 ( \7278 , \7276 , \7277 );
xnor \U$7026 ( \7279 , \7278 , \7163 );
xor \U$7027 ( \7280 , \7275 , \7279 );
and \U$7028 ( \7281 , \5986 , \7175 );
and \U$7029 ( \7282 , \5998 , \7173 );
nor \U$7030 ( \7283 , \7281 , \7282 );
xnor \U$7031 ( \7284 , \7283 , \7181 );
xor \U$7032 ( \7285 , \7280 , \7284 );
and \U$7033 ( \7286 , \5881 , \7082 );
and \U$7034 ( \7287 , \5893 , \7080 );
nor \U$7035 ( \7288 , \7286 , \7287 );
xnor \U$7036 ( \7289 , \7288 , \7088 );
and \U$7037 ( \7290 , \5906 , \7099 );
and \U$7038 ( \7291 , \5918 , \7097 );
nor \U$7039 ( \7292 , \7290 , \7291 );
xnor \U$7040 ( \7293 , \7292 , \7105 );
xor \U$7041 ( \7294 , \7289 , \7293 );
and \U$7042 ( \7295 , \5925 , \7117 );
and \U$7043 ( \7296 , \5937 , \7115 );
nor \U$7044 ( \7297 , \7295 , \7296 );
xnor \U$7045 ( \7298 , \7297 , \7123 );
xor \U$7046 ( \7299 , \7294 , \7298 );
xor \U$7047 ( \7300 , \7285 , \7299 );
and \U$7048 ( \7301 , \5819 , \7026 );
and \U$7049 ( \7302 , \5831 , \7024 );
nor \U$7050 ( \7303 , \7301 , \7302 );
xnor \U$7051 ( \7304 , \7303 , \7032 );
and \U$7052 ( \7305 , \5842 , \7043 );
and \U$7053 ( \7306 , \5854 , \7041 );
nor \U$7054 ( \7307 , \7305 , \7306 );
xnor \U$7055 ( \7308 , \7307 , \7049 );
xor \U$7056 ( \7309 , \7304 , \7308 );
and \U$7057 ( \7310 , \5861 , \7061 );
and \U$7058 ( \7311 , \5873 , \7059 );
nor \U$7059 ( \7312 , \7310 , \7311 );
xnor \U$7060 ( \7313 , \7312 , \7067 );
xor \U$7061 ( \7314 , \7309 , \7313 );
xor \U$7062 ( \7315 , \7300 , \7314 );
and \U$7063 ( \7316 , \7271 , \7315 );
and \U$7064 ( \7317 , \7230 , \7234 );
and \U$7065 ( \7318 , \7234 , \7239 );
and \U$7066 ( \7319 , \7230 , \7239 );
or \U$7067 ( \7320 , \7317 , \7318 , \7319 );
nand \U$7068 ( \7321 , \6065 , \5766 );
xnor \U$7069 ( \7322 , \7321 , \5775 );
xor \U$7070 ( \7323 , \7320 , \7322 );
and \U$7071 ( \7324 , \6006 , \7192 );
and \U$7072 ( \7325 , \6018 , \7190 );
nor \U$7073 ( \7326 , \7324 , \7325 );
xnor \U$7074 ( \7327 , \7326 , \7198 );
and \U$7075 ( \7328 , \6029 , \7203 );
and \U$7076 ( \7329 , \6041 , \7201 );
nor \U$7077 ( \7330 , \7328 , \7329 );
xnor \U$7078 ( \7331 , \7330 , \6824 );
xor \U$7079 ( \7332 , \7327 , \7331 );
and \U$7080 ( \7333 , \6048 , \5750 );
and \U$7081 ( \7334 , \6057 , \5748 );
nor \U$7082 ( \7335 , \7333 , \7334 );
xnor \U$7083 ( \7336 , \7335 , \5755 );
xor \U$7084 ( \7337 , \7332 , \7336 );
xor \U$7085 ( \7338 , \7323 , \7337 );
and \U$7086 ( \7339 , \7315 , \7338 );
and \U$7087 ( \7340 , \7271 , \7338 );
or \U$7088 ( \7341 , \7316 , \7339 , \7340 );
and \U$7089 ( \7342 , \7261 , \7341 );
and \U$7090 ( \7343 , \5775 , \7265 );
and \U$7091 ( \7344 , \7265 , \7270 );
and \U$7092 ( \7345 , \5775 , \7270 );
or \U$7093 ( \7346 , \7343 , \7344 , \7345 );
and \U$7094 ( \7347 , \7304 , \7308 );
and \U$7095 ( \7348 , \7308 , \7313 );
and \U$7096 ( \7349 , \7304 , \7313 );
or \U$7097 ( \7350 , \7347 , \7348 , \7349 );
xor \U$7098 ( \7351 , \7346 , \7350 );
and \U$7099 ( \7352 , \7289 , \7293 );
and \U$7100 ( \7353 , \7293 , \7298 );
and \U$7101 ( \7354 , \7289 , \7298 );
or \U$7102 ( \7355 , \7352 , \7353 , \7354 );
xor \U$7103 ( \7356 , \7351 , \7355 );
and \U$7104 ( \7357 , \7341 , \7356 );
and \U$7105 ( \7358 , \7261 , \7356 );
or \U$7106 ( \7359 , \7342 , \7357 , \7358 );
and \U$7107 ( \7360 , \5792 , \6991 );
and \U$7108 ( \7361 , \5758 , \6988 );
nor \U$7109 ( \7362 , \7360 , \7361 );
xnor \U$7110 ( \7363 , \7362 , \6985 );
and \U$7111 ( \7364 , \5811 , \7006 );
and \U$7112 ( \7365 , \5780 , \7004 );
nor \U$7113 ( \7366 , \7364 , \7365 );
xnor \U$7114 ( \7367 , \7366 , \7012 );
xor \U$7115 ( \7368 , \7363 , \7367 );
and \U$7116 ( \7369 , \5831 , \7026 );
and \U$7117 ( \7370 , \5799 , \7024 );
nor \U$7118 ( \7371 , \7369 , \7370 );
xnor \U$7119 ( \7372 , \7371 , \7032 );
xor \U$7120 ( \7373 , \7368 , \7372 );
and \U$7121 ( \7374 , \5979 , \7157 );
and \U$7122 ( \7375 , \5945 , \7155 );
nor \U$7123 ( \7376 , \7374 , \7375 );
xnor \U$7124 ( \7377 , \7376 , \7163 );
and \U$7125 ( \7378 , \5998 , \7175 );
and \U$7126 ( \7379 , \5967 , \7173 );
nor \U$7127 ( \7380 , \7378 , \7379 );
xnor \U$7128 ( \7381 , \7380 , \7181 );
xor \U$7129 ( \7382 , \7377 , \7381 );
and \U$7130 ( \7383 , \6018 , \7192 );
and \U$7131 ( \7384 , \5986 , \7190 );
nor \U$7132 ( \7385 , \7383 , \7384 );
xnor \U$7133 ( \7386 , \7385 , \7198 );
xor \U$7134 ( \7387 , \7382 , \7386 );
and \U$7135 ( \7388 , \5918 , \7099 );
and \U$7136 ( \7389 , \5881 , \7097 );
nor \U$7137 ( \7390 , \7388 , \7389 );
xnor \U$7138 ( \7391 , \7390 , \7105 );
and \U$7139 ( \7392 , \5937 , \7117 );
and \U$7140 ( \7393 , \5906 , \7115 );
nor \U$7141 ( \7394 , \7392 , \7393 );
xnor \U$7142 ( \7395 , \7394 , \7123 );
xor \U$7143 ( \7396 , \7391 , \7395 );
and \U$7144 ( \7397 , \5957 , \7140 );
and \U$7145 ( \7398 , \5925 , \7138 );
nor \U$7146 ( \7399 , \7397 , \7398 );
xnor \U$7147 ( \7400 , \7399 , \7146 );
xor \U$7148 ( \7401 , \7396 , \7400 );
xor \U$7149 ( \7402 , \7387 , \7401 );
and \U$7150 ( \7403 , \5854 , \7043 );
and \U$7151 ( \7404 , \5819 , \7041 );
nor \U$7152 ( \7405 , \7403 , \7404 );
xnor \U$7153 ( \7406 , \7405 , \7049 );
and \U$7154 ( \7407 , \5873 , \7061 );
and \U$7155 ( \7408 , \5842 , \7059 );
nor \U$7156 ( \7409 , \7407 , \7408 );
xnor \U$7157 ( \7410 , \7409 , \7067 );
xor \U$7158 ( \7411 , \7406 , \7410 );
and \U$7159 ( \7412 , \5893 , \7082 );
and \U$7160 ( \7413 , \5861 , \7080 );
nor \U$7161 ( \7414 , \7412 , \7413 );
xnor \U$7162 ( \7415 , \7414 , \7088 );
xor \U$7163 ( \7416 , \7411 , \7415 );
xor \U$7164 ( \7417 , \7402 , \7416 );
xor \U$7165 ( \7418 , \7373 , \7417 );
and \U$7166 ( \7419 , \7275 , \7279 );
and \U$7167 ( \7420 , \7279 , \7284 );
and \U$7168 ( \7421 , \7275 , \7284 );
or \U$7169 ( \7422 , \7419 , \7420 , \7421 );
and \U$7170 ( \7423 , \7327 , \7331 );
and \U$7171 ( \7424 , \7331 , \7336 );
and \U$7172 ( \7425 , \7327 , \7336 );
or \U$7173 ( \7426 , \7423 , \7424 , \7425 );
xor \U$7174 ( \7427 , \7422 , \7426 );
and \U$7175 ( \7428 , \6041 , \7203 );
and \U$7176 ( \7429 , \6006 , \7201 );
nor \U$7177 ( \7430 , \7428 , \7429 );
xnor \U$7178 ( \7431 , \7430 , \6824 );
and \U$7179 ( \7432 , \6057 , \5750 );
and \U$7180 ( \7433 , \6029 , \5748 );
nor \U$7181 ( \7434 , \7432 , \7433 );
xnor \U$7182 ( \7435 , \7434 , \5755 );
xor \U$7183 ( \7436 , \7431 , \7435 );
and \U$7184 ( \7437 , \6065 , \5768 );
and \U$7185 ( \7438 , \6048 , \5766 );
nor \U$7186 ( \7439 , \7437 , \7438 );
xnor \U$7187 ( \7440 , \7439 , \5775 );
xor \U$7188 ( \7441 , \7436 , \7440 );
xor \U$7189 ( \7442 , \7427 , \7441 );
xor \U$7190 ( \7443 , \7418 , \7442 );
and \U$7191 ( \7444 , \5811 , \6991 );
and \U$7192 ( \7445 , \5780 , \6988 );
nor \U$7193 ( \7446 , \7444 , \7445 );
xnor \U$7194 ( \7447 , \7446 , \6985 );
and \U$7195 ( \7448 , \5831 , \7006 );
and \U$7196 ( \7449 , \5799 , \7004 );
nor \U$7197 ( \7450 , \7448 , \7449 );
xnor \U$7198 ( \7451 , \7450 , \7012 );
and \U$7199 ( \7452 , \7447 , \7451 );
and \U$7200 ( \7453 , \5854 , \7026 );
and \U$7201 ( \7454 , \5819 , \7024 );
nor \U$7202 ( \7455 , \7453 , \7454 );
xnor \U$7203 ( \7456 , \7455 , \7032 );
and \U$7204 ( \7457 , \7451 , \7456 );
and \U$7205 ( \7458 , \7447 , \7456 );
or \U$7206 ( \7459 , \7452 , \7457 , \7458 );
and \U$7207 ( \7460 , \5873 , \7043 );
and \U$7208 ( \7461 , \5842 , \7041 );
nor \U$7209 ( \7462 , \7460 , \7461 );
xnor \U$7210 ( \7463 , \7462 , \7049 );
and \U$7211 ( \7464 , \5893 , \7061 );
and \U$7212 ( \7465 , \5861 , \7059 );
nor \U$7213 ( \7466 , \7464 , \7465 );
xnor \U$7214 ( \7467 , \7466 , \7067 );
and \U$7215 ( \7468 , \7463 , \7467 );
and \U$7216 ( \7469 , \5918 , \7082 );
and \U$7217 ( \7470 , \5881 , \7080 );
nor \U$7218 ( \7471 , \7469 , \7470 );
xnor \U$7219 ( \7472 , \7471 , \7088 );
and \U$7220 ( \7473 , \7467 , \7472 );
and \U$7221 ( \7474 , \7463 , \7472 );
or \U$7222 ( \7475 , \7468 , \7473 , \7474 );
and \U$7223 ( \7476 , \7459 , \7475 );
and \U$7224 ( \7477 , \7245 , \7249 );
and \U$7225 ( \7478 , \7249 , \7254 );
and \U$7226 ( \7479 , \7245 , \7254 );
or \U$7227 ( \7480 , \7477 , \7478 , \7479 );
and \U$7228 ( \7481 , \7475 , \7480 );
and \U$7229 ( \7482 , \7459 , \7480 );
or \U$7230 ( \7483 , \7476 , \7481 , \7482 );
and \U$7231 ( \7484 , \7320 , \7322 );
and \U$7232 ( \7485 , \7322 , \7337 );
and \U$7233 ( \7486 , \7320 , \7337 );
or \U$7234 ( \7487 , \7484 , \7485 , \7486 );
xor \U$7235 ( \7488 , \7483 , \7487 );
and \U$7236 ( \7489 , \7285 , \7299 );
and \U$7237 ( \7490 , \7299 , \7314 );
and \U$7238 ( \7491 , \7285 , \7314 );
or \U$7239 ( \7492 , \7489 , \7490 , \7491 );
xor \U$7240 ( \7493 , \7488 , \7492 );
and \U$7241 ( \7494 , \7443 , \7493 );
and \U$7242 ( \7495 , \7359 , \7494 );
and \U$7243 ( \7496 , \5861 , \7082 );
and \U$7244 ( \7497 , \5873 , \7080 );
nor \U$7245 ( \7498 , \7496 , \7497 );
xnor \U$7246 ( \7499 , \7498 , \7088 );
and \U$7247 ( \7500 , \5881 , \7099 );
and \U$7248 ( \7501 , \5893 , \7097 );
nor \U$7249 ( \7502 , \7500 , \7501 );
xnor \U$7250 ( \7503 , \7502 , \7105 );
xor \U$7251 ( \7504 , \7499 , \7503 );
and \U$7252 ( \7505 , \5906 , \7117 );
and \U$7253 ( \7506 , \5918 , \7115 );
nor \U$7254 ( \7507 , \7505 , \7506 );
xnor \U$7255 ( \7508 , \7507 , \7123 );
xor \U$7256 ( \7509 , \7504 , \7508 );
and \U$7257 ( \7510 , \5799 , \7026 );
and \U$7258 ( \7511 , \5811 , \7024 );
nor \U$7259 ( \7512 , \7510 , \7511 );
xnor \U$7260 ( \7513 , \7512 , \7032 );
and \U$7261 ( \7514 , \5819 , \7043 );
and \U$7262 ( \7515 , \5831 , \7041 );
nor \U$7263 ( \7516 , \7514 , \7515 );
xnor \U$7264 ( \7517 , \7516 , \7049 );
xor \U$7265 ( \7518 , \7513 , \7517 );
and \U$7266 ( \7519 , \5842 , \7061 );
and \U$7267 ( \7520 , \5854 , \7059 );
nor \U$7268 ( \7521 , \7519 , \7520 );
xnor \U$7269 ( \7522 , \7521 , \7067 );
xor \U$7270 ( \7523 , \7518 , \7522 );
xor \U$7271 ( \7524 , \7509 , \7523 );
and \U$7272 ( \7525 , \5758 , \6991 );
and \U$7273 ( \7526 , \5770 , \6988 );
nor \U$7274 ( \7527 , \7525 , \7526 );
xnor \U$7275 ( \7528 , \7527 , \6985 );
xor \U$7276 ( \7529 , \5797 , \7528 );
and \U$7277 ( \7530 , \5780 , \7006 );
and \U$7278 ( \7531 , \5792 , \7004 );
nor \U$7279 ( \7532 , \7530 , \7531 );
xnor \U$7280 ( \7533 , \7532 , \7012 );
xor \U$7281 ( \7534 , \7529 , \7533 );
xor \U$7282 ( \7535 , \7524 , \7534 );
nand \U$7283 ( \7536 , \6065 , \5788 );
xnor \U$7284 ( \7537 , \7536 , \5797 );
and \U$7285 ( \7538 , \5986 , \7192 );
and \U$7286 ( \7539 , \5998 , \7190 );
nor \U$7287 ( \7540 , \7538 , \7539 );
xnor \U$7288 ( \7541 , \7540 , \7198 );
and \U$7289 ( \7542 , \6006 , \7203 );
and \U$7290 ( \7543 , \6018 , \7201 );
nor \U$7291 ( \7544 , \7542 , \7543 );
xnor \U$7292 ( \7545 , \7544 , \6824 );
xor \U$7293 ( \7546 , \7541 , \7545 );
and \U$7294 ( \7547 , \6029 , \5750 );
and \U$7295 ( \7548 , \6041 , \5748 );
nor \U$7296 ( \7549 , \7547 , \7548 );
xnor \U$7297 ( \7550 , \7549 , \5755 );
xor \U$7298 ( \7551 , \7546 , \7550 );
xor \U$7299 ( \7552 , \7537 , \7551 );
and \U$7300 ( \7553 , \5925 , \7140 );
and \U$7301 ( \7554 , \5937 , \7138 );
nor \U$7302 ( \7555 , \7553 , \7554 );
xnor \U$7303 ( \7556 , \7555 , \7146 );
and \U$7304 ( \7557 , \5945 , \7157 );
and \U$7305 ( \7558 , \5957 , \7155 );
nor \U$7306 ( \7559 , \7557 , \7558 );
xnor \U$7307 ( \7560 , \7559 , \7163 );
xor \U$7308 ( \7561 , \7556 , \7560 );
and \U$7309 ( \7562 , \5967 , \7175 );
and \U$7310 ( \7563 , \5979 , \7173 );
nor \U$7311 ( \7564 , \7562 , \7563 );
xnor \U$7312 ( \7565 , \7564 , \7181 );
xor \U$7313 ( \7566 , \7561 , \7565 );
xor \U$7314 ( \7567 , \7552 , \7566 );
xor \U$7315 ( \7568 , \7535 , \7567 );
and \U$7316 ( \7569 , \7377 , \7381 );
and \U$7317 ( \7570 , \7381 , \7386 );
and \U$7318 ( \7571 , \7377 , \7386 );
or \U$7319 ( \7572 , \7569 , \7570 , \7571 );
and \U$7320 ( \7573 , \7431 , \7435 );
and \U$7321 ( \7574 , \7435 , \7440 );
and \U$7322 ( \7575 , \7431 , \7440 );
or \U$7323 ( \7576 , \7573 , \7574 , \7575 );
xor \U$7324 ( \7577 , \7572 , \7576 );
and \U$7325 ( \7578 , \6048 , \5768 );
and \U$7326 ( \7579 , \6057 , \5766 );
nor \U$7327 ( \7580 , \7578 , \7579 );
xnor \U$7328 ( \7581 , \7580 , \5775 );
xor \U$7329 ( \7582 , \7577 , \7581 );
xor \U$7330 ( \7583 , \7568 , \7582 );
and \U$7331 ( \7584 , \7494 , \7583 );
and \U$7332 ( \7585 , \7359 , \7583 );
or \U$7333 ( \7586 , \7495 , \7584 , \7585 );
and \U$7334 ( \7587 , \7346 , \7350 );
and \U$7335 ( \7588 , \7350 , \7355 );
and \U$7336 ( \7589 , \7346 , \7355 );
or \U$7337 ( \7590 , \7587 , \7588 , \7589 );
and \U$7338 ( \7591 , \7422 , \7426 );
and \U$7339 ( \7592 , \7426 , \7441 );
and \U$7340 ( \7593 , \7422 , \7441 );
or \U$7341 ( \7594 , \7591 , \7592 , \7593 );
xor \U$7342 ( \7595 , \7590 , \7594 );
and \U$7343 ( \7596 , \7387 , \7401 );
and \U$7344 ( \7597 , \7401 , \7416 );
and \U$7345 ( \7598 , \7387 , \7416 );
or \U$7346 ( \7599 , \7596 , \7597 , \7598 );
xor \U$7347 ( \7600 , \7595 , \7599 );
and \U$7348 ( \7601 , \7483 , \7487 );
and \U$7349 ( \7602 , \7487 , \7492 );
and \U$7350 ( \7603 , \7483 , \7492 );
or \U$7351 ( \7604 , \7601 , \7602 , \7603 );
and \U$7352 ( \7605 , \7373 , \7417 );
and \U$7353 ( \7606 , \7417 , \7442 );
and \U$7354 ( \7607 , \7373 , \7442 );
or \U$7355 ( \7608 , \7605 , \7606 , \7607 );
xor \U$7356 ( \7609 , \7604 , \7608 );
and \U$7357 ( \7610 , \7363 , \7367 );
and \U$7358 ( \7611 , \7367 , \7372 );
and \U$7359 ( \7612 , \7363 , \7372 );
or \U$7360 ( \7613 , \7610 , \7611 , \7612 );
and \U$7361 ( \7614 , \7406 , \7410 );
and \U$7362 ( \7615 , \7410 , \7415 );
and \U$7363 ( \7616 , \7406 , \7415 );
or \U$7364 ( \7617 , \7614 , \7615 , \7616 );
xor \U$7365 ( \7618 , \7613 , \7617 );
and \U$7366 ( \7619 , \7391 , \7395 );
and \U$7367 ( \7620 , \7395 , \7400 );
and \U$7368 ( \7621 , \7391 , \7400 );
or \U$7369 ( \7622 , \7619 , \7620 , \7621 );
xor \U$7370 ( \7623 , \7618 , \7622 );
xor \U$7371 ( \7624 , \7609 , \7623 );
and \U$7372 ( \7625 , \7600 , \7624 );
xor \U$7373 ( \7626 , \7586 , \7625 );
and \U$7374 ( \7627 , \7604 , \7608 );
and \U$7375 ( \7628 , \7608 , \7623 );
and \U$7376 ( \7629 , \7604 , \7623 );
or \U$7377 ( \7630 , \7627 , \7628 , \7629 );
and \U$7378 ( \7631 , \7509 , \7523 );
and \U$7379 ( \7632 , \7523 , \7534 );
and \U$7380 ( \7633 , \7509 , \7534 );
or \U$7381 ( \7634 , \7631 , \7632 , \7633 );
and \U$7382 ( \7635 , \5831 , \7043 );
and \U$7383 ( \7636 , \5799 , \7041 );
nor \U$7384 ( \7637 , \7635 , \7636 );
xnor \U$7385 ( \7638 , \7637 , \7049 );
and \U$7386 ( \7639 , \5854 , \7061 );
and \U$7387 ( \7640 , \5819 , \7059 );
nor \U$7388 ( \7641 , \7639 , \7640 );
xnor \U$7389 ( \7642 , \7641 , \7067 );
xor \U$7390 ( \7643 , \7638 , \7642 );
and \U$7391 ( \7644 , \5873 , \7082 );
and \U$7392 ( \7645 , \5842 , \7080 );
nor \U$7393 ( \7646 , \7644 , \7645 );
xnor \U$7394 ( \7647 , \7646 , \7088 );
xor \U$7395 ( \7648 , \7643 , \7647 );
xor \U$7396 ( \7649 , \7634 , \7648 );
and \U$7397 ( \7650 , \5770 , \6991 );
and \U$7398 ( \7651 , \5737 , \6988 );
nor \U$7399 ( \7652 , \7650 , \7651 );
xnor \U$7400 ( \7653 , \7652 , \6985 );
and \U$7401 ( \7654 , \5792 , \7006 );
and \U$7402 ( \7655 , \5758 , \7004 );
nor \U$7403 ( \7656 , \7654 , \7655 );
xnor \U$7404 ( \7657 , \7656 , \7012 );
xor \U$7405 ( \7658 , \7653 , \7657 );
and \U$7406 ( \7659 , \5811 , \7026 );
and \U$7407 ( \7660 , \5780 , \7024 );
nor \U$7408 ( \7661 , \7659 , \7660 );
xnor \U$7409 ( \7662 , \7661 , \7032 );
xor \U$7410 ( \7663 , \7658 , \7662 );
xor \U$7411 ( \7664 , \7649 , \7663 );
and \U$7412 ( \7665 , \7613 , \7617 );
and \U$7413 ( \7666 , \7617 , \7622 );
and \U$7414 ( \7667 , \7613 , \7622 );
or \U$7415 ( \7668 , \7665 , \7666 , \7667 );
and \U$7416 ( \7669 , \7572 , \7576 );
and \U$7417 ( \7670 , \7576 , \7581 );
and \U$7418 ( \7671 , \7572 , \7581 );
or \U$7419 ( \7672 , \7669 , \7670 , \7671 );
xor \U$7420 ( \7673 , \7668 , \7672 );
and \U$7421 ( \7674 , \7537 , \7551 );
and \U$7422 ( \7675 , \7551 , \7566 );
and \U$7423 ( \7676 , \7537 , \7566 );
or \U$7424 ( \7677 , \7674 , \7675 , \7676 );
xor \U$7425 ( \7678 , \7673 , \7677 );
xor \U$7426 ( \7679 , \7664 , \7678 );
xor \U$7427 ( \7680 , \7630 , \7679 );
and \U$7428 ( \7681 , \7590 , \7594 );
and \U$7429 ( \7682 , \7594 , \7599 );
and \U$7430 ( \7683 , \7590 , \7599 );
or \U$7431 ( \7684 , \7681 , \7682 , \7683 );
and \U$7432 ( \7685 , \7535 , \7567 );
and \U$7433 ( \7686 , \7567 , \7582 );
and \U$7434 ( \7687 , \7535 , \7582 );
or \U$7435 ( \7688 , \7685 , \7686 , \7687 );
xor \U$7436 ( \7689 , \7684 , \7688 );
and \U$7437 ( \7690 , \6018 , \7203 );
and \U$7438 ( \7691 , \5986 , \7201 );
nor \U$7439 ( \7692 , \7690 , \7691 );
xnor \U$7440 ( \7693 , \7692 , \6824 );
and \U$7441 ( \7694 , \6041 , \5750 );
and \U$7442 ( \7695 , \6006 , \5748 );
nor \U$7443 ( \7696 , \7694 , \7695 );
xnor \U$7444 ( \7697 , \7696 , \5755 );
xor \U$7445 ( \7698 , \7693 , \7697 );
and \U$7446 ( \7699 , \6057 , \5768 );
and \U$7447 ( \7700 , \6029 , \5766 );
nor \U$7448 ( \7701 , \7699 , \7700 );
xnor \U$7449 ( \7702 , \7701 , \5775 );
xor \U$7450 ( \7703 , \7698 , \7702 );
and \U$7451 ( \7704 , \5957 , \7157 );
and \U$7452 ( \7705 , \5925 , \7155 );
nor \U$7453 ( \7706 , \7704 , \7705 );
xnor \U$7454 ( \7707 , \7706 , \7163 );
and \U$7455 ( \7708 , \5979 , \7175 );
and \U$7456 ( \7709 , \5945 , \7173 );
nor \U$7457 ( \7710 , \7708 , \7709 );
xnor \U$7458 ( \7711 , \7710 , \7181 );
xor \U$7459 ( \7712 , \7707 , \7711 );
and \U$7460 ( \7713 , \5998 , \7192 );
and \U$7461 ( \7714 , \5967 , \7190 );
nor \U$7462 ( \7715 , \7713 , \7714 );
xnor \U$7463 ( \7716 , \7715 , \7198 );
xor \U$7464 ( \7717 , \7712 , \7716 );
xor \U$7465 ( \7718 , \7703 , \7717 );
and \U$7466 ( \7719 , \5893 , \7099 );
and \U$7467 ( \7720 , \5861 , \7097 );
nor \U$7468 ( \7721 , \7719 , \7720 );
xnor \U$7469 ( \7722 , \7721 , \7105 );
and \U$7470 ( \7723 , \5918 , \7117 );
and \U$7471 ( \7724 , \5881 , \7115 );
nor \U$7472 ( \7725 , \7723 , \7724 );
xnor \U$7473 ( \7726 , \7725 , \7123 );
xor \U$7474 ( \7727 , \7722 , \7726 );
and \U$7475 ( \7728 , \5937 , \7140 );
and \U$7476 ( \7729 , \5906 , \7138 );
nor \U$7477 ( \7730 , \7728 , \7729 );
xnor \U$7478 ( \7731 , \7730 , \7146 );
xor \U$7479 ( \7732 , \7727 , \7731 );
xor \U$7480 ( \7733 , \7718 , \7732 );
and \U$7481 ( \7734 , \7556 , \7560 );
and \U$7482 ( \7735 , \7560 , \7565 );
and \U$7483 ( \7736 , \7556 , \7565 );
or \U$7484 ( \7737 , \7734 , \7735 , \7736 );
and \U$7485 ( \7738 , \7541 , \7545 );
and \U$7486 ( \7739 , \7545 , \7550 );
and \U$7487 ( \7740 , \7541 , \7550 );
or \U$7488 ( \7741 , \7738 , \7739 , \7740 );
xor \U$7489 ( \7742 , \7737 , \7741 );
and \U$7490 ( \7743 , \6065 , \5790 );
and \U$7491 ( \7744 , \6048 , \5788 );
nor \U$7492 ( \7745 , \7743 , \7744 );
xnor \U$7493 ( \7746 , \7745 , \5797 );
xor \U$7494 ( \7747 , \7742 , \7746 );
xor \U$7495 ( \7748 , \7733 , \7747 );
and \U$7496 ( \7749 , \5797 , \7528 );
and \U$7497 ( \7750 , \7528 , \7533 );
and \U$7498 ( \7751 , \5797 , \7533 );
or \U$7499 ( \7752 , \7749 , \7750 , \7751 );
and \U$7500 ( \7753 , \7513 , \7517 );
and \U$7501 ( \7754 , \7517 , \7522 );
and \U$7502 ( \7755 , \7513 , \7522 );
or \U$7503 ( \7756 , \7753 , \7754 , \7755 );
xor \U$7504 ( \7757 , \7752 , \7756 );
and \U$7505 ( \7758 , \7499 , \7503 );
and \U$7506 ( \7759 , \7503 , \7508 );
and \U$7507 ( \7760 , \7499 , \7508 );
or \U$7508 ( \7761 , \7758 , \7759 , \7760 );
xor \U$7509 ( \7762 , \7757 , \7761 );
xor \U$7510 ( \7763 , \7748 , \7762 );
xor \U$7511 ( \7764 , \7689 , \7763 );
xor \U$7512 ( \7765 , \7680 , \7764 );
xor \U$7513 ( \7766 , \7626 , \7765 );
and \U$7514 ( \7767 , \5831 , \6991 );
and \U$7515 ( \7768 , \5799 , \6988 );
nor \U$7516 ( \7769 , \7767 , \7768 );
xnor \U$7517 ( \7770 , \7769 , \6985 );
and \U$7518 ( \7771 , \5854 , \7006 );
and \U$7519 ( \7772 , \5819 , \7004 );
nor \U$7520 ( \7773 , \7771 , \7772 );
xnor \U$7521 ( \7774 , \7773 , \7012 );
and \U$7522 ( \7775 , \7770 , \7774 );
and \U$7523 ( \7776 , \5873 , \7026 );
and \U$7524 ( \7777 , \5842 , \7024 );
nor \U$7525 ( \7778 , \7776 , \7777 );
xnor \U$7526 ( \7779 , \7778 , \7032 );
and \U$7527 ( \7780 , \7774 , \7779 );
and \U$7528 ( \7781 , \7770 , \7779 );
or \U$7529 ( \7782 , \7775 , \7780 , \7781 );
and \U$7530 ( \7783 , \5893 , \7043 );
and \U$7531 ( \7784 , \5861 , \7041 );
nor \U$7532 ( \7785 , \7783 , \7784 );
xnor \U$7533 ( \7786 , \7785 , \7049 );
and \U$7534 ( \7787 , \5918 , \7061 );
and \U$7535 ( \7788 , \5881 , \7059 );
nor \U$7536 ( \7789 , \7787 , \7788 );
xnor \U$7537 ( \7790 , \7789 , \7067 );
and \U$7538 ( \7791 , \7786 , \7790 );
and \U$7539 ( \7792 , \5937 , \7082 );
and \U$7540 ( \7793 , \5906 , \7080 );
nor \U$7541 ( \7794 , \7792 , \7793 );
xnor \U$7542 ( \7795 , \7794 , \7088 );
and \U$7543 ( \7796 , \7790 , \7795 );
and \U$7544 ( \7797 , \7786 , \7795 );
or \U$7545 ( \7798 , \7791 , \7796 , \7797 );
and \U$7546 ( \7799 , \7782 , \7798 );
and \U$7547 ( \7800 , \5957 , \7099 );
and \U$7548 ( \7801 , \5925 , \7097 );
nor \U$7549 ( \7802 , \7800 , \7801 );
xnor \U$7550 ( \7803 , \7802 , \7105 );
and \U$7551 ( \7804 , \5979 , \7117 );
and \U$7552 ( \7805 , \5945 , \7115 );
nor \U$7553 ( \7806 , \7804 , \7805 );
xnor \U$7554 ( \7807 , \7806 , \7123 );
and \U$7555 ( \7808 , \7803 , \7807 );
and \U$7556 ( \7809 , \5998 , \7140 );
and \U$7557 ( \7810 , \5967 , \7138 );
nor \U$7558 ( \7811 , \7809 , \7810 );
xnor \U$7559 ( \7812 , \7811 , \7146 );
and \U$7560 ( \7813 , \7807 , \7812 );
and \U$7561 ( \7814 , \7803 , \7812 );
or \U$7562 ( \7815 , \7808 , \7813 , \7814 );
and \U$7563 ( \7816 , \7798 , \7815 );
and \U$7564 ( \7817 , \7782 , \7815 );
or \U$7565 ( \7818 , \7799 , \7816 , \7817 );
and \U$7566 ( \7819 , \6018 , \7157 );
and \U$7567 ( \7820 , \5986 , \7155 );
nor \U$7568 ( \7821 , \7819 , \7820 );
xnor \U$7569 ( \7822 , \7821 , \7163 );
and \U$7570 ( \7823 , \6041 , \7175 );
and \U$7571 ( \7824 , \6006 , \7173 );
nor \U$7572 ( \7825 , \7823 , \7824 );
xnor \U$7573 ( \7826 , \7825 , \7181 );
and \U$7574 ( \7827 , \7822 , \7826 );
and \U$7575 ( \7828 , \6057 , \7192 );
and \U$7576 ( \7829 , \6029 , \7190 );
nor \U$7577 ( \7830 , \7828 , \7829 );
xnor \U$7578 ( \7831 , \7830 , \7198 );
and \U$7579 ( \7832 , \7826 , \7831 );
and \U$7580 ( \7833 , \7822 , \7831 );
or \U$7581 ( \7834 , \7827 , \7832 , \7833 );
xor \U$7582 ( \7835 , \7199 , \7207 );
xor \U$7583 ( \7836 , \7835 , \7210 );
and \U$7584 ( \7837 , \7834 , \7836 );
xor \U$7585 ( \7838 , \7147 , \7164 );
xor \U$7586 ( \7839 , \7838 , \7182 );
and \U$7587 ( \7840 , \7836 , \7839 );
and \U$7588 ( \7841 , \7834 , \7839 );
or \U$7589 ( \7842 , \7837 , \7840 , \7841 );
and \U$7590 ( \7843 , \7818 , \7842 );
xor \U$7591 ( \7844 , \7089 , \7106 );
xor \U$7592 ( \7845 , \7844 , \7124 );
xor \U$7593 ( \7846 , \7033 , \7050 );
xor \U$7594 ( \7847 , \7846 , \7068 );
and \U$7595 ( \7848 , \7845 , \7847 );
xor \U$7596 ( \7849 , \5755 , \6995 );
xor \U$7597 ( \7850 , \7849 , \7013 );
and \U$7598 ( \7851 , \7847 , \7850 );
and \U$7599 ( \7852 , \7845 , \7850 );
or \U$7600 ( \7853 , \7848 , \7851 , \7852 );
and \U$7601 ( \7854 , \7842 , \7853 );
and \U$7602 ( \7855 , \7818 , \7853 );
or \U$7603 ( \7856 , \7843 , \7854 , \7855 );
xor \U$7604 ( \7857 , \7463 , \7467 );
xor \U$7605 ( \7858 , \7857 , \7472 );
xor \U$7606 ( \7859 , \7447 , \7451 );
xor \U$7607 ( \7860 , \7859 , \7456 );
and \U$7608 ( \7861 , \7858 , \7860 );
xor \U$7609 ( \7862 , \7226 , \7240 );
xor \U$7610 ( \7863 , \7862 , \7255 );
and \U$7611 ( \7864 , \7860 , \7863 );
and \U$7612 ( \7865 , \7858 , \7863 );
or \U$7613 ( \7866 , \7861 , \7864 , \7865 );
and \U$7614 ( \7867 , \7856 , \7866 );
xor \U$7615 ( \7868 , \7459 , \7475 );
xor \U$7616 ( \7869 , \7868 , \7480 );
and \U$7617 ( \7870 , \7866 , \7869 );
and \U$7618 ( \7871 , \7856 , \7869 );
or \U$7619 ( \7872 , \7867 , \7870 , \7871 );
xor \U$7620 ( \7873 , \7443 , \7493 );
and \U$7621 ( \7874 , \7872 , \7873 );
xor \U$7622 ( \7875 , \7261 , \7341 );
xor \U$7623 ( \7876 , \7875 , \7356 );
and \U$7624 ( \7877 , \7873 , \7876 );
and \U$7625 ( \7878 , \7872 , \7876 );
or \U$7626 ( \7879 , \7874 , \7877 , \7878 );
xor \U$7627 ( \7880 , \7600 , \7624 );
and \U$7628 ( \7881 , \7879 , \7880 );
xor \U$7629 ( \7882 , \7359 , \7494 );
xor \U$7630 ( \7883 , \7882 , \7583 );
and \U$7631 ( \7884 , \7880 , \7883 );
and \U$7632 ( \7885 , \7879 , \7883 );
or \U$7633 ( \7886 , \7881 , \7884 , \7885 );
nor \U$7634 ( \7887 , \7766 , \7886 );
and \U$7635 ( \7888 , \7630 , \7679 );
and \U$7636 ( \7889 , \7679 , \7764 );
and \U$7637 ( \7890 , \7630 , \7764 );
or \U$7638 ( \7891 , \7888 , \7889 , \7890 );
and \U$7639 ( \7892 , \7668 , \7672 );
and \U$7640 ( \7893 , \7672 , \7677 );
and \U$7641 ( \7894 , \7668 , \7677 );
or \U$7642 ( \7895 , \7892 , \7893 , \7894 );
and \U$7643 ( \7896 , \7634 , \7648 );
and \U$7644 ( \7897 , \7648 , \7663 );
and \U$7645 ( \7898 , \7634 , \7663 );
or \U$7646 ( \7899 , \7896 , \7897 , \7898 );
xor \U$7647 ( \7900 , \7895 , \7899 );
and \U$7648 ( \7901 , \7733 , \7747 );
and \U$7649 ( \7902 , \7747 , \7762 );
and \U$7650 ( \7903 , \7733 , \7762 );
or \U$7651 ( \7904 , \7901 , \7902 , \7903 );
xor \U$7652 ( \7905 , \7900 , \7904 );
xor \U$7653 ( \7906 , \7891 , \7905 );
and \U$7654 ( \7907 , \7684 , \7688 );
and \U$7655 ( \7908 , \7688 , \7763 );
and \U$7656 ( \7909 , \7684 , \7763 );
or \U$7657 ( \7910 , \7907 , \7908 , \7909 );
and \U$7658 ( \7911 , \7664 , \7678 );
xor \U$7659 ( \7912 , \7910 , \7911 );
and \U$7660 ( \7913 , \7707 , \7711 );
and \U$7661 ( \7914 , \7711 , \7716 );
and \U$7662 ( \7915 , \7707 , \7716 );
or \U$7663 ( \7916 , \7913 , \7914 , \7915 );
and \U$7664 ( \7917 , \7693 , \7697 );
and \U$7665 ( \7918 , \7697 , \7702 );
and \U$7666 ( \7919 , \7693 , \7702 );
or \U$7667 ( \7920 , \7917 , \7918 , \7919 );
xor \U$7668 ( \7921 , \7916 , \7920 );
and \U$7669 ( \7922 , \6029 , \5768 );
and \U$7670 ( \7923 , \6041 , \5766 );
nor \U$7671 ( \7924 , \7922 , \7923 );
xnor \U$7672 ( \7925 , \7924 , \5775 );
and \U$7673 ( \7926 , \6048 , \5790 );
and \U$7674 ( \7927 , \6057 , \5788 );
nor \U$7675 ( \7928 , \7926 , \7927 );
xnor \U$7676 ( \7929 , \7928 , \5797 );
xor \U$7677 ( \7930 , \7925 , \7929 );
nand \U$7678 ( \7931 , \6065 , \5807 );
xnor \U$7679 ( \7932 , \7931 , \5816 );
xor \U$7680 ( \7933 , \7930 , \7932 );
xor \U$7681 ( \7934 , \7921 , \7933 );
and \U$7682 ( \7935 , \7653 , \7657 );
and \U$7683 ( \7936 , \7657 , \7662 );
and \U$7684 ( \7937 , \7653 , \7662 );
or \U$7685 ( \7938 , \7935 , \7936 , \7937 );
and \U$7686 ( \7939 , \7638 , \7642 );
and \U$7687 ( \7940 , \7642 , \7647 );
and \U$7688 ( \7941 , \7638 , \7647 );
or \U$7689 ( \7942 , \7939 , \7940 , \7941 );
xor \U$7690 ( \7943 , \7938 , \7942 );
and \U$7691 ( \7944 , \7722 , \7726 );
and \U$7692 ( \7945 , \7726 , \7731 );
and \U$7693 ( \7946 , \7722 , \7731 );
or \U$7694 ( \7947 , \7944 , \7945 , \7946 );
xor \U$7695 ( \7948 , \7943 , \7947 );
xor \U$7696 ( \7949 , \7934 , \7948 );
and \U$7697 ( \7950 , \5780 , \7026 );
and \U$7698 ( \7951 , \5792 , \7024 );
nor \U$7699 ( \7952 , \7950 , \7951 );
xnor \U$7700 ( \7953 , \7952 , \7032 );
and \U$7701 ( \7954 , \5799 , \7043 );
and \U$7702 ( \7955 , \5811 , \7041 );
nor \U$7703 ( \7956 , \7954 , \7955 );
xnor \U$7704 ( \7957 , \7956 , \7049 );
xor \U$7705 ( \7958 , \7953 , \7957 );
and \U$7706 ( \7959 , \5819 , \7061 );
and \U$7707 ( \7960 , \5831 , \7059 );
nor \U$7708 ( \7961 , \7959 , \7960 );
xnor \U$7709 ( \7962 , \7961 , \7067 );
xor \U$7710 ( \7963 , \7958 , \7962 );
and \U$7711 ( \7964 , \5737 , \6991 );
not \U$7712 ( \7965 , \7964 );
xnor \U$7713 ( \7966 , \7965 , \6985 );
xor \U$7714 ( \7967 , \5816 , \7966 );
and \U$7715 ( \7968 , \5758 , \7006 );
and \U$7716 ( \7969 , \5770 , \7004 );
nor \U$7717 ( \7970 , \7968 , \7969 );
xnor \U$7718 ( \7971 , \7970 , \7012 );
xor \U$7719 ( \7972 , \7967 , \7971 );
xor \U$7720 ( \7973 , \7963 , \7972 );
and \U$7721 ( \7974 , \5967 , \7192 );
and \U$7722 ( \7975 , \5979 , \7190 );
nor \U$7723 ( \7976 , \7974 , \7975 );
xnor \U$7724 ( \7977 , \7976 , \7198 );
and \U$7725 ( \7978 , \5986 , \7203 );
and \U$7726 ( \7979 , \5998 , \7201 );
nor \U$7727 ( \7980 , \7978 , \7979 );
xnor \U$7728 ( \7981 , \7980 , \6824 );
xor \U$7729 ( \7982 , \7977 , \7981 );
and \U$7730 ( \7983 , \6006 , \5750 );
and \U$7731 ( \7984 , \6018 , \5748 );
nor \U$7732 ( \7985 , \7983 , \7984 );
xnor \U$7733 ( \7986 , \7985 , \5755 );
xor \U$7734 ( \7987 , \7982 , \7986 );
and \U$7735 ( \7988 , \5906 , \7140 );
and \U$7736 ( \7989 , \5918 , \7138 );
nor \U$7737 ( \7990 , \7988 , \7989 );
xnor \U$7738 ( \7991 , \7990 , \7146 );
and \U$7739 ( \7992 , \5925 , \7157 );
and \U$7740 ( \7993 , \5937 , \7155 );
nor \U$7741 ( \7994 , \7992 , \7993 );
xnor \U$7742 ( \7995 , \7994 , \7163 );
xor \U$7743 ( \7996 , \7991 , \7995 );
and \U$7744 ( \7997 , \5945 , \7175 );
and \U$7745 ( \7998 , \5957 , \7173 );
nor \U$7746 ( \7999 , \7997 , \7998 );
xnor \U$7747 ( \8000 , \7999 , \7181 );
xor \U$7748 ( \8001 , \7996 , \8000 );
xor \U$7749 ( \8002 , \7987 , \8001 );
and \U$7750 ( \8003 , \5842 , \7082 );
and \U$7751 ( \8004 , \5854 , \7080 );
nor \U$7752 ( \8005 , \8003 , \8004 );
xnor \U$7753 ( \8006 , \8005 , \7088 );
and \U$7754 ( \8007 , \5861 , \7099 );
and \U$7755 ( \8008 , \5873 , \7097 );
nor \U$7756 ( \8009 , \8007 , \8008 );
xnor \U$7757 ( \8010 , \8009 , \7105 );
xor \U$7758 ( \8011 , \8006 , \8010 );
and \U$7759 ( \8012 , \5881 , \7117 );
and \U$7760 ( \8013 , \5893 , \7115 );
nor \U$7761 ( \8014 , \8012 , \8013 );
xnor \U$7762 ( \8015 , \8014 , \7123 );
xor \U$7763 ( \8016 , \8011 , \8015 );
xor \U$7764 ( \8017 , \8002 , \8016 );
xor \U$7765 ( \8018 , \7973 , \8017 );
xor \U$7766 ( \8019 , \7949 , \8018 );
and \U$7767 ( \8020 , \7752 , \7756 );
and \U$7768 ( \8021 , \7756 , \7761 );
and \U$7769 ( \8022 , \7752 , \7761 );
or \U$7770 ( \8023 , \8020 , \8021 , \8022 );
and \U$7771 ( \8024 , \7737 , \7741 );
and \U$7772 ( \8025 , \7741 , \7746 );
and \U$7773 ( \8026 , \7737 , \7746 );
or \U$7774 ( \8027 , \8024 , \8025 , \8026 );
xor \U$7775 ( \8028 , \8023 , \8027 );
and \U$7776 ( \8029 , \7703 , \7717 );
and \U$7777 ( \8030 , \7717 , \7732 );
and \U$7778 ( \8031 , \7703 , \7732 );
or \U$7779 ( \8032 , \8029 , \8030 , \8031 );
xor \U$7780 ( \8033 , \8028 , \8032 );
xor \U$7781 ( \8034 , \8019 , \8033 );
xor \U$7782 ( \8035 , \7912 , \8034 );
xor \U$7783 ( \8036 , \7906 , \8035 );
and \U$7784 ( \8037 , \7586 , \7625 );
and \U$7785 ( \8038 , \7625 , \7765 );
and \U$7786 ( \8039 , \7586 , \7765 );
or \U$7787 ( \8040 , \8037 , \8038 , \8039 );
nor \U$7788 ( \8041 , \8036 , \8040 );
nor \U$7789 ( \8042 , \7887 , \8041 );
and \U$7790 ( \8043 , \7910 , \7911 );
and \U$7791 ( \8044 , \7911 , \8034 );
and \U$7792 ( \8045 , \7910 , \8034 );
or \U$7793 ( \8046 , \8043 , \8044 , \8045 );
and \U$7794 ( \8047 , \8023 , \8027 );
and \U$7795 ( \8048 , \8027 , \8032 );
and \U$7796 ( \8049 , \8023 , \8032 );
or \U$7797 ( \8050 , \8047 , \8048 , \8049 );
and \U$7798 ( \8051 , \7963 , \7972 );
and \U$7799 ( \8052 , \7972 , \8017 );
and \U$7800 ( \8053 , \7963 , \8017 );
or \U$7801 ( \8054 , \8051 , \8052 , \8053 );
xor \U$7802 ( \8055 , \8050 , \8054 );
and \U$7803 ( \8056 , \7934 , \7948 );
xor \U$7804 ( \8057 , \8055 , \8056 );
xor \U$7805 ( \8058 , \8046 , \8057 );
and \U$7806 ( \8059 , \7895 , \7899 );
and \U$7807 ( \8060 , \7899 , \7904 );
and \U$7808 ( \8061 , \7895 , \7904 );
or \U$7809 ( \8062 , \8059 , \8060 , \8061 );
and \U$7810 ( \8063 , \7949 , \8018 );
and \U$7811 ( \8064 , \8018 , \8033 );
and \U$7812 ( \8065 , \7949 , \8033 );
or \U$7813 ( \8066 , \8063 , \8064 , \8065 );
xor \U$7814 ( \8067 , \8062 , \8066 );
and \U$7815 ( \8068 , \5816 , \7966 );
and \U$7816 ( \8069 , \7966 , \7971 );
and \U$7817 ( \8070 , \5816 , \7971 );
or \U$7818 ( \8071 , \8068 , \8069 , \8070 );
and \U$7819 ( \8072 , \7953 , \7957 );
and \U$7820 ( \8073 , \7957 , \7962 );
and \U$7821 ( \8074 , \7953 , \7962 );
or \U$7822 ( \8075 , \8072 , \8073 , \8074 );
xor \U$7823 ( \8076 , \8071 , \8075 );
and \U$7824 ( \8077 , \8006 , \8010 );
and \U$7825 ( \8078 , \8010 , \8015 );
and \U$7826 ( \8079 , \8006 , \8015 );
or \U$7827 ( \8080 , \8077 , \8078 , \8079 );
xor \U$7828 ( \8081 , \8076 , \8080 );
and \U$7829 ( \8082 , \5873 , \7099 );
and \U$7830 ( \8083 , \5842 , \7097 );
nor \U$7831 ( \8084 , \8082 , \8083 );
xnor \U$7832 ( \8085 , \8084 , \7105 );
and \U$7833 ( \8086 , \5893 , \7117 );
and \U$7834 ( \8087 , \5861 , \7115 );
nor \U$7835 ( \8088 , \8086 , \8087 );
xnor \U$7836 ( \8089 , \8088 , \7123 );
xor \U$7837 ( \8090 , \8085 , \8089 );
and \U$7838 ( \8091 , \5918 , \7140 );
and \U$7839 ( \8092 , \5881 , \7138 );
nor \U$7840 ( \8093 , \8091 , \8092 );
xnor \U$7841 ( \8094 , \8093 , \7146 );
xor \U$7842 ( \8095 , \8090 , \8094 );
and \U$7843 ( \8096 , \5811 , \7043 );
and \U$7844 ( \8097 , \5780 , \7041 );
nor \U$7845 ( \8098 , \8096 , \8097 );
xnor \U$7846 ( \8099 , \8098 , \7049 );
and \U$7847 ( \8100 , \5831 , \7061 );
and \U$7848 ( \8101 , \5799 , \7059 );
nor \U$7849 ( \8102 , \8100 , \8101 );
xnor \U$7850 ( \8103 , \8102 , \7067 );
xor \U$7851 ( \8104 , \8099 , \8103 );
and \U$7852 ( \8105 , \5854 , \7082 );
and \U$7853 ( \8106 , \5819 , \7080 );
nor \U$7854 ( \8107 , \8105 , \8106 );
xnor \U$7855 ( \8108 , \8107 , \7088 );
xor \U$7856 ( \8109 , \8104 , \8108 );
xor \U$7857 ( \8110 , \8095 , \8109 );
not \U$7858 ( \8111 , \6985 );
and \U$7859 ( \8112 , \5770 , \7006 );
and \U$7860 ( \8113 , \5737 , \7004 );
nor \U$7861 ( \8114 , \8112 , \8113 );
xnor \U$7862 ( \8115 , \8114 , \7012 );
xor \U$7863 ( \8116 , \8111 , \8115 );
and \U$7864 ( \8117 , \5792 , \7026 );
and \U$7865 ( \8118 , \5758 , \7024 );
nor \U$7866 ( \8119 , \8117 , \8118 );
xnor \U$7867 ( \8120 , \8119 , \7032 );
xor \U$7868 ( \8121 , \8116 , \8120 );
xor \U$7869 ( \8122 , \8110 , \8121 );
and \U$7870 ( \8123 , \6057 , \5790 );
and \U$7871 ( \8124 , \6029 , \5788 );
nor \U$7872 ( \8125 , \8123 , \8124 );
xnor \U$7873 ( \8126 , \8125 , \5797 );
and \U$7874 ( \8127 , \6065 , \5809 );
and \U$7875 ( \8128 , \6048 , \5807 );
nor \U$7876 ( \8129 , \8127 , \8128 );
xnor \U$7877 ( \8130 , \8129 , \5816 );
xnor \U$7878 ( \8131 , \8126 , \8130 );
and \U$7879 ( \8132 , \5998 , \7203 );
and \U$7880 ( \8133 , \5967 , \7201 );
nor \U$7881 ( \8134 , \8132 , \8133 );
xnor \U$7882 ( \8135 , \8134 , \6824 );
and \U$7883 ( \8136 , \6018 , \5750 );
and \U$7884 ( \8137 , \5986 , \5748 );
nor \U$7885 ( \8138 , \8136 , \8137 );
xnor \U$7886 ( \8139 , \8138 , \5755 );
xor \U$7887 ( \8140 , \8135 , \8139 );
and \U$7888 ( \8141 , \6041 , \5768 );
and \U$7889 ( \8142 , \6006 , \5766 );
nor \U$7890 ( \8143 , \8141 , \8142 );
xnor \U$7891 ( \8144 , \8143 , \5775 );
xor \U$7892 ( \8145 , \8140 , \8144 );
xor \U$7893 ( \8146 , \8131 , \8145 );
and \U$7894 ( \8147 , \5937 , \7157 );
and \U$7895 ( \8148 , \5906 , \7155 );
nor \U$7896 ( \8149 , \8147 , \8148 );
xnor \U$7897 ( \8150 , \8149 , \7163 );
and \U$7898 ( \8151 , \5957 , \7175 );
and \U$7899 ( \8152 , \5925 , \7173 );
nor \U$7900 ( \8153 , \8151 , \8152 );
xnor \U$7901 ( \8154 , \8153 , \7181 );
xor \U$7902 ( \8155 , \8150 , \8154 );
and \U$7903 ( \8156 , \5979 , \7192 );
and \U$7904 ( \8157 , \5945 , \7190 );
nor \U$7905 ( \8158 , \8156 , \8157 );
xnor \U$7906 ( \8159 , \8158 , \7198 );
xor \U$7907 ( \8160 , \8155 , \8159 );
xor \U$7908 ( \8161 , \8146 , \8160 );
xor \U$7909 ( \8162 , \8122 , \8161 );
and \U$7910 ( \8163 , \7991 , \7995 );
and \U$7911 ( \8164 , \7995 , \8000 );
and \U$7912 ( \8165 , \7991 , \8000 );
or \U$7913 ( \8166 , \8163 , \8164 , \8165 );
and \U$7914 ( \8167 , \7977 , \7981 );
and \U$7915 ( \8168 , \7981 , \7986 );
and \U$7916 ( \8169 , \7977 , \7986 );
or \U$7917 ( \8170 , \8167 , \8168 , \8169 );
xor \U$7918 ( \8171 , \8166 , \8170 );
and \U$7919 ( \8172 , \7925 , \7929 );
and \U$7920 ( \8173 , \7929 , \7932 );
and \U$7921 ( \8174 , \7925 , \7932 );
or \U$7922 ( \8175 , \8172 , \8173 , \8174 );
xor \U$7923 ( \8176 , \8171 , \8175 );
xor \U$7924 ( \8177 , \8162 , \8176 );
xor \U$7925 ( \8178 , \8081 , \8177 );
and \U$7926 ( \8179 , \7938 , \7942 );
and \U$7927 ( \8180 , \7942 , \7947 );
and \U$7928 ( \8181 , \7938 , \7947 );
or \U$7929 ( \8182 , \8179 , \8180 , \8181 );
and \U$7930 ( \8183 , \7916 , \7920 );
and \U$7931 ( \8184 , \7920 , \7933 );
and \U$7932 ( \8185 , \7916 , \7933 );
or \U$7933 ( \8186 , \8183 , \8184 , \8185 );
xor \U$7934 ( \8187 , \8182 , \8186 );
and \U$7935 ( \8188 , \7987 , \8001 );
and \U$7936 ( \8189 , \8001 , \8016 );
and \U$7937 ( \8190 , \7987 , \8016 );
or \U$7938 ( \8191 , \8188 , \8189 , \8190 );
xor \U$7939 ( \8192 , \8187 , \8191 );
xor \U$7940 ( \8193 , \8178 , \8192 );
xor \U$7941 ( \8194 , \8067 , \8193 );
xor \U$7942 ( \8195 , \8058 , \8194 );
and \U$7943 ( \8196 , \7891 , \7905 );
and \U$7944 ( \8197 , \7905 , \8035 );
and \U$7945 ( \8198 , \7891 , \8035 );
or \U$7946 ( \8199 , \8196 , \8197 , \8198 );
nor \U$7947 ( \8200 , \8195 , \8199 );
and \U$7948 ( \8201 , \8062 , \8066 );
and \U$7949 ( \8202 , \8066 , \8193 );
and \U$7950 ( \8203 , \8062 , \8193 );
or \U$7951 ( \8204 , \8201 , \8202 , \8203 );
and \U$7952 ( \8205 , \8071 , \8075 );
and \U$7953 ( \8206 , \8075 , \8080 );
and \U$7954 ( \8207 , \8071 , \8080 );
or \U$7955 ( \8208 , \8205 , \8206 , \8207 );
and \U$7956 ( \8209 , \8166 , \8170 );
and \U$7957 ( \8210 , \8170 , \8175 );
and \U$7958 ( \8211 , \8166 , \8175 );
or \U$7959 ( \8212 , \8209 , \8210 , \8211 );
xor \U$7960 ( \8213 , \8208 , \8212 );
and \U$7961 ( \8214 , \8131 , \8145 );
and \U$7962 ( \8215 , \8145 , \8160 );
and \U$7963 ( \8216 , \8131 , \8160 );
or \U$7964 ( \8217 , \8214 , \8215 , \8216 );
xor \U$7965 ( \8218 , \8213 , \8217 );
and \U$7966 ( \8219 , \8182 , \8186 );
and \U$7967 ( \8220 , \8186 , \8191 );
and \U$7968 ( \8221 , \8182 , \8191 );
or \U$7969 ( \8222 , \8219 , \8220 , \8221 );
and \U$7970 ( \8223 , \8122 , \8161 );
and \U$7971 ( \8224 , \8161 , \8176 );
and \U$7972 ( \8225 , \8122 , \8176 );
or \U$7973 ( \8226 , \8223 , \8224 , \8225 );
xor \U$7974 ( \8227 , \8222 , \8226 );
and \U$7975 ( \8228 , \6029 , \5790 );
and \U$7976 ( \8229 , \6041 , \5788 );
nor \U$7977 ( \8230 , \8228 , \8229 );
xnor \U$7978 ( \8231 , \8230 , \5797 );
and \U$7979 ( \8232 , \6048 , \5809 );
and \U$7980 ( \8233 , \6057 , \5807 );
nor \U$7981 ( \8234 , \8232 , \8233 );
xnor \U$7982 ( \8235 , \8234 , \5816 );
xor \U$7983 ( \8236 , \8231 , \8235 );
nand \U$7984 ( \8237 , \6065 , \5827 );
xnor \U$7985 ( \8238 , \8237 , \5836 );
xor \U$7986 ( \8239 , \8236 , \8238 );
and \U$7987 ( \8240 , \5967 , \7203 );
and \U$7988 ( \8241 , \5979 , \7201 );
nor \U$7989 ( \8242 , \8240 , \8241 );
xnor \U$7990 ( \8243 , \8242 , \6824 );
and \U$7991 ( \8244 , \5986 , \5750 );
and \U$7992 ( \8245 , \5998 , \5748 );
nor \U$7993 ( \8246 , \8244 , \8245 );
xnor \U$7994 ( \8247 , \8246 , \5755 );
xor \U$7995 ( \8248 , \8243 , \8247 );
and \U$7996 ( \8249 , \6006 , \5768 );
and \U$7997 ( \8250 , \6018 , \5766 );
nor \U$7998 ( \8251 , \8249 , \8250 );
xnor \U$7999 ( \8252 , \8251 , \5775 );
xor \U$8000 ( \8253 , \8248 , \8252 );
xnor \U$8001 ( \8254 , \8239 , \8253 );
and \U$8002 ( \8255 , \8150 , \8154 );
and \U$8003 ( \8256 , \8154 , \8159 );
and \U$8004 ( \8257 , \8150 , \8159 );
or \U$8005 ( \8258 , \8255 , \8256 , \8257 );
and \U$8006 ( \8259 , \8135 , \8139 );
and \U$8007 ( \8260 , \8139 , \8144 );
and \U$8008 ( \8261 , \8135 , \8144 );
or \U$8009 ( \8262 , \8259 , \8260 , \8261 );
xor \U$8010 ( \8263 , \8258 , \8262 );
or \U$8011 ( \8264 , \8126 , \8130 );
xor \U$8012 ( \8265 , \8263 , \8264 );
xor \U$8013 ( \8266 , \8254 , \8265 );
and \U$8014 ( \8267 , \8111 , \8115 );
and \U$8015 ( \8268 , \8115 , \8120 );
and \U$8016 ( \8269 , \8111 , \8120 );
or \U$8017 ( \8270 , \8267 , \8268 , \8269 );
and \U$8018 ( \8271 , \8099 , \8103 );
and \U$8019 ( \8272 , \8103 , \8108 );
and \U$8020 ( \8273 , \8099 , \8108 );
or \U$8021 ( \8274 , \8271 , \8272 , \8273 );
xor \U$8022 ( \8275 , \8270 , \8274 );
and \U$8023 ( \8276 , \8085 , \8089 );
and \U$8024 ( \8277 , \8089 , \8094 );
and \U$8025 ( \8278 , \8085 , \8094 );
or \U$8026 ( \8279 , \8276 , \8277 , \8278 );
xor \U$8027 ( \8280 , \8275 , \8279 );
xor \U$8028 ( \8281 , \8266 , \8280 );
xor \U$8029 ( \8282 , \8227 , \8281 );
xor \U$8030 ( \8283 , \8218 , \8282 );
xor \U$8031 ( \8284 , \8204 , \8283 );
and \U$8032 ( \8285 , \8050 , \8054 );
and \U$8033 ( \8286 , \8054 , \8056 );
and \U$8034 ( \8287 , \8050 , \8056 );
or \U$8035 ( \8288 , \8285 , \8286 , \8287 );
and \U$8036 ( \8289 , \8081 , \8177 );
and \U$8037 ( \8290 , \8177 , \8192 );
and \U$8038 ( \8291 , \8081 , \8192 );
or \U$8039 ( \8292 , \8289 , \8290 , \8291 );
xor \U$8040 ( \8293 , \8288 , \8292 );
and \U$8041 ( \8294 , \8095 , \8109 );
and \U$8042 ( \8295 , \8109 , \8121 );
and \U$8043 ( \8296 , \8095 , \8121 );
or \U$8044 ( \8297 , \8294 , \8295 , \8296 );
and \U$8045 ( \8298 , \5737 , \7006 );
not \U$8046 ( \8299 , \8298 );
xnor \U$8047 ( \8300 , \8299 , \7012 );
xor \U$8048 ( \8301 , \5836 , \8300 );
and \U$8049 ( \8302 , \5758 , \7026 );
and \U$8050 ( \8303 , \5770 , \7024 );
nor \U$8051 ( \8304 , \8302 , \8303 );
xnor \U$8052 ( \8305 , \8304 , \7032 );
xor \U$8053 ( \8306 , \8301 , \8305 );
xor \U$8054 ( \8307 , \8297 , \8306 );
and \U$8055 ( \8308 , \5906 , \7157 );
and \U$8056 ( \8309 , \5918 , \7155 );
nor \U$8057 ( \8310 , \8308 , \8309 );
xnor \U$8058 ( \8311 , \8310 , \7163 );
and \U$8059 ( \8312 , \5925 , \7175 );
and \U$8060 ( \8313 , \5937 , \7173 );
nor \U$8061 ( \8314 , \8312 , \8313 );
xnor \U$8062 ( \8315 , \8314 , \7181 );
xor \U$8063 ( \8316 , \8311 , \8315 );
and \U$8064 ( \8317 , \5945 , \7192 );
and \U$8065 ( \8318 , \5957 , \7190 );
nor \U$8066 ( \8319 , \8317 , \8318 );
xnor \U$8067 ( \8320 , \8319 , \7198 );
xor \U$8068 ( \8321 , \8316 , \8320 );
and \U$8069 ( \8322 , \5842 , \7099 );
and \U$8070 ( \8323 , \5854 , \7097 );
nor \U$8071 ( \8324 , \8322 , \8323 );
xnor \U$8072 ( \8325 , \8324 , \7105 );
and \U$8073 ( \8326 , \5861 , \7117 );
and \U$8074 ( \8327 , \5873 , \7115 );
nor \U$8075 ( \8328 , \8326 , \8327 );
xnor \U$8076 ( \8329 , \8328 , \7123 );
xor \U$8077 ( \8330 , \8325 , \8329 );
and \U$8078 ( \8331 , \5881 , \7140 );
and \U$8079 ( \8332 , \5893 , \7138 );
nor \U$8080 ( \8333 , \8331 , \8332 );
xnor \U$8081 ( \8334 , \8333 , \7146 );
xor \U$8082 ( \8335 , \8330 , \8334 );
xor \U$8083 ( \8336 , \8321 , \8335 );
and \U$8084 ( \8337 , \5780 , \7043 );
and \U$8085 ( \8338 , \5792 , \7041 );
nor \U$8086 ( \8339 , \8337 , \8338 );
xnor \U$8087 ( \8340 , \8339 , \7049 );
and \U$8088 ( \8341 , \5799 , \7061 );
and \U$8089 ( \8342 , \5811 , \7059 );
nor \U$8090 ( \8343 , \8341 , \8342 );
xnor \U$8091 ( \8344 , \8343 , \7067 );
xor \U$8092 ( \8345 , \8340 , \8344 );
and \U$8093 ( \8346 , \5819 , \7082 );
and \U$8094 ( \8347 , \5831 , \7080 );
nor \U$8095 ( \8348 , \8346 , \8347 );
xnor \U$8096 ( \8349 , \8348 , \7088 );
xor \U$8097 ( \8350 , \8345 , \8349 );
xor \U$8098 ( \8351 , \8336 , \8350 );
xor \U$8099 ( \8352 , \8307 , \8351 );
xor \U$8100 ( \8353 , \8293 , \8352 );
xor \U$8101 ( \8354 , \8284 , \8353 );
and \U$8102 ( \8355 , \8046 , \8057 );
and \U$8103 ( \8356 , \8057 , \8194 );
and \U$8104 ( \8357 , \8046 , \8194 );
or \U$8105 ( \8358 , \8355 , \8356 , \8357 );
nor \U$8106 ( \8359 , \8354 , \8358 );
nor \U$8107 ( \8360 , \8200 , \8359 );
nand \U$8108 ( \8361 , \8042 , \8360 );
and \U$8109 ( \8362 , \8288 , \8292 );
and \U$8110 ( \8363 , \8292 , \8352 );
and \U$8111 ( \8364 , \8288 , \8352 );
or \U$8112 ( \8365 , \8362 , \8363 , \8364 );
and \U$8113 ( \8366 , \8218 , \8282 );
xor \U$8114 ( \8367 , \8365 , \8366 );
and \U$8115 ( \8368 , \8222 , \8226 );
and \U$8116 ( \8369 , \8226 , \8281 );
and \U$8117 ( \8370 , \8222 , \8281 );
or \U$8118 ( \8371 , \8368 , \8369 , \8370 );
and \U$8119 ( \8372 , \8311 , \8315 );
and \U$8120 ( \8373 , \8315 , \8320 );
and \U$8121 ( \8374 , \8311 , \8320 );
or \U$8122 ( \8375 , \8372 , \8373 , \8374 );
and \U$8123 ( \8376 , \8243 , \8247 );
and \U$8124 ( \8377 , \8247 , \8252 );
and \U$8125 ( \8378 , \8243 , \8252 );
or \U$8126 ( \8379 , \8376 , \8377 , \8378 );
xor \U$8127 ( \8380 , \8375 , \8379 );
and \U$8128 ( \8381 , \8231 , \8235 );
and \U$8129 ( \8382 , \8235 , \8238 );
and \U$8130 ( \8383 , \8231 , \8238 );
or \U$8131 ( \8384 , \8381 , \8382 , \8383 );
xor \U$8132 ( \8385 , \8380 , \8384 );
and \U$8133 ( \8386 , \5836 , \8300 );
and \U$8134 ( \8387 , \8300 , \8305 );
and \U$8135 ( \8388 , \5836 , \8305 );
or \U$8136 ( \8389 , \8386 , \8387 , \8388 );
and \U$8137 ( \8390 , \8340 , \8344 );
and \U$8138 ( \8391 , \8344 , \8349 );
and \U$8139 ( \8392 , \8340 , \8349 );
or \U$8140 ( \8393 , \8390 , \8391 , \8392 );
xor \U$8141 ( \8394 , \8389 , \8393 );
and \U$8142 ( \8395 , \8325 , \8329 );
and \U$8143 ( \8396 , \8329 , \8334 );
and \U$8144 ( \8397 , \8325 , \8334 );
or \U$8145 ( \8398 , \8395 , \8396 , \8397 );
xor \U$8146 ( \8399 , \8394 , \8398 );
xor \U$8147 ( \8400 , \8385 , \8399 );
and \U$8148 ( \8401 , \8321 , \8335 );
and \U$8149 ( \8402 , \8335 , \8350 );
and \U$8150 ( \8403 , \8321 , \8350 );
or \U$8151 ( \8404 , \8401 , \8402 , \8403 );
and \U$8152 ( \8405 , \5873 , \7117 );
and \U$8153 ( \8406 , \5842 , \7115 );
nor \U$8154 ( \8407 , \8405 , \8406 );
xnor \U$8155 ( \8408 , \8407 , \7123 );
and \U$8156 ( \8409 , \5893 , \7140 );
and \U$8157 ( \8410 , \5861 , \7138 );
nor \U$8158 ( \8411 , \8409 , \8410 );
xnor \U$8159 ( \8412 , \8411 , \7146 );
xor \U$8160 ( \8413 , \8408 , \8412 );
and \U$8161 ( \8414 , \5918 , \7157 );
and \U$8162 ( \8415 , \5881 , \7155 );
nor \U$8163 ( \8416 , \8414 , \8415 );
xnor \U$8164 ( \8417 , \8416 , \7163 );
xor \U$8165 ( \8418 , \8413 , \8417 );
and \U$8166 ( \8419 , \5811 , \7061 );
and \U$8167 ( \8420 , \5780 , \7059 );
nor \U$8168 ( \8421 , \8419 , \8420 );
xnor \U$8169 ( \8422 , \8421 , \7067 );
and \U$8170 ( \8423 , \5831 , \7082 );
and \U$8171 ( \8424 , \5799 , \7080 );
nor \U$8172 ( \8425 , \8423 , \8424 );
xnor \U$8173 ( \8426 , \8425 , \7088 );
xor \U$8174 ( \8427 , \8422 , \8426 );
and \U$8175 ( \8428 , \5854 , \7099 );
and \U$8176 ( \8429 , \5819 , \7097 );
nor \U$8177 ( \8430 , \8428 , \8429 );
xnor \U$8178 ( \8431 , \8430 , \7105 );
xor \U$8179 ( \8432 , \8427 , \8431 );
xor \U$8180 ( \8433 , \8418 , \8432 );
not \U$8181 ( \8434 , \7012 );
and \U$8182 ( \8435 , \5770 , \7026 );
and \U$8183 ( \8436 , \5737 , \7024 );
nor \U$8184 ( \8437 , \8435 , \8436 );
xnor \U$8185 ( \8438 , \8437 , \7032 );
xor \U$8186 ( \8439 , \8434 , \8438 );
and \U$8187 ( \8440 , \5792 , \7043 );
and \U$8188 ( \8441 , \5758 , \7041 );
nor \U$8189 ( \8442 , \8440 , \8441 );
xnor \U$8190 ( \8443 , \8442 , \7049 );
xor \U$8191 ( \8444 , \8439 , \8443 );
xor \U$8192 ( \8445 , \8433 , \8444 );
xor \U$8193 ( \8446 , \8404 , \8445 );
and \U$8194 ( \8447 , \6057 , \5809 );
and \U$8195 ( \8448 , \6029 , \5807 );
nor \U$8196 ( \8449 , \8447 , \8448 );
xnor \U$8197 ( \8450 , \8449 , \5816 );
and \U$8198 ( \8451 , \6065 , \5829 );
and \U$8199 ( \8452 , \6048 , \5827 );
nor \U$8200 ( \8453 , \8451 , \8452 );
xnor \U$8201 ( \8454 , \8453 , \5836 );
xor \U$8202 ( \8455 , \8450 , \8454 );
and \U$8203 ( \8456 , \5998 , \5750 );
and \U$8204 ( \8457 , \5967 , \5748 );
nor \U$8205 ( \8458 , \8456 , \8457 );
xnor \U$8206 ( \8459 , \8458 , \5755 );
and \U$8207 ( \8460 , \6018 , \5768 );
and \U$8208 ( \8461 , \5986 , \5766 );
nor \U$8209 ( \8462 , \8460 , \8461 );
xnor \U$8210 ( \8463 , \8462 , \5775 );
xor \U$8211 ( \8464 , \8459 , \8463 );
and \U$8212 ( \8465 , \6041 , \5790 );
and \U$8213 ( \8466 , \6006 , \5788 );
nor \U$8214 ( \8467 , \8465 , \8466 );
xnor \U$8215 ( \8468 , \8467 , \5797 );
xor \U$8216 ( \8469 , \8464 , \8468 );
xor \U$8217 ( \8470 , \8455 , \8469 );
and \U$8218 ( \8471 , \5937 , \7175 );
and \U$8219 ( \8472 , \5906 , \7173 );
nor \U$8220 ( \8473 , \8471 , \8472 );
xnor \U$8221 ( \8474 , \8473 , \7181 );
and \U$8222 ( \8475 , \5957 , \7192 );
and \U$8223 ( \8476 , \5925 , \7190 );
nor \U$8224 ( \8477 , \8475 , \8476 );
xnor \U$8225 ( \8478 , \8477 , \7198 );
xor \U$8226 ( \8479 , \8474 , \8478 );
and \U$8227 ( \8480 , \5979 , \7203 );
and \U$8228 ( \8481 , \5945 , \7201 );
nor \U$8229 ( \8482 , \8480 , \8481 );
xnor \U$8230 ( \8483 , \8482 , \6824 );
xor \U$8231 ( \8484 , \8479 , \8483 );
xor \U$8232 ( \8485 , \8470 , \8484 );
xor \U$8233 ( \8486 , \8446 , \8485 );
xor \U$8234 ( \8487 , \8400 , \8486 );
and \U$8235 ( \8488 , \8270 , \8274 );
and \U$8236 ( \8489 , \8274 , \8279 );
and \U$8237 ( \8490 , \8270 , \8279 );
or \U$8238 ( \8491 , \8488 , \8489 , \8490 );
and \U$8239 ( \8492 , \8258 , \8262 );
and \U$8240 ( \8493 , \8262 , \8264 );
and \U$8241 ( \8494 , \8258 , \8264 );
or \U$8242 ( \8495 , \8492 , \8493 , \8494 );
xor \U$8243 ( \8496 , \8491 , \8495 );
or \U$8244 ( \8497 , \8239 , \8253 );
xor \U$8245 ( \8498 , \8496 , \8497 );
xor \U$8246 ( \8499 , \8487 , \8498 );
xor \U$8247 ( \8500 , \8371 , \8499 );
and \U$8248 ( \8501 , \8208 , \8212 );
and \U$8249 ( \8502 , \8212 , \8217 );
and \U$8250 ( \8503 , \8208 , \8217 );
or \U$8251 ( \8504 , \8501 , \8502 , \8503 );
and \U$8252 ( \8505 , \8297 , \8306 );
and \U$8253 ( \8506 , \8306 , \8351 );
and \U$8254 ( \8507 , \8297 , \8351 );
or \U$8255 ( \8508 , \8505 , \8506 , \8507 );
xor \U$8256 ( \8509 , \8504 , \8508 );
and \U$8257 ( \8510 , \8254 , \8265 );
and \U$8258 ( \8511 , \8265 , \8280 );
and \U$8259 ( \8512 , \8254 , \8280 );
or \U$8260 ( \8513 , \8510 , \8511 , \8512 );
xor \U$8261 ( \8514 , \8509 , \8513 );
xor \U$8262 ( \8515 , \8500 , \8514 );
xor \U$8263 ( \8516 , \8367 , \8515 );
and \U$8264 ( \8517 , \8204 , \8283 );
and \U$8265 ( \8518 , \8283 , \8353 );
and \U$8266 ( \8519 , \8204 , \8353 );
or \U$8267 ( \8520 , \8517 , \8518 , \8519 );
nor \U$8268 ( \8521 , \8516 , \8520 );
and \U$8269 ( \8522 , \8371 , \8499 );
and \U$8270 ( \8523 , \8499 , \8514 );
and \U$8271 ( \8524 , \8371 , \8514 );
or \U$8272 ( \8525 , \8522 , \8523 , \8524 );
and \U$8273 ( \8526 , \8491 , \8495 );
and \U$8274 ( \8527 , \8495 , \8497 );
and \U$8275 ( \8528 , \8491 , \8497 );
or \U$8276 ( \8529 , \8526 , \8527 , \8528 );
and \U$8277 ( \8530 , \8404 , \8445 );
and \U$8278 ( \8531 , \8445 , \8485 );
and \U$8279 ( \8532 , \8404 , \8485 );
or \U$8280 ( \8533 , \8530 , \8531 , \8532 );
xor \U$8281 ( \8534 , \8529 , \8533 );
and \U$8282 ( \8535 , \8385 , \8399 );
xor \U$8283 ( \8536 , \8534 , \8535 );
xor \U$8284 ( \8537 , \8525 , \8536 );
and \U$8285 ( \8538 , \8504 , \8508 );
and \U$8286 ( \8539 , \8508 , \8513 );
and \U$8287 ( \8540 , \8504 , \8513 );
or \U$8288 ( \8541 , \8538 , \8539 , \8540 );
and \U$8289 ( \8542 , \8400 , \8486 );
and \U$8290 ( \8543 , \8486 , \8498 );
and \U$8291 ( \8544 , \8400 , \8498 );
or \U$8292 ( \8545 , \8542 , \8543 , \8544 );
xor \U$8293 ( \8546 , \8541 , \8545 );
and \U$8294 ( \8547 , \6029 , \5809 );
and \U$8295 ( \8548 , \6041 , \5807 );
nor \U$8296 ( \8549 , \8547 , \8548 );
xnor \U$8297 ( \8550 , \8549 , \5816 );
and \U$8298 ( \8551 , \6048 , \5829 );
and \U$8299 ( \8552 , \6057 , \5827 );
nor \U$8300 ( \8553 , \8551 , \8552 );
xnor \U$8301 ( \8554 , \8553 , \5836 );
xor \U$8302 ( \8555 , \8550 , \8554 );
nand \U$8303 ( \8556 , \6065 , \5850 );
xnor \U$8304 ( \8557 , \8556 , \5859 );
xor \U$8305 ( \8558 , \8555 , \8557 );
and \U$8306 ( \8559 , \5967 , \5750 );
and \U$8307 ( \8560 , \5979 , \5748 );
nor \U$8308 ( \8561 , \8559 , \8560 );
xnor \U$8309 ( \8562 , \8561 , \5755 );
and \U$8310 ( \8563 , \5986 , \5768 );
and \U$8311 ( \8564 , \5998 , \5766 );
nor \U$8312 ( \8565 , \8563 , \8564 );
xnor \U$8313 ( \8566 , \8565 , \5775 );
xor \U$8314 ( \8567 , \8562 , \8566 );
and \U$8315 ( \8568 , \6006 , \5790 );
and \U$8316 ( \8569 , \6018 , \5788 );
nor \U$8317 ( \8570 , \8568 , \8569 );
xnor \U$8318 ( \8571 , \8570 , \5797 );
xor \U$8319 ( \8572 , \8567 , \8571 );
xnor \U$8320 ( \8573 , \8558 , \8572 );
and \U$8321 ( \8574 , \8474 , \8478 );
and \U$8322 ( \8575 , \8478 , \8483 );
and \U$8323 ( \8576 , \8474 , \8483 );
or \U$8324 ( \8577 , \8574 , \8575 , \8576 );
and \U$8325 ( \8578 , \8459 , \8463 );
and \U$8326 ( \8579 , \8463 , \8468 );
and \U$8327 ( \8580 , \8459 , \8468 );
or \U$8328 ( \8581 , \8578 , \8579 , \8580 );
xor \U$8329 ( \8582 , \8577 , \8581 );
and \U$8330 ( \8583 , \8450 , \8454 );
xor \U$8331 ( \8584 , \8582 , \8583 );
xor \U$8332 ( \8585 , \8573 , \8584 );
and \U$8333 ( \8586 , \8434 , \8438 );
and \U$8334 ( \8587 , \8438 , \8443 );
and \U$8335 ( \8588 , \8434 , \8443 );
or \U$8336 ( \8589 , \8586 , \8587 , \8588 );
and \U$8337 ( \8590 , \8422 , \8426 );
and \U$8338 ( \8591 , \8426 , \8431 );
and \U$8339 ( \8592 , \8422 , \8431 );
or \U$8340 ( \8593 , \8590 , \8591 , \8592 );
xor \U$8341 ( \8594 , \8589 , \8593 );
and \U$8342 ( \8595 , \8408 , \8412 );
and \U$8343 ( \8596 , \8412 , \8417 );
and \U$8344 ( \8597 , \8408 , \8417 );
or \U$8345 ( \8598 , \8595 , \8596 , \8597 );
xor \U$8346 ( \8599 , \8594 , \8598 );
xor \U$8347 ( \8600 , \8585 , \8599 );
and \U$8348 ( \8601 , \8418 , \8432 );
and \U$8349 ( \8602 , \8432 , \8444 );
and \U$8350 ( \8603 , \8418 , \8444 );
or \U$8351 ( \8604 , \8601 , \8602 , \8603 );
and \U$8352 ( \8605 , \5737 , \7026 );
not \U$8353 ( \8606 , \8605 );
xnor \U$8354 ( \8607 , \8606 , \7032 );
xor \U$8355 ( \8608 , \5859 , \8607 );
and \U$8356 ( \8609 , \5758 , \7043 );
and \U$8357 ( \8610 , \5770 , \7041 );
nor \U$8358 ( \8611 , \8609 , \8610 );
xnor \U$8359 ( \8612 , \8611 , \7049 );
xor \U$8360 ( \8613 , \8608 , \8612 );
xor \U$8361 ( \8614 , \8604 , \8613 );
and \U$8362 ( \8615 , \5906 , \7175 );
and \U$8363 ( \8616 , \5918 , \7173 );
nor \U$8364 ( \8617 , \8615 , \8616 );
xnor \U$8365 ( \8618 , \8617 , \7181 );
and \U$8366 ( \8619 , \5925 , \7192 );
and \U$8367 ( \8620 , \5937 , \7190 );
nor \U$8368 ( \8621 , \8619 , \8620 );
xnor \U$8369 ( \8622 , \8621 , \7198 );
xor \U$8370 ( \8623 , \8618 , \8622 );
and \U$8371 ( \8624 , \5945 , \7203 );
and \U$8372 ( \8625 , \5957 , \7201 );
nor \U$8373 ( \8626 , \8624 , \8625 );
xnor \U$8374 ( \8627 , \8626 , \6824 );
xor \U$8375 ( \8628 , \8623 , \8627 );
and \U$8376 ( \8629 , \5842 , \7117 );
and \U$8377 ( \8630 , \5854 , \7115 );
nor \U$8378 ( \8631 , \8629 , \8630 );
xnor \U$8379 ( \8632 , \8631 , \7123 );
and \U$8380 ( \8633 , \5861 , \7140 );
and \U$8381 ( \8634 , \5873 , \7138 );
nor \U$8382 ( \8635 , \8633 , \8634 );
xnor \U$8383 ( \8636 , \8635 , \7146 );
xor \U$8384 ( \8637 , \8632 , \8636 );
and \U$8385 ( \8638 , \5881 , \7157 );
and \U$8386 ( \8639 , \5893 , \7155 );
nor \U$8387 ( \8640 , \8638 , \8639 );
xnor \U$8388 ( \8641 , \8640 , \7163 );
xor \U$8389 ( \8642 , \8637 , \8641 );
xor \U$8390 ( \8643 , \8628 , \8642 );
and \U$8391 ( \8644 , \5780 , \7061 );
and \U$8392 ( \8645 , \5792 , \7059 );
nor \U$8393 ( \8646 , \8644 , \8645 );
xnor \U$8394 ( \8647 , \8646 , \7067 );
and \U$8395 ( \8648 , \5799 , \7082 );
and \U$8396 ( \8649 , \5811 , \7080 );
nor \U$8397 ( \8650 , \8648 , \8649 );
xnor \U$8398 ( \8651 , \8650 , \7088 );
xor \U$8399 ( \8652 , \8647 , \8651 );
and \U$8400 ( \8653 , \5819 , \7099 );
and \U$8401 ( \8654 , \5831 , \7097 );
nor \U$8402 ( \8655 , \8653 , \8654 );
xnor \U$8403 ( \8656 , \8655 , \7105 );
xor \U$8404 ( \8657 , \8652 , \8656 );
xor \U$8405 ( \8658 , \8643 , \8657 );
xor \U$8406 ( \8659 , \8614 , \8658 );
xor \U$8407 ( \8660 , \8600 , \8659 );
and \U$8408 ( \8661 , \8389 , \8393 );
and \U$8409 ( \8662 , \8393 , \8398 );
and \U$8410 ( \8663 , \8389 , \8398 );
or \U$8411 ( \8664 , \8661 , \8662 , \8663 );
and \U$8412 ( \8665 , \8375 , \8379 );
and \U$8413 ( \8666 , \8379 , \8384 );
and \U$8414 ( \8667 , \8375 , \8384 );
or \U$8415 ( \8668 , \8665 , \8666 , \8667 );
xor \U$8416 ( \8669 , \8664 , \8668 );
and \U$8417 ( \8670 , \8455 , \8469 );
and \U$8418 ( \8671 , \8469 , \8484 );
and \U$8419 ( \8672 , \8455 , \8484 );
or \U$8420 ( \8673 , \8670 , \8671 , \8672 );
xor \U$8421 ( \8674 , \8669 , \8673 );
xor \U$8422 ( \8675 , \8660 , \8674 );
xor \U$8423 ( \8676 , \8546 , \8675 );
xor \U$8424 ( \8677 , \8537 , \8676 );
and \U$8425 ( \8678 , \8365 , \8366 );
and \U$8426 ( \8679 , \8366 , \8515 );
and \U$8427 ( \8680 , \8365 , \8515 );
or \U$8428 ( \8681 , \8678 , \8679 , \8680 );
nor \U$8429 ( \8682 , \8677 , \8681 );
nor \U$8430 ( \8683 , \8521 , \8682 );
and \U$8431 ( \8684 , \8541 , \8545 );
and \U$8432 ( \8685 , \8545 , \8675 );
and \U$8433 ( \8686 , \8541 , \8675 );
or \U$8434 ( \8687 , \8684 , \8685 , \8686 );
and \U$8435 ( \8688 , \8664 , \8668 );
and \U$8436 ( \8689 , \8668 , \8673 );
and \U$8437 ( \8690 , \8664 , \8673 );
or \U$8438 ( \8691 , \8688 , \8689 , \8690 );
and \U$8439 ( \8692 , \8604 , \8613 );
and \U$8440 ( \8693 , \8613 , \8658 );
and \U$8441 ( \8694 , \8604 , \8658 );
or \U$8442 ( \8695 , \8692 , \8693 , \8694 );
xor \U$8443 ( \8696 , \8691 , \8695 );
and \U$8444 ( \8697 , \8573 , \8584 );
and \U$8445 ( \8698 , \8584 , \8599 );
and \U$8446 ( \8699 , \8573 , \8599 );
or \U$8447 ( \8700 , \8697 , \8698 , \8699 );
xor \U$8448 ( \8701 , \8696 , \8700 );
xor \U$8449 ( \8702 , \8687 , \8701 );
and \U$8450 ( \8703 , \8529 , \8533 );
and \U$8451 ( \8704 , \8533 , \8535 );
and \U$8452 ( \8705 , \8529 , \8535 );
or \U$8453 ( \8706 , \8703 , \8704 , \8705 );
and \U$8454 ( \8707 , \8600 , \8659 );
and \U$8455 ( \8708 , \8659 , \8674 );
and \U$8456 ( \8709 , \8600 , \8674 );
or \U$8457 ( \8710 , \8707 , \8708 , \8709 );
xor \U$8458 ( \8711 , \8706 , \8710 );
and \U$8459 ( \8712 , \8618 , \8622 );
and \U$8460 ( \8713 , \8622 , \8627 );
and \U$8461 ( \8714 , \8618 , \8627 );
or \U$8462 ( \8715 , \8712 , \8713 , \8714 );
and \U$8463 ( \8716 , \8562 , \8566 );
and \U$8464 ( \8717 , \8566 , \8571 );
and \U$8465 ( \8718 , \8562 , \8571 );
or \U$8466 ( \8719 , \8716 , \8717 , \8718 );
xor \U$8467 ( \8720 , \8715 , \8719 );
and \U$8468 ( \8721 , \8550 , \8554 );
and \U$8469 ( \8722 , \8554 , \8557 );
and \U$8470 ( \8723 , \8550 , \8557 );
or \U$8471 ( \8724 , \8721 , \8722 , \8723 );
xor \U$8472 ( \8725 , \8720 , \8724 );
and \U$8473 ( \8726 , \5859 , \8607 );
and \U$8474 ( \8727 , \8607 , \8612 );
and \U$8475 ( \8728 , \5859 , \8612 );
or \U$8476 ( \8729 , \8726 , \8727 , \8728 );
and \U$8477 ( \8730 , \8647 , \8651 );
and \U$8478 ( \8731 , \8651 , \8656 );
and \U$8479 ( \8732 , \8647 , \8656 );
or \U$8480 ( \8733 , \8730 , \8731 , \8732 );
xor \U$8481 ( \8734 , \8729 , \8733 );
and \U$8482 ( \8735 , \8632 , \8636 );
and \U$8483 ( \8736 , \8636 , \8641 );
and \U$8484 ( \8737 , \8632 , \8641 );
or \U$8485 ( \8738 , \8735 , \8736 , \8737 );
xor \U$8486 ( \8739 , \8734 , \8738 );
xor \U$8487 ( \8740 , \8725 , \8739 );
and \U$8488 ( \8741 , \8628 , \8642 );
and \U$8489 ( \8742 , \8642 , \8657 );
and \U$8490 ( \8743 , \8628 , \8657 );
or \U$8491 ( \8744 , \8741 , \8742 , \8743 );
and \U$8492 ( \8745 , \5873 , \7140 );
and \U$8493 ( \8746 , \5842 , \7138 );
nor \U$8494 ( \8747 , \8745 , \8746 );
xnor \U$8495 ( \8748 , \8747 , \7146 );
and \U$8496 ( \8749 , \5893 , \7157 );
and \U$8497 ( \8750 , \5861 , \7155 );
nor \U$8498 ( \8751 , \8749 , \8750 );
xnor \U$8499 ( \8752 , \8751 , \7163 );
xor \U$8500 ( \8753 , \8748 , \8752 );
and \U$8501 ( \8754 , \5918 , \7175 );
and \U$8502 ( \8755 , \5881 , \7173 );
nor \U$8503 ( \8756 , \8754 , \8755 );
xnor \U$8504 ( \8757 , \8756 , \7181 );
xor \U$8505 ( \8758 , \8753 , \8757 );
and \U$8506 ( \8759 , \5811 , \7082 );
and \U$8507 ( \8760 , \5780 , \7080 );
nor \U$8508 ( \8761 , \8759 , \8760 );
xnor \U$8509 ( \8762 , \8761 , \7088 );
and \U$8510 ( \8763 , \5831 , \7099 );
and \U$8511 ( \8764 , \5799 , \7097 );
nor \U$8512 ( \8765 , \8763 , \8764 );
xnor \U$8513 ( \8766 , \8765 , \7105 );
xor \U$8514 ( \8767 , \8762 , \8766 );
and \U$8515 ( \8768 , \5854 , \7117 );
and \U$8516 ( \8769 , \5819 , \7115 );
nor \U$8517 ( \8770 , \8768 , \8769 );
xnor \U$8518 ( \8771 , \8770 , \7123 );
xor \U$8519 ( \8772 , \8767 , \8771 );
xor \U$8520 ( \8773 , \8758 , \8772 );
not \U$8521 ( \8774 , \7032 );
and \U$8522 ( \8775 , \5770 , \7043 );
and \U$8523 ( \8776 , \5737 , \7041 );
nor \U$8524 ( \8777 , \8775 , \8776 );
xnor \U$8525 ( \8778 , \8777 , \7049 );
xor \U$8526 ( \8779 , \8774 , \8778 );
and \U$8527 ( \8780 , \5792 , \7061 );
and \U$8528 ( \8781 , \5758 , \7059 );
nor \U$8529 ( \8782 , \8780 , \8781 );
xnor \U$8530 ( \8783 , \8782 , \7067 );
xor \U$8531 ( \8784 , \8779 , \8783 );
xor \U$8532 ( \8785 , \8773 , \8784 );
xor \U$8533 ( \8786 , \8744 , \8785 );
and \U$8534 ( \8787 , \6057 , \5829 );
and \U$8535 ( \8788 , \6029 , \5827 );
nor \U$8536 ( \8789 , \8787 , \8788 );
xnor \U$8537 ( \8790 , \8789 , \5836 );
and \U$8538 ( \8791 , \6065 , \5852 );
and \U$8539 ( \8792 , \6048 , \5850 );
nor \U$8540 ( \8793 , \8791 , \8792 );
xnor \U$8541 ( \8794 , \8793 , \5859 );
xor \U$8542 ( \8795 , \8790 , \8794 );
and \U$8543 ( \8796 , \5998 , \5768 );
and \U$8544 ( \8797 , \5967 , \5766 );
nor \U$8545 ( \8798 , \8796 , \8797 );
xnor \U$8546 ( \8799 , \8798 , \5775 );
and \U$8547 ( \8800 , \6018 , \5790 );
and \U$8548 ( \8801 , \5986 , \5788 );
nor \U$8549 ( \8802 , \8800 , \8801 );
xnor \U$8550 ( \8803 , \8802 , \5797 );
xor \U$8551 ( \8804 , \8799 , \8803 );
and \U$8552 ( \8805 , \6041 , \5809 );
and \U$8553 ( \8806 , \6006 , \5807 );
nor \U$8554 ( \8807 , \8805 , \8806 );
xnor \U$8555 ( \8808 , \8807 , \5816 );
xor \U$8556 ( \8809 , \8804 , \8808 );
xor \U$8557 ( \8810 , \8795 , \8809 );
and \U$8558 ( \8811 , \5937 , \7192 );
and \U$8559 ( \8812 , \5906 , \7190 );
nor \U$8560 ( \8813 , \8811 , \8812 );
xnor \U$8561 ( \8814 , \8813 , \7198 );
and \U$8562 ( \8815 , \5957 , \7203 );
and \U$8563 ( \8816 , \5925 , \7201 );
nor \U$8564 ( \8817 , \8815 , \8816 );
xnor \U$8565 ( \8818 , \8817 , \6824 );
xor \U$8566 ( \8819 , \8814 , \8818 );
and \U$8567 ( \8820 , \5979 , \5750 );
and \U$8568 ( \8821 , \5945 , \5748 );
nor \U$8569 ( \8822 , \8820 , \8821 );
xnor \U$8570 ( \8823 , \8822 , \5755 );
xor \U$8571 ( \8824 , \8819 , \8823 );
xor \U$8572 ( \8825 , \8810 , \8824 );
xor \U$8573 ( \8826 , \8786 , \8825 );
xor \U$8574 ( \8827 , \8740 , \8826 );
and \U$8575 ( \8828 , \8589 , \8593 );
and \U$8576 ( \8829 , \8593 , \8598 );
and \U$8577 ( \8830 , \8589 , \8598 );
or \U$8578 ( \8831 , \8828 , \8829 , \8830 );
and \U$8579 ( \8832 , \8577 , \8581 );
and \U$8580 ( \8833 , \8581 , \8583 );
and \U$8581 ( \8834 , \8577 , \8583 );
or \U$8582 ( \8835 , \8832 , \8833 , \8834 );
xor \U$8583 ( \8836 , \8831 , \8835 );
or \U$8584 ( \8837 , \8558 , \8572 );
xor \U$8585 ( \8838 , \8836 , \8837 );
xor \U$8586 ( \8839 , \8827 , \8838 );
xor \U$8587 ( \8840 , \8711 , \8839 );
xor \U$8588 ( \8841 , \8702 , \8840 );
and \U$8589 ( \8842 , \8525 , \8536 );
and \U$8590 ( \8843 , \8536 , \8676 );
and \U$8591 ( \8844 , \8525 , \8676 );
or \U$8592 ( \8845 , \8842 , \8843 , \8844 );
nor \U$8593 ( \8846 , \8841 , \8845 );
and \U$8594 ( \8847 , \8706 , \8710 );
and \U$8595 ( \8848 , \8710 , \8839 );
and \U$8596 ( \8849 , \8706 , \8839 );
or \U$8597 ( \8850 , \8847 , \8848 , \8849 );
and \U$8598 ( \8851 , \8831 , \8835 );
and \U$8599 ( \8852 , \8835 , \8837 );
and \U$8600 ( \8853 , \8831 , \8837 );
or \U$8601 ( \8854 , \8851 , \8852 , \8853 );
and \U$8602 ( \8855 , \8744 , \8785 );
and \U$8603 ( \8856 , \8785 , \8825 );
and \U$8604 ( \8857 , \8744 , \8825 );
or \U$8605 ( \8858 , \8855 , \8856 , \8857 );
xor \U$8606 ( \8859 , \8854 , \8858 );
and \U$8607 ( \8860 , \8725 , \8739 );
xor \U$8608 ( \8861 , \8859 , \8860 );
xor \U$8609 ( \8862 , \8850 , \8861 );
and \U$8610 ( \8863 , \8691 , \8695 );
and \U$8611 ( \8864 , \8695 , \8700 );
and \U$8612 ( \8865 , \8691 , \8700 );
or \U$8613 ( \8866 , \8863 , \8864 , \8865 );
and \U$8614 ( \8867 , \8740 , \8826 );
and \U$8615 ( \8868 , \8826 , \8838 );
and \U$8616 ( \8869 , \8740 , \8838 );
or \U$8617 ( \8870 , \8867 , \8868 , \8869 );
xor \U$8618 ( \8871 , \8866 , \8870 );
and \U$8619 ( \8872 , \6029 , \5829 );
and \U$8620 ( \8873 , \6041 , \5827 );
nor \U$8621 ( \8874 , \8872 , \8873 );
xnor \U$8622 ( \8875 , \8874 , \5836 );
and \U$8623 ( \8876 , \6048 , \5852 );
and \U$8624 ( \8877 , \6057 , \5850 );
nor \U$8625 ( \8878 , \8876 , \8877 );
xnor \U$8626 ( \8879 , \8878 , \5859 );
xor \U$8627 ( \8880 , \8875 , \8879 );
nand \U$8628 ( \8881 , \6065 , \5869 );
xnor \U$8629 ( \8882 , \8881 , \5878 );
xor \U$8630 ( \8883 , \8880 , \8882 );
and \U$8631 ( \8884 , \5967 , \5768 );
and \U$8632 ( \8885 , \5979 , \5766 );
nor \U$8633 ( \8886 , \8884 , \8885 );
xnor \U$8634 ( \8887 , \8886 , \5775 );
and \U$8635 ( \8888 , \5986 , \5790 );
and \U$8636 ( \8889 , \5998 , \5788 );
nor \U$8637 ( \8890 , \8888 , \8889 );
xnor \U$8638 ( \8891 , \8890 , \5797 );
xor \U$8639 ( \8892 , \8887 , \8891 );
and \U$8640 ( \8893 , \6006 , \5809 );
and \U$8641 ( \8894 , \6018 , \5807 );
nor \U$8642 ( \8895 , \8893 , \8894 );
xnor \U$8643 ( \8896 , \8895 , \5816 );
xor \U$8644 ( \8897 , \8892 , \8896 );
xnor \U$8645 ( \8898 , \8883 , \8897 );
and \U$8646 ( \8899 , \8814 , \8818 );
and \U$8647 ( \8900 , \8818 , \8823 );
and \U$8648 ( \8901 , \8814 , \8823 );
or \U$8649 ( \8902 , \8899 , \8900 , \8901 );
and \U$8650 ( \8903 , \8799 , \8803 );
and \U$8651 ( \8904 , \8803 , \8808 );
and \U$8652 ( \8905 , \8799 , \8808 );
or \U$8653 ( \8906 , \8903 , \8904 , \8905 );
xor \U$8654 ( \8907 , \8902 , \8906 );
and \U$8655 ( \8908 , \8790 , \8794 );
xor \U$8656 ( \8909 , \8907 , \8908 );
xor \U$8657 ( \8910 , \8898 , \8909 );
and \U$8658 ( \8911 , \8774 , \8778 );
and \U$8659 ( \8912 , \8778 , \8783 );
and \U$8660 ( \8913 , \8774 , \8783 );
or \U$8661 ( \8914 , \8911 , \8912 , \8913 );
and \U$8662 ( \8915 , \8762 , \8766 );
and \U$8663 ( \8916 , \8766 , \8771 );
and \U$8664 ( \8917 , \8762 , \8771 );
or \U$8665 ( \8918 , \8915 , \8916 , \8917 );
xor \U$8666 ( \8919 , \8914 , \8918 );
and \U$8667 ( \8920 , \8748 , \8752 );
and \U$8668 ( \8921 , \8752 , \8757 );
and \U$8669 ( \8922 , \8748 , \8757 );
or \U$8670 ( \8923 , \8920 , \8921 , \8922 );
xor \U$8671 ( \8924 , \8919 , \8923 );
xor \U$8672 ( \8925 , \8910 , \8924 );
and \U$8673 ( \8926 , \8758 , \8772 );
and \U$8674 ( \8927 , \8772 , \8784 );
and \U$8675 ( \8928 , \8758 , \8784 );
or \U$8676 ( \8929 , \8926 , \8927 , \8928 );
and \U$8677 ( \8930 , \5737 , \7043 );
not \U$8678 ( \8931 , \8930 );
xnor \U$8679 ( \8932 , \8931 , \7049 );
xor \U$8680 ( \8933 , \5878 , \8932 );
and \U$8681 ( \8934 , \5758 , \7061 );
and \U$8682 ( \8935 , \5770 , \7059 );
nor \U$8683 ( \8936 , \8934 , \8935 );
xnor \U$8684 ( \8937 , \8936 , \7067 );
xor \U$8685 ( \8938 , \8933 , \8937 );
xor \U$8686 ( \8939 , \8929 , \8938 );
and \U$8687 ( \8940 , \5906 , \7192 );
and \U$8688 ( \8941 , \5918 , \7190 );
nor \U$8689 ( \8942 , \8940 , \8941 );
xnor \U$8690 ( \8943 , \8942 , \7198 );
and \U$8691 ( \8944 , \5925 , \7203 );
and \U$8692 ( \8945 , \5937 , \7201 );
nor \U$8693 ( \8946 , \8944 , \8945 );
xnor \U$8694 ( \8947 , \8946 , \6824 );
xor \U$8695 ( \8948 , \8943 , \8947 );
and \U$8696 ( \8949 , \5945 , \5750 );
and \U$8697 ( \8950 , \5957 , \5748 );
nor \U$8698 ( \8951 , \8949 , \8950 );
xnor \U$8699 ( \8952 , \8951 , \5755 );
xor \U$8700 ( \8953 , \8948 , \8952 );
and \U$8701 ( \8954 , \5842 , \7140 );
and \U$8702 ( \8955 , \5854 , \7138 );
nor \U$8703 ( \8956 , \8954 , \8955 );
xnor \U$8704 ( \8957 , \8956 , \7146 );
and \U$8705 ( \8958 , \5861 , \7157 );
and \U$8706 ( \8959 , \5873 , \7155 );
nor \U$8707 ( \8960 , \8958 , \8959 );
xnor \U$8708 ( \8961 , \8960 , \7163 );
xor \U$8709 ( \8962 , \8957 , \8961 );
and \U$8710 ( \8963 , \5881 , \7175 );
and \U$8711 ( \8964 , \5893 , \7173 );
nor \U$8712 ( \8965 , \8963 , \8964 );
xnor \U$8713 ( \8966 , \8965 , \7181 );
xor \U$8714 ( \8967 , \8962 , \8966 );
xor \U$8715 ( \8968 , \8953 , \8967 );
and \U$8716 ( \8969 , \5780 , \7082 );
and \U$8717 ( \8970 , \5792 , \7080 );
nor \U$8718 ( \8971 , \8969 , \8970 );
xnor \U$8719 ( \8972 , \8971 , \7088 );
and \U$8720 ( \8973 , \5799 , \7099 );
and \U$8721 ( \8974 , \5811 , \7097 );
nor \U$8722 ( \8975 , \8973 , \8974 );
xnor \U$8723 ( \8976 , \8975 , \7105 );
xor \U$8724 ( \8977 , \8972 , \8976 );
and \U$8725 ( \8978 , \5819 , \7117 );
and \U$8726 ( \8979 , \5831 , \7115 );
nor \U$8727 ( \8980 , \8978 , \8979 );
xnor \U$8728 ( \8981 , \8980 , \7123 );
xor \U$8729 ( \8982 , \8977 , \8981 );
xor \U$8730 ( \8983 , \8968 , \8982 );
xor \U$8731 ( \8984 , \8939 , \8983 );
xor \U$8732 ( \8985 , \8925 , \8984 );
and \U$8733 ( \8986 , \8729 , \8733 );
and \U$8734 ( \8987 , \8733 , \8738 );
and \U$8735 ( \8988 , \8729 , \8738 );
or \U$8736 ( \8989 , \8986 , \8987 , \8988 );
and \U$8737 ( \8990 , \8715 , \8719 );
and \U$8738 ( \8991 , \8719 , \8724 );
and \U$8739 ( \8992 , \8715 , \8724 );
or \U$8740 ( \8993 , \8990 , \8991 , \8992 );
xor \U$8741 ( \8994 , \8989 , \8993 );
and \U$8742 ( \8995 , \8795 , \8809 );
and \U$8743 ( \8996 , \8809 , \8824 );
and \U$8744 ( \8997 , \8795 , \8824 );
or \U$8745 ( \8998 , \8995 , \8996 , \8997 );
xor \U$8746 ( \8999 , \8994 , \8998 );
xor \U$8747 ( \9000 , \8985 , \8999 );
xor \U$8748 ( \9001 , \8871 , \9000 );
xor \U$8749 ( \9002 , \8862 , \9001 );
and \U$8750 ( \9003 , \8687 , \8701 );
and \U$8751 ( \9004 , \8701 , \8840 );
and \U$8752 ( \9005 , \8687 , \8840 );
or \U$8753 ( \9006 , \9003 , \9004 , \9005 );
nor \U$8754 ( \9007 , \9002 , \9006 );
nor \U$8755 ( \9008 , \8846 , \9007 );
nand \U$8756 ( \9009 , \8683 , \9008 );
nor \U$8757 ( \9010 , \8361 , \9009 );
and \U$8758 ( \9011 , \8866 , \8870 );
and \U$8759 ( \9012 , \8870 , \9000 );
and \U$8760 ( \9013 , \8866 , \9000 );
or \U$8761 ( \9014 , \9011 , \9012 , \9013 );
and \U$8762 ( \9015 , \8989 , \8993 );
and \U$8763 ( \9016 , \8993 , \8998 );
and \U$8764 ( \9017 , \8989 , \8998 );
or \U$8765 ( \9018 , \9015 , \9016 , \9017 );
and \U$8766 ( \9019 , \8929 , \8938 );
and \U$8767 ( \9020 , \8938 , \8983 );
and \U$8768 ( \9021 , \8929 , \8983 );
or \U$8769 ( \9022 , \9019 , \9020 , \9021 );
xor \U$8770 ( \9023 , \9018 , \9022 );
and \U$8771 ( \9024 , \8898 , \8909 );
and \U$8772 ( \9025 , \8909 , \8924 );
and \U$8773 ( \9026 , \8898 , \8924 );
or \U$8774 ( \9027 , \9024 , \9025 , \9026 );
xor \U$8775 ( \9028 , \9023 , \9027 );
xor \U$8776 ( \9029 , \9014 , \9028 );
and \U$8777 ( \9030 , \8854 , \8858 );
and \U$8778 ( \9031 , \8858 , \8860 );
and \U$8779 ( \9032 , \8854 , \8860 );
or \U$8780 ( \9033 , \9030 , \9031 , \9032 );
and \U$8781 ( \9034 , \8925 , \8984 );
and \U$8782 ( \9035 , \8984 , \8999 );
and \U$8783 ( \9036 , \8925 , \8999 );
or \U$8784 ( \9037 , \9034 , \9035 , \9036 );
xor \U$8785 ( \9038 , \9033 , \9037 );
and \U$8786 ( \9039 , \8943 , \8947 );
and \U$8787 ( \9040 , \8947 , \8952 );
and \U$8788 ( \9041 , \8943 , \8952 );
or \U$8789 ( \9042 , \9039 , \9040 , \9041 );
and \U$8790 ( \9043 , \8887 , \8891 );
and \U$8791 ( \9044 , \8891 , \8896 );
and \U$8792 ( \9045 , \8887 , \8896 );
or \U$8793 ( \9046 , \9043 , \9044 , \9045 );
xor \U$8794 ( \9047 , \9042 , \9046 );
and \U$8795 ( \9048 , \8875 , \8879 );
and \U$8796 ( \9049 , \8879 , \8882 );
and \U$8797 ( \9050 , \8875 , \8882 );
or \U$8798 ( \9051 , \9048 , \9049 , \9050 );
xor \U$8799 ( \9052 , \9047 , \9051 );
and \U$8800 ( \9053 , \5878 , \8932 );
and \U$8801 ( \9054 , \8932 , \8937 );
and \U$8802 ( \9055 , \5878 , \8937 );
or \U$8803 ( \9056 , \9053 , \9054 , \9055 );
and \U$8804 ( \9057 , \8972 , \8976 );
and \U$8805 ( \9058 , \8976 , \8981 );
and \U$8806 ( \9059 , \8972 , \8981 );
or \U$8807 ( \9060 , \9057 , \9058 , \9059 );
xor \U$8808 ( \9061 , \9056 , \9060 );
and \U$8809 ( \9062 , \8957 , \8961 );
and \U$8810 ( \9063 , \8961 , \8966 );
and \U$8811 ( \9064 , \8957 , \8966 );
or \U$8812 ( \9065 , \9062 , \9063 , \9064 );
xor \U$8813 ( \9066 , \9061 , \9065 );
xor \U$8814 ( \9067 , \9052 , \9066 );
and \U$8815 ( \9068 , \8953 , \8967 );
and \U$8816 ( \9069 , \8967 , \8982 );
and \U$8817 ( \9070 , \8953 , \8982 );
or \U$8818 ( \9071 , \9068 , \9069 , \9070 );
and \U$8819 ( \9072 , \5873 , \7157 );
and \U$8820 ( \9073 , \5842 , \7155 );
nor \U$8821 ( \9074 , \9072 , \9073 );
xnor \U$8822 ( \9075 , \9074 , \7163 );
and \U$8823 ( \9076 , \5893 , \7175 );
and \U$8824 ( \9077 , \5861 , \7173 );
nor \U$8825 ( \9078 , \9076 , \9077 );
xnor \U$8826 ( \9079 , \9078 , \7181 );
xor \U$8827 ( \9080 , \9075 , \9079 );
and \U$8828 ( \9081 , \5918 , \7192 );
and \U$8829 ( \9082 , \5881 , \7190 );
nor \U$8830 ( \9083 , \9081 , \9082 );
xnor \U$8831 ( \9084 , \9083 , \7198 );
xor \U$8832 ( \9085 , \9080 , \9084 );
and \U$8833 ( \9086 , \5811 , \7099 );
and \U$8834 ( \9087 , \5780 , \7097 );
nor \U$8835 ( \9088 , \9086 , \9087 );
xnor \U$8836 ( \9089 , \9088 , \7105 );
and \U$8837 ( \9090 , \5831 , \7117 );
and \U$8838 ( \9091 , \5799 , \7115 );
nor \U$8839 ( \9092 , \9090 , \9091 );
xnor \U$8840 ( \9093 , \9092 , \7123 );
xor \U$8841 ( \9094 , \9089 , \9093 );
and \U$8842 ( \9095 , \5854 , \7140 );
and \U$8843 ( \9096 , \5819 , \7138 );
nor \U$8844 ( \9097 , \9095 , \9096 );
xnor \U$8845 ( \9098 , \9097 , \7146 );
xor \U$8846 ( \9099 , \9094 , \9098 );
xor \U$8847 ( \9100 , \9085 , \9099 );
not \U$8848 ( \9101 , \7049 );
and \U$8849 ( \9102 , \5770 , \7061 );
and \U$8850 ( \9103 , \5737 , \7059 );
nor \U$8851 ( \9104 , \9102 , \9103 );
xnor \U$8852 ( \9105 , \9104 , \7067 );
xor \U$8853 ( \9106 , \9101 , \9105 );
and \U$8854 ( \9107 , \5792 , \7082 );
and \U$8855 ( \9108 , \5758 , \7080 );
nor \U$8856 ( \9109 , \9107 , \9108 );
xnor \U$8857 ( \9110 , \9109 , \7088 );
xor \U$8858 ( \9111 , \9106 , \9110 );
xor \U$8859 ( \9112 , \9100 , \9111 );
xor \U$8860 ( \9113 , \9071 , \9112 );
and \U$8861 ( \9114 , \6057 , \5852 );
and \U$8862 ( \9115 , \6029 , \5850 );
nor \U$8863 ( \9116 , \9114 , \9115 );
xnor \U$8864 ( \9117 , \9116 , \5859 );
and \U$8865 ( \9118 , \6065 , \5871 );
and \U$8866 ( \9119 , \6048 , \5869 );
nor \U$8867 ( \9120 , \9118 , \9119 );
xnor \U$8868 ( \9121 , \9120 , \5878 );
xor \U$8869 ( \9122 , \9117 , \9121 );
and \U$8870 ( \9123 , \5998 , \5790 );
and \U$8871 ( \9124 , \5967 , \5788 );
nor \U$8872 ( \9125 , \9123 , \9124 );
xnor \U$8873 ( \9126 , \9125 , \5797 );
and \U$8874 ( \9127 , \6018 , \5809 );
and \U$8875 ( \9128 , \5986 , \5807 );
nor \U$8876 ( \9129 , \9127 , \9128 );
xnor \U$8877 ( \9130 , \9129 , \5816 );
xor \U$8878 ( \9131 , \9126 , \9130 );
and \U$8879 ( \9132 , \6041 , \5829 );
and \U$8880 ( \9133 , \6006 , \5827 );
nor \U$8881 ( \9134 , \9132 , \9133 );
xnor \U$8882 ( \9135 , \9134 , \5836 );
xor \U$8883 ( \9136 , \9131 , \9135 );
xor \U$8884 ( \9137 , \9122 , \9136 );
and \U$8885 ( \9138 , \5937 , \7203 );
and \U$8886 ( \9139 , \5906 , \7201 );
nor \U$8887 ( \9140 , \9138 , \9139 );
xnor \U$8888 ( \9141 , \9140 , \6824 );
and \U$8889 ( \9142 , \5957 , \5750 );
and \U$8890 ( \9143 , \5925 , \5748 );
nor \U$8891 ( \9144 , \9142 , \9143 );
xnor \U$8892 ( \9145 , \9144 , \5755 );
xor \U$8893 ( \9146 , \9141 , \9145 );
and \U$8894 ( \9147 , \5979 , \5768 );
and \U$8895 ( \9148 , \5945 , \5766 );
nor \U$8896 ( \9149 , \9147 , \9148 );
xnor \U$8897 ( \9150 , \9149 , \5775 );
xor \U$8898 ( \9151 , \9146 , \9150 );
xor \U$8899 ( \9152 , \9137 , \9151 );
xor \U$8900 ( \9153 , \9113 , \9152 );
xor \U$8901 ( \9154 , \9067 , \9153 );
and \U$8902 ( \9155 , \8914 , \8918 );
and \U$8903 ( \9156 , \8918 , \8923 );
and \U$8904 ( \9157 , \8914 , \8923 );
or \U$8905 ( \9158 , \9155 , \9156 , \9157 );
and \U$8906 ( \9159 , \8902 , \8906 );
and \U$8907 ( \9160 , \8906 , \8908 );
and \U$8908 ( \9161 , \8902 , \8908 );
or \U$8909 ( \9162 , \9159 , \9160 , \9161 );
xor \U$8910 ( \9163 , \9158 , \9162 );
or \U$8911 ( \9164 , \8883 , \8897 );
xor \U$8912 ( \9165 , \9163 , \9164 );
xor \U$8913 ( \9166 , \9154 , \9165 );
xor \U$8914 ( \9167 , \9038 , \9166 );
xor \U$8915 ( \9168 , \9029 , \9167 );
and \U$8916 ( \9169 , \8850 , \8861 );
and \U$8917 ( \9170 , \8861 , \9001 );
and \U$8918 ( \9171 , \8850 , \9001 );
or \U$8919 ( \9172 , \9169 , \9170 , \9171 );
nor \U$8920 ( \9173 , \9168 , \9172 );
and \U$8921 ( \9174 , \9033 , \9037 );
and \U$8922 ( \9175 , \9037 , \9166 );
and \U$8923 ( \9176 , \9033 , \9166 );
or \U$8924 ( \9177 , \9174 , \9175 , \9176 );
and \U$8925 ( \9178 , \9158 , \9162 );
and \U$8926 ( \9179 , \9162 , \9164 );
and \U$8927 ( \9180 , \9158 , \9164 );
or \U$8928 ( \9181 , \9178 , \9179 , \9180 );
and \U$8929 ( \9182 , \9071 , \9112 );
and \U$8930 ( \9183 , \9112 , \9152 );
and \U$8931 ( \9184 , \9071 , \9152 );
or \U$8932 ( \9185 , \9182 , \9183 , \9184 );
xor \U$8933 ( \9186 , \9181 , \9185 );
and \U$8934 ( \9187 , \9052 , \9066 );
xor \U$8935 ( \9188 , \9186 , \9187 );
xor \U$8936 ( \9189 , \9177 , \9188 );
and \U$8937 ( \9190 , \9018 , \9022 );
and \U$8938 ( \9191 , \9022 , \9027 );
and \U$8939 ( \9192 , \9018 , \9027 );
or \U$8940 ( \9193 , \9190 , \9191 , \9192 );
and \U$8941 ( \9194 , \9067 , \9153 );
and \U$8942 ( \9195 , \9153 , \9165 );
and \U$8943 ( \9196 , \9067 , \9165 );
or \U$8944 ( \9197 , \9194 , \9195 , \9196 );
xor \U$8945 ( \9198 , \9193 , \9197 );
and \U$8946 ( \9199 , \6029 , \5852 );
and \U$8947 ( \9200 , \6041 , \5850 );
nor \U$8948 ( \9201 , \9199 , \9200 );
xnor \U$8949 ( \9202 , \9201 , \5859 );
and \U$8950 ( \9203 , \6048 , \5871 );
and \U$8951 ( \9204 , \6057 , \5869 );
nor \U$8952 ( \9205 , \9203 , \9204 );
xnor \U$8953 ( \9206 , \9205 , \5878 );
xor \U$8954 ( \9207 , \9202 , \9206 );
nand \U$8955 ( \9208 , \6065 , \5889 );
xnor \U$8956 ( \9209 , \9208 , \5898 );
xor \U$8957 ( \9210 , \9207 , \9209 );
and \U$8958 ( \9211 , \5967 , \5790 );
and \U$8959 ( \9212 , \5979 , \5788 );
nor \U$8960 ( \9213 , \9211 , \9212 );
xnor \U$8961 ( \9214 , \9213 , \5797 );
and \U$8962 ( \9215 , \5986 , \5809 );
and \U$8963 ( \9216 , \5998 , \5807 );
nor \U$8964 ( \9217 , \9215 , \9216 );
xnor \U$8965 ( \9218 , \9217 , \5816 );
xor \U$8966 ( \9219 , \9214 , \9218 );
and \U$8967 ( \9220 , \6006 , \5829 );
and \U$8968 ( \9221 , \6018 , \5827 );
nor \U$8969 ( \9222 , \9220 , \9221 );
xnor \U$8970 ( \9223 , \9222 , \5836 );
xor \U$8971 ( \9224 , \9219 , \9223 );
xnor \U$8972 ( \9225 , \9210 , \9224 );
and \U$8973 ( \9226 , \9141 , \9145 );
and \U$8974 ( \9227 , \9145 , \9150 );
and \U$8975 ( \9228 , \9141 , \9150 );
or \U$8976 ( \9229 , \9226 , \9227 , \9228 );
and \U$8977 ( \9230 , \9126 , \9130 );
and \U$8978 ( \9231 , \9130 , \9135 );
and \U$8979 ( \9232 , \9126 , \9135 );
or \U$8980 ( \9233 , \9230 , \9231 , \9232 );
xor \U$8981 ( \9234 , \9229 , \9233 );
and \U$8982 ( \9235 , \9117 , \9121 );
xor \U$8983 ( \9236 , \9234 , \9235 );
xor \U$8984 ( \9237 , \9225 , \9236 );
and \U$8985 ( \9238 , \9101 , \9105 );
and \U$8986 ( \9239 , \9105 , \9110 );
and \U$8987 ( \9240 , \9101 , \9110 );
or \U$8988 ( \9241 , \9238 , \9239 , \9240 );
and \U$8989 ( \9242 , \9089 , \9093 );
and \U$8990 ( \9243 , \9093 , \9098 );
and \U$8991 ( \9244 , \9089 , \9098 );
or \U$8992 ( \9245 , \9242 , \9243 , \9244 );
xor \U$8993 ( \9246 , \9241 , \9245 );
and \U$8994 ( \9247 , \9075 , \9079 );
and \U$8995 ( \9248 , \9079 , \9084 );
and \U$8996 ( \9249 , \9075 , \9084 );
or \U$8997 ( \9250 , \9247 , \9248 , \9249 );
xor \U$8998 ( \9251 , \9246 , \9250 );
xor \U$8999 ( \9252 , \9237 , \9251 );
and \U$9000 ( \9253 , \9085 , \9099 );
and \U$9001 ( \9254 , \9099 , \9111 );
and \U$9002 ( \9255 , \9085 , \9111 );
or \U$9003 ( \9256 , \9253 , \9254 , \9255 );
and \U$9004 ( \9257 , \5737 , \7061 );
not \U$9005 ( \9258 , \9257 );
xnor \U$9006 ( \9259 , \9258 , \7067 );
xor \U$9007 ( \9260 , \5898 , \9259 );
and \U$9008 ( \9261 , \5758 , \7082 );
and \U$9009 ( \9262 , \5770 , \7080 );
nor \U$9010 ( \9263 , \9261 , \9262 );
xnor \U$9011 ( \9264 , \9263 , \7088 );
xor \U$9012 ( \9265 , \9260 , \9264 );
xor \U$9013 ( \9266 , \9256 , \9265 );
and \U$9014 ( \9267 , \5906 , \7203 );
and \U$9015 ( \9268 , \5918 , \7201 );
nor \U$9016 ( \9269 , \9267 , \9268 );
xnor \U$9017 ( \9270 , \9269 , \6824 );
and \U$9018 ( \9271 , \5925 , \5750 );
and \U$9019 ( \9272 , \5937 , \5748 );
nor \U$9020 ( \9273 , \9271 , \9272 );
xnor \U$9021 ( \9274 , \9273 , \5755 );
xor \U$9022 ( \9275 , \9270 , \9274 );
and \U$9023 ( \9276 , \5945 , \5768 );
and \U$9024 ( \9277 , \5957 , \5766 );
nor \U$9025 ( \9278 , \9276 , \9277 );
xnor \U$9026 ( \9279 , \9278 , \5775 );
xor \U$9027 ( \9280 , \9275 , \9279 );
and \U$9028 ( \9281 , \5842 , \7157 );
and \U$9029 ( \9282 , \5854 , \7155 );
nor \U$9030 ( \9283 , \9281 , \9282 );
xnor \U$9031 ( \9284 , \9283 , \7163 );
and \U$9032 ( \9285 , \5861 , \7175 );
and \U$9033 ( \9286 , \5873 , \7173 );
nor \U$9034 ( \9287 , \9285 , \9286 );
xnor \U$9035 ( \9288 , \9287 , \7181 );
xor \U$9036 ( \9289 , \9284 , \9288 );
and \U$9037 ( \9290 , \5881 , \7192 );
and \U$9038 ( \9291 , \5893 , \7190 );
nor \U$9039 ( \9292 , \9290 , \9291 );
xnor \U$9040 ( \9293 , \9292 , \7198 );
xor \U$9041 ( \9294 , \9289 , \9293 );
xor \U$9042 ( \9295 , \9280 , \9294 );
and \U$9043 ( \9296 , \5780 , \7099 );
and \U$9044 ( \9297 , \5792 , \7097 );
nor \U$9045 ( \9298 , \9296 , \9297 );
xnor \U$9046 ( \9299 , \9298 , \7105 );
and \U$9047 ( \9300 , \5799 , \7117 );
and \U$9048 ( \9301 , \5811 , \7115 );
nor \U$9049 ( \9302 , \9300 , \9301 );
xnor \U$9050 ( \9303 , \9302 , \7123 );
xor \U$9051 ( \9304 , \9299 , \9303 );
and \U$9052 ( \9305 , \5819 , \7140 );
and \U$9053 ( \9306 , \5831 , \7138 );
nor \U$9054 ( \9307 , \9305 , \9306 );
xnor \U$9055 ( \9308 , \9307 , \7146 );
xor \U$9056 ( \9309 , \9304 , \9308 );
xor \U$9057 ( \9310 , \9295 , \9309 );
xor \U$9058 ( \9311 , \9266 , \9310 );
xor \U$9059 ( \9312 , \9252 , \9311 );
and \U$9060 ( \9313 , \9056 , \9060 );
and \U$9061 ( \9314 , \9060 , \9065 );
and \U$9062 ( \9315 , \9056 , \9065 );
or \U$9063 ( \9316 , \9313 , \9314 , \9315 );
and \U$9064 ( \9317 , \9042 , \9046 );
and \U$9065 ( \9318 , \9046 , \9051 );
and \U$9066 ( \9319 , \9042 , \9051 );
or \U$9067 ( \9320 , \9317 , \9318 , \9319 );
xor \U$9068 ( \9321 , \9316 , \9320 );
and \U$9069 ( \9322 , \9122 , \9136 );
and \U$9070 ( \9323 , \9136 , \9151 );
and \U$9071 ( \9324 , \9122 , \9151 );
or \U$9072 ( \9325 , \9322 , \9323 , \9324 );
xor \U$9073 ( \9326 , \9321 , \9325 );
xor \U$9074 ( \9327 , \9312 , \9326 );
xor \U$9075 ( \9328 , \9198 , \9327 );
xor \U$9076 ( \9329 , \9189 , \9328 );
and \U$9077 ( \9330 , \9014 , \9028 );
and \U$9078 ( \9331 , \9028 , \9167 );
and \U$9079 ( \9332 , \9014 , \9167 );
or \U$9080 ( \9333 , \9330 , \9331 , \9332 );
nor \U$9081 ( \9334 , \9329 , \9333 );
nor \U$9082 ( \9335 , \9173 , \9334 );
and \U$9083 ( \9336 , \9193 , \9197 );
and \U$9084 ( \9337 , \9197 , \9327 );
and \U$9085 ( \9338 , \9193 , \9327 );
or \U$9086 ( \9339 , \9336 , \9337 , \9338 );
and \U$9087 ( \9340 , \9316 , \9320 );
and \U$9088 ( \9341 , \9320 , \9325 );
and \U$9089 ( \9342 , \9316 , \9325 );
or \U$9090 ( \9343 , \9340 , \9341 , \9342 );
and \U$9091 ( \9344 , \9256 , \9265 );
and \U$9092 ( \9345 , \9265 , \9310 );
and \U$9093 ( \9346 , \9256 , \9310 );
or \U$9094 ( \9347 , \9344 , \9345 , \9346 );
xor \U$9095 ( \9348 , \9343 , \9347 );
and \U$9096 ( \9349 , \9225 , \9236 );
and \U$9097 ( \9350 , \9236 , \9251 );
and \U$9098 ( \9351 , \9225 , \9251 );
or \U$9099 ( \9352 , \9349 , \9350 , \9351 );
xor \U$9100 ( \9353 , \9348 , \9352 );
xor \U$9101 ( \9354 , \9339 , \9353 );
and \U$9102 ( \9355 , \9181 , \9185 );
and \U$9103 ( \9356 , \9185 , \9187 );
and \U$9104 ( \9357 , \9181 , \9187 );
or \U$9105 ( \9358 , \9355 , \9356 , \9357 );
and \U$9106 ( \9359 , \9252 , \9311 );
and \U$9107 ( \9360 , \9311 , \9326 );
and \U$9108 ( \9361 , \9252 , \9326 );
or \U$9109 ( \9362 , \9359 , \9360 , \9361 );
xor \U$9110 ( \9363 , \9358 , \9362 );
and \U$9111 ( \9364 , \9270 , \9274 );
and \U$9112 ( \9365 , \9274 , \9279 );
and \U$9113 ( \9366 , \9270 , \9279 );
or \U$9114 ( \9367 , \9364 , \9365 , \9366 );
and \U$9115 ( \9368 , \9214 , \9218 );
and \U$9116 ( \9369 , \9218 , \9223 );
and \U$9117 ( \9370 , \9214 , \9223 );
or \U$9118 ( \9371 , \9368 , \9369 , \9370 );
xor \U$9119 ( \9372 , \9367 , \9371 );
and \U$9120 ( \9373 , \9202 , \9206 );
and \U$9121 ( \9374 , \9206 , \9209 );
and \U$9122 ( \9375 , \9202 , \9209 );
or \U$9123 ( \9376 , \9373 , \9374 , \9375 );
xor \U$9124 ( \9377 , \9372 , \9376 );
and \U$9125 ( \9378 , \5898 , \9259 );
and \U$9126 ( \9379 , \9259 , \9264 );
and \U$9127 ( \9380 , \5898 , \9264 );
or \U$9128 ( \9381 , \9378 , \9379 , \9380 );
and \U$9129 ( \9382 , \9299 , \9303 );
and \U$9130 ( \9383 , \9303 , \9308 );
and \U$9131 ( \9384 , \9299 , \9308 );
or \U$9132 ( \9385 , \9382 , \9383 , \9384 );
xor \U$9133 ( \9386 , \9381 , \9385 );
and \U$9134 ( \9387 , \9284 , \9288 );
and \U$9135 ( \9388 , \9288 , \9293 );
and \U$9136 ( \9389 , \9284 , \9293 );
or \U$9137 ( \9390 , \9387 , \9388 , \9389 );
xor \U$9138 ( \9391 , \9386 , \9390 );
xor \U$9139 ( \9392 , \9377 , \9391 );
and \U$9140 ( \9393 , \9280 , \9294 );
and \U$9141 ( \9394 , \9294 , \9309 );
and \U$9142 ( \9395 , \9280 , \9309 );
or \U$9143 ( \9396 , \9393 , \9394 , \9395 );
and \U$9144 ( \9397 , \5873 , \7175 );
and \U$9145 ( \9398 , \5842 , \7173 );
nor \U$9146 ( \9399 , \9397 , \9398 );
xnor \U$9147 ( \9400 , \9399 , \7181 );
and \U$9148 ( \9401 , \5893 , \7192 );
and \U$9149 ( \9402 , \5861 , \7190 );
nor \U$9150 ( \9403 , \9401 , \9402 );
xnor \U$9151 ( \9404 , \9403 , \7198 );
xor \U$9152 ( \9405 , \9400 , \9404 );
and \U$9153 ( \9406 , \5918 , \7203 );
and \U$9154 ( \9407 , \5881 , \7201 );
nor \U$9155 ( \9408 , \9406 , \9407 );
xnor \U$9156 ( \9409 , \9408 , \6824 );
xor \U$9157 ( \9410 , \9405 , \9409 );
and \U$9158 ( \9411 , \5811 , \7117 );
and \U$9159 ( \9412 , \5780 , \7115 );
nor \U$9160 ( \9413 , \9411 , \9412 );
xnor \U$9161 ( \9414 , \9413 , \7123 );
and \U$9162 ( \9415 , \5831 , \7140 );
and \U$9163 ( \9416 , \5799 , \7138 );
nor \U$9164 ( \9417 , \9415 , \9416 );
xnor \U$9165 ( \9418 , \9417 , \7146 );
xor \U$9166 ( \9419 , \9414 , \9418 );
and \U$9167 ( \9420 , \5854 , \7157 );
and \U$9168 ( \9421 , \5819 , \7155 );
nor \U$9169 ( \9422 , \9420 , \9421 );
xnor \U$9170 ( \9423 , \9422 , \7163 );
xor \U$9171 ( \9424 , \9419 , \9423 );
xor \U$9172 ( \9425 , \9410 , \9424 );
not \U$9173 ( \9426 , \7067 );
and \U$9174 ( \9427 , \5770 , \7082 );
and \U$9175 ( \9428 , \5737 , \7080 );
nor \U$9176 ( \9429 , \9427 , \9428 );
xnor \U$9177 ( \9430 , \9429 , \7088 );
xor \U$9178 ( \9431 , \9426 , \9430 );
and \U$9179 ( \9432 , \5792 , \7099 );
and \U$9180 ( \9433 , \5758 , \7097 );
nor \U$9181 ( \9434 , \9432 , \9433 );
xnor \U$9182 ( \9435 , \9434 , \7105 );
xor \U$9183 ( \9436 , \9431 , \9435 );
xor \U$9184 ( \9437 , \9425 , \9436 );
xor \U$9185 ( \9438 , \9396 , \9437 );
and \U$9186 ( \9439 , \6057 , \5871 );
and \U$9187 ( \9440 , \6029 , \5869 );
nor \U$9188 ( \9441 , \9439 , \9440 );
xnor \U$9189 ( \9442 , \9441 , \5878 );
and \U$9190 ( \9443 , \6065 , \5891 );
and \U$9191 ( \9444 , \6048 , \5889 );
nor \U$9192 ( \9445 , \9443 , \9444 );
xnor \U$9193 ( \9446 , \9445 , \5898 );
xor \U$9194 ( \9447 , \9442 , \9446 );
and \U$9195 ( \9448 , \5998 , \5809 );
and \U$9196 ( \9449 , \5967 , \5807 );
nor \U$9197 ( \9450 , \9448 , \9449 );
xnor \U$9198 ( \9451 , \9450 , \5816 );
and \U$9199 ( \9452 , \6018 , \5829 );
and \U$9200 ( \9453 , \5986 , \5827 );
nor \U$9201 ( \9454 , \9452 , \9453 );
xnor \U$9202 ( \9455 , \9454 , \5836 );
xor \U$9203 ( \9456 , \9451 , \9455 );
and \U$9204 ( \9457 , \6041 , \5852 );
and \U$9205 ( \9458 , \6006 , \5850 );
nor \U$9206 ( \9459 , \9457 , \9458 );
xnor \U$9207 ( \9460 , \9459 , \5859 );
xor \U$9208 ( \9461 , \9456 , \9460 );
xor \U$9209 ( \9462 , \9447 , \9461 );
and \U$9210 ( \9463 , \5937 , \5750 );
and \U$9211 ( \9464 , \5906 , \5748 );
nor \U$9212 ( \9465 , \9463 , \9464 );
xnor \U$9213 ( \9466 , \9465 , \5755 );
and \U$9214 ( \9467 , \5957 , \5768 );
and \U$9215 ( \9468 , \5925 , \5766 );
nor \U$9216 ( \9469 , \9467 , \9468 );
xnor \U$9217 ( \9470 , \9469 , \5775 );
xor \U$9218 ( \9471 , \9466 , \9470 );
and \U$9219 ( \9472 , \5979 , \5790 );
and \U$9220 ( \9473 , \5945 , \5788 );
nor \U$9221 ( \9474 , \9472 , \9473 );
xnor \U$9222 ( \9475 , \9474 , \5797 );
xor \U$9223 ( \9476 , \9471 , \9475 );
xor \U$9224 ( \9477 , \9462 , \9476 );
xor \U$9225 ( \9478 , \9438 , \9477 );
xor \U$9226 ( \9479 , \9392 , \9478 );
and \U$9227 ( \9480 , \9241 , \9245 );
and \U$9228 ( \9481 , \9245 , \9250 );
and \U$9229 ( \9482 , \9241 , \9250 );
or \U$9230 ( \9483 , \9480 , \9481 , \9482 );
and \U$9231 ( \9484 , \9229 , \9233 );
and \U$9232 ( \9485 , \9233 , \9235 );
and \U$9233 ( \9486 , \9229 , \9235 );
or \U$9234 ( \9487 , \9484 , \9485 , \9486 );
xor \U$9235 ( \9488 , \9483 , \9487 );
or \U$9236 ( \9489 , \9210 , \9224 );
xor \U$9237 ( \9490 , \9488 , \9489 );
xor \U$9238 ( \9491 , \9479 , \9490 );
xor \U$9239 ( \9492 , \9363 , \9491 );
xor \U$9240 ( \9493 , \9354 , \9492 );
and \U$9241 ( \9494 , \9177 , \9188 );
and \U$9242 ( \9495 , \9188 , \9328 );
and \U$9243 ( \9496 , \9177 , \9328 );
or \U$9244 ( \9497 , \9494 , \9495 , \9496 );
nor \U$9245 ( \9498 , \9493 , \9497 );
and \U$9246 ( \9499 , \9358 , \9362 );
and \U$9247 ( \9500 , \9362 , \9491 );
and \U$9248 ( \9501 , \9358 , \9491 );
or \U$9249 ( \9502 , \9499 , \9500 , \9501 );
and \U$9250 ( \9503 , \9483 , \9487 );
and \U$9251 ( \9504 , \9487 , \9489 );
and \U$9252 ( \9505 , \9483 , \9489 );
or \U$9253 ( \9506 , \9503 , \9504 , \9505 );
and \U$9254 ( \9507 , \9396 , \9437 );
and \U$9255 ( \9508 , \9437 , \9477 );
and \U$9256 ( \9509 , \9396 , \9477 );
or \U$9257 ( \9510 , \9507 , \9508 , \9509 );
xor \U$9258 ( \9511 , \9506 , \9510 );
and \U$9259 ( \9512 , \9377 , \9391 );
xor \U$9260 ( \9513 , \9511 , \9512 );
xor \U$9261 ( \9514 , \9502 , \9513 );
and \U$9262 ( \9515 , \9343 , \9347 );
and \U$9263 ( \9516 , \9347 , \9352 );
and \U$9264 ( \9517 , \9343 , \9352 );
or \U$9265 ( \9518 , \9515 , \9516 , \9517 );
and \U$9266 ( \9519 , \9392 , \9478 );
and \U$9267 ( \9520 , \9478 , \9490 );
and \U$9268 ( \9521 , \9392 , \9490 );
or \U$9269 ( \9522 , \9519 , \9520 , \9521 );
xor \U$9270 ( \9523 , \9518 , \9522 );
and \U$9271 ( \9524 , \6029 , \5871 );
and \U$9272 ( \9525 , \6041 , \5869 );
nor \U$9273 ( \9526 , \9524 , \9525 );
xnor \U$9274 ( \9527 , \9526 , \5878 );
and \U$9275 ( \9528 , \6048 , \5891 );
and \U$9276 ( \9529 , \6057 , \5889 );
nor \U$9277 ( \9530 , \9528 , \9529 );
xnor \U$9278 ( \9531 , \9530 , \5898 );
xor \U$9279 ( \9532 , \9527 , \9531 );
nand \U$9280 ( \9533 , \6065 , \5914 );
xnor \U$9281 ( \9534 , \9533 , \5923 );
xor \U$9282 ( \9535 , \9532 , \9534 );
and \U$9283 ( \9536 , \5967 , \5809 );
and \U$9284 ( \9537 , \5979 , \5807 );
nor \U$9285 ( \9538 , \9536 , \9537 );
xnor \U$9286 ( \9539 , \9538 , \5816 );
and \U$9287 ( \9540 , \5986 , \5829 );
and \U$9288 ( \9541 , \5998 , \5827 );
nor \U$9289 ( \9542 , \9540 , \9541 );
xnor \U$9290 ( \9543 , \9542 , \5836 );
xor \U$9291 ( \9544 , \9539 , \9543 );
and \U$9292 ( \9545 , \6006 , \5852 );
and \U$9293 ( \9546 , \6018 , \5850 );
nor \U$9294 ( \9547 , \9545 , \9546 );
xnor \U$9295 ( \9548 , \9547 , \5859 );
xor \U$9296 ( \9549 , \9544 , \9548 );
xnor \U$9297 ( \9550 , \9535 , \9549 );
and \U$9298 ( \9551 , \9466 , \9470 );
and \U$9299 ( \9552 , \9470 , \9475 );
and \U$9300 ( \9553 , \9466 , \9475 );
or \U$9301 ( \9554 , \9551 , \9552 , \9553 );
and \U$9302 ( \9555 , \9451 , \9455 );
and \U$9303 ( \9556 , \9455 , \9460 );
and \U$9304 ( \9557 , \9451 , \9460 );
or \U$9305 ( \9558 , \9555 , \9556 , \9557 );
xor \U$9306 ( \9559 , \9554 , \9558 );
and \U$9307 ( \9560 , \9442 , \9446 );
xor \U$9308 ( \9561 , \9559 , \9560 );
xor \U$9309 ( \9562 , \9550 , \9561 );
and \U$9310 ( \9563 , \9426 , \9430 );
and \U$9311 ( \9564 , \9430 , \9435 );
and \U$9312 ( \9565 , \9426 , \9435 );
or \U$9313 ( \9566 , \9563 , \9564 , \9565 );
and \U$9314 ( \9567 , \9414 , \9418 );
and \U$9315 ( \9568 , \9418 , \9423 );
and \U$9316 ( \9569 , \9414 , \9423 );
or \U$9317 ( \9570 , \9567 , \9568 , \9569 );
xor \U$9318 ( \9571 , \9566 , \9570 );
and \U$9319 ( \9572 , \9400 , \9404 );
and \U$9320 ( \9573 , \9404 , \9409 );
and \U$9321 ( \9574 , \9400 , \9409 );
or \U$9322 ( \9575 , \9572 , \9573 , \9574 );
xor \U$9323 ( \9576 , \9571 , \9575 );
xor \U$9324 ( \9577 , \9562 , \9576 );
and \U$9325 ( \9578 , \9410 , \9424 );
and \U$9326 ( \9579 , \9424 , \9436 );
and \U$9327 ( \9580 , \9410 , \9436 );
or \U$9328 ( \9581 , \9578 , \9579 , \9580 );
and \U$9329 ( \9582 , \5737 , \7082 );
not \U$9330 ( \9583 , \9582 );
xnor \U$9331 ( \9584 , \9583 , \7088 );
xor \U$9332 ( \9585 , \5923 , \9584 );
and \U$9333 ( \9586 , \5758 , \7099 );
and \U$9334 ( \9587 , \5770 , \7097 );
nor \U$9335 ( \9588 , \9586 , \9587 );
xnor \U$9336 ( \9589 , \9588 , \7105 );
xor \U$9337 ( \9590 , \9585 , \9589 );
xor \U$9338 ( \9591 , \9581 , \9590 );
and \U$9339 ( \9592 , \5906 , \5750 );
and \U$9340 ( \9593 , \5918 , \5748 );
nor \U$9341 ( \9594 , \9592 , \9593 );
xnor \U$9342 ( \9595 , \9594 , \5755 );
and \U$9343 ( \9596 , \5925 , \5768 );
and \U$9344 ( \9597 , \5937 , \5766 );
nor \U$9345 ( \9598 , \9596 , \9597 );
xnor \U$9346 ( \9599 , \9598 , \5775 );
xor \U$9347 ( \9600 , \9595 , \9599 );
and \U$9348 ( \9601 , \5945 , \5790 );
and \U$9349 ( \9602 , \5957 , \5788 );
nor \U$9350 ( \9603 , \9601 , \9602 );
xnor \U$9351 ( \9604 , \9603 , \5797 );
xor \U$9352 ( \9605 , \9600 , \9604 );
and \U$9353 ( \9606 , \5842 , \7175 );
and \U$9354 ( \9607 , \5854 , \7173 );
nor \U$9355 ( \9608 , \9606 , \9607 );
xnor \U$9356 ( \9609 , \9608 , \7181 );
and \U$9357 ( \9610 , \5861 , \7192 );
and \U$9358 ( \9611 , \5873 , \7190 );
nor \U$9359 ( \9612 , \9610 , \9611 );
xnor \U$9360 ( \9613 , \9612 , \7198 );
xor \U$9361 ( \9614 , \9609 , \9613 );
and \U$9362 ( \9615 , \5881 , \7203 );
and \U$9363 ( \9616 , \5893 , \7201 );
nor \U$9364 ( \9617 , \9615 , \9616 );
xnor \U$9365 ( \9618 , \9617 , \6824 );
xor \U$9366 ( \9619 , \9614 , \9618 );
xor \U$9367 ( \9620 , \9605 , \9619 );
and \U$9368 ( \9621 , \5780 , \7117 );
and \U$9369 ( \9622 , \5792 , \7115 );
nor \U$9370 ( \9623 , \9621 , \9622 );
xnor \U$9371 ( \9624 , \9623 , \7123 );
and \U$9372 ( \9625 , \5799 , \7140 );
and \U$9373 ( \9626 , \5811 , \7138 );
nor \U$9374 ( \9627 , \9625 , \9626 );
xnor \U$9375 ( \9628 , \9627 , \7146 );
xor \U$9376 ( \9629 , \9624 , \9628 );
and \U$9377 ( \9630 , \5819 , \7157 );
and \U$9378 ( \9631 , \5831 , \7155 );
nor \U$9379 ( \9632 , \9630 , \9631 );
xnor \U$9380 ( \9633 , \9632 , \7163 );
xor \U$9381 ( \9634 , \9629 , \9633 );
xor \U$9382 ( \9635 , \9620 , \9634 );
xor \U$9383 ( \9636 , \9591 , \9635 );
xor \U$9384 ( \9637 , \9577 , \9636 );
and \U$9385 ( \9638 , \9381 , \9385 );
and \U$9386 ( \9639 , \9385 , \9390 );
and \U$9387 ( \9640 , \9381 , \9390 );
or \U$9388 ( \9641 , \9638 , \9639 , \9640 );
and \U$9389 ( \9642 , \9367 , \9371 );
and \U$9390 ( \9643 , \9371 , \9376 );
and \U$9391 ( \9644 , \9367 , \9376 );
or \U$9392 ( \9645 , \9642 , \9643 , \9644 );
xor \U$9393 ( \9646 , \9641 , \9645 );
and \U$9394 ( \9647 , \9447 , \9461 );
and \U$9395 ( \9648 , \9461 , \9476 );
and \U$9396 ( \9649 , \9447 , \9476 );
or \U$9397 ( \9650 , \9647 , \9648 , \9649 );
xor \U$9398 ( \9651 , \9646 , \9650 );
xor \U$9399 ( \9652 , \9637 , \9651 );
xor \U$9400 ( \9653 , \9523 , \9652 );
xor \U$9401 ( \9654 , \9514 , \9653 );
and \U$9402 ( \9655 , \9339 , \9353 );
and \U$9403 ( \9656 , \9353 , \9492 );
and \U$9404 ( \9657 , \9339 , \9492 );
or \U$9405 ( \9658 , \9655 , \9656 , \9657 );
nor \U$9406 ( \9659 , \9654 , \9658 );
nor \U$9407 ( \9660 , \9498 , \9659 );
nand \U$9408 ( \9661 , \9335 , \9660 );
and \U$9409 ( \9662 , \9518 , \9522 );
and \U$9410 ( \9663 , \9522 , \9652 );
and \U$9411 ( \9664 , \9518 , \9652 );
or \U$9412 ( \9665 , \9662 , \9663 , \9664 );
and \U$9413 ( \9666 , \9641 , \9645 );
and \U$9414 ( \9667 , \9645 , \9650 );
and \U$9415 ( \9668 , \9641 , \9650 );
or \U$9416 ( \9669 , \9666 , \9667 , \9668 );
and \U$9417 ( \9670 , \9581 , \9590 );
and \U$9418 ( \9671 , \9590 , \9635 );
and \U$9419 ( \9672 , \9581 , \9635 );
or \U$9420 ( \9673 , \9670 , \9671 , \9672 );
xor \U$9421 ( \9674 , \9669 , \9673 );
and \U$9422 ( \9675 , \9550 , \9561 );
and \U$9423 ( \9676 , \9561 , \9576 );
and \U$9424 ( \9677 , \9550 , \9576 );
or \U$9425 ( \9678 , \9675 , \9676 , \9677 );
xor \U$9426 ( \9679 , \9674 , \9678 );
xor \U$9427 ( \9680 , \9665 , \9679 );
and \U$9428 ( \9681 , \9506 , \9510 );
and \U$9429 ( \9682 , \9510 , \9512 );
and \U$9430 ( \9683 , \9506 , \9512 );
or \U$9431 ( \9684 , \9681 , \9682 , \9683 );
and \U$9432 ( \9685 , \9577 , \9636 );
and \U$9433 ( \9686 , \9636 , \9651 );
and \U$9434 ( \9687 , \9577 , \9651 );
or \U$9435 ( \9688 , \9685 , \9686 , \9687 );
xor \U$9436 ( \9689 , \9684 , \9688 );
and \U$9437 ( \9690 , \9595 , \9599 );
and \U$9438 ( \9691 , \9599 , \9604 );
and \U$9439 ( \9692 , \9595 , \9604 );
or \U$9440 ( \9693 , \9690 , \9691 , \9692 );
and \U$9441 ( \9694 , \9539 , \9543 );
and \U$9442 ( \9695 , \9543 , \9548 );
and \U$9443 ( \9696 , \9539 , \9548 );
or \U$9444 ( \9697 , \9694 , \9695 , \9696 );
xor \U$9445 ( \9698 , \9693 , \9697 );
and \U$9446 ( \9699 , \9527 , \9531 );
and \U$9447 ( \9700 , \9531 , \9534 );
and \U$9448 ( \9701 , \9527 , \9534 );
or \U$9449 ( \9702 , \9699 , \9700 , \9701 );
xor \U$9450 ( \9703 , \9698 , \9702 );
and \U$9451 ( \9704 , \5923 , \9584 );
and \U$9452 ( \9705 , \9584 , \9589 );
and \U$9453 ( \9706 , \5923 , \9589 );
or \U$9454 ( \9707 , \9704 , \9705 , \9706 );
and \U$9455 ( \9708 , \9624 , \9628 );
and \U$9456 ( \9709 , \9628 , \9633 );
and \U$9457 ( \9710 , \9624 , \9633 );
or \U$9458 ( \9711 , \9708 , \9709 , \9710 );
xor \U$9459 ( \9712 , \9707 , \9711 );
and \U$9460 ( \9713 , \9609 , \9613 );
and \U$9461 ( \9714 , \9613 , \9618 );
and \U$9462 ( \9715 , \9609 , \9618 );
or \U$9463 ( \9716 , \9713 , \9714 , \9715 );
xor \U$9464 ( \9717 , \9712 , \9716 );
xor \U$9465 ( \9718 , \9703 , \9717 );
and \U$9466 ( \9719 , \9605 , \9619 );
and \U$9467 ( \9720 , \9619 , \9634 );
and \U$9468 ( \9721 , \9605 , \9634 );
or \U$9469 ( \9722 , \9719 , \9720 , \9721 );
and \U$9470 ( \9723 , \5873 , \7192 );
and \U$9471 ( \9724 , \5842 , \7190 );
nor \U$9472 ( \9725 , \9723 , \9724 );
xnor \U$9473 ( \9726 , \9725 , \7198 );
and \U$9474 ( \9727 , \5893 , \7203 );
and \U$9475 ( \9728 , \5861 , \7201 );
nor \U$9476 ( \9729 , \9727 , \9728 );
xnor \U$9477 ( \9730 , \9729 , \6824 );
xor \U$9478 ( \9731 , \9726 , \9730 );
and \U$9479 ( \9732 , \5918 , \5750 );
and \U$9480 ( \9733 , \5881 , \5748 );
nor \U$9481 ( \9734 , \9732 , \9733 );
xnor \U$9482 ( \9735 , \9734 , \5755 );
xor \U$9483 ( \9736 , \9731 , \9735 );
and \U$9484 ( \9737 , \5811 , \7140 );
and \U$9485 ( \9738 , \5780 , \7138 );
nor \U$9486 ( \9739 , \9737 , \9738 );
xnor \U$9487 ( \9740 , \9739 , \7146 );
and \U$9488 ( \9741 , \5831 , \7157 );
and \U$9489 ( \9742 , \5799 , \7155 );
nor \U$9490 ( \9743 , \9741 , \9742 );
xnor \U$9491 ( \9744 , \9743 , \7163 );
xor \U$9492 ( \9745 , \9740 , \9744 );
and \U$9493 ( \9746 , \5854 , \7175 );
and \U$9494 ( \9747 , \5819 , \7173 );
nor \U$9495 ( \9748 , \9746 , \9747 );
xnor \U$9496 ( \9749 , \9748 , \7181 );
xor \U$9497 ( \9750 , \9745 , \9749 );
xor \U$9498 ( \9751 , \9736 , \9750 );
not \U$9499 ( \9752 , \7088 );
and \U$9500 ( \9753 , \5770 , \7099 );
and \U$9501 ( \9754 , \5737 , \7097 );
nor \U$9502 ( \9755 , \9753 , \9754 );
xnor \U$9503 ( \9756 , \9755 , \7105 );
xor \U$9504 ( \9757 , \9752 , \9756 );
and \U$9505 ( \9758 , \5792 , \7117 );
and \U$9506 ( \9759 , \5758 , \7115 );
nor \U$9507 ( \9760 , \9758 , \9759 );
xnor \U$9508 ( \9761 , \9760 , \7123 );
xor \U$9509 ( \9762 , \9757 , \9761 );
xor \U$9510 ( \9763 , \9751 , \9762 );
xor \U$9511 ( \9764 , \9722 , \9763 );
and \U$9512 ( \9765 , \6057 , \5891 );
and \U$9513 ( \9766 , \6029 , \5889 );
nor \U$9514 ( \9767 , \9765 , \9766 );
xnor \U$9515 ( \9768 , \9767 , \5898 );
and \U$9516 ( \9769 , \6065 , \5916 );
and \U$9517 ( \9770 , \6048 , \5914 );
nor \U$9518 ( \9771 , \9769 , \9770 );
xnor \U$9519 ( \9772 , \9771 , \5923 );
xor \U$9520 ( \9773 , \9768 , \9772 );
and \U$9521 ( \9774 , \5998 , \5829 );
and \U$9522 ( \9775 , \5967 , \5827 );
nor \U$9523 ( \9776 , \9774 , \9775 );
xnor \U$9524 ( \9777 , \9776 , \5836 );
and \U$9525 ( \9778 , \6018 , \5852 );
and \U$9526 ( \9779 , \5986 , \5850 );
nor \U$9527 ( \9780 , \9778 , \9779 );
xnor \U$9528 ( \9781 , \9780 , \5859 );
xor \U$9529 ( \9782 , \9777 , \9781 );
and \U$9530 ( \9783 , \6041 , \5871 );
and \U$9531 ( \9784 , \6006 , \5869 );
nor \U$9532 ( \9785 , \9783 , \9784 );
xnor \U$9533 ( \9786 , \9785 , \5878 );
xor \U$9534 ( \9787 , \9782 , \9786 );
xor \U$9535 ( \9788 , \9773 , \9787 );
and \U$9536 ( \9789 , \5937 , \5768 );
and \U$9537 ( \9790 , \5906 , \5766 );
nor \U$9538 ( \9791 , \9789 , \9790 );
xnor \U$9539 ( \9792 , \9791 , \5775 );
and \U$9540 ( \9793 , \5957 , \5790 );
and \U$9541 ( \9794 , \5925 , \5788 );
nor \U$9542 ( \9795 , \9793 , \9794 );
xnor \U$9543 ( \9796 , \9795 , \5797 );
xor \U$9544 ( \9797 , \9792 , \9796 );
and \U$9545 ( \9798 , \5979 , \5809 );
and \U$9546 ( \9799 , \5945 , \5807 );
nor \U$9547 ( \9800 , \9798 , \9799 );
xnor \U$9548 ( \9801 , \9800 , \5816 );
xor \U$9549 ( \9802 , \9797 , \9801 );
xor \U$9550 ( \9803 , \9788 , \9802 );
xor \U$9551 ( \9804 , \9764 , \9803 );
xor \U$9552 ( \9805 , \9718 , \9804 );
and \U$9553 ( \9806 , \9566 , \9570 );
and \U$9554 ( \9807 , \9570 , \9575 );
and \U$9555 ( \9808 , \9566 , \9575 );
or \U$9556 ( \9809 , \9806 , \9807 , \9808 );
and \U$9557 ( \9810 , \9554 , \9558 );
and \U$9558 ( \9811 , \9558 , \9560 );
and \U$9559 ( \9812 , \9554 , \9560 );
or \U$9560 ( \9813 , \9810 , \9811 , \9812 );
xor \U$9561 ( \9814 , \9809 , \9813 );
or \U$9562 ( \9815 , \9535 , \9549 );
xor \U$9563 ( \9816 , \9814 , \9815 );
xor \U$9564 ( \9817 , \9805 , \9816 );
xor \U$9565 ( \9818 , \9689 , \9817 );
xor \U$9566 ( \9819 , \9680 , \9818 );
and \U$9567 ( \9820 , \9502 , \9513 );
and \U$9568 ( \9821 , \9513 , \9653 );
and \U$9569 ( \9822 , \9502 , \9653 );
or \U$9570 ( \9823 , \9820 , \9821 , \9822 );
nor \U$9571 ( \9824 , \9819 , \9823 );
and \U$9572 ( \9825 , \9684 , \9688 );
and \U$9573 ( \9826 , \9688 , \9817 );
and \U$9574 ( \9827 , \9684 , \9817 );
or \U$9575 ( \9828 , \9825 , \9826 , \9827 );
and \U$9576 ( \9829 , \9809 , \9813 );
and \U$9577 ( \9830 , \9813 , \9815 );
and \U$9578 ( \9831 , \9809 , \9815 );
or \U$9579 ( \9832 , \9829 , \9830 , \9831 );
and \U$9580 ( \9833 , \9722 , \9763 );
and \U$9581 ( \9834 , \9763 , \9803 );
and \U$9582 ( \9835 , \9722 , \9803 );
or \U$9583 ( \9836 , \9833 , \9834 , \9835 );
xor \U$9584 ( \9837 , \9832 , \9836 );
and \U$9585 ( \9838 , \9703 , \9717 );
xor \U$9586 ( \9839 , \9837 , \9838 );
xor \U$9587 ( \9840 , \9828 , \9839 );
and \U$9588 ( \9841 , \9669 , \9673 );
and \U$9589 ( \9842 , \9673 , \9678 );
and \U$9590 ( \9843 , \9669 , \9678 );
or \U$9591 ( \9844 , \9841 , \9842 , \9843 );
and \U$9592 ( \9845 , \9718 , \9804 );
and \U$9593 ( \9846 , \9804 , \9816 );
and \U$9594 ( \9847 , \9718 , \9816 );
or \U$9595 ( \9848 , \9845 , \9846 , \9847 );
xor \U$9596 ( \9849 , \9844 , \9848 );
and \U$9597 ( \9850 , \6029 , \5891 );
and \U$9598 ( \9851 , \6041 , \5889 );
nor \U$9599 ( \9852 , \9850 , \9851 );
xnor \U$9600 ( \9853 , \9852 , \5898 );
and \U$9601 ( \9854 , \6048 , \5916 );
and \U$9602 ( \9855 , \6057 , \5914 );
nor \U$9603 ( \9856 , \9854 , \9855 );
xnor \U$9604 ( \9857 , \9856 , \5923 );
xor \U$9605 ( \9858 , \9853 , \9857 );
nand \U$9606 ( \9859 , \6065 , \5933 );
xnor \U$9607 ( \9860 , \9859 , \5942 );
xor \U$9608 ( \9861 , \9858 , \9860 );
and \U$9609 ( \9862 , \5967 , \5829 );
and \U$9610 ( \9863 , \5979 , \5827 );
nor \U$9611 ( \9864 , \9862 , \9863 );
xnor \U$9612 ( \9865 , \9864 , \5836 );
and \U$9613 ( \9866 , \5986 , \5852 );
and \U$9614 ( \9867 , \5998 , \5850 );
nor \U$9615 ( \9868 , \9866 , \9867 );
xnor \U$9616 ( \9869 , \9868 , \5859 );
xor \U$9617 ( \9870 , \9865 , \9869 );
and \U$9618 ( \9871 , \6006 , \5871 );
and \U$9619 ( \9872 , \6018 , \5869 );
nor \U$9620 ( \9873 , \9871 , \9872 );
xnor \U$9621 ( \9874 , \9873 , \5878 );
xor \U$9622 ( \9875 , \9870 , \9874 );
xnor \U$9623 ( \9876 , \9861 , \9875 );
and \U$9624 ( \9877 , \9792 , \9796 );
and \U$9625 ( \9878 , \9796 , \9801 );
and \U$9626 ( \9879 , \9792 , \9801 );
or \U$9627 ( \9880 , \9877 , \9878 , \9879 );
and \U$9628 ( \9881 , \9777 , \9781 );
and \U$9629 ( \9882 , \9781 , \9786 );
and \U$9630 ( \9883 , \9777 , \9786 );
or \U$9631 ( \9884 , \9881 , \9882 , \9883 );
xor \U$9632 ( \9885 , \9880 , \9884 );
and \U$9633 ( \9886 , \9768 , \9772 );
xor \U$9634 ( \9887 , \9885 , \9886 );
xor \U$9635 ( \9888 , \9876 , \9887 );
and \U$9636 ( \9889 , \9752 , \9756 );
and \U$9637 ( \9890 , \9756 , \9761 );
and \U$9638 ( \9891 , \9752 , \9761 );
or \U$9639 ( \9892 , \9889 , \9890 , \9891 );
and \U$9640 ( \9893 , \9740 , \9744 );
and \U$9641 ( \9894 , \9744 , \9749 );
and \U$9642 ( \9895 , \9740 , \9749 );
or \U$9643 ( \9896 , \9893 , \9894 , \9895 );
xor \U$9644 ( \9897 , \9892 , \9896 );
and \U$9645 ( \9898 , \9726 , \9730 );
and \U$9646 ( \9899 , \9730 , \9735 );
and \U$9647 ( \9900 , \9726 , \9735 );
or \U$9648 ( \9901 , \9898 , \9899 , \9900 );
xor \U$9649 ( \9902 , \9897 , \9901 );
xor \U$9650 ( \9903 , \9888 , \9902 );
and \U$9651 ( \9904 , \9736 , \9750 );
and \U$9652 ( \9905 , \9750 , \9762 );
and \U$9653 ( \9906 , \9736 , \9762 );
or \U$9654 ( \9907 , \9904 , \9905 , \9906 );
and \U$9655 ( \9908 , \5737 , \7099 );
not \U$9656 ( \9909 , \9908 );
xnor \U$9657 ( \9910 , \9909 , \7105 );
xor \U$9658 ( \9911 , \5942 , \9910 );
and \U$9659 ( \9912 , \5758 , \7117 );
and \U$9660 ( \9913 , \5770 , \7115 );
nor \U$9661 ( \9914 , \9912 , \9913 );
xnor \U$9662 ( \9915 , \9914 , \7123 );
xor \U$9663 ( \9916 , \9911 , \9915 );
xor \U$9664 ( \9917 , \9907 , \9916 );
and \U$9665 ( \9918 , \5906 , \5768 );
and \U$9666 ( \9919 , \5918 , \5766 );
nor \U$9667 ( \9920 , \9918 , \9919 );
xnor \U$9668 ( \9921 , \9920 , \5775 );
and \U$9669 ( \9922 , \5925 , \5790 );
and \U$9670 ( \9923 , \5937 , \5788 );
nor \U$9671 ( \9924 , \9922 , \9923 );
xnor \U$9672 ( \9925 , \9924 , \5797 );
xor \U$9673 ( \9926 , \9921 , \9925 );
and \U$9674 ( \9927 , \5945 , \5809 );
and \U$9675 ( \9928 , \5957 , \5807 );
nor \U$9676 ( \9929 , \9927 , \9928 );
xnor \U$9677 ( \9930 , \9929 , \5816 );
xor \U$9678 ( \9931 , \9926 , \9930 );
and \U$9679 ( \9932 , \5842 , \7192 );
and \U$9680 ( \9933 , \5854 , \7190 );
nor \U$9681 ( \9934 , \9932 , \9933 );
xnor \U$9682 ( \9935 , \9934 , \7198 );
and \U$9683 ( \9936 , \5861 , \7203 );
and \U$9684 ( \9937 , \5873 , \7201 );
nor \U$9685 ( \9938 , \9936 , \9937 );
xnor \U$9686 ( \9939 , \9938 , \6824 );
xor \U$9687 ( \9940 , \9935 , \9939 );
and \U$9688 ( \9941 , \5881 , \5750 );
and \U$9689 ( \9942 , \5893 , \5748 );
nor \U$9690 ( \9943 , \9941 , \9942 );
xnor \U$9691 ( \9944 , \9943 , \5755 );
xor \U$9692 ( \9945 , \9940 , \9944 );
xor \U$9693 ( \9946 , \9931 , \9945 );
and \U$9694 ( \9947 , \5780 , \7140 );
and \U$9695 ( \9948 , \5792 , \7138 );
nor \U$9696 ( \9949 , \9947 , \9948 );
xnor \U$9697 ( \9950 , \9949 , \7146 );
and \U$9698 ( \9951 , \5799 , \7157 );
and \U$9699 ( \9952 , \5811 , \7155 );
nor \U$9700 ( \9953 , \9951 , \9952 );
xnor \U$9701 ( \9954 , \9953 , \7163 );
xor \U$9702 ( \9955 , \9950 , \9954 );
and \U$9703 ( \9956 , \5819 , \7175 );
and \U$9704 ( \9957 , \5831 , \7173 );
nor \U$9705 ( \9958 , \9956 , \9957 );
xnor \U$9706 ( \9959 , \9958 , \7181 );
xor \U$9707 ( \9960 , \9955 , \9959 );
xor \U$9708 ( \9961 , \9946 , \9960 );
xor \U$9709 ( \9962 , \9917 , \9961 );
xor \U$9710 ( \9963 , \9903 , \9962 );
and \U$9711 ( \9964 , \9707 , \9711 );
and \U$9712 ( \9965 , \9711 , \9716 );
and \U$9713 ( \9966 , \9707 , \9716 );
or \U$9714 ( \9967 , \9964 , \9965 , \9966 );
and \U$9715 ( \9968 , \9693 , \9697 );
and \U$9716 ( \9969 , \9697 , \9702 );
and \U$9717 ( \9970 , \9693 , \9702 );
or \U$9718 ( \9971 , \9968 , \9969 , \9970 );
xor \U$9719 ( \9972 , \9967 , \9971 );
and \U$9720 ( \9973 , \9773 , \9787 );
and \U$9721 ( \9974 , \9787 , \9802 );
and \U$9722 ( \9975 , \9773 , \9802 );
or \U$9723 ( \9976 , \9973 , \9974 , \9975 );
xor \U$9724 ( \9977 , \9972 , \9976 );
xor \U$9725 ( \9978 , \9963 , \9977 );
xor \U$9726 ( \9979 , \9849 , \9978 );
xor \U$9727 ( \9980 , \9840 , \9979 );
and \U$9728 ( \9981 , \9665 , \9679 );
and \U$9729 ( \9982 , \9679 , \9818 );
and \U$9730 ( \9983 , \9665 , \9818 );
or \U$9731 ( \9984 , \9981 , \9982 , \9983 );
nor \U$9732 ( \9985 , \9980 , \9984 );
nor \U$9733 ( \9986 , \9824 , \9985 );
and \U$9734 ( \9987 , \9844 , \9848 );
and \U$9735 ( \9988 , \9848 , \9978 );
and \U$9736 ( \9989 , \9844 , \9978 );
or \U$9737 ( \9990 , \9987 , \9988 , \9989 );
and \U$9738 ( \9991 , \9967 , \9971 );
and \U$9739 ( \9992 , \9971 , \9976 );
and \U$9740 ( \9993 , \9967 , \9976 );
or \U$9741 ( \9994 , \9991 , \9992 , \9993 );
and \U$9742 ( \9995 , \9907 , \9916 );
and \U$9743 ( \9996 , \9916 , \9961 );
and \U$9744 ( \9997 , \9907 , \9961 );
or \U$9745 ( \9998 , \9995 , \9996 , \9997 );
xor \U$9746 ( \9999 , \9994 , \9998 );
and \U$9747 ( \10000 , \9876 , \9887 );
and \U$9748 ( \10001 , \9887 , \9902 );
and \U$9749 ( \10002 , \9876 , \9902 );
or \U$9750 ( \10003 , \10000 , \10001 , \10002 );
xor \U$9751 ( \10004 , \9999 , \10003 );
xor \U$9752 ( \10005 , \9990 , \10004 );
and \U$9753 ( \10006 , \9832 , \9836 );
and \U$9754 ( \10007 , \9836 , \9838 );
and \U$9755 ( \10008 , \9832 , \9838 );
or \U$9756 ( \10009 , \10006 , \10007 , \10008 );
and \U$9757 ( \10010 , \9903 , \9962 );
and \U$9758 ( \10011 , \9962 , \9977 );
and \U$9759 ( \10012 , \9903 , \9977 );
or \U$9760 ( \10013 , \10010 , \10011 , \10012 );
xor \U$9761 ( \10014 , \10009 , \10013 );
and \U$9762 ( \10015 , \9921 , \9925 );
and \U$9763 ( \10016 , \9925 , \9930 );
and \U$9764 ( \10017 , \9921 , \9930 );
or \U$9765 ( \10018 , \10015 , \10016 , \10017 );
and \U$9766 ( \10019 , \9865 , \9869 );
and \U$9767 ( \10020 , \9869 , \9874 );
and \U$9768 ( \10021 , \9865 , \9874 );
or \U$9769 ( \10022 , \10019 , \10020 , \10021 );
xor \U$9770 ( \10023 , \10018 , \10022 );
and \U$9771 ( \10024 , \9853 , \9857 );
and \U$9772 ( \10025 , \9857 , \9860 );
and \U$9773 ( \10026 , \9853 , \9860 );
or \U$9774 ( \10027 , \10024 , \10025 , \10026 );
xor \U$9775 ( \10028 , \10023 , \10027 );
and \U$9776 ( \10029 , \5942 , \9910 );
and \U$9777 ( \10030 , \9910 , \9915 );
and \U$9778 ( \10031 , \5942 , \9915 );
or \U$9779 ( \10032 , \10029 , \10030 , \10031 );
and \U$9780 ( \10033 , \9950 , \9954 );
and \U$9781 ( \10034 , \9954 , \9959 );
and \U$9782 ( \10035 , \9950 , \9959 );
or \U$9783 ( \10036 , \10033 , \10034 , \10035 );
xor \U$9784 ( \10037 , \10032 , \10036 );
and \U$9785 ( \10038 , \9935 , \9939 );
and \U$9786 ( \10039 , \9939 , \9944 );
and \U$9787 ( \10040 , \9935 , \9944 );
or \U$9788 ( \10041 , \10038 , \10039 , \10040 );
xor \U$9789 ( \10042 , \10037 , \10041 );
xor \U$9790 ( \10043 , \10028 , \10042 );
and \U$9791 ( \10044 , \9931 , \9945 );
and \U$9792 ( \10045 , \9945 , \9960 );
and \U$9793 ( \10046 , \9931 , \9960 );
or \U$9794 ( \10047 , \10044 , \10045 , \10046 );
and \U$9795 ( \10048 , \5873 , \7203 );
and \U$9796 ( \10049 , \5842 , \7201 );
nor \U$9797 ( \10050 , \10048 , \10049 );
xnor \U$9798 ( \10051 , \10050 , \6824 );
and \U$9799 ( \10052 , \5893 , \5750 );
and \U$9800 ( \10053 , \5861 , \5748 );
nor \U$9801 ( \10054 , \10052 , \10053 );
xnor \U$9802 ( \10055 , \10054 , \5755 );
xor \U$9803 ( \10056 , \10051 , \10055 );
and \U$9804 ( \10057 , \5918 , \5768 );
and \U$9805 ( \10058 , \5881 , \5766 );
nor \U$9806 ( \10059 , \10057 , \10058 );
xnor \U$9807 ( \10060 , \10059 , \5775 );
xor \U$9808 ( \10061 , \10056 , \10060 );
and \U$9809 ( \10062 , \5811 , \7157 );
and \U$9810 ( \10063 , \5780 , \7155 );
nor \U$9811 ( \10064 , \10062 , \10063 );
xnor \U$9812 ( \10065 , \10064 , \7163 );
and \U$9813 ( \10066 , \5831 , \7175 );
and \U$9814 ( \10067 , \5799 , \7173 );
nor \U$9815 ( \10068 , \10066 , \10067 );
xnor \U$9816 ( \10069 , \10068 , \7181 );
xor \U$9817 ( \10070 , \10065 , \10069 );
and \U$9818 ( \10071 , \5854 , \7192 );
and \U$9819 ( \10072 , \5819 , \7190 );
nor \U$9820 ( \10073 , \10071 , \10072 );
xnor \U$9821 ( \10074 , \10073 , \7198 );
xor \U$9822 ( \10075 , \10070 , \10074 );
xor \U$9823 ( \10076 , \10061 , \10075 );
not \U$9824 ( \10077 , \7105 );
and \U$9825 ( \10078 , \5770 , \7117 );
and \U$9826 ( \10079 , \5737 , \7115 );
nor \U$9827 ( \10080 , \10078 , \10079 );
xnor \U$9828 ( \10081 , \10080 , \7123 );
xor \U$9829 ( \10082 , \10077 , \10081 );
and \U$9830 ( \10083 , \5792 , \7140 );
and \U$9831 ( \10084 , \5758 , \7138 );
nor \U$9832 ( \10085 , \10083 , \10084 );
xnor \U$9833 ( \10086 , \10085 , \7146 );
xor \U$9834 ( \10087 , \10082 , \10086 );
xor \U$9835 ( \10088 , \10076 , \10087 );
xor \U$9836 ( \10089 , \10047 , \10088 );
and \U$9837 ( \10090 , \6057 , \5916 );
and \U$9838 ( \10091 , \6029 , \5914 );
nor \U$9839 ( \10092 , \10090 , \10091 );
xnor \U$9840 ( \10093 , \10092 , \5923 );
and \U$9841 ( \10094 , \6065 , \5935 );
and \U$9842 ( \10095 , \6048 , \5933 );
nor \U$9843 ( \10096 , \10094 , \10095 );
xnor \U$9844 ( \10097 , \10096 , \5942 );
xor \U$9845 ( \10098 , \10093 , \10097 );
and \U$9846 ( \10099 , \5998 , \5852 );
and \U$9847 ( \10100 , \5967 , \5850 );
nor \U$9848 ( \10101 , \10099 , \10100 );
xnor \U$9849 ( \10102 , \10101 , \5859 );
and \U$9850 ( \10103 , \6018 , \5871 );
and \U$9851 ( \10104 , \5986 , \5869 );
nor \U$9852 ( \10105 , \10103 , \10104 );
xnor \U$9853 ( \10106 , \10105 , \5878 );
xor \U$9854 ( \10107 , \10102 , \10106 );
and \U$9855 ( \10108 , \6041 , \5891 );
and \U$9856 ( \10109 , \6006 , \5889 );
nor \U$9857 ( \10110 , \10108 , \10109 );
xnor \U$9858 ( \10111 , \10110 , \5898 );
xor \U$9859 ( \10112 , \10107 , \10111 );
xor \U$9860 ( \10113 , \10098 , \10112 );
and \U$9861 ( \10114 , \5937 , \5790 );
and \U$9862 ( \10115 , \5906 , \5788 );
nor \U$9863 ( \10116 , \10114 , \10115 );
xnor \U$9864 ( \10117 , \10116 , \5797 );
and \U$9865 ( \10118 , \5957 , \5809 );
and \U$9866 ( \10119 , \5925 , \5807 );
nor \U$9867 ( \10120 , \10118 , \10119 );
xnor \U$9868 ( \10121 , \10120 , \5816 );
xor \U$9869 ( \10122 , \10117 , \10121 );
and \U$9870 ( \10123 , \5979 , \5829 );
and \U$9871 ( \10124 , \5945 , \5827 );
nor \U$9872 ( \10125 , \10123 , \10124 );
xnor \U$9873 ( \10126 , \10125 , \5836 );
xor \U$9874 ( \10127 , \10122 , \10126 );
xor \U$9875 ( \10128 , \10113 , \10127 );
xor \U$9876 ( \10129 , \10089 , \10128 );
xor \U$9877 ( \10130 , \10043 , \10129 );
and \U$9878 ( \10131 , \9892 , \9896 );
and \U$9879 ( \10132 , \9896 , \9901 );
and \U$9880 ( \10133 , \9892 , \9901 );
or \U$9881 ( \10134 , \10131 , \10132 , \10133 );
and \U$9882 ( \10135 , \9880 , \9884 );
and \U$9883 ( \10136 , \9884 , \9886 );
and \U$9884 ( \10137 , \9880 , \9886 );
or \U$9885 ( \10138 , \10135 , \10136 , \10137 );
xor \U$9886 ( \10139 , \10134 , \10138 );
or \U$9887 ( \10140 , \9861 , \9875 );
xor \U$9888 ( \10141 , \10139 , \10140 );
xor \U$9889 ( \10142 , \10130 , \10141 );
xor \U$9890 ( \10143 , \10014 , \10142 );
xor \U$9891 ( \10144 , \10005 , \10143 );
and \U$9892 ( \10145 , \9828 , \9839 );
and \U$9893 ( \10146 , \9839 , \9979 );
and \U$9894 ( \10147 , \9828 , \9979 );
or \U$9895 ( \10148 , \10145 , \10146 , \10147 );
nor \U$9896 ( \10149 , \10144 , \10148 );
and \U$9897 ( \10150 , \10009 , \10013 );
and \U$9898 ( \10151 , \10013 , \10142 );
and \U$9899 ( \10152 , \10009 , \10142 );
or \U$9900 ( \10153 , \10150 , \10151 , \10152 );
and \U$9901 ( \10154 , \10134 , \10138 );
and \U$9902 ( \10155 , \10138 , \10140 );
and \U$9903 ( \10156 , \10134 , \10140 );
or \U$9904 ( \10157 , \10154 , \10155 , \10156 );
and \U$9905 ( \10158 , \10047 , \10088 );
and \U$9906 ( \10159 , \10088 , \10128 );
and \U$9907 ( \10160 , \10047 , \10128 );
or \U$9908 ( \10161 , \10158 , \10159 , \10160 );
xor \U$9909 ( \10162 , \10157 , \10161 );
and \U$9910 ( \10163 , \10028 , \10042 );
xor \U$9911 ( \10164 , \10162 , \10163 );
xor \U$9912 ( \10165 , \10153 , \10164 );
and \U$9913 ( \10166 , \9994 , \9998 );
and \U$9914 ( \10167 , \9998 , \10003 );
and \U$9915 ( \10168 , \9994 , \10003 );
or \U$9916 ( \10169 , \10166 , \10167 , \10168 );
and \U$9917 ( \10170 , \10043 , \10129 );
and \U$9918 ( \10171 , \10129 , \10141 );
and \U$9919 ( \10172 , \10043 , \10141 );
or \U$9920 ( \10173 , \10170 , \10171 , \10172 );
xor \U$9921 ( \10174 , \10169 , \10173 );
and \U$9922 ( \10175 , \6029 , \5916 );
and \U$9923 ( \10176 , \6041 , \5914 );
nor \U$9924 ( \10177 , \10175 , \10176 );
xnor \U$9925 ( \10178 , \10177 , \5923 );
and \U$9926 ( \10179 , \6048 , \5935 );
and \U$9927 ( \10180 , \6057 , \5933 );
nor \U$9928 ( \10181 , \10179 , \10180 );
xnor \U$9929 ( \10182 , \10181 , \5942 );
xor \U$9930 ( \10183 , \10178 , \10182 );
nand \U$9931 ( \10184 , \6065 , \5953 );
xnor \U$9932 ( \10185 , \10184 , \5962 );
xor \U$9933 ( \10186 , \10183 , \10185 );
and \U$9934 ( \10187 , \5967 , \5852 );
and \U$9935 ( \10188 , \5979 , \5850 );
nor \U$9936 ( \10189 , \10187 , \10188 );
xnor \U$9937 ( \10190 , \10189 , \5859 );
and \U$9938 ( \10191 , \5986 , \5871 );
and \U$9939 ( \10192 , \5998 , \5869 );
nor \U$9940 ( \10193 , \10191 , \10192 );
xnor \U$9941 ( \10194 , \10193 , \5878 );
xor \U$9942 ( \10195 , \10190 , \10194 );
and \U$9943 ( \10196 , \6006 , \5891 );
and \U$9944 ( \10197 , \6018 , \5889 );
nor \U$9945 ( \10198 , \10196 , \10197 );
xnor \U$9946 ( \10199 , \10198 , \5898 );
xor \U$9947 ( \10200 , \10195 , \10199 );
xnor \U$9948 ( \10201 , \10186 , \10200 );
and \U$9949 ( \10202 , \10117 , \10121 );
and \U$9950 ( \10203 , \10121 , \10126 );
and \U$9951 ( \10204 , \10117 , \10126 );
or \U$9952 ( \10205 , \10202 , \10203 , \10204 );
and \U$9953 ( \10206 , \10102 , \10106 );
and \U$9954 ( \10207 , \10106 , \10111 );
and \U$9955 ( \10208 , \10102 , \10111 );
or \U$9956 ( \10209 , \10206 , \10207 , \10208 );
xor \U$9957 ( \10210 , \10205 , \10209 );
and \U$9958 ( \10211 , \10093 , \10097 );
xor \U$9959 ( \10212 , \10210 , \10211 );
xor \U$9960 ( \10213 , \10201 , \10212 );
and \U$9961 ( \10214 , \10077 , \10081 );
and \U$9962 ( \10215 , \10081 , \10086 );
and \U$9963 ( \10216 , \10077 , \10086 );
or \U$9964 ( \10217 , \10214 , \10215 , \10216 );
and \U$9965 ( \10218 , \10065 , \10069 );
and \U$9966 ( \10219 , \10069 , \10074 );
and \U$9967 ( \10220 , \10065 , \10074 );
or \U$9968 ( \10221 , \10218 , \10219 , \10220 );
xor \U$9969 ( \10222 , \10217 , \10221 );
and \U$9970 ( \10223 , \10051 , \10055 );
and \U$9971 ( \10224 , \10055 , \10060 );
and \U$9972 ( \10225 , \10051 , \10060 );
or \U$9973 ( \10226 , \10223 , \10224 , \10225 );
xor \U$9974 ( \10227 , \10222 , \10226 );
xor \U$9975 ( \10228 , \10213 , \10227 );
and \U$9976 ( \10229 , \10061 , \10075 );
and \U$9977 ( \10230 , \10075 , \10087 );
and \U$9978 ( \10231 , \10061 , \10087 );
or \U$9979 ( \10232 , \10229 , \10230 , \10231 );
and \U$9980 ( \10233 , \5737 , \7117 );
not \U$9981 ( \10234 , \10233 );
xnor \U$9982 ( \10235 , \10234 , \7123 );
xor \U$9983 ( \10236 , \5962 , \10235 );
and \U$9984 ( \10237 , \5758 , \7140 );
and \U$9985 ( \10238 , \5770 , \7138 );
nor \U$9986 ( \10239 , \10237 , \10238 );
xnor \U$9987 ( \10240 , \10239 , \7146 );
xor \U$9988 ( \10241 , \10236 , \10240 );
xor \U$9989 ( \10242 , \10232 , \10241 );
and \U$9990 ( \10243 , \5906 , \5790 );
and \U$9991 ( \10244 , \5918 , \5788 );
nor \U$9992 ( \10245 , \10243 , \10244 );
xnor \U$9993 ( \10246 , \10245 , \5797 );
and \U$9994 ( \10247 , \5925 , \5809 );
and \U$9995 ( \10248 , \5937 , \5807 );
nor \U$9996 ( \10249 , \10247 , \10248 );
xnor \U$9997 ( \10250 , \10249 , \5816 );
xor \U$9998 ( \10251 , \10246 , \10250 );
and \U$9999 ( \10252 , \5945 , \5829 );
and \U$10000 ( \10253 , \5957 , \5827 );
nor \U$10001 ( \10254 , \10252 , \10253 );
xnor \U$10002 ( \10255 , \10254 , \5836 );
xor \U$10003 ( \10256 , \10251 , \10255 );
and \U$10004 ( \10257 , \5842 , \7203 );
and \U$10005 ( \10258 , \5854 , \7201 );
nor \U$10006 ( \10259 , \10257 , \10258 );
xnor \U$10007 ( \10260 , \10259 , \6824 );
and \U$10008 ( \10261 , \5861 , \5750 );
and \U$10009 ( \10262 , \5873 , \5748 );
nor \U$10010 ( \10263 , \10261 , \10262 );
xnor \U$10011 ( \10264 , \10263 , \5755 );
xor \U$10012 ( \10265 , \10260 , \10264 );
and \U$10013 ( \10266 , \5881 , \5768 );
and \U$10014 ( \10267 , \5893 , \5766 );
nor \U$10015 ( \10268 , \10266 , \10267 );
xnor \U$10016 ( \10269 , \10268 , \5775 );
xor \U$10017 ( \10270 , \10265 , \10269 );
xor \U$10018 ( \10271 , \10256 , \10270 );
and \U$10019 ( \10272 , \5780 , \7157 );
and \U$10020 ( \10273 , \5792 , \7155 );
nor \U$10021 ( \10274 , \10272 , \10273 );
xnor \U$10022 ( \10275 , \10274 , \7163 );
and \U$10023 ( \10276 , \5799 , \7175 );
and \U$10024 ( \10277 , \5811 , \7173 );
nor \U$10025 ( \10278 , \10276 , \10277 );
xnor \U$10026 ( \10279 , \10278 , \7181 );
xor \U$10027 ( \10280 , \10275 , \10279 );
and \U$10028 ( \10281 , \5819 , \7192 );
and \U$10029 ( \10282 , \5831 , \7190 );
nor \U$10030 ( \10283 , \10281 , \10282 );
xnor \U$10031 ( \10284 , \10283 , \7198 );
xor \U$10032 ( \10285 , \10280 , \10284 );
xor \U$10033 ( \10286 , \10271 , \10285 );
xor \U$10034 ( \10287 , \10242 , \10286 );
xor \U$10035 ( \10288 , \10228 , \10287 );
and \U$10036 ( \10289 , \10032 , \10036 );
and \U$10037 ( \10290 , \10036 , \10041 );
and \U$10038 ( \10291 , \10032 , \10041 );
or \U$10039 ( \10292 , \10289 , \10290 , \10291 );
and \U$10040 ( \10293 , \10018 , \10022 );
and \U$10041 ( \10294 , \10022 , \10027 );
and \U$10042 ( \10295 , \10018 , \10027 );
or \U$10043 ( \10296 , \10293 , \10294 , \10295 );
xor \U$10044 ( \10297 , \10292 , \10296 );
and \U$10045 ( \10298 , \10098 , \10112 );
and \U$10046 ( \10299 , \10112 , \10127 );
and \U$10047 ( \10300 , \10098 , \10127 );
or \U$10048 ( \10301 , \10298 , \10299 , \10300 );
xor \U$10049 ( \10302 , \10297 , \10301 );
xor \U$10050 ( \10303 , \10288 , \10302 );
xor \U$10051 ( \10304 , \10174 , \10303 );
xor \U$10052 ( \10305 , \10165 , \10304 );
and \U$10053 ( \10306 , \9990 , \10004 );
and \U$10054 ( \10307 , \10004 , \10143 );
and \U$10055 ( \10308 , \9990 , \10143 );
or \U$10056 ( \10309 , \10306 , \10307 , \10308 );
nor \U$10057 ( \10310 , \10305 , \10309 );
nor \U$10058 ( \10311 , \10149 , \10310 );
nand \U$10059 ( \10312 , \9986 , \10311 );
nor \U$10060 ( \10313 , \9661 , \10312 );
nand \U$10061 ( \10314 , \9010 , \10313 );
and \U$10062 ( \10315 , \10169 , \10173 );
and \U$10063 ( \10316 , \10173 , \10303 );
and \U$10064 ( \10317 , \10169 , \10303 );
or \U$10065 ( \10318 , \10315 , \10316 , \10317 );
and \U$10066 ( \10319 , \10292 , \10296 );
and \U$10067 ( \10320 , \10296 , \10301 );
and \U$10068 ( \10321 , \10292 , \10301 );
or \U$10069 ( \10322 , \10319 , \10320 , \10321 );
and \U$10070 ( \10323 , \10232 , \10241 );
and \U$10071 ( \10324 , \10241 , \10286 );
and \U$10072 ( \10325 , \10232 , \10286 );
or \U$10073 ( \10326 , \10323 , \10324 , \10325 );
xor \U$10074 ( \10327 , \10322 , \10326 );
and \U$10075 ( \10328 , \10201 , \10212 );
and \U$10076 ( \10329 , \10212 , \10227 );
and \U$10077 ( \10330 , \10201 , \10227 );
or \U$10078 ( \10331 , \10328 , \10329 , \10330 );
xor \U$10079 ( \10332 , \10327 , \10331 );
xor \U$10080 ( \10333 , \10318 , \10332 );
and \U$10081 ( \10334 , \10157 , \10161 );
and \U$10082 ( \10335 , \10161 , \10163 );
and \U$10083 ( \10336 , \10157 , \10163 );
or \U$10084 ( \10337 , \10334 , \10335 , \10336 );
and \U$10085 ( \10338 , \10228 , \10287 );
and \U$10086 ( \10339 , \10287 , \10302 );
and \U$10087 ( \10340 , \10228 , \10302 );
or \U$10088 ( \10341 , \10338 , \10339 , \10340 );
xor \U$10089 ( \10342 , \10337 , \10341 );
and \U$10090 ( \10343 , \10246 , \10250 );
and \U$10091 ( \10344 , \10250 , \10255 );
and \U$10092 ( \10345 , \10246 , \10255 );
or \U$10093 ( \10346 , \10343 , \10344 , \10345 );
and \U$10094 ( \10347 , \10190 , \10194 );
and \U$10095 ( \10348 , \10194 , \10199 );
and \U$10096 ( \10349 , \10190 , \10199 );
or \U$10097 ( \10350 , \10347 , \10348 , \10349 );
xor \U$10098 ( \10351 , \10346 , \10350 );
and \U$10099 ( \10352 , \10178 , \10182 );
and \U$10100 ( \10353 , \10182 , \10185 );
and \U$10101 ( \10354 , \10178 , \10185 );
or \U$10102 ( \10355 , \10352 , \10353 , \10354 );
xor \U$10103 ( \10356 , \10351 , \10355 );
and \U$10104 ( \10357 , \5962 , \10235 );
and \U$10105 ( \10358 , \10235 , \10240 );
and \U$10106 ( \10359 , \5962 , \10240 );
or \U$10107 ( \10360 , \10357 , \10358 , \10359 );
and \U$10108 ( \10361 , \10275 , \10279 );
and \U$10109 ( \10362 , \10279 , \10284 );
and \U$10110 ( \10363 , \10275 , \10284 );
or \U$10111 ( \10364 , \10361 , \10362 , \10363 );
xor \U$10112 ( \10365 , \10360 , \10364 );
and \U$10113 ( \10366 , \10260 , \10264 );
and \U$10114 ( \10367 , \10264 , \10269 );
and \U$10115 ( \10368 , \10260 , \10269 );
or \U$10116 ( \10369 , \10366 , \10367 , \10368 );
xor \U$10117 ( \10370 , \10365 , \10369 );
xor \U$10118 ( \10371 , \10356 , \10370 );
and \U$10119 ( \10372 , \10256 , \10270 );
and \U$10120 ( \10373 , \10270 , \10285 );
and \U$10121 ( \10374 , \10256 , \10285 );
or \U$10122 ( \10375 , \10372 , \10373 , \10374 );
and \U$10123 ( \10376 , \5873 , \5750 );
and \U$10124 ( \10377 , \5842 , \5748 );
nor \U$10125 ( \10378 , \10376 , \10377 );
xnor \U$10126 ( \10379 , \10378 , \5755 );
and \U$10127 ( \10380 , \5893 , \5768 );
and \U$10128 ( \10381 , \5861 , \5766 );
nor \U$10129 ( \10382 , \10380 , \10381 );
xnor \U$10130 ( \10383 , \10382 , \5775 );
xor \U$10131 ( \10384 , \10379 , \10383 );
and \U$10132 ( \10385 , \5918 , \5790 );
and \U$10133 ( \10386 , \5881 , \5788 );
nor \U$10134 ( \10387 , \10385 , \10386 );
xnor \U$10135 ( \10388 , \10387 , \5797 );
xor \U$10136 ( \10389 , \10384 , \10388 );
and \U$10137 ( \10390 , \5811 , \7175 );
and \U$10138 ( \10391 , \5780 , \7173 );
nor \U$10139 ( \10392 , \10390 , \10391 );
xnor \U$10140 ( \10393 , \10392 , \7181 );
and \U$10141 ( \10394 , \5831 , \7192 );
and \U$10142 ( \10395 , \5799 , \7190 );
nor \U$10143 ( \10396 , \10394 , \10395 );
xnor \U$10144 ( \10397 , \10396 , \7198 );
xor \U$10145 ( \10398 , \10393 , \10397 );
and \U$10146 ( \10399 , \5854 , \7203 );
and \U$10147 ( \10400 , \5819 , \7201 );
nor \U$10148 ( \10401 , \10399 , \10400 );
xnor \U$10149 ( \10402 , \10401 , \6824 );
xor \U$10150 ( \10403 , \10398 , \10402 );
xor \U$10151 ( \10404 , \10389 , \10403 );
not \U$10152 ( \10405 , \7123 );
and \U$10153 ( \10406 , \5770 , \7140 );
and \U$10154 ( \10407 , \5737 , \7138 );
nor \U$10155 ( \10408 , \10406 , \10407 );
xnor \U$10156 ( \10409 , \10408 , \7146 );
xor \U$10157 ( \10410 , \10405 , \10409 );
and \U$10158 ( \10411 , \5792 , \7157 );
and \U$10159 ( \10412 , \5758 , \7155 );
nor \U$10160 ( \10413 , \10411 , \10412 );
xnor \U$10161 ( \10414 , \10413 , \7163 );
xor \U$10162 ( \10415 , \10410 , \10414 );
xor \U$10163 ( \10416 , \10404 , \10415 );
xor \U$10164 ( \10417 , \10375 , \10416 );
and \U$10165 ( \10418 , \6057 , \5935 );
and \U$10166 ( \10419 , \6029 , \5933 );
nor \U$10167 ( \10420 , \10418 , \10419 );
xnor \U$10168 ( \10421 , \10420 , \5942 );
and \U$10169 ( \10422 , \6065 , \5955 );
and \U$10170 ( \10423 , \6048 , \5953 );
nor \U$10171 ( \10424 , \10422 , \10423 );
xnor \U$10172 ( \10425 , \10424 , \5962 );
xor \U$10173 ( \10426 , \10421 , \10425 );
and \U$10174 ( \10427 , \5998 , \5871 );
and \U$10175 ( \10428 , \5967 , \5869 );
nor \U$10176 ( \10429 , \10427 , \10428 );
xnor \U$10177 ( \10430 , \10429 , \5878 );
and \U$10178 ( \10431 , \6018 , \5891 );
and \U$10179 ( \10432 , \5986 , \5889 );
nor \U$10180 ( \10433 , \10431 , \10432 );
xnor \U$10181 ( \10434 , \10433 , \5898 );
xor \U$10182 ( \10435 , \10430 , \10434 );
and \U$10183 ( \10436 , \6041 , \5916 );
and \U$10184 ( \10437 , \6006 , \5914 );
nor \U$10185 ( \10438 , \10436 , \10437 );
xnor \U$10186 ( \10439 , \10438 , \5923 );
xor \U$10187 ( \10440 , \10435 , \10439 );
xor \U$10188 ( \10441 , \10426 , \10440 );
and \U$10189 ( \10442 , \5937 , \5809 );
and \U$10190 ( \10443 , \5906 , \5807 );
nor \U$10191 ( \10444 , \10442 , \10443 );
xnor \U$10192 ( \10445 , \10444 , \5816 );
and \U$10193 ( \10446 , \5957 , \5829 );
and \U$10194 ( \10447 , \5925 , \5827 );
nor \U$10195 ( \10448 , \10446 , \10447 );
xnor \U$10196 ( \10449 , \10448 , \5836 );
xor \U$10197 ( \10450 , \10445 , \10449 );
and \U$10198 ( \10451 , \5979 , \5852 );
and \U$10199 ( \10452 , \5945 , \5850 );
nor \U$10200 ( \10453 , \10451 , \10452 );
xnor \U$10201 ( \10454 , \10453 , \5859 );
xor \U$10202 ( \10455 , \10450 , \10454 );
xor \U$10203 ( \10456 , \10441 , \10455 );
xor \U$10204 ( \10457 , \10417 , \10456 );
xor \U$10205 ( \10458 , \10371 , \10457 );
and \U$10206 ( \10459 , \10217 , \10221 );
and \U$10207 ( \10460 , \10221 , \10226 );
and \U$10208 ( \10461 , \10217 , \10226 );
or \U$10209 ( \10462 , \10459 , \10460 , \10461 );
and \U$10210 ( \10463 , \10205 , \10209 );
and \U$10211 ( \10464 , \10209 , \10211 );
and \U$10212 ( \10465 , \10205 , \10211 );
or \U$10213 ( \10466 , \10463 , \10464 , \10465 );
xor \U$10214 ( \10467 , \10462 , \10466 );
or \U$10215 ( \10468 , \10186 , \10200 );
xor \U$10216 ( \10469 , \10467 , \10468 );
xor \U$10217 ( \10470 , \10458 , \10469 );
xor \U$10218 ( \10471 , \10342 , \10470 );
xor \U$10219 ( \10472 , \10333 , \10471 );
and \U$10220 ( \10473 , \10153 , \10164 );
and \U$10221 ( \10474 , \10164 , \10304 );
and \U$10222 ( \10475 , \10153 , \10304 );
or \U$10223 ( \10476 , \10473 , \10474 , \10475 );
nor \U$10224 ( \10477 , \10472 , \10476 );
and \U$10225 ( \10478 , \10337 , \10341 );
and \U$10226 ( \10479 , \10341 , \10470 );
and \U$10227 ( \10480 , \10337 , \10470 );
or \U$10228 ( \10481 , \10478 , \10479 , \10480 );
and \U$10229 ( \10482 , \10462 , \10466 );
and \U$10230 ( \10483 , \10466 , \10468 );
and \U$10231 ( \10484 , \10462 , \10468 );
or \U$10232 ( \10485 , \10482 , \10483 , \10484 );
and \U$10233 ( \10486 , \10375 , \10416 );
and \U$10234 ( \10487 , \10416 , \10456 );
and \U$10235 ( \10488 , \10375 , \10456 );
or \U$10236 ( \10489 , \10486 , \10487 , \10488 );
xor \U$10237 ( \10490 , \10485 , \10489 );
and \U$10238 ( \10491 , \10356 , \10370 );
xor \U$10239 ( \10492 , \10490 , \10491 );
xor \U$10240 ( \10493 , \10481 , \10492 );
and \U$10241 ( \10494 , \10322 , \10326 );
and \U$10242 ( \10495 , \10326 , \10331 );
and \U$10243 ( \10496 , \10322 , \10331 );
or \U$10244 ( \10497 , \10494 , \10495 , \10496 );
and \U$10245 ( \10498 , \10371 , \10457 );
and \U$10246 ( \10499 , \10457 , \10469 );
and \U$10247 ( \10500 , \10371 , \10469 );
or \U$10248 ( \10501 , \10498 , \10499 , \10500 );
xor \U$10249 ( \10502 , \10497 , \10501 );
and \U$10250 ( \10503 , \6029 , \5935 );
and \U$10251 ( \10504 , \6041 , \5933 );
nor \U$10252 ( \10505 , \10503 , \10504 );
xnor \U$10253 ( \10506 , \10505 , \5942 );
and \U$10254 ( \10507 , \6048 , \5955 );
and \U$10255 ( \10508 , \6057 , \5953 );
nor \U$10256 ( \10509 , \10507 , \10508 );
xnor \U$10257 ( \10510 , \10509 , \5962 );
xor \U$10258 ( \10511 , \10506 , \10510 );
nand \U$10259 ( \10512 , \6065 , \5975 );
xnor \U$10260 ( \10513 , \10512 , \5984 );
xor \U$10261 ( \10514 , \10511 , \10513 );
and \U$10262 ( \10515 , \5967 , \5871 );
and \U$10263 ( \10516 , \5979 , \5869 );
nor \U$10264 ( \10517 , \10515 , \10516 );
xnor \U$10265 ( \10518 , \10517 , \5878 );
and \U$10266 ( \10519 , \5986 , \5891 );
and \U$10267 ( \10520 , \5998 , \5889 );
nor \U$10268 ( \10521 , \10519 , \10520 );
xnor \U$10269 ( \10522 , \10521 , \5898 );
xor \U$10270 ( \10523 , \10518 , \10522 );
and \U$10271 ( \10524 , \6006 , \5916 );
and \U$10272 ( \10525 , \6018 , \5914 );
nor \U$10273 ( \10526 , \10524 , \10525 );
xnor \U$10274 ( \10527 , \10526 , \5923 );
xor \U$10275 ( \10528 , \10523 , \10527 );
xnor \U$10276 ( \10529 , \10514 , \10528 );
and \U$10277 ( \10530 , \10445 , \10449 );
and \U$10278 ( \10531 , \10449 , \10454 );
and \U$10279 ( \10532 , \10445 , \10454 );
or \U$10280 ( \10533 , \10530 , \10531 , \10532 );
and \U$10281 ( \10534 , \10430 , \10434 );
and \U$10282 ( \10535 , \10434 , \10439 );
and \U$10283 ( \10536 , \10430 , \10439 );
or \U$10284 ( \10537 , \10534 , \10535 , \10536 );
xor \U$10285 ( \10538 , \10533 , \10537 );
and \U$10286 ( \10539 , \10421 , \10425 );
xor \U$10287 ( \10540 , \10538 , \10539 );
xor \U$10288 ( \10541 , \10529 , \10540 );
and \U$10289 ( \10542 , \10405 , \10409 );
and \U$10290 ( \10543 , \10409 , \10414 );
and \U$10291 ( \10544 , \10405 , \10414 );
or \U$10292 ( \10545 , \10542 , \10543 , \10544 );
and \U$10293 ( \10546 , \10393 , \10397 );
and \U$10294 ( \10547 , \10397 , \10402 );
and \U$10295 ( \10548 , \10393 , \10402 );
or \U$10296 ( \10549 , \10546 , \10547 , \10548 );
xor \U$10297 ( \10550 , \10545 , \10549 );
and \U$10298 ( \10551 , \10379 , \10383 );
and \U$10299 ( \10552 , \10383 , \10388 );
and \U$10300 ( \10553 , \10379 , \10388 );
or \U$10301 ( \10554 , \10551 , \10552 , \10553 );
xor \U$10302 ( \10555 , \10550 , \10554 );
xor \U$10303 ( \10556 , \10541 , \10555 );
and \U$10304 ( \10557 , \10389 , \10403 );
and \U$10305 ( \10558 , \10403 , \10415 );
and \U$10306 ( \10559 , \10389 , \10415 );
or \U$10307 ( \10560 , \10557 , \10558 , \10559 );
and \U$10308 ( \10561 , \5737 , \7140 );
not \U$10309 ( \10562 , \10561 );
xnor \U$10310 ( \10563 , \10562 , \7146 );
xor \U$10311 ( \10564 , \5984 , \10563 );
and \U$10312 ( \10565 , \5758 , \7157 );
and \U$10313 ( \10566 , \5770 , \7155 );
nor \U$10314 ( \10567 , \10565 , \10566 );
xnor \U$10315 ( \10568 , \10567 , \7163 );
xor \U$10316 ( \10569 , \10564 , \10568 );
xor \U$10317 ( \10570 , \10560 , \10569 );
and \U$10318 ( \10571 , \5906 , \5809 );
and \U$10319 ( \10572 , \5918 , \5807 );
nor \U$10320 ( \10573 , \10571 , \10572 );
xnor \U$10321 ( \10574 , \10573 , \5816 );
and \U$10322 ( \10575 , \5925 , \5829 );
and \U$10323 ( \10576 , \5937 , \5827 );
nor \U$10324 ( \10577 , \10575 , \10576 );
xnor \U$10325 ( \10578 , \10577 , \5836 );
xor \U$10326 ( \10579 , \10574 , \10578 );
and \U$10327 ( \10580 , \5945 , \5852 );
and \U$10328 ( \10581 , \5957 , \5850 );
nor \U$10329 ( \10582 , \10580 , \10581 );
xnor \U$10330 ( \10583 , \10582 , \5859 );
xor \U$10331 ( \10584 , \10579 , \10583 );
and \U$10332 ( \10585 , \5842 , \5750 );
and \U$10333 ( \10586 , \5854 , \5748 );
nor \U$10334 ( \10587 , \10585 , \10586 );
xnor \U$10335 ( \10588 , \10587 , \5755 );
and \U$10336 ( \10589 , \5861 , \5768 );
and \U$10337 ( \10590 , \5873 , \5766 );
nor \U$10338 ( \10591 , \10589 , \10590 );
xnor \U$10339 ( \10592 , \10591 , \5775 );
xor \U$10340 ( \10593 , \10588 , \10592 );
and \U$10341 ( \10594 , \5881 , \5790 );
and \U$10342 ( \10595 , \5893 , \5788 );
nor \U$10343 ( \10596 , \10594 , \10595 );
xnor \U$10344 ( \10597 , \10596 , \5797 );
xor \U$10345 ( \10598 , \10593 , \10597 );
xor \U$10346 ( \10599 , \10584 , \10598 );
and \U$10347 ( \10600 , \5780 , \7175 );
and \U$10348 ( \10601 , \5792 , \7173 );
nor \U$10349 ( \10602 , \10600 , \10601 );
xnor \U$10350 ( \10603 , \10602 , \7181 );
and \U$10351 ( \10604 , \5799 , \7192 );
and \U$10352 ( \10605 , \5811 , \7190 );
nor \U$10353 ( \10606 , \10604 , \10605 );
xnor \U$10354 ( \10607 , \10606 , \7198 );
xor \U$10355 ( \10608 , \10603 , \10607 );
and \U$10356 ( \10609 , \5819 , \7203 );
and \U$10357 ( \10610 , \5831 , \7201 );
nor \U$10358 ( \10611 , \10609 , \10610 );
xnor \U$10359 ( \10612 , \10611 , \6824 );
xor \U$10360 ( \10613 , \10608 , \10612 );
xor \U$10361 ( \10614 , \10599 , \10613 );
xor \U$10362 ( \10615 , \10570 , \10614 );
xor \U$10363 ( \10616 , \10556 , \10615 );
and \U$10364 ( \10617 , \10360 , \10364 );
and \U$10365 ( \10618 , \10364 , \10369 );
and \U$10366 ( \10619 , \10360 , \10369 );
or \U$10367 ( \10620 , \10617 , \10618 , \10619 );
and \U$10368 ( \10621 , \10346 , \10350 );
and \U$10369 ( \10622 , \10350 , \10355 );
and \U$10370 ( \10623 , \10346 , \10355 );
or \U$10371 ( \10624 , \10621 , \10622 , \10623 );
xor \U$10372 ( \10625 , \10620 , \10624 );
and \U$10373 ( \10626 , \10426 , \10440 );
and \U$10374 ( \10627 , \10440 , \10455 );
and \U$10375 ( \10628 , \10426 , \10455 );
or \U$10376 ( \10629 , \10626 , \10627 , \10628 );
xor \U$10377 ( \10630 , \10625 , \10629 );
xor \U$10378 ( \10631 , \10616 , \10630 );
xor \U$10379 ( \10632 , \10502 , \10631 );
xor \U$10380 ( \10633 , \10493 , \10632 );
and \U$10381 ( \10634 , \10318 , \10332 );
and \U$10382 ( \10635 , \10332 , \10471 );
and \U$10383 ( \10636 , \10318 , \10471 );
or \U$10384 ( \10637 , \10634 , \10635 , \10636 );
nor \U$10385 ( \10638 , \10633 , \10637 );
nor \U$10386 ( \10639 , \10477 , \10638 );
and \U$10387 ( \10640 , \10497 , \10501 );
and \U$10388 ( \10641 , \10501 , \10631 );
and \U$10389 ( \10642 , \10497 , \10631 );
or \U$10390 ( \10643 , \10640 , \10641 , \10642 );
and \U$10391 ( \10644 , \10620 , \10624 );
and \U$10392 ( \10645 , \10624 , \10629 );
and \U$10393 ( \10646 , \10620 , \10629 );
or \U$10394 ( \10647 , \10644 , \10645 , \10646 );
and \U$10395 ( \10648 , \10560 , \10569 );
and \U$10396 ( \10649 , \10569 , \10614 );
and \U$10397 ( \10650 , \10560 , \10614 );
or \U$10398 ( \10651 , \10648 , \10649 , \10650 );
xor \U$10399 ( \10652 , \10647 , \10651 );
and \U$10400 ( \10653 , \10529 , \10540 );
and \U$10401 ( \10654 , \10540 , \10555 );
and \U$10402 ( \10655 , \10529 , \10555 );
or \U$10403 ( \10656 , \10653 , \10654 , \10655 );
xor \U$10404 ( \10657 , \10652 , \10656 );
xor \U$10405 ( \10658 , \10643 , \10657 );
and \U$10406 ( \10659 , \10485 , \10489 );
and \U$10407 ( \10660 , \10489 , \10491 );
and \U$10408 ( \10661 , \10485 , \10491 );
or \U$10409 ( \10662 , \10659 , \10660 , \10661 );
and \U$10410 ( \10663 , \10556 , \10615 );
and \U$10411 ( \10664 , \10615 , \10630 );
and \U$10412 ( \10665 , \10556 , \10630 );
or \U$10413 ( \10666 , \10663 , \10664 , \10665 );
xor \U$10414 ( \10667 , \10662 , \10666 );
and \U$10415 ( \10668 , \10574 , \10578 );
and \U$10416 ( \10669 , \10578 , \10583 );
and \U$10417 ( \10670 , \10574 , \10583 );
or \U$10418 ( \10671 , \10668 , \10669 , \10670 );
and \U$10419 ( \10672 , \10518 , \10522 );
and \U$10420 ( \10673 , \10522 , \10527 );
and \U$10421 ( \10674 , \10518 , \10527 );
or \U$10422 ( \10675 , \10672 , \10673 , \10674 );
xor \U$10423 ( \10676 , \10671 , \10675 );
and \U$10424 ( \10677 , \10506 , \10510 );
and \U$10425 ( \10678 , \10510 , \10513 );
and \U$10426 ( \10679 , \10506 , \10513 );
or \U$10427 ( \10680 , \10677 , \10678 , \10679 );
xor \U$10428 ( \10681 , \10676 , \10680 );
and \U$10429 ( \10682 , \5984 , \10563 );
and \U$10430 ( \10683 , \10563 , \10568 );
and \U$10431 ( \10684 , \5984 , \10568 );
or \U$10432 ( \10685 , \10682 , \10683 , \10684 );
and \U$10433 ( \10686 , \10603 , \10607 );
and \U$10434 ( \10687 , \10607 , \10612 );
and \U$10435 ( \10688 , \10603 , \10612 );
or \U$10436 ( \10689 , \10686 , \10687 , \10688 );
xor \U$10437 ( \10690 , \10685 , \10689 );
and \U$10438 ( \10691 , \10588 , \10592 );
and \U$10439 ( \10692 , \10592 , \10597 );
and \U$10440 ( \10693 , \10588 , \10597 );
or \U$10441 ( \10694 , \10691 , \10692 , \10693 );
xor \U$10442 ( \10695 , \10690 , \10694 );
xor \U$10443 ( \10696 , \10681 , \10695 );
and \U$10444 ( \10697 , \10584 , \10598 );
and \U$10445 ( \10698 , \10598 , \10613 );
and \U$10446 ( \10699 , \10584 , \10613 );
or \U$10447 ( \10700 , \10697 , \10698 , \10699 );
and \U$10448 ( \10701 , \5873 , \5768 );
and \U$10449 ( \10702 , \5842 , \5766 );
nor \U$10450 ( \10703 , \10701 , \10702 );
xnor \U$10451 ( \10704 , \10703 , \5775 );
and \U$10452 ( \10705 , \5893 , \5790 );
and \U$10453 ( \10706 , \5861 , \5788 );
nor \U$10454 ( \10707 , \10705 , \10706 );
xnor \U$10455 ( \10708 , \10707 , \5797 );
xor \U$10456 ( \10709 , \10704 , \10708 );
and \U$10457 ( \10710 , \5918 , \5809 );
and \U$10458 ( \10711 , \5881 , \5807 );
nor \U$10459 ( \10712 , \10710 , \10711 );
xnor \U$10460 ( \10713 , \10712 , \5816 );
xor \U$10461 ( \10714 , \10709 , \10713 );
and \U$10462 ( \10715 , \5811 , \7192 );
and \U$10463 ( \10716 , \5780 , \7190 );
nor \U$10464 ( \10717 , \10715 , \10716 );
xnor \U$10465 ( \10718 , \10717 , \7198 );
and \U$10466 ( \10719 , \5831 , \7203 );
and \U$10467 ( \10720 , \5799 , \7201 );
nor \U$10468 ( \10721 , \10719 , \10720 );
xnor \U$10469 ( \10722 , \10721 , \6824 );
xor \U$10470 ( \10723 , \10718 , \10722 );
and \U$10471 ( \10724 , \5854 , \5750 );
and \U$10472 ( \10725 , \5819 , \5748 );
nor \U$10473 ( \10726 , \10724 , \10725 );
xnor \U$10474 ( \10727 , \10726 , \5755 );
xor \U$10475 ( \10728 , \10723 , \10727 );
xor \U$10476 ( \10729 , \10714 , \10728 );
not \U$10477 ( \10730 , \7146 );
and \U$10478 ( \10731 , \5770 , \7157 );
and \U$10479 ( \10732 , \5737 , \7155 );
nor \U$10480 ( \10733 , \10731 , \10732 );
xnor \U$10481 ( \10734 , \10733 , \7163 );
xor \U$10482 ( \10735 , \10730 , \10734 );
and \U$10483 ( \10736 , \5792 , \7175 );
and \U$10484 ( \10737 , \5758 , \7173 );
nor \U$10485 ( \10738 , \10736 , \10737 );
xnor \U$10486 ( \10739 , \10738 , \7181 );
xor \U$10487 ( \10740 , \10735 , \10739 );
xor \U$10488 ( \10741 , \10729 , \10740 );
xor \U$10489 ( \10742 , \10700 , \10741 );
and \U$10490 ( \10743 , \6057 , \5955 );
and \U$10491 ( \10744 , \6029 , \5953 );
nor \U$10492 ( \10745 , \10743 , \10744 );
xnor \U$10493 ( \10746 , \10745 , \5962 );
and \U$10494 ( \10747 , \6065 , \5977 );
and \U$10495 ( \10748 , \6048 , \5975 );
nor \U$10496 ( \10749 , \10747 , \10748 );
xnor \U$10497 ( \10750 , \10749 , \5984 );
xor \U$10498 ( \10751 , \10746 , \10750 );
and \U$10499 ( \10752 , \5998 , \5891 );
and \U$10500 ( \10753 , \5967 , \5889 );
nor \U$10501 ( \10754 , \10752 , \10753 );
xnor \U$10502 ( \10755 , \10754 , \5898 );
and \U$10503 ( \10756 , \6018 , \5916 );
and \U$10504 ( \10757 , \5986 , \5914 );
nor \U$10505 ( \10758 , \10756 , \10757 );
xnor \U$10506 ( \10759 , \10758 , \5923 );
xor \U$10507 ( \10760 , \10755 , \10759 );
and \U$10508 ( \10761 , \6041 , \5935 );
and \U$10509 ( \10762 , \6006 , \5933 );
nor \U$10510 ( \10763 , \10761 , \10762 );
xnor \U$10511 ( \10764 , \10763 , \5942 );
xor \U$10512 ( \10765 , \10760 , \10764 );
xor \U$10513 ( \10766 , \10751 , \10765 );
and \U$10514 ( \10767 , \5937 , \5829 );
and \U$10515 ( \10768 , \5906 , \5827 );
nor \U$10516 ( \10769 , \10767 , \10768 );
xnor \U$10517 ( \10770 , \10769 , \5836 );
and \U$10518 ( \10771 , \5957 , \5852 );
and \U$10519 ( \10772 , \5925 , \5850 );
nor \U$10520 ( \10773 , \10771 , \10772 );
xnor \U$10521 ( \10774 , \10773 , \5859 );
xor \U$10522 ( \10775 , \10770 , \10774 );
and \U$10523 ( \10776 , \5979 , \5871 );
and \U$10524 ( \10777 , \5945 , \5869 );
nor \U$10525 ( \10778 , \10776 , \10777 );
xnor \U$10526 ( \10779 , \10778 , \5878 );
xor \U$10527 ( \10780 , \10775 , \10779 );
xor \U$10528 ( \10781 , \10766 , \10780 );
xor \U$10529 ( \10782 , \10742 , \10781 );
xor \U$10530 ( \10783 , \10696 , \10782 );
and \U$10531 ( \10784 , \10545 , \10549 );
and \U$10532 ( \10785 , \10549 , \10554 );
and \U$10533 ( \10786 , \10545 , \10554 );
or \U$10534 ( \10787 , \10784 , \10785 , \10786 );
and \U$10535 ( \10788 , \10533 , \10537 );
and \U$10536 ( \10789 , \10537 , \10539 );
and \U$10537 ( \10790 , \10533 , \10539 );
or \U$10538 ( \10791 , \10788 , \10789 , \10790 );
xor \U$10539 ( \10792 , \10787 , \10791 );
or \U$10540 ( \10793 , \10514 , \10528 );
xor \U$10541 ( \10794 , \10792 , \10793 );
xor \U$10542 ( \10795 , \10783 , \10794 );
xor \U$10543 ( \10796 , \10667 , \10795 );
xor \U$10544 ( \10797 , \10658 , \10796 );
and \U$10545 ( \10798 , \10481 , \10492 );
and \U$10546 ( \10799 , \10492 , \10632 );
and \U$10547 ( \10800 , \10481 , \10632 );
or \U$10548 ( \10801 , \10798 , \10799 , \10800 );
nor \U$10549 ( \10802 , \10797 , \10801 );
and \U$10550 ( \10803 , \10662 , \10666 );
and \U$10551 ( \10804 , \10666 , \10795 );
and \U$10552 ( \10805 , \10662 , \10795 );
or \U$10553 ( \10806 , \10803 , \10804 , \10805 );
and \U$10554 ( \10807 , \10787 , \10791 );
and \U$10555 ( \10808 , \10791 , \10793 );
and \U$10556 ( \10809 , \10787 , \10793 );
or \U$10557 ( \10810 , \10807 , \10808 , \10809 );
and \U$10558 ( \10811 , \10700 , \10741 );
and \U$10559 ( \10812 , \10741 , \10781 );
and \U$10560 ( \10813 , \10700 , \10781 );
or \U$10561 ( \10814 , \10811 , \10812 , \10813 );
xor \U$10562 ( \10815 , \10810 , \10814 );
and \U$10563 ( \10816 , \10681 , \10695 );
xor \U$10564 ( \10817 , \10815 , \10816 );
xor \U$10565 ( \10818 , \10806 , \10817 );
and \U$10566 ( \10819 , \10647 , \10651 );
and \U$10567 ( \10820 , \10651 , \10656 );
and \U$10568 ( \10821 , \10647 , \10656 );
or \U$10569 ( \10822 , \10819 , \10820 , \10821 );
and \U$10570 ( \10823 , \10696 , \10782 );
and \U$10571 ( \10824 , \10782 , \10794 );
and \U$10572 ( \10825 , \10696 , \10794 );
or \U$10573 ( \10826 , \10823 , \10824 , \10825 );
xor \U$10574 ( \10827 , \10822 , \10826 );
and \U$10575 ( \10828 , \6029 , \5955 );
and \U$10576 ( \10829 , \6041 , \5953 );
nor \U$10577 ( \10830 , \10828 , \10829 );
xnor \U$10578 ( \10831 , \10830 , \5962 );
and \U$10579 ( \10832 , \6048 , \5977 );
and \U$10580 ( \10833 , \6057 , \5975 );
nor \U$10581 ( \10834 , \10832 , \10833 );
xnor \U$10582 ( \10835 , \10834 , \5984 );
xor \U$10583 ( \10836 , \10831 , \10835 );
nand \U$10584 ( \10837 , \6065 , \5994 );
xnor \U$10585 ( \10838 , \10837 , \6003 );
xor \U$10586 ( \10839 , \10836 , \10838 );
and \U$10587 ( \10840 , \5967 , \5891 );
and \U$10588 ( \10841 , \5979 , \5889 );
nor \U$10589 ( \10842 , \10840 , \10841 );
xnor \U$10590 ( \10843 , \10842 , \5898 );
and \U$10591 ( \10844 , \5986 , \5916 );
and \U$10592 ( \10845 , \5998 , \5914 );
nor \U$10593 ( \10846 , \10844 , \10845 );
xnor \U$10594 ( \10847 , \10846 , \5923 );
xor \U$10595 ( \10848 , \10843 , \10847 );
and \U$10596 ( \10849 , \6006 , \5935 );
and \U$10597 ( \10850 , \6018 , \5933 );
nor \U$10598 ( \10851 , \10849 , \10850 );
xnor \U$10599 ( \10852 , \10851 , \5942 );
xor \U$10600 ( \10853 , \10848 , \10852 );
xnor \U$10601 ( \10854 , \10839 , \10853 );
and \U$10602 ( \10855 , \10770 , \10774 );
and \U$10603 ( \10856 , \10774 , \10779 );
and \U$10604 ( \10857 , \10770 , \10779 );
or \U$10605 ( \10858 , \10855 , \10856 , \10857 );
and \U$10606 ( \10859 , \10755 , \10759 );
and \U$10607 ( \10860 , \10759 , \10764 );
and \U$10608 ( \10861 , \10755 , \10764 );
or \U$10609 ( \10862 , \10859 , \10860 , \10861 );
xor \U$10610 ( \10863 , \10858 , \10862 );
and \U$10611 ( \10864 , \10746 , \10750 );
xor \U$10612 ( \10865 , \10863 , \10864 );
xor \U$10613 ( \10866 , \10854 , \10865 );
and \U$10614 ( \10867 , \10730 , \10734 );
and \U$10615 ( \10868 , \10734 , \10739 );
and \U$10616 ( \10869 , \10730 , \10739 );
or \U$10617 ( \10870 , \10867 , \10868 , \10869 );
and \U$10618 ( \10871 , \10718 , \10722 );
and \U$10619 ( \10872 , \10722 , \10727 );
and \U$10620 ( \10873 , \10718 , \10727 );
or \U$10621 ( \10874 , \10871 , \10872 , \10873 );
xor \U$10622 ( \10875 , \10870 , \10874 );
and \U$10623 ( \10876 , \10704 , \10708 );
and \U$10624 ( \10877 , \10708 , \10713 );
and \U$10625 ( \10878 , \10704 , \10713 );
or \U$10626 ( \10879 , \10876 , \10877 , \10878 );
xor \U$10627 ( \10880 , \10875 , \10879 );
xor \U$10628 ( \10881 , \10866 , \10880 );
and \U$10629 ( \10882 , \10714 , \10728 );
and \U$10630 ( \10883 , \10728 , \10740 );
and \U$10631 ( \10884 , \10714 , \10740 );
or \U$10632 ( \10885 , \10882 , \10883 , \10884 );
and \U$10633 ( \10886 , \5737 , \7157 );
not \U$10634 ( \10887 , \10886 );
xnor \U$10635 ( \10888 , \10887 , \7163 );
xor \U$10636 ( \10889 , \6003 , \10888 );
and \U$10637 ( \10890 , \5758 , \7175 );
and \U$10638 ( \10891 , \5770 , \7173 );
nor \U$10639 ( \10892 , \10890 , \10891 );
xnor \U$10640 ( \10893 , \10892 , \7181 );
xor \U$10641 ( \10894 , \10889 , \10893 );
xor \U$10642 ( \10895 , \10885 , \10894 );
and \U$10643 ( \10896 , \5906 , \5829 );
and \U$10644 ( \10897 , \5918 , \5827 );
nor \U$10645 ( \10898 , \10896 , \10897 );
xnor \U$10646 ( \10899 , \10898 , \5836 );
and \U$10647 ( \10900 , \5925 , \5852 );
and \U$10648 ( \10901 , \5937 , \5850 );
nor \U$10649 ( \10902 , \10900 , \10901 );
xnor \U$10650 ( \10903 , \10902 , \5859 );
xor \U$10651 ( \10904 , \10899 , \10903 );
and \U$10652 ( \10905 , \5945 , \5871 );
and \U$10653 ( \10906 , \5957 , \5869 );
nor \U$10654 ( \10907 , \10905 , \10906 );
xnor \U$10655 ( \10908 , \10907 , \5878 );
xor \U$10656 ( \10909 , \10904 , \10908 );
and \U$10657 ( \10910 , \5842 , \5768 );
and \U$10658 ( \10911 , \5854 , \5766 );
nor \U$10659 ( \10912 , \10910 , \10911 );
xnor \U$10660 ( \10913 , \10912 , \5775 );
and \U$10661 ( \10914 , \5861 , \5790 );
and \U$10662 ( \10915 , \5873 , \5788 );
nor \U$10663 ( \10916 , \10914 , \10915 );
xnor \U$10664 ( \10917 , \10916 , \5797 );
xor \U$10665 ( \10918 , \10913 , \10917 );
and \U$10666 ( \10919 , \5881 , \5809 );
and \U$10667 ( \10920 , \5893 , \5807 );
nor \U$10668 ( \10921 , \10919 , \10920 );
xnor \U$10669 ( \10922 , \10921 , \5816 );
xor \U$10670 ( \10923 , \10918 , \10922 );
xor \U$10671 ( \10924 , \10909 , \10923 );
and \U$10672 ( \10925 , \5780 , \7192 );
and \U$10673 ( \10926 , \5792 , \7190 );
nor \U$10674 ( \10927 , \10925 , \10926 );
xnor \U$10675 ( \10928 , \10927 , \7198 );
and \U$10676 ( \10929 , \5799 , \7203 );
and \U$10677 ( \10930 , \5811 , \7201 );
nor \U$10678 ( \10931 , \10929 , \10930 );
xnor \U$10679 ( \10932 , \10931 , \6824 );
xor \U$10680 ( \10933 , \10928 , \10932 );
and \U$10681 ( \10934 , \5819 , \5750 );
and \U$10682 ( \10935 , \5831 , \5748 );
nor \U$10683 ( \10936 , \10934 , \10935 );
xnor \U$10684 ( \10937 , \10936 , \5755 );
xor \U$10685 ( \10938 , \10933 , \10937 );
xor \U$10686 ( \10939 , \10924 , \10938 );
xor \U$10687 ( \10940 , \10895 , \10939 );
xor \U$10688 ( \10941 , \10881 , \10940 );
and \U$10689 ( \10942 , \10685 , \10689 );
and \U$10690 ( \10943 , \10689 , \10694 );
and \U$10691 ( \10944 , \10685 , \10694 );
or \U$10692 ( \10945 , \10942 , \10943 , \10944 );
and \U$10693 ( \10946 , \10671 , \10675 );
and \U$10694 ( \10947 , \10675 , \10680 );
and \U$10695 ( \10948 , \10671 , \10680 );
or \U$10696 ( \10949 , \10946 , \10947 , \10948 );
xor \U$10697 ( \10950 , \10945 , \10949 );
and \U$10698 ( \10951 , \10751 , \10765 );
and \U$10699 ( \10952 , \10765 , \10780 );
and \U$10700 ( \10953 , \10751 , \10780 );
or \U$10701 ( \10954 , \10951 , \10952 , \10953 );
xor \U$10702 ( \10955 , \10950 , \10954 );
xor \U$10703 ( \10956 , \10941 , \10955 );
xor \U$10704 ( \10957 , \10827 , \10956 );
xor \U$10705 ( \10958 , \10818 , \10957 );
and \U$10706 ( \10959 , \10643 , \10657 );
and \U$10707 ( \10960 , \10657 , \10796 );
and \U$10708 ( \10961 , \10643 , \10796 );
or \U$10709 ( \10962 , \10959 , \10960 , \10961 );
nor \U$10710 ( \10963 , \10958 , \10962 );
nor \U$10711 ( \10964 , \10802 , \10963 );
nand \U$10712 ( \10965 , \10639 , \10964 );
and \U$10713 ( \10966 , \10822 , \10826 );
and \U$10714 ( \10967 , \10826 , \10956 );
and \U$10715 ( \10968 , \10822 , \10956 );
or \U$10716 ( \10969 , \10966 , \10967 , \10968 );
and \U$10717 ( \10970 , \10945 , \10949 );
and \U$10718 ( \10971 , \10949 , \10954 );
and \U$10719 ( \10972 , \10945 , \10954 );
or \U$10720 ( \10973 , \10970 , \10971 , \10972 );
and \U$10721 ( \10974 , \10885 , \10894 );
and \U$10722 ( \10975 , \10894 , \10939 );
and \U$10723 ( \10976 , \10885 , \10939 );
or \U$10724 ( \10977 , \10974 , \10975 , \10976 );
xor \U$10725 ( \10978 , \10973 , \10977 );
and \U$10726 ( \10979 , \10854 , \10865 );
and \U$10727 ( \10980 , \10865 , \10880 );
and \U$10728 ( \10981 , \10854 , \10880 );
or \U$10729 ( \10982 , \10979 , \10980 , \10981 );
xor \U$10730 ( \10983 , \10978 , \10982 );
xor \U$10731 ( \10984 , \10969 , \10983 );
and \U$10732 ( \10985 , \10810 , \10814 );
and \U$10733 ( \10986 , \10814 , \10816 );
and \U$10734 ( \10987 , \10810 , \10816 );
or \U$10735 ( \10988 , \10985 , \10986 , \10987 );
and \U$10736 ( \10989 , \10881 , \10940 );
and \U$10737 ( \10990 , \10940 , \10955 );
and \U$10738 ( \10991 , \10881 , \10955 );
or \U$10739 ( \10992 , \10989 , \10990 , \10991 );
xor \U$10740 ( \10993 , \10988 , \10992 );
and \U$10741 ( \10994 , \10899 , \10903 );
and \U$10742 ( \10995 , \10903 , \10908 );
and \U$10743 ( \10996 , \10899 , \10908 );
or \U$10744 ( \10997 , \10994 , \10995 , \10996 );
and \U$10745 ( \10998 , \10843 , \10847 );
and \U$10746 ( \10999 , \10847 , \10852 );
and \U$10747 ( \11000 , \10843 , \10852 );
or \U$10748 ( \11001 , \10998 , \10999 , \11000 );
xor \U$10749 ( \11002 , \10997 , \11001 );
and \U$10750 ( \11003 , \10831 , \10835 );
and \U$10751 ( \11004 , \10835 , \10838 );
and \U$10752 ( \11005 , \10831 , \10838 );
or \U$10753 ( \11006 , \11003 , \11004 , \11005 );
xor \U$10754 ( \11007 , \11002 , \11006 );
and \U$10755 ( \11008 , \6003 , \10888 );
and \U$10756 ( \11009 , \10888 , \10893 );
and \U$10757 ( \11010 , \6003 , \10893 );
or \U$10758 ( \11011 , \11008 , \11009 , \11010 );
and \U$10759 ( \11012 , \10928 , \10932 );
and \U$10760 ( \11013 , \10932 , \10937 );
and \U$10761 ( \11014 , \10928 , \10937 );
or \U$10762 ( \11015 , \11012 , \11013 , \11014 );
xor \U$10763 ( \11016 , \11011 , \11015 );
and \U$10764 ( \11017 , \10913 , \10917 );
and \U$10765 ( \11018 , \10917 , \10922 );
and \U$10766 ( \11019 , \10913 , \10922 );
or \U$10767 ( \11020 , \11017 , \11018 , \11019 );
xor \U$10768 ( \11021 , \11016 , \11020 );
xor \U$10769 ( \11022 , \11007 , \11021 );
and \U$10770 ( \11023 , \10909 , \10923 );
and \U$10771 ( \11024 , \10923 , \10938 );
and \U$10772 ( \11025 , \10909 , \10938 );
or \U$10773 ( \11026 , \11023 , \11024 , \11025 );
and \U$10774 ( \11027 , \5873 , \5790 );
and \U$10775 ( \11028 , \5842 , \5788 );
nor \U$10776 ( \11029 , \11027 , \11028 );
xnor \U$10777 ( \11030 , \11029 , \5797 );
and \U$10778 ( \11031 , \5893 , \5809 );
and \U$10779 ( \11032 , \5861 , \5807 );
nor \U$10780 ( \11033 , \11031 , \11032 );
xnor \U$10781 ( \11034 , \11033 , \5816 );
xor \U$10782 ( \11035 , \11030 , \11034 );
and \U$10783 ( \11036 , \5918 , \5829 );
and \U$10784 ( \11037 , \5881 , \5827 );
nor \U$10785 ( \11038 , \11036 , \11037 );
xnor \U$10786 ( \11039 , \11038 , \5836 );
xor \U$10787 ( \11040 , \11035 , \11039 );
and \U$10788 ( \11041 , \5811 , \7203 );
and \U$10789 ( \11042 , \5780 , \7201 );
nor \U$10790 ( \11043 , \11041 , \11042 );
xnor \U$10791 ( \11044 , \11043 , \6824 );
and \U$10792 ( \11045 , \5831 , \5750 );
and \U$10793 ( \11046 , \5799 , \5748 );
nor \U$10794 ( \11047 , \11045 , \11046 );
xnor \U$10795 ( \11048 , \11047 , \5755 );
xor \U$10796 ( \11049 , \11044 , \11048 );
and \U$10797 ( \11050 , \5854 , \5768 );
and \U$10798 ( \11051 , \5819 , \5766 );
nor \U$10799 ( \11052 , \11050 , \11051 );
xnor \U$10800 ( \11053 , \11052 , \5775 );
xor \U$10801 ( \11054 , \11049 , \11053 );
xor \U$10802 ( \11055 , \11040 , \11054 );
not \U$10803 ( \11056 , \7163 );
and \U$10804 ( \11057 , \5770 , \7175 );
and \U$10805 ( \11058 , \5737 , \7173 );
nor \U$10806 ( \11059 , \11057 , \11058 );
xnor \U$10807 ( \11060 , \11059 , \7181 );
xor \U$10808 ( \11061 , \11056 , \11060 );
and \U$10809 ( \11062 , \5792 , \7192 );
and \U$10810 ( \11063 , \5758 , \7190 );
nor \U$10811 ( \11064 , \11062 , \11063 );
xnor \U$10812 ( \11065 , \11064 , \7198 );
xor \U$10813 ( \11066 , \11061 , \11065 );
xor \U$10814 ( \11067 , \11055 , \11066 );
xor \U$10815 ( \11068 , \11026 , \11067 );
and \U$10816 ( \11069 , \6057 , \5977 );
and \U$10817 ( \11070 , \6029 , \5975 );
nor \U$10818 ( \11071 , \11069 , \11070 );
xnor \U$10819 ( \11072 , \11071 , \5984 );
and \U$10820 ( \11073 , \6065 , \5996 );
and \U$10821 ( \11074 , \6048 , \5994 );
nor \U$10822 ( \11075 , \11073 , \11074 );
xnor \U$10823 ( \11076 , \11075 , \6003 );
xor \U$10824 ( \11077 , \11072 , \11076 );
and \U$10825 ( \11078 , \5998 , \5916 );
and \U$10826 ( \11079 , \5967 , \5914 );
nor \U$10827 ( \11080 , \11078 , \11079 );
xnor \U$10828 ( \11081 , \11080 , \5923 );
and \U$10829 ( \11082 , \6018 , \5935 );
and \U$10830 ( \11083 , \5986 , \5933 );
nor \U$10831 ( \11084 , \11082 , \11083 );
xnor \U$10832 ( \11085 , \11084 , \5942 );
xor \U$10833 ( \11086 , \11081 , \11085 );
and \U$10834 ( \11087 , \6041 , \5955 );
and \U$10835 ( \11088 , \6006 , \5953 );
nor \U$10836 ( \11089 , \11087 , \11088 );
xnor \U$10837 ( \11090 , \11089 , \5962 );
xor \U$10838 ( \11091 , \11086 , \11090 );
xor \U$10839 ( \11092 , \11077 , \11091 );
and \U$10840 ( \11093 , \5937 , \5852 );
and \U$10841 ( \11094 , \5906 , \5850 );
nor \U$10842 ( \11095 , \11093 , \11094 );
xnor \U$10843 ( \11096 , \11095 , \5859 );
and \U$10844 ( \11097 , \5957 , \5871 );
and \U$10845 ( \11098 , \5925 , \5869 );
nor \U$10846 ( \11099 , \11097 , \11098 );
xnor \U$10847 ( \11100 , \11099 , \5878 );
xor \U$10848 ( \11101 , \11096 , \11100 );
and \U$10849 ( \11102 , \5979 , \5891 );
and \U$10850 ( \11103 , \5945 , \5889 );
nor \U$10851 ( \11104 , \11102 , \11103 );
xnor \U$10852 ( \11105 , \11104 , \5898 );
xor \U$10853 ( \11106 , \11101 , \11105 );
xor \U$10854 ( \11107 , \11092 , \11106 );
xor \U$10855 ( \11108 , \11068 , \11107 );
xor \U$10856 ( \11109 , \11022 , \11108 );
and \U$10857 ( \11110 , \10870 , \10874 );
and \U$10858 ( \11111 , \10874 , \10879 );
and \U$10859 ( \11112 , \10870 , \10879 );
or \U$10860 ( \11113 , \11110 , \11111 , \11112 );
and \U$10861 ( \11114 , \10858 , \10862 );
and \U$10862 ( \11115 , \10862 , \10864 );
and \U$10863 ( \11116 , \10858 , \10864 );
or \U$10864 ( \11117 , \11114 , \11115 , \11116 );
xor \U$10865 ( \11118 , \11113 , \11117 );
or \U$10866 ( \11119 , \10839 , \10853 );
xor \U$10867 ( \11120 , \11118 , \11119 );
xor \U$10868 ( \11121 , \11109 , \11120 );
xor \U$10869 ( \11122 , \10993 , \11121 );
xor \U$10870 ( \11123 , \10984 , \11122 );
and \U$10871 ( \11124 , \10806 , \10817 );
and \U$10872 ( \11125 , \10817 , \10957 );
and \U$10873 ( \11126 , \10806 , \10957 );
or \U$10874 ( \11127 , \11124 , \11125 , \11126 );
nor \U$10875 ( \11128 , \11123 , \11127 );
and \U$10876 ( \11129 , \10988 , \10992 );
and \U$10877 ( \11130 , \10992 , \11121 );
and \U$10878 ( \11131 , \10988 , \11121 );
or \U$10879 ( \11132 , \11129 , \11130 , \11131 );
and \U$10880 ( \11133 , \11113 , \11117 );
and \U$10881 ( \11134 , \11117 , \11119 );
and \U$10882 ( \11135 , \11113 , \11119 );
or \U$10883 ( \11136 , \11133 , \11134 , \11135 );
and \U$10884 ( \11137 , \11026 , \11067 );
and \U$10885 ( \11138 , \11067 , \11107 );
and \U$10886 ( \11139 , \11026 , \11107 );
or \U$10887 ( \11140 , \11137 , \11138 , \11139 );
xor \U$10888 ( \11141 , \11136 , \11140 );
and \U$10889 ( \11142 , \11007 , \11021 );
xor \U$10890 ( \11143 , \11141 , \11142 );
xor \U$10891 ( \11144 , \11132 , \11143 );
and \U$10892 ( \11145 , \10973 , \10977 );
and \U$10893 ( \11146 , \10977 , \10982 );
and \U$10894 ( \11147 , \10973 , \10982 );
or \U$10895 ( \11148 , \11145 , \11146 , \11147 );
and \U$10896 ( \11149 , \11022 , \11108 );
and \U$10897 ( \11150 , \11108 , \11120 );
and \U$10898 ( \11151 , \11022 , \11120 );
or \U$10899 ( \11152 , \11149 , \11150 , \11151 );
xor \U$10900 ( \11153 , \11148 , \11152 );
and \U$10901 ( \11154 , \6029 , \5977 );
and \U$10902 ( \11155 , \6041 , \5975 );
nor \U$10903 ( \11156 , \11154 , \11155 );
xnor \U$10904 ( \11157 , \11156 , \5984 );
and \U$10905 ( \11158 , \6048 , \5996 );
and \U$10906 ( \11159 , \6057 , \5994 );
nor \U$10907 ( \11160 , \11158 , \11159 );
xnor \U$10908 ( \11161 , \11160 , \6003 );
xor \U$10909 ( \11162 , \11157 , \11161 );
nand \U$10910 ( \11163 , \6065 , \6014 );
xnor \U$10911 ( \11164 , \11163 , \6023 );
xor \U$10912 ( \11165 , \11162 , \11164 );
and \U$10913 ( \11166 , \5967 , \5916 );
and \U$10914 ( \11167 , \5979 , \5914 );
nor \U$10915 ( \11168 , \11166 , \11167 );
xnor \U$10916 ( \11169 , \11168 , \5923 );
and \U$10917 ( \11170 , \5986 , \5935 );
and \U$10918 ( \11171 , \5998 , \5933 );
nor \U$10919 ( \11172 , \11170 , \11171 );
xnor \U$10920 ( \11173 , \11172 , \5942 );
xor \U$10921 ( \11174 , \11169 , \11173 );
and \U$10922 ( \11175 , \6006 , \5955 );
and \U$10923 ( \11176 , \6018 , \5953 );
nor \U$10924 ( \11177 , \11175 , \11176 );
xnor \U$10925 ( \11178 , \11177 , \5962 );
xor \U$10926 ( \11179 , \11174 , \11178 );
xnor \U$10927 ( \11180 , \11165 , \11179 );
and \U$10928 ( \11181 , \11096 , \11100 );
and \U$10929 ( \11182 , \11100 , \11105 );
and \U$10930 ( \11183 , \11096 , \11105 );
or \U$10931 ( \11184 , \11181 , \11182 , \11183 );
and \U$10932 ( \11185 , \11081 , \11085 );
and \U$10933 ( \11186 , \11085 , \11090 );
and \U$10934 ( \11187 , \11081 , \11090 );
or \U$10935 ( \11188 , \11185 , \11186 , \11187 );
xor \U$10936 ( \11189 , \11184 , \11188 );
and \U$10937 ( \11190 , \11072 , \11076 );
xor \U$10938 ( \11191 , \11189 , \11190 );
xor \U$10939 ( \11192 , \11180 , \11191 );
and \U$10940 ( \11193 , \11056 , \11060 );
and \U$10941 ( \11194 , \11060 , \11065 );
and \U$10942 ( \11195 , \11056 , \11065 );
or \U$10943 ( \11196 , \11193 , \11194 , \11195 );
and \U$10944 ( \11197 , \11044 , \11048 );
and \U$10945 ( \11198 , \11048 , \11053 );
and \U$10946 ( \11199 , \11044 , \11053 );
or \U$10947 ( \11200 , \11197 , \11198 , \11199 );
xor \U$10948 ( \11201 , \11196 , \11200 );
and \U$10949 ( \11202 , \11030 , \11034 );
and \U$10950 ( \11203 , \11034 , \11039 );
and \U$10951 ( \11204 , \11030 , \11039 );
or \U$10952 ( \11205 , \11202 , \11203 , \11204 );
xor \U$10953 ( \11206 , \11201 , \11205 );
xor \U$10954 ( \11207 , \11192 , \11206 );
and \U$10955 ( \11208 , \11040 , \11054 );
and \U$10956 ( \11209 , \11054 , \11066 );
and \U$10957 ( \11210 , \11040 , \11066 );
or \U$10958 ( \11211 , \11208 , \11209 , \11210 );
and \U$10959 ( \11212 , \5737 , \7175 );
not \U$10960 ( \11213 , \11212 );
xnor \U$10961 ( \11214 , \11213 , \7181 );
xor \U$10962 ( \11215 , \6023 , \11214 );
and \U$10963 ( \11216 , \5758 , \7192 );
and \U$10964 ( \11217 , \5770 , \7190 );
nor \U$10965 ( \11218 , \11216 , \11217 );
xnor \U$10966 ( \11219 , \11218 , \7198 );
xor \U$10967 ( \11220 , \11215 , \11219 );
xor \U$10968 ( \11221 , \11211 , \11220 );
and \U$10969 ( \11222 , \5906 , \5852 );
and \U$10970 ( \11223 , \5918 , \5850 );
nor \U$10971 ( \11224 , \11222 , \11223 );
xnor \U$10972 ( \11225 , \11224 , \5859 );
and \U$10973 ( \11226 , \5925 , \5871 );
and \U$10974 ( \11227 , \5937 , \5869 );
nor \U$10975 ( \11228 , \11226 , \11227 );
xnor \U$10976 ( \11229 , \11228 , \5878 );
xor \U$10977 ( \11230 , \11225 , \11229 );
and \U$10978 ( \11231 , \5945 , \5891 );
and \U$10979 ( \11232 , \5957 , \5889 );
nor \U$10980 ( \11233 , \11231 , \11232 );
xnor \U$10981 ( \11234 , \11233 , \5898 );
xor \U$10982 ( \11235 , \11230 , \11234 );
and \U$10983 ( \11236 , \5842 , \5790 );
and \U$10984 ( \11237 , \5854 , \5788 );
nor \U$10985 ( \11238 , \11236 , \11237 );
xnor \U$10986 ( \11239 , \11238 , \5797 );
and \U$10987 ( \11240 , \5861 , \5809 );
and \U$10988 ( \11241 , \5873 , \5807 );
nor \U$10989 ( \11242 , \11240 , \11241 );
xnor \U$10990 ( \11243 , \11242 , \5816 );
xor \U$10991 ( \11244 , \11239 , \11243 );
and \U$10992 ( \11245 , \5881 , \5829 );
and \U$10993 ( \11246 , \5893 , \5827 );
nor \U$10994 ( \11247 , \11245 , \11246 );
xnor \U$10995 ( \11248 , \11247 , \5836 );
xor \U$10996 ( \11249 , \11244 , \11248 );
xor \U$10997 ( \11250 , \11235 , \11249 );
and \U$10998 ( \11251 , \5780 , \7203 );
and \U$10999 ( \11252 , \5792 , \7201 );
nor \U$11000 ( \11253 , \11251 , \11252 );
xnor \U$11001 ( \11254 , \11253 , \6824 );
and \U$11002 ( \11255 , \5799 , \5750 );
and \U$11003 ( \11256 , \5811 , \5748 );
nor \U$11004 ( \11257 , \11255 , \11256 );
xnor \U$11005 ( \11258 , \11257 , \5755 );
xor \U$11006 ( \11259 , \11254 , \11258 );
and \U$11007 ( \11260 , \5819 , \5768 );
and \U$11008 ( \11261 , \5831 , \5766 );
nor \U$11009 ( \11262 , \11260 , \11261 );
xnor \U$11010 ( \11263 , \11262 , \5775 );
xor \U$11011 ( \11264 , \11259 , \11263 );
xor \U$11012 ( \11265 , \11250 , \11264 );
xor \U$11013 ( \11266 , \11221 , \11265 );
xor \U$11014 ( \11267 , \11207 , \11266 );
and \U$11015 ( \11268 , \11011 , \11015 );
and \U$11016 ( \11269 , \11015 , \11020 );
and \U$11017 ( \11270 , \11011 , \11020 );
or \U$11018 ( \11271 , \11268 , \11269 , \11270 );
and \U$11019 ( \11272 , \10997 , \11001 );
and \U$11020 ( \11273 , \11001 , \11006 );
and \U$11021 ( \11274 , \10997 , \11006 );
or \U$11022 ( \11275 , \11272 , \11273 , \11274 );
xor \U$11023 ( \11276 , \11271 , \11275 );
and \U$11024 ( \11277 , \11077 , \11091 );
and \U$11025 ( \11278 , \11091 , \11106 );
and \U$11026 ( \11279 , \11077 , \11106 );
or \U$11027 ( \11280 , \11277 , \11278 , \11279 );
xor \U$11028 ( \11281 , \11276 , \11280 );
xor \U$11029 ( \11282 , \11267 , \11281 );
xor \U$11030 ( \11283 , \11153 , \11282 );
xor \U$11031 ( \11284 , \11144 , \11283 );
and \U$11032 ( \11285 , \10969 , \10983 );
and \U$11033 ( \11286 , \10983 , \11122 );
and \U$11034 ( \11287 , \10969 , \11122 );
or \U$11035 ( \11288 , \11285 , \11286 , \11287 );
nor \U$11036 ( \11289 , \11284 , \11288 );
nor \U$11037 ( \11290 , \11128 , \11289 );
and \U$11038 ( \11291 , \11148 , \11152 );
and \U$11039 ( \11292 , \11152 , \11282 );
and \U$11040 ( \11293 , \11148 , \11282 );
or \U$11041 ( \11294 , \11291 , \11292 , \11293 );
and \U$11042 ( \11295 , \11271 , \11275 );
and \U$11043 ( \11296 , \11275 , \11280 );
and \U$11044 ( \11297 , \11271 , \11280 );
or \U$11045 ( \11298 , \11295 , \11296 , \11297 );
and \U$11046 ( \11299 , \11211 , \11220 );
and \U$11047 ( \11300 , \11220 , \11265 );
and \U$11048 ( \11301 , \11211 , \11265 );
or \U$11049 ( \11302 , \11299 , \11300 , \11301 );
xor \U$11050 ( \11303 , \11298 , \11302 );
and \U$11051 ( \11304 , \11180 , \11191 );
and \U$11052 ( \11305 , \11191 , \11206 );
and \U$11053 ( \11306 , \11180 , \11206 );
or \U$11054 ( \11307 , \11304 , \11305 , \11306 );
xor \U$11055 ( \11308 , \11303 , \11307 );
xor \U$11056 ( \11309 , \11294 , \11308 );
and \U$11057 ( \11310 , \11136 , \11140 );
and \U$11058 ( \11311 , \11140 , \11142 );
and \U$11059 ( \11312 , \11136 , \11142 );
or \U$11060 ( \11313 , \11310 , \11311 , \11312 );
and \U$11061 ( \11314 , \11207 , \11266 );
and \U$11062 ( \11315 , \11266 , \11281 );
and \U$11063 ( \11316 , \11207 , \11281 );
or \U$11064 ( \11317 , \11314 , \11315 , \11316 );
xor \U$11065 ( \11318 , \11313 , \11317 );
and \U$11066 ( \11319 , \11225 , \11229 );
and \U$11067 ( \11320 , \11229 , \11234 );
and \U$11068 ( \11321 , \11225 , \11234 );
or \U$11069 ( \11322 , \11319 , \11320 , \11321 );
and \U$11070 ( \11323 , \11169 , \11173 );
and \U$11071 ( \11324 , \11173 , \11178 );
and \U$11072 ( \11325 , \11169 , \11178 );
or \U$11073 ( \11326 , \11323 , \11324 , \11325 );
xor \U$11074 ( \11327 , \11322 , \11326 );
and \U$11075 ( \11328 , \11157 , \11161 );
and \U$11076 ( \11329 , \11161 , \11164 );
and \U$11077 ( \11330 , \11157 , \11164 );
or \U$11078 ( \11331 , \11328 , \11329 , \11330 );
xor \U$11079 ( \11332 , \11327 , \11331 );
and \U$11080 ( \11333 , \6023 , \11214 );
and \U$11081 ( \11334 , \11214 , \11219 );
and \U$11082 ( \11335 , \6023 , \11219 );
or \U$11083 ( \11336 , \11333 , \11334 , \11335 );
and \U$11084 ( \11337 , \11254 , \11258 );
and \U$11085 ( \11338 , \11258 , \11263 );
and \U$11086 ( \11339 , \11254 , \11263 );
or \U$11087 ( \11340 , \11337 , \11338 , \11339 );
xor \U$11088 ( \11341 , \11336 , \11340 );
and \U$11089 ( \11342 , \11239 , \11243 );
and \U$11090 ( \11343 , \11243 , \11248 );
and \U$11091 ( \11344 , \11239 , \11248 );
or \U$11092 ( \11345 , \11342 , \11343 , \11344 );
xor \U$11093 ( \11346 , \11341 , \11345 );
xor \U$11094 ( \11347 , \11332 , \11346 );
and \U$11095 ( \11348 , \11235 , \11249 );
and \U$11096 ( \11349 , \11249 , \11264 );
and \U$11097 ( \11350 , \11235 , \11264 );
or \U$11098 ( \11351 , \11348 , \11349 , \11350 );
and \U$11099 ( \11352 , \5873 , \5809 );
and \U$11100 ( \11353 , \5842 , \5807 );
nor \U$11101 ( \11354 , \11352 , \11353 );
xnor \U$11102 ( \11355 , \11354 , \5816 );
and \U$11103 ( \11356 , \5893 , \5829 );
and \U$11104 ( \11357 , \5861 , \5827 );
nor \U$11105 ( \11358 , \11356 , \11357 );
xnor \U$11106 ( \11359 , \11358 , \5836 );
xor \U$11107 ( \11360 , \11355 , \11359 );
and \U$11108 ( \11361 , \5918 , \5852 );
and \U$11109 ( \11362 , \5881 , \5850 );
nor \U$11110 ( \11363 , \11361 , \11362 );
xnor \U$11111 ( \11364 , \11363 , \5859 );
xor \U$11112 ( \11365 , \11360 , \11364 );
and \U$11113 ( \11366 , \5811 , \5750 );
and \U$11114 ( \11367 , \5780 , \5748 );
nor \U$11115 ( \11368 , \11366 , \11367 );
xnor \U$11116 ( \11369 , \11368 , \5755 );
and \U$11117 ( \11370 , \5831 , \5768 );
and \U$11118 ( \11371 , \5799 , \5766 );
nor \U$11119 ( \11372 , \11370 , \11371 );
xnor \U$11120 ( \11373 , \11372 , \5775 );
xor \U$11121 ( \11374 , \11369 , \11373 );
and \U$11122 ( \11375 , \5854 , \5790 );
and \U$11123 ( \11376 , \5819 , \5788 );
nor \U$11124 ( \11377 , \11375 , \11376 );
xnor \U$11125 ( \11378 , \11377 , \5797 );
xor \U$11126 ( \11379 , \11374 , \11378 );
xor \U$11127 ( \11380 , \11365 , \11379 );
not \U$11128 ( \11381 , \7181 );
and \U$11129 ( \11382 , \5770 , \7192 );
and \U$11130 ( \11383 , \5737 , \7190 );
nor \U$11131 ( \11384 , \11382 , \11383 );
xnor \U$11132 ( \11385 , \11384 , \7198 );
xor \U$11133 ( \11386 , \11381 , \11385 );
and \U$11134 ( \11387 , \5792 , \7203 );
and \U$11135 ( \11388 , \5758 , \7201 );
nor \U$11136 ( \11389 , \11387 , \11388 );
xnor \U$11137 ( \11390 , \11389 , \6824 );
xor \U$11138 ( \11391 , \11386 , \11390 );
xor \U$11139 ( \11392 , \11380 , \11391 );
xor \U$11140 ( \11393 , \11351 , \11392 );
and \U$11141 ( \11394 , \6057 , \5996 );
and \U$11142 ( \11395 , \6029 , \5994 );
nor \U$11143 ( \11396 , \11394 , \11395 );
xnor \U$11144 ( \11397 , \11396 , \6003 );
and \U$11145 ( \11398 , \6065 , \6016 );
and \U$11146 ( \11399 , \6048 , \6014 );
nor \U$11147 ( \11400 , \11398 , \11399 );
xnor \U$11148 ( \11401 , \11400 , \6023 );
xor \U$11149 ( \11402 , \11397 , \11401 );
and \U$11150 ( \11403 , \5998 , \5935 );
and \U$11151 ( \11404 , \5967 , \5933 );
nor \U$11152 ( \11405 , \11403 , \11404 );
xnor \U$11153 ( \11406 , \11405 , \5942 );
and \U$11154 ( \11407 , \6018 , \5955 );
and \U$11155 ( \11408 , \5986 , \5953 );
nor \U$11156 ( \11409 , \11407 , \11408 );
xnor \U$11157 ( \11410 , \11409 , \5962 );
xor \U$11158 ( \11411 , \11406 , \11410 );
and \U$11159 ( \11412 , \6041 , \5977 );
and \U$11160 ( \11413 , \6006 , \5975 );
nor \U$11161 ( \11414 , \11412 , \11413 );
xnor \U$11162 ( \11415 , \11414 , \5984 );
xor \U$11163 ( \11416 , \11411 , \11415 );
xor \U$11164 ( \11417 , \11402 , \11416 );
and \U$11165 ( \11418 , \5937 , \5871 );
and \U$11166 ( \11419 , \5906 , \5869 );
nor \U$11167 ( \11420 , \11418 , \11419 );
xnor \U$11168 ( \11421 , \11420 , \5878 );
and \U$11169 ( \11422 , \5957 , \5891 );
and \U$11170 ( \11423 , \5925 , \5889 );
nor \U$11171 ( \11424 , \11422 , \11423 );
xnor \U$11172 ( \11425 , \11424 , \5898 );
xor \U$11173 ( \11426 , \11421 , \11425 );
and \U$11174 ( \11427 , \5979 , \5916 );
and \U$11175 ( \11428 , \5945 , \5914 );
nor \U$11176 ( \11429 , \11427 , \11428 );
xnor \U$11177 ( \11430 , \11429 , \5923 );
xor \U$11178 ( \11431 , \11426 , \11430 );
xor \U$11179 ( \11432 , \11417 , \11431 );
xor \U$11180 ( \11433 , \11393 , \11432 );
xor \U$11181 ( \11434 , \11347 , \11433 );
and \U$11182 ( \11435 , \11196 , \11200 );
and \U$11183 ( \11436 , \11200 , \11205 );
and \U$11184 ( \11437 , \11196 , \11205 );
or \U$11185 ( \11438 , \11435 , \11436 , \11437 );
and \U$11186 ( \11439 , \11184 , \11188 );
and \U$11187 ( \11440 , \11188 , \11190 );
and \U$11188 ( \11441 , \11184 , \11190 );
or \U$11189 ( \11442 , \11439 , \11440 , \11441 );
xor \U$11190 ( \11443 , \11438 , \11442 );
or \U$11191 ( \11444 , \11165 , \11179 );
xor \U$11192 ( \11445 , \11443 , \11444 );
xor \U$11193 ( \11446 , \11434 , \11445 );
xor \U$11194 ( \11447 , \11318 , \11446 );
xor \U$11195 ( \11448 , \11309 , \11447 );
and \U$11196 ( \11449 , \11132 , \11143 );
and \U$11197 ( \11450 , \11143 , \11283 );
and \U$11198 ( \11451 , \11132 , \11283 );
or \U$11199 ( \11452 , \11449 , \11450 , \11451 );
nor \U$11200 ( \11453 , \11448 , \11452 );
and \U$11201 ( \11454 , \11313 , \11317 );
and \U$11202 ( \11455 , \11317 , \11446 );
and \U$11203 ( \11456 , \11313 , \11446 );
or \U$11204 ( \11457 , \11454 , \11455 , \11456 );
and \U$11205 ( \11458 , \11438 , \11442 );
and \U$11206 ( \11459 , \11442 , \11444 );
and \U$11207 ( \11460 , \11438 , \11444 );
or \U$11208 ( \11461 , \11458 , \11459 , \11460 );
and \U$11209 ( \11462 , \11351 , \11392 );
and \U$11210 ( \11463 , \11392 , \11432 );
and \U$11211 ( \11464 , \11351 , \11432 );
or \U$11212 ( \11465 , \11462 , \11463 , \11464 );
xor \U$11213 ( \11466 , \11461 , \11465 );
and \U$11214 ( \11467 , \11332 , \11346 );
xor \U$11215 ( \11468 , \11466 , \11467 );
xor \U$11216 ( \11469 , \11457 , \11468 );
and \U$11217 ( \11470 , \11298 , \11302 );
and \U$11218 ( \11471 , \11302 , \11307 );
and \U$11219 ( \11472 , \11298 , \11307 );
or \U$11220 ( \11473 , \11470 , \11471 , \11472 );
and \U$11221 ( \11474 , \11347 , \11433 );
and \U$11222 ( \11475 , \11433 , \11445 );
and \U$11223 ( \11476 , \11347 , \11445 );
or \U$11224 ( \11477 , \11474 , \11475 , \11476 );
xor \U$11225 ( \11478 , \11473 , \11477 );
and \U$11226 ( \11479 , \6029 , \5996 );
and \U$11227 ( \11480 , \6041 , \5994 );
nor \U$11228 ( \11481 , \11479 , \11480 );
xnor \U$11229 ( \11482 , \11481 , \6003 );
and \U$11230 ( \11483 , \6048 , \6016 );
and \U$11231 ( \11484 , \6057 , \6014 );
nor \U$11232 ( \11485 , \11483 , \11484 );
xnor \U$11233 ( \11486 , \11485 , \6023 );
xor \U$11234 ( \11487 , \11482 , \11486 );
nand \U$11235 ( \11488 , \6065 , \6037 );
xnor \U$11236 ( \11489 , \11488 , \6046 );
xor \U$11237 ( \11490 , \11487 , \11489 );
and \U$11238 ( \11491 , \5967 , \5935 );
and \U$11239 ( \11492 , \5979 , \5933 );
nor \U$11240 ( \11493 , \11491 , \11492 );
xnor \U$11241 ( \11494 , \11493 , \5942 );
and \U$11242 ( \11495 , \5986 , \5955 );
and \U$11243 ( \11496 , \5998 , \5953 );
nor \U$11244 ( \11497 , \11495 , \11496 );
xnor \U$11245 ( \11498 , \11497 , \5962 );
xor \U$11246 ( \11499 , \11494 , \11498 );
and \U$11247 ( \11500 , \6006 , \5977 );
and \U$11248 ( \11501 , \6018 , \5975 );
nor \U$11249 ( \11502 , \11500 , \11501 );
xnor \U$11250 ( \11503 , \11502 , \5984 );
xor \U$11251 ( \11504 , \11499 , \11503 );
xnor \U$11252 ( \11505 , \11490 , \11504 );
and \U$11253 ( \11506 , \11421 , \11425 );
and \U$11254 ( \11507 , \11425 , \11430 );
and \U$11255 ( \11508 , \11421 , \11430 );
or \U$11256 ( \11509 , \11506 , \11507 , \11508 );
and \U$11257 ( \11510 , \11406 , \11410 );
and \U$11258 ( \11511 , \11410 , \11415 );
and \U$11259 ( \11512 , \11406 , \11415 );
or \U$11260 ( \11513 , \11510 , \11511 , \11512 );
xor \U$11261 ( \11514 , \11509 , \11513 );
and \U$11262 ( \11515 , \11397 , \11401 );
xor \U$11263 ( \11516 , \11514 , \11515 );
xor \U$11264 ( \11517 , \11505 , \11516 );
and \U$11265 ( \11518 , \11381 , \11385 );
and \U$11266 ( \11519 , \11385 , \11390 );
and \U$11267 ( \11520 , \11381 , \11390 );
or \U$11268 ( \11521 , \11518 , \11519 , \11520 );
and \U$11269 ( \11522 , \11369 , \11373 );
and \U$11270 ( \11523 , \11373 , \11378 );
and \U$11271 ( \11524 , \11369 , \11378 );
or \U$11272 ( \11525 , \11522 , \11523 , \11524 );
xor \U$11273 ( \11526 , \11521 , \11525 );
and \U$11274 ( \11527 , \11355 , \11359 );
and \U$11275 ( \11528 , \11359 , \11364 );
and \U$11276 ( \11529 , \11355 , \11364 );
or \U$11277 ( \11530 , \11527 , \11528 , \11529 );
xor \U$11278 ( \11531 , \11526 , \11530 );
xor \U$11279 ( \11532 , \11517 , \11531 );
and \U$11280 ( \11533 , \11365 , \11379 );
and \U$11281 ( \11534 , \11379 , \11391 );
and \U$11282 ( \11535 , \11365 , \11391 );
or \U$11283 ( \11536 , \11533 , \11534 , \11535 );
and \U$11284 ( \11537 , \5737 , \7192 );
not \U$11285 ( \11538 , \11537 );
xnor \U$11286 ( \11539 , \11538 , \7198 );
xor \U$11287 ( \11540 , \6046 , \11539 );
and \U$11288 ( \11541 , \5758 , \7203 );
and \U$11289 ( \11542 , \5770 , \7201 );
nor \U$11290 ( \11543 , \11541 , \11542 );
xnor \U$11291 ( \11544 , \11543 , \6824 );
xor \U$11292 ( \11545 , \11540 , \11544 );
xor \U$11293 ( \11546 , \11536 , \11545 );
and \U$11294 ( \11547 , \5906 , \5871 );
and \U$11295 ( \11548 , \5918 , \5869 );
nor \U$11296 ( \11549 , \11547 , \11548 );
xnor \U$11297 ( \11550 , \11549 , \5878 );
and \U$11298 ( \11551 , \5925 , \5891 );
and \U$11299 ( \11552 , \5937 , \5889 );
nor \U$11300 ( \11553 , \11551 , \11552 );
xnor \U$11301 ( \11554 , \11553 , \5898 );
xor \U$11302 ( \11555 , \11550 , \11554 );
and \U$11303 ( \11556 , \5945 , \5916 );
and \U$11304 ( \11557 , \5957 , \5914 );
nor \U$11305 ( \11558 , \11556 , \11557 );
xnor \U$11306 ( \11559 , \11558 , \5923 );
xor \U$11307 ( \11560 , \11555 , \11559 );
and \U$11308 ( \11561 , \5842 , \5809 );
and \U$11309 ( \11562 , \5854 , \5807 );
nor \U$11310 ( \11563 , \11561 , \11562 );
xnor \U$11311 ( \11564 , \11563 , \5816 );
and \U$11312 ( \11565 , \5861 , \5829 );
and \U$11313 ( \11566 , \5873 , \5827 );
nor \U$11314 ( \11567 , \11565 , \11566 );
xnor \U$11315 ( \11568 , \11567 , \5836 );
xor \U$11316 ( \11569 , \11564 , \11568 );
and \U$11317 ( \11570 , \5881 , \5852 );
and \U$11318 ( \11571 , \5893 , \5850 );
nor \U$11319 ( \11572 , \11570 , \11571 );
xnor \U$11320 ( \11573 , \11572 , \5859 );
xor \U$11321 ( \11574 , \11569 , \11573 );
xor \U$11322 ( \11575 , \11560 , \11574 );
and \U$11323 ( \11576 , \5780 , \5750 );
and \U$11324 ( \11577 , \5792 , \5748 );
nor \U$11325 ( \11578 , \11576 , \11577 );
xnor \U$11326 ( \11579 , \11578 , \5755 );
and \U$11327 ( \11580 , \5799 , \5768 );
and \U$11328 ( \11581 , \5811 , \5766 );
nor \U$11329 ( \11582 , \11580 , \11581 );
xnor \U$11330 ( \11583 , \11582 , \5775 );
xor \U$11331 ( \11584 , \11579 , \11583 );
and \U$11332 ( \11585 , \5819 , \5790 );
and \U$11333 ( \11586 , \5831 , \5788 );
nor \U$11334 ( \11587 , \11585 , \11586 );
xnor \U$11335 ( \11588 , \11587 , \5797 );
xor \U$11336 ( \11589 , \11584 , \11588 );
xor \U$11337 ( \11590 , \11575 , \11589 );
xor \U$11338 ( \11591 , \11546 , \11590 );
xor \U$11339 ( \11592 , \11532 , \11591 );
and \U$11340 ( \11593 , \11336 , \11340 );
and \U$11341 ( \11594 , \11340 , \11345 );
and \U$11342 ( \11595 , \11336 , \11345 );
or \U$11343 ( \11596 , \11593 , \11594 , \11595 );
and \U$11344 ( \11597 , \11322 , \11326 );
and \U$11345 ( \11598 , \11326 , \11331 );
and \U$11346 ( \11599 , \11322 , \11331 );
or \U$11347 ( \11600 , \11597 , \11598 , \11599 );
xor \U$11348 ( \11601 , \11596 , \11600 );
and \U$11349 ( \11602 , \11402 , \11416 );
and \U$11350 ( \11603 , \11416 , \11431 );
and \U$11351 ( \11604 , \11402 , \11431 );
or \U$11352 ( \11605 , \11602 , \11603 , \11604 );
xor \U$11353 ( \11606 , \11601 , \11605 );
xor \U$11354 ( \11607 , \11592 , \11606 );
xor \U$11355 ( \11608 , \11478 , \11607 );
xor \U$11356 ( \11609 , \11469 , \11608 );
and \U$11357 ( \11610 , \11294 , \11308 );
and \U$11358 ( \11611 , \11308 , \11447 );
and \U$11359 ( \11612 , \11294 , \11447 );
or \U$11360 ( \11613 , \11610 , \11611 , \11612 );
nor \U$11361 ( \11614 , \11609 , \11613 );
nor \U$11362 ( \11615 , \11453 , \11614 );
nand \U$11363 ( \11616 , \11290 , \11615 );
nor \U$11364 ( \11617 , \10965 , \11616 );
and \U$11365 ( \11618 , \11473 , \11477 );
and \U$11366 ( \11619 , \11477 , \11607 );
and \U$11367 ( \11620 , \11473 , \11607 );
or \U$11368 ( \11621 , \11618 , \11619 , \11620 );
and \U$11369 ( \11622 , \11596 , \11600 );
and \U$11370 ( \11623 , \11600 , \11605 );
and \U$11371 ( \11624 , \11596 , \11605 );
or \U$11372 ( \11625 , \11622 , \11623 , \11624 );
and \U$11373 ( \11626 , \11536 , \11545 );
and \U$11374 ( \11627 , \11545 , \11590 );
and \U$11375 ( \11628 , \11536 , \11590 );
or \U$11376 ( \11629 , \11626 , \11627 , \11628 );
xor \U$11377 ( \11630 , \11625 , \11629 );
and \U$11378 ( \11631 , \11505 , \11516 );
and \U$11379 ( \11632 , \11516 , \11531 );
and \U$11380 ( \11633 , \11505 , \11531 );
or \U$11381 ( \11634 , \11631 , \11632 , \11633 );
xor \U$11382 ( \11635 , \11630 , \11634 );
xor \U$11383 ( \11636 , \11621 , \11635 );
and \U$11384 ( \11637 , \11461 , \11465 );
and \U$11385 ( \11638 , \11465 , \11467 );
and \U$11386 ( \11639 , \11461 , \11467 );
or \U$11387 ( \11640 , \11637 , \11638 , \11639 );
and \U$11388 ( \11641 , \11532 , \11591 );
and \U$11389 ( \11642 , \11591 , \11606 );
and \U$11390 ( \11643 , \11532 , \11606 );
or \U$11391 ( \11644 , \11641 , \11642 , \11643 );
xor \U$11392 ( \11645 , \11640 , \11644 );
and \U$11393 ( \11646 , \11550 , \11554 );
and \U$11394 ( \11647 , \11554 , \11559 );
and \U$11395 ( \11648 , \11550 , \11559 );
or \U$11396 ( \11649 , \11646 , \11647 , \11648 );
and \U$11397 ( \11650 , \11494 , \11498 );
and \U$11398 ( \11651 , \11498 , \11503 );
and \U$11399 ( \11652 , \11494 , \11503 );
or \U$11400 ( \11653 , \11650 , \11651 , \11652 );
xor \U$11401 ( \11654 , \11649 , \11653 );
and \U$11402 ( \11655 , \11482 , \11486 );
and \U$11403 ( \11656 , \11486 , \11489 );
and \U$11404 ( \11657 , \11482 , \11489 );
or \U$11405 ( \11658 , \11655 , \11656 , \11657 );
xor \U$11406 ( \11659 , \11654 , \11658 );
and \U$11407 ( \11660 , \6046 , \11539 );
and \U$11408 ( \11661 , \11539 , \11544 );
and \U$11409 ( \11662 , \6046 , \11544 );
or \U$11410 ( \11663 , \11660 , \11661 , \11662 );
and \U$11411 ( \11664 , \11579 , \11583 );
and \U$11412 ( \11665 , \11583 , \11588 );
and \U$11413 ( \11666 , \11579 , \11588 );
or \U$11414 ( \11667 , \11664 , \11665 , \11666 );
xor \U$11415 ( \11668 , \11663 , \11667 );
and \U$11416 ( \11669 , \11564 , \11568 );
and \U$11417 ( \11670 , \11568 , \11573 );
and \U$11418 ( \11671 , \11564 , \11573 );
or \U$11419 ( \11672 , \11669 , \11670 , \11671 );
xor \U$11420 ( \11673 , \11668 , \11672 );
xor \U$11421 ( \11674 , \11659 , \11673 );
and \U$11422 ( \11675 , \11560 , \11574 );
and \U$11423 ( \11676 , \11574 , \11589 );
and \U$11424 ( \11677 , \11560 , \11589 );
or \U$11425 ( \11678 , \11675 , \11676 , \11677 );
and \U$11426 ( \11679 , \5873 , \5829 );
and \U$11427 ( \11680 , \5842 , \5827 );
nor \U$11428 ( \11681 , \11679 , \11680 );
xnor \U$11429 ( \11682 , \11681 , \5836 );
and \U$11430 ( \11683 , \5893 , \5852 );
and \U$11431 ( \11684 , \5861 , \5850 );
nor \U$11432 ( \11685 , \11683 , \11684 );
xnor \U$11433 ( \11686 , \11685 , \5859 );
xor \U$11434 ( \11687 , \11682 , \11686 );
and \U$11435 ( \11688 , \5918 , \5871 );
and \U$11436 ( \11689 , \5881 , \5869 );
nor \U$11437 ( \11690 , \11688 , \11689 );
xnor \U$11438 ( \11691 , \11690 , \5878 );
xor \U$11439 ( \11692 , \11687 , \11691 );
and \U$11440 ( \11693 , \5811 , \5768 );
and \U$11441 ( \11694 , \5780 , \5766 );
nor \U$11442 ( \11695 , \11693 , \11694 );
xnor \U$11443 ( \11696 , \11695 , \5775 );
and \U$11444 ( \11697 , \5831 , \5790 );
and \U$11445 ( \11698 , \5799 , \5788 );
nor \U$11446 ( \11699 , \11697 , \11698 );
xnor \U$11447 ( \11700 , \11699 , \5797 );
xor \U$11448 ( \11701 , \11696 , \11700 );
and \U$11449 ( \11702 , \5854 , \5809 );
and \U$11450 ( \11703 , \5819 , \5807 );
nor \U$11451 ( \11704 , \11702 , \11703 );
xnor \U$11452 ( \11705 , \11704 , \5816 );
xor \U$11453 ( \11706 , \11701 , \11705 );
xor \U$11454 ( \11707 , \11692 , \11706 );
not \U$11455 ( \11708 , \7198 );
and \U$11456 ( \11709 , \5770 , \7203 );
and \U$11457 ( \11710 , \5737 , \7201 );
nor \U$11458 ( \11711 , \11709 , \11710 );
xnor \U$11459 ( \11712 , \11711 , \6824 );
xor \U$11460 ( \11713 , \11708 , \11712 );
and \U$11461 ( \11714 , \5792 , \5750 );
and \U$11462 ( \11715 , \5758 , \5748 );
nor \U$11463 ( \11716 , \11714 , \11715 );
xnor \U$11464 ( \11717 , \11716 , \5755 );
xor \U$11465 ( \11718 , \11713 , \11717 );
xor \U$11466 ( \11719 , \11707 , \11718 );
xor \U$11467 ( \11720 , \11678 , \11719 );
and \U$11468 ( \11721 , \6057 , \6016 );
and \U$11469 ( \11722 , \6029 , \6014 );
nor \U$11470 ( \11723 , \11721 , \11722 );
xnor \U$11471 ( \11724 , \11723 , \6023 );
and \U$11472 ( \11725 , \6065 , \6039 );
and \U$11473 ( \11726 , \6048 , \6037 );
nor \U$11474 ( \11727 , \11725 , \11726 );
xnor \U$11475 ( \11728 , \11727 , \6046 );
xor \U$11476 ( \11729 , \11724 , \11728 );
and \U$11477 ( \11730 , \5998 , \5955 );
and \U$11478 ( \11731 , \5967 , \5953 );
nor \U$11479 ( \11732 , \11730 , \11731 );
xnor \U$11480 ( \11733 , \11732 , \5962 );
and \U$11481 ( \11734 , \6018 , \5977 );
and \U$11482 ( \11735 , \5986 , \5975 );
nor \U$11483 ( \11736 , \11734 , \11735 );
xnor \U$11484 ( \11737 , \11736 , \5984 );
xor \U$11485 ( \11738 , \11733 , \11737 );
and \U$11486 ( \11739 , \6041 , \5996 );
and \U$11487 ( \11740 , \6006 , \5994 );
nor \U$11488 ( \11741 , \11739 , \11740 );
xnor \U$11489 ( \11742 , \11741 , \6003 );
xor \U$11490 ( \11743 , \11738 , \11742 );
xor \U$11491 ( \11744 , \11729 , \11743 );
and \U$11492 ( \11745 , \5937 , \5891 );
and \U$11493 ( \11746 , \5906 , \5889 );
nor \U$11494 ( \11747 , \11745 , \11746 );
xnor \U$11495 ( \11748 , \11747 , \5898 );
and \U$11496 ( \11749 , \5957 , \5916 );
and \U$11497 ( \11750 , \5925 , \5914 );
nor \U$11498 ( \11751 , \11749 , \11750 );
xnor \U$11499 ( \11752 , \11751 , \5923 );
xor \U$11500 ( \11753 , \11748 , \11752 );
and \U$11501 ( \11754 , \5979 , \5935 );
and \U$11502 ( \11755 , \5945 , \5933 );
nor \U$11503 ( \11756 , \11754 , \11755 );
xnor \U$11504 ( \11757 , \11756 , \5942 );
xor \U$11505 ( \11758 , \11753 , \11757 );
xor \U$11506 ( \11759 , \11744 , \11758 );
xor \U$11507 ( \11760 , \11720 , \11759 );
xor \U$11508 ( \11761 , \11674 , \11760 );
and \U$11509 ( \11762 , \11521 , \11525 );
and \U$11510 ( \11763 , \11525 , \11530 );
and \U$11511 ( \11764 , \11521 , \11530 );
or \U$11512 ( \11765 , \11762 , \11763 , \11764 );
and \U$11513 ( \11766 , \11509 , \11513 );
and \U$11514 ( \11767 , \11513 , \11515 );
and \U$11515 ( \11768 , \11509 , \11515 );
or \U$11516 ( \11769 , \11766 , \11767 , \11768 );
xor \U$11517 ( \11770 , \11765 , \11769 );
or \U$11518 ( \11771 , \11490 , \11504 );
xor \U$11519 ( \11772 , \11770 , \11771 );
xor \U$11520 ( \11773 , \11761 , \11772 );
xor \U$11521 ( \11774 , \11645 , \11773 );
xor \U$11522 ( \11775 , \11636 , \11774 );
and \U$11523 ( \11776 , \11457 , \11468 );
and \U$11524 ( \11777 , \11468 , \11608 );
and \U$11525 ( \11778 , \11457 , \11608 );
or \U$11526 ( \11779 , \11776 , \11777 , \11778 );
nor \U$11527 ( \11780 , \11775 , \11779 );
and \U$11528 ( \11781 , \11640 , \11644 );
and \U$11529 ( \11782 , \11644 , \11773 );
and \U$11530 ( \11783 , \11640 , \11773 );
or \U$11531 ( \11784 , \11781 , \11782 , \11783 );
and \U$11532 ( \11785 , \11765 , \11769 );
and \U$11533 ( \11786 , \11769 , \11771 );
and \U$11534 ( \11787 , \11765 , \11771 );
or \U$11535 ( \11788 , \11785 , \11786 , \11787 );
and \U$11536 ( \11789 , \11678 , \11719 );
and \U$11537 ( \11790 , \11719 , \11759 );
and \U$11538 ( \11791 , \11678 , \11759 );
or \U$11539 ( \11792 , \11789 , \11790 , \11791 );
xor \U$11540 ( \11793 , \11788 , \11792 );
and \U$11541 ( \11794 , \11659 , \11673 );
xor \U$11542 ( \11795 , \11793 , \11794 );
xor \U$11543 ( \11796 , \11784 , \11795 );
and \U$11544 ( \11797 , \11625 , \11629 );
and \U$11545 ( \11798 , \11629 , \11634 );
and \U$11546 ( \11799 , \11625 , \11634 );
or \U$11547 ( \11800 , \11797 , \11798 , \11799 );
and \U$11548 ( \11801 , \11674 , \11760 );
and \U$11549 ( \11802 , \11760 , \11772 );
and \U$11550 ( \11803 , \11674 , \11772 );
or \U$11551 ( \11804 , \11801 , \11802 , \11803 );
xor \U$11552 ( \11805 , \11800 , \11804 );
and \U$11553 ( \11806 , \6029 , \6016 );
and \U$11554 ( \11807 , \6041 , \6014 );
nor \U$11555 ( \11808 , \11806 , \11807 );
xnor \U$11556 ( \11809 , \11808 , \6023 );
and \U$11557 ( \11810 , \6048 , \6039 );
and \U$11558 ( \11811 , \6057 , \6037 );
nor \U$11559 ( \11812 , \11810 , \11811 );
xnor \U$11560 ( \11813 , \11812 , \6046 );
xor \U$11561 ( \11814 , \11809 , \11813 );
nand \U$11562 ( \11815 , \6065 , \6053 );
xnor \U$11563 ( \11816 , \11815 , \6062 );
xor \U$11564 ( \11817 , \11814 , \11816 );
and \U$11565 ( \11818 , \5967 , \5955 );
and \U$11566 ( \11819 , \5979 , \5953 );
nor \U$11567 ( \11820 , \11818 , \11819 );
xnor \U$11568 ( \11821 , \11820 , \5962 );
and \U$11569 ( \11822 , \5986 , \5977 );
and \U$11570 ( \11823 , \5998 , \5975 );
nor \U$11571 ( \11824 , \11822 , \11823 );
xnor \U$11572 ( \11825 , \11824 , \5984 );
xor \U$11573 ( \11826 , \11821 , \11825 );
and \U$11574 ( \11827 , \6006 , \5996 );
and \U$11575 ( \11828 , \6018 , \5994 );
nor \U$11576 ( \11829 , \11827 , \11828 );
xnor \U$11577 ( \11830 , \11829 , \6003 );
xor \U$11578 ( \11831 , \11826 , \11830 );
xnor \U$11579 ( \11832 , \11817 , \11831 );
and \U$11580 ( \11833 , \11748 , \11752 );
and \U$11581 ( \11834 , \11752 , \11757 );
and \U$11582 ( \11835 , \11748 , \11757 );
or \U$11583 ( \11836 , \11833 , \11834 , \11835 );
and \U$11584 ( \11837 , \11733 , \11737 );
and \U$11585 ( \11838 , \11737 , \11742 );
and \U$11586 ( \11839 , \11733 , \11742 );
or \U$11587 ( \11840 , \11837 , \11838 , \11839 );
xor \U$11588 ( \11841 , \11836 , \11840 );
and \U$11589 ( \11842 , \11724 , \11728 );
xor \U$11590 ( \11843 , \11841 , \11842 );
xor \U$11591 ( \11844 , \11832 , \11843 );
and \U$11592 ( \11845 , \11708 , \11712 );
and \U$11593 ( \11846 , \11712 , \11717 );
and \U$11594 ( \11847 , \11708 , \11717 );
or \U$11595 ( \11848 , \11845 , \11846 , \11847 );
and \U$11596 ( \11849 , \11696 , \11700 );
and \U$11597 ( \11850 , \11700 , \11705 );
and \U$11598 ( \11851 , \11696 , \11705 );
or \U$11599 ( \11852 , \11849 , \11850 , \11851 );
xor \U$11600 ( \11853 , \11848 , \11852 );
and \U$11601 ( \11854 , \11682 , \11686 );
and \U$11602 ( \11855 , \11686 , \11691 );
and \U$11603 ( \11856 , \11682 , \11691 );
or \U$11604 ( \11857 , \11854 , \11855 , \11856 );
xor \U$11605 ( \11858 , \11853 , \11857 );
xor \U$11606 ( \11859 , \11844 , \11858 );
and \U$11607 ( \11860 , \11692 , \11706 );
and \U$11608 ( \11861 , \11706 , \11718 );
and \U$11609 ( \11862 , \11692 , \11718 );
or \U$11610 ( \11863 , \11860 , \11861 , \11862 );
and \U$11611 ( \11864 , \5737 , \7203 );
not \U$11612 ( \11865 , \11864 );
xnor \U$11613 ( \11866 , \11865 , \6824 );
xor \U$11614 ( \11867 , \6062 , \11866 );
and \U$11615 ( \11868 , \5758 , \5750 );
and \U$11616 ( \11869 , \5770 , \5748 );
nor \U$11617 ( \11870 , \11868 , \11869 );
xnor \U$11618 ( \11871 , \11870 , \5755 );
xor \U$11619 ( \11872 , \11867 , \11871 );
xor \U$11620 ( \11873 , \11863 , \11872 );
and \U$11621 ( \11874 , \5906 , \5891 );
and \U$11622 ( \11875 , \5918 , \5889 );
nor \U$11623 ( \11876 , \11874 , \11875 );
xnor \U$11624 ( \11877 , \11876 , \5898 );
and \U$11625 ( \11878 , \5925 , \5916 );
and \U$11626 ( \11879 , \5937 , \5914 );
nor \U$11627 ( \11880 , \11878 , \11879 );
xnor \U$11628 ( \11881 , \11880 , \5923 );
xor \U$11629 ( \11882 , \11877 , \11881 );
and \U$11630 ( \11883 , \5945 , \5935 );
and \U$11631 ( \11884 , \5957 , \5933 );
nor \U$11632 ( \11885 , \11883 , \11884 );
xnor \U$11633 ( \11886 , \11885 , \5942 );
xor \U$11634 ( \11887 , \11882 , \11886 );
and \U$11635 ( \11888 , \5842 , \5829 );
and \U$11636 ( \11889 , \5854 , \5827 );
nor \U$11637 ( \11890 , \11888 , \11889 );
xnor \U$11638 ( \11891 , \11890 , \5836 );
and \U$11639 ( \11892 , \5861 , \5852 );
and \U$11640 ( \11893 , \5873 , \5850 );
nor \U$11641 ( \11894 , \11892 , \11893 );
xnor \U$11642 ( \11895 , \11894 , \5859 );
xor \U$11643 ( \11896 , \11891 , \11895 );
and \U$11644 ( \11897 , \5881 , \5871 );
and \U$11645 ( \11898 , \5893 , \5869 );
nor \U$11646 ( \11899 , \11897 , \11898 );
xnor \U$11647 ( \11900 , \11899 , \5878 );
xor \U$11648 ( \11901 , \11896 , \11900 );
xor \U$11649 ( \11902 , \11887 , \11901 );
and \U$11650 ( \11903 , \5780 , \5768 );
and \U$11651 ( \11904 , \5792 , \5766 );
nor \U$11652 ( \11905 , \11903 , \11904 );
xnor \U$11653 ( \11906 , \11905 , \5775 );
and \U$11654 ( \11907 , \5799 , \5790 );
and \U$11655 ( \11908 , \5811 , \5788 );
nor \U$11656 ( \11909 , \11907 , \11908 );
xnor \U$11657 ( \11910 , \11909 , \5797 );
xor \U$11658 ( \11911 , \11906 , \11910 );
and \U$11659 ( \11912 , \5819 , \5809 );
and \U$11660 ( \11913 , \5831 , \5807 );
nor \U$11661 ( \11914 , \11912 , \11913 );
xnor \U$11662 ( \11915 , \11914 , \5816 );
xor \U$11663 ( \11916 , \11911 , \11915 );
xor \U$11664 ( \11917 , \11902 , \11916 );
xor \U$11665 ( \11918 , \11873 , \11917 );
xor \U$11666 ( \11919 , \11859 , \11918 );
and \U$11667 ( \11920 , \11663 , \11667 );
and \U$11668 ( \11921 , \11667 , \11672 );
and \U$11669 ( \11922 , \11663 , \11672 );
or \U$11670 ( \11923 , \11920 , \11921 , \11922 );
and \U$11671 ( \11924 , \11649 , \11653 );
and \U$11672 ( \11925 , \11653 , \11658 );
and \U$11673 ( \11926 , \11649 , \11658 );
or \U$11674 ( \11927 , \11924 , \11925 , \11926 );
xor \U$11675 ( \11928 , \11923 , \11927 );
and \U$11676 ( \11929 , \11729 , \11743 );
and \U$11677 ( \11930 , \11743 , \11758 );
and \U$11678 ( \11931 , \11729 , \11758 );
or \U$11679 ( \11932 , \11929 , \11930 , \11931 );
xor \U$11680 ( \11933 , \11928 , \11932 );
xor \U$11681 ( \11934 , \11919 , \11933 );
xor \U$11682 ( \11935 , \11805 , \11934 );
xor \U$11683 ( \11936 , \11796 , \11935 );
and \U$11684 ( \11937 , \11621 , \11635 );
and \U$11685 ( \11938 , \11635 , \11774 );
and \U$11686 ( \11939 , \11621 , \11774 );
or \U$11687 ( \11940 , \11937 , \11938 , \11939 );
nor \U$11688 ( \11941 , \11936 , \11940 );
nor \U$11689 ( \11942 , \11780 , \11941 );
and \U$11690 ( \11943 , \11800 , \11804 );
and \U$11691 ( \11944 , \11804 , \11934 );
and \U$11692 ( \11945 , \11800 , \11934 );
or \U$11693 ( \11946 , \11943 , \11944 , \11945 );
and \U$11694 ( \11947 , \11923 , \11927 );
and \U$11695 ( \11948 , \11927 , \11932 );
and \U$11696 ( \11949 , \11923 , \11932 );
or \U$11697 ( \11950 , \11947 , \11948 , \11949 );
and \U$11698 ( \11951 , \11863 , \11872 );
and \U$11699 ( \11952 , \11872 , \11917 );
and \U$11700 ( \11953 , \11863 , \11917 );
or \U$11701 ( \11954 , \11951 , \11952 , \11953 );
xor \U$11702 ( \11955 , \11950 , \11954 );
and \U$11703 ( \11956 , \11832 , \11843 );
and \U$11704 ( \11957 , \11843 , \11858 );
and \U$11705 ( \11958 , \11832 , \11858 );
or \U$11706 ( \11959 , \11956 , \11957 , \11958 );
xor \U$11707 ( \11960 , \11955 , \11959 );
xor \U$11708 ( \11961 , \11946 , \11960 );
and \U$11709 ( \11962 , \11788 , \11792 );
and \U$11710 ( \11963 , \11792 , \11794 );
and \U$11711 ( \11964 , \11788 , \11794 );
or \U$11712 ( \11965 , \11962 , \11963 , \11964 );
and \U$11713 ( \11966 , \11859 , \11918 );
and \U$11714 ( \11967 , \11918 , \11933 );
and \U$11715 ( \11968 , \11859 , \11933 );
or \U$11716 ( \11969 , \11966 , \11967 , \11968 );
xor \U$11717 ( \11970 , \11965 , \11969 );
and \U$11718 ( \11971 , \11877 , \11881 );
and \U$11719 ( \11972 , \11881 , \11886 );
and \U$11720 ( \11973 , \11877 , \11886 );
or \U$11721 ( \11974 , \11971 , \11972 , \11973 );
and \U$11722 ( \11975 , \11821 , \11825 );
and \U$11723 ( \11976 , \11825 , \11830 );
and \U$11724 ( \11977 , \11821 , \11830 );
or \U$11725 ( \11978 , \11975 , \11976 , \11977 );
xor \U$11726 ( \11979 , \11974 , \11978 );
and \U$11727 ( \11980 , \11809 , \11813 );
and \U$11728 ( \11981 , \11813 , \11816 );
and \U$11729 ( \11982 , \11809 , \11816 );
or \U$11730 ( \11983 , \11980 , \11981 , \11982 );
xor \U$11731 ( \11984 , \11979 , \11983 );
and \U$11732 ( \11985 , \6062 , \11866 );
and \U$11733 ( \11986 , \11866 , \11871 );
and \U$11734 ( \11987 , \6062 , \11871 );
or \U$11735 ( \11988 , \11985 , \11986 , \11987 );
and \U$11736 ( \11989 , \11906 , \11910 );
and \U$11737 ( \11990 , \11910 , \11915 );
and \U$11738 ( \11991 , \11906 , \11915 );
or \U$11739 ( \11992 , \11989 , \11990 , \11991 );
xor \U$11740 ( \11993 , \11988 , \11992 );
and \U$11741 ( \11994 , \11891 , \11895 );
and \U$11742 ( \11995 , \11895 , \11900 );
and \U$11743 ( \11996 , \11891 , \11900 );
or \U$11744 ( \11997 , \11994 , \11995 , \11996 );
xor \U$11745 ( \11998 , \11993 , \11997 );
xor \U$11746 ( \11999 , \11984 , \11998 );
and \U$11747 ( \12000 , \11887 , \11901 );
and \U$11748 ( \12001 , \11901 , \11916 );
and \U$11749 ( \12002 , \11887 , \11916 );
or \U$11750 ( \12003 , \12000 , \12001 , \12002 );
xor \U$11751 ( \12004 , \6858 , \6862 );
xor \U$11752 ( \12005 , \12004 , \6867 );
xor \U$11753 ( \12006 , \6841 , \6845 );
xor \U$11754 ( \12007 , \12006 , \6850 );
xor \U$11755 ( \12008 , \12005 , \12007 );
xor \U$11756 ( \12009 , \6825 , \6829 );
xor \U$11757 ( \12010 , \12009 , \6834 );
xor \U$11758 ( \12011 , \12008 , \12010 );
xor \U$11759 ( \12012 , \12003 , \12011 );
xor \U$11760 ( \12013 , \6910 , \6914 );
xor \U$11761 ( \12014 , \6893 , \6897 );
xor \U$11762 ( \12015 , \12014 , \6902 );
xor \U$11763 ( \12016 , \12013 , \12015 );
xor \U$11764 ( \12017 , \6877 , \6881 );
xor \U$11765 ( \12018 , \12017 , \6886 );
xor \U$11766 ( \12019 , \12016 , \12018 );
xor \U$11767 ( \12020 , \12012 , \12019 );
xor \U$11768 ( \12021 , \11999 , \12020 );
and \U$11769 ( \12022 , \11848 , \11852 );
and \U$11770 ( \12023 , \11852 , \11857 );
and \U$11771 ( \12024 , \11848 , \11857 );
or \U$11772 ( \12025 , \12022 , \12023 , \12024 );
and \U$11773 ( \12026 , \11836 , \11840 );
and \U$11774 ( \12027 , \11840 , \11842 );
and \U$11775 ( \12028 , \11836 , \11842 );
or \U$11776 ( \12029 , \12026 , \12027 , \12028 );
xor \U$11777 ( \12030 , \12025 , \12029 );
or \U$11778 ( \12031 , \11817 , \11831 );
xor \U$11779 ( \12032 , \12030 , \12031 );
xor \U$11780 ( \12033 , \12021 , \12032 );
xor \U$11781 ( \12034 , \11970 , \12033 );
xor \U$11782 ( \12035 , \11961 , \12034 );
and \U$11783 ( \12036 , \11784 , \11795 );
and \U$11784 ( \12037 , \11795 , \11935 );
and \U$11785 ( \12038 , \11784 , \11935 );
or \U$11786 ( \12039 , \12036 , \12037 , \12038 );
nor \U$11787 ( \12040 , \12035 , \12039 );
and \U$11788 ( \12041 , \11965 , \11969 );
and \U$11789 ( \12042 , \11969 , \12033 );
and \U$11790 ( \12043 , \11965 , \12033 );
or \U$11791 ( \12044 , \12041 , \12042 , \12043 );
and \U$11792 ( \12045 , \12025 , \12029 );
and \U$11793 ( \12046 , \12029 , \12031 );
and \U$11794 ( \12047 , \12025 , \12031 );
or \U$11795 ( \12048 , \12045 , \12046 , \12047 );
and \U$11796 ( \12049 , \12003 , \12011 );
and \U$11797 ( \12050 , \12011 , \12019 );
and \U$11798 ( \12051 , \12003 , \12019 );
or \U$11799 ( \12052 , \12049 , \12050 , \12051 );
xor \U$11800 ( \12053 , \12048 , \12052 );
and \U$11801 ( \12054 , \11984 , \11998 );
xor \U$11802 ( \12055 , \12053 , \12054 );
xor \U$11803 ( \12056 , \12044 , \12055 );
and \U$11804 ( \12057 , \11950 , \11954 );
and \U$11805 ( \12058 , \11954 , \11959 );
and \U$11806 ( \12059 , \11950 , \11959 );
or \U$11807 ( \12060 , \12057 , \12058 , \12059 );
and \U$11808 ( \12061 , \11999 , \12020 );
and \U$11809 ( \12062 , \12020 , \12032 );
and \U$11810 ( \12063 , \11999 , \12032 );
or \U$11811 ( \12064 , \12061 , \12062 , \12063 );
xor \U$11812 ( \12065 , \12060 , \12064 );
xnor \U$11813 ( \12066 , \6921 , \6923 );
xor \U$11814 ( \12067 , \6889 , \6905 );
xor \U$11815 ( \12068 , \12067 , \6915 );
xor \U$11816 ( \12069 , \12066 , \12068 );
xor \U$11817 ( \12070 , \6837 , \6853 );
xor \U$11818 ( \12071 , \12070 , \6870 );
xor \U$11819 ( \12072 , \12069 , \12071 );
and \U$11820 ( \12073 , \12005 , \12007 );
and \U$11821 ( \12074 , \12007 , \12010 );
and \U$11822 ( \12075 , \12005 , \12010 );
or \U$11823 ( \12076 , \12073 , \12074 , \12075 );
xor \U$11824 ( \12077 , \5736 , \5756 );
xor \U$11825 ( \12078 , \12077 , \5776 );
xor \U$11826 ( \12079 , \12076 , \12078 );
xor \U$11827 ( \12080 , \6929 , \6931 );
xor \U$11828 ( \12081 , \12080 , \6934 );
xor \U$11829 ( \12082 , \12079 , \12081 );
xor \U$11830 ( \12083 , \12072 , \12082 );
and \U$11831 ( \12084 , \11988 , \11992 );
and \U$11832 ( \12085 , \11992 , \11997 );
and \U$11833 ( \12086 , \11988 , \11997 );
or \U$11834 ( \12087 , \12084 , \12085 , \12086 );
and \U$11835 ( \12088 , \11974 , \11978 );
and \U$11836 ( \12089 , \11978 , \11983 );
and \U$11837 ( \12090 , \11974 , \11983 );
or \U$11838 ( \12091 , \12088 , \12089 , \12090 );
xor \U$11839 ( \12092 , \12087 , \12091 );
and \U$11840 ( \12093 , \12013 , \12015 );
and \U$11841 ( \12094 , \12015 , \12018 );
and \U$11842 ( \12095 , \12013 , \12018 );
or \U$11843 ( \12096 , \12093 , \12094 , \12095 );
xor \U$11844 ( \12097 , \12092 , \12096 );
xor \U$11845 ( \12098 , \12083 , \12097 );
xor \U$11846 ( \12099 , \12065 , \12098 );
xor \U$11847 ( \12100 , \12056 , \12099 );
and \U$11848 ( \12101 , \11946 , \11960 );
and \U$11849 ( \12102 , \11960 , \12034 );
and \U$11850 ( \12103 , \11946 , \12034 );
or \U$11851 ( \12104 , \12101 , \12102 , \12103 );
nor \U$11852 ( \12105 , \12100 , \12104 );
nor \U$11853 ( \12106 , \12040 , \12105 );
nand \U$11854 ( \12107 , \11942 , \12106 );
and \U$11855 ( \12108 , \12060 , \12064 );
and \U$11856 ( \12109 , \12064 , \12098 );
and \U$11857 ( \12110 , \12060 , \12098 );
or \U$11858 ( \12111 , \12108 , \12109 , \12110 );
and \U$11859 ( \12112 , \12087 , \12091 );
and \U$11860 ( \12113 , \12091 , \12096 );
and \U$11861 ( \12114 , \12087 , \12096 );
or \U$11862 ( \12115 , \12112 , \12113 , \12114 );
and \U$11863 ( \12116 , \12076 , \12078 );
and \U$11864 ( \12117 , \12078 , \12081 );
and \U$11865 ( \12118 , \12076 , \12081 );
or \U$11866 ( \12119 , \12116 , \12117 , \12118 );
xor \U$11867 ( \12120 , \12115 , \12119 );
and \U$11868 ( \12121 , \12066 , \12068 );
and \U$11869 ( \12122 , \12068 , \12071 );
and \U$11870 ( \12123 , \12066 , \12071 );
or \U$11871 ( \12124 , \12121 , \12122 , \12123 );
xor \U$11872 ( \12125 , \12120 , \12124 );
xor \U$11873 ( \12126 , \12111 , \12125 );
and \U$11874 ( \12127 , \12048 , \12052 );
and \U$11875 ( \12128 , \12052 , \12054 );
and \U$11876 ( \12129 , \12048 , \12054 );
or \U$11877 ( \12130 , \12127 , \12128 , \12129 );
and \U$11878 ( \12131 , \12072 , \12082 );
and \U$11879 ( \12132 , \12082 , \12097 );
and \U$11880 ( \12133 , \12072 , \12097 );
or \U$11881 ( \12134 , \12131 , \12132 , \12133 );
xor \U$11882 ( \12135 , \12130 , \12134 );
xor \U$11883 ( \12136 , \6948 , \6950 );
xor \U$11884 ( \12137 , \6937 , \6939 );
xor \U$11885 ( \12138 , \12137 , \6942 );
xor \U$11886 ( \12139 , \12136 , \12138 );
xor \U$11887 ( \12140 , \6873 , \6918 );
xor \U$11888 ( \12141 , \12140 , \6924 );
xor \U$11889 ( \12142 , \12139 , \12141 );
xor \U$11890 ( \12143 , \12135 , \12142 );
xor \U$11891 ( \12144 , \12126 , \12143 );
and \U$11892 ( \12145 , \12044 , \12055 );
and \U$11893 ( \12146 , \12055 , \12099 );
and \U$11894 ( \12147 , \12044 , \12099 );
or \U$11895 ( \12148 , \12145 , \12146 , \12147 );
nor \U$11896 ( \12149 , \12144 , \12148 );
and \U$11897 ( \12150 , \12130 , \12134 );
and \U$11898 ( \12151 , \12134 , \12142 );
and \U$11899 ( \12152 , \12130 , \12142 );
or \U$11900 ( \12153 , \12150 , \12151 , \12152 );
xor \U$11901 ( \12154 , \6927 , \6945 );
xor \U$11902 ( \12155 , \12154 , \6951 );
xor \U$11903 ( \12156 , \12153 , \12155 );
and \U$11904 ( \12157 , \12115 , \12119 );
and \U$11905 ( \12158 , \12119 , \12124 );
and \U$11906 ( \12159 , \12115 , \12124 );
or \U$11907 ( \12160 , \12157 , \12158 , \12159 );
and \U$11908 ( \12161 , \12136 , \12138 );
and \U$11909 ( \12162 , \12138 , \12141 );
and \U$11910 ( \12163 , \12136 , \12141 );
or \U$11911 ( \12164 , \12161 , \12162 , \12163 );
xor \U$11912 ( \12165 , \12160 , \12164 );
xor \U$11913 ( \12166 , \6956 , \6958 );
xor \U$11914 ( \12167 , \12166 , \6961 );
xor \U$11915 ( \12168 , \12165 , \12167 );
xor \U$11916 ( \12169 , \12156 , \12168 );
and \U$11917 ( \12170 , \12111 , \12125 );
and \U$11918 ( \12171 , \12125 , \12143 );
and \U$11919 ( \12172 , \12111 , \12143 );
or \U$11920 ( \12173 , \12170 , \12171 , \12172 );
nor \U$11921 ( \12174 , \12169 , \12173 );
nor \U$11922 ( \12175 , \12149 , \12174 );
and \U$11923 ( \12176 , \12160 , \12164 );
and \U$11924 ( \12177 , \12164 , \12167 );
and \U$11925 ( \12178 , \12160 , \12167 );
or \U$11926 ( \12179 , \12176 , \12177 , \12178 );
xor \U$11927 ( \12180 , \6122 , \6284 );
xor \U$11928 ( \12181 , \12180 , \6342 );
xor \U$11929 ( \12182 , \12179 , \12181 );
xor \U$11930 ( \12183 , \6954 , \6964 );
xor \U$11931 ( \12184 , \12183 , \6967 );
xor \U$11932 ( \12185 , \12182 , \12184 );
and \U$11933 ( \12186 , \12153 , \12155 );
and \U$11934 ( \12187 , \12155 , \12168 );
and \U$11935 ( \12188 , \12153 , \12168 );
or \U$11936 ( \12189 , \12186 , \12187 , \12188 );
nor \U$11937 ( \12190 , \12185 , \12189 );
xor \U$11938 ( \12191 , \6970 , \6972 );
xor \U$11939 ( \12192 , \12191 , \6975 );
and \U$11940 ( \12193 , \12179 , \12181 );
and \U$11941 ( \12194 , \12181 , \12184 );
and \U$11942 ( \12195 , \12179 , \12184 );
or \U$11943 ( \12196 , \12193 , \12194 , \12195 );
nor \U$11944 ( \12197 , \12192 , \12196 );
nor \U$11945 ( \12198 , \12190 , \12197 );
nand \U$11946 ( \12199 , \12175 , \12198 );
nor \U$11947 ( \12200 , \12107 , \12199 );
nand \U$11948 ( \12201 , \11617 , \12200 );
nor \U$11949 ( \12202 , \10314 , \12201 );
and \U$11950 ( \12203 , \5945 , \6991 );
and \U$11951 ( \12204 , \5957 , \6988 );
nor \U$11952 ( \12205 , \12203 , \12204 );
xnor \U$11953 ( \12206 , \12205 , \6985 );
and \U$11954 ( \12207 , \7105 , \12206 );
and \U$11955 ( \12208 , \5967 , \7006 );
and \U$11956 ( \12209 , \5979 , \7004 );
nor \U$11957 ( \12210 , \12208 , \12209 );
xnor \U$11958 ( \12211 , \12210 , \7012 );
and \U$11959 ( \12212 , \12206 , \12211 );
and \U$11960 ( \12213 , \7105 , \12211 );
or \U$11961 ( \12214 , \12207 , \12212 , \12213 );
and \U$11962 ( \12215 , \5986 , \7026 );
and \U$11963 ( \12216 , \5998 , \7024 );
nor \U$11964 ( \12217 , \12215 , \12216 );
xnor \U$11965 ( \12218 , \12217 , \7032 );
and \U$11966 ( \12219 , \6006 , \7043 );
and \U$11967 ( \12220 , \6018 , \7041 );
nor \U$11968 ( \12221 , \12219 , \12220 );
xnor \U$11969 ( \12222 , \12221 , \7049 );
and \U$11970 ( \12223 , \12218 , \12222 );
and \U$11971 ( \12224 , \6029 , \7061 );
and \U$11972 ( \12225 , \6041 , \7059 );
nor \U$11973 ( \12226 , \12224 , \12225 );
xnor \U$11974 ( \12227 , \12226 , \7067 );
and \U$11975 ( \12228 , \12222 , \12227 );
and \U$11976 ( \12229 , \12218 , \12227 );
or \U$11977 ( \12230 , \12223 , \12228 , \12229 );
and \U$11978 ( \12231 , \12214 , \12230 );
and \U$11979 ( \12232 , \6065 , \7099 );
and \U$11980 ( \12233 , \6048 , \7097 );
nor \U$11981 ( \12234 , \12232 , \12233 );
xnor \U$11982 ( \12235 , \12234 , \7105 );
and \U$11983 ( \12236 , \12230 , \12235 );
and \U$11984 ( \12237 , \12214 , \12235 );
or \U$11985 ( \12238 , \12231 , \12236 , \12237 );
and \U$11986 ( \12239 , \5967 , \7026 );
and \U$11987 ( \12240 , \5979 , \7024 );
nor \U$11988 ( \12241 , \12239 , \12240 );
xnor \U$11989 ( \12242 , \12241 , \7032 );
and \U$11990 ( \12243 , \5986 , \7043 );
and \U$11991 ( \12244 , \5998 , \7041 );
nor \U$11992 ( \12245 , \12243 , \12244 );
xnor \U$11993 ( \12246 , \12245 , \7049 );
xor \U$11994 ( \12247 , \12242 , \12246 );
and \U$11995 ( \12248 , \6006 , \7061 );
and \U$11996 ( \12249 , \6018 , \7059 );
nor \U$11997 ( \12250 , \12248 , \12249 );
xnor \U$11998 ( \12251 , \12250 , \7067 );
xor \U$11999 ( \12252 , \12247 , \12251 );
and \U$12000 ( \12253 , \5925 , \6991 );
and \U$12001 ( \12254 , \5937 , \6988 );
nor \U$12002 ( \12255 , \12253 , \12254 );
xnor \U$12003 ( \12256 , \12255 , \6985 );
xor \U$12004 ( \12257 , \7123 , \12256 );
and \U$12005 ( \12258 , \5945 , \7006 );
and \U$12006 ( \12259 , \5957 , \7004 );
nor \U$12007 ( \12260 , \12258 , \12259 );
xnor \U$12008 ( \12261 , \12260 , \7012 );
xor \U$12009 ( \12262 , \12257 , \12261 );
xor \U$12010 ( \12263 , \12252 , \12262 );
and \U$12011 ( \12264 , \12238 , \12263 );
and \U$12012 ( \12265 , \5957 , \6991 );
and \U$12013 ( \12266 , \5925 , \6988 );
nor \U$12014 ( \12267 , \12265 , \12266 );
xnor \U$12015 ( \12268 , \12267 , \6985 );
and \U$12016 ( \12269 , \5979 , \7006 );
and \U$12017 ( \12270 , \5945 , \7004 );
nor \U$12018 ( \12271 , \12269 , \12270 );
xnor \U$12019 ( \12272 , \12271 , \7012 );
and \U$12020 ( \12273 , \12268 , \12272 );
and \U$12021 ( \12274 , \5998 , \7026 );
and \U$12022 ( \12275 , \5967 , \7024 );
nor \U$12023 ( \12276 , \12274 , \12275 );
xnor \U$12024 ( \12277 , \12276 , \7032 );
and \U$12025 ( \12278 , \12272 , \12277 );
and \U$12026 ( \12279 , \12268 , \12277 );
or \U$12027 ( \12280 , \12273 , \12278 , \12279 );
and \U$12028 ( \12281 , \6018 , \7043 );
and \U$12029 ( \12282 , \5986 , \7041 );
nor \U$12030 ( \12283 , \12281 , \12282 );
xnor \U$12031 ( \12284 , \12283 , \7049 );
and \U$12032 ( \12285 , \6041 , \7061 );
and \U$12033 ( \12286 , \6006 , \7059 );
nor \U$12034 ( \12287 , \12285 , \12286 );
xnor \U$12035 ( \12288 , \12287 , \7067 );
and \U$12036 ( \12289 , \12284 , \12288 );
and \U$12037 ( \12290 , \6057 , \7082 );
and \U$12038 ( \12291 , \6029 , \7080 );
nor \U$12039 ( \12292 , \12290 , \12291 );
xnor \U$12040 ( \12293 , \12292 , \7088 );
and \U$12041 ( \12294 , \12288 , \12293 );
and \U$12042 ( \12295 , \12284 , \12293 );
or \U$12043 ( \12296 , \12289 , \12294 , \12295 );
xor \U$12044 ( \12297 , \12280 , \12296 );
and \U$12045 ( \12298 , \6029 , \7082 );
and \U$12046 ( \12299 , \6041 , \7080 );
nor \U$12047 ( \12300 , \12298 , \12299 );
xnor \U$12048 ( \12301 , \12300 , \7088 );
and \U$12049 ( \12302 , \6048 , \7099 );
and \U$12050 ( \12303 , \6057 , \7097 );
nor \U$12051 ( \12304 , \12302 , \12303 );
xnor \U$12052 ( \12305 , \12304 , \7105 );
xor \U$12053 ( \12306 , \12301 , \12305 );
nand \U$12054 ( \12307 , \6065 , \7115 );
xnor \U$12055 ( \12308 , \12307 , \7123 );
xor \U$12056 ( \12309 , \12306 , \12308 );
xor \U$12057 ( \12310 , \12297 , \12309 );
and \U$12058 ( \12311 , \12263 , \12310 );
and \U$12059 ( \12312 , \12238 , \12310 );
or \U$12060 ( \12313 , \12264 , \12311 , \12312 );
and \U$12061 ( \12314 , \7123 , \12256 );
and \U$12062 ( \12315 , \12256 , \12261 );
and \U$12063 ( \12316 , \7123 , \12261 );
or \U$12064 ( \12317 , \12314 , \12315 , \12316 );
and \U$12065 ( \12318 , \12242 , \12246 );
and \U$12066 ( \12319 , \12246 , \12251 );
and \U$12067 ( \12320 , \12242 , \12251 );
or \U$12068 ( \12321 , \12318 , \12319 , \12320 );
xor \U$12069 ( \12322 , \12317 , \12321 );
and \U$12070 ( \12323 , \12301 , \12305 );
and \U$12071 ( \12324 , \12305 , \12308 );
and \U$12072 ( \12325 , \12301 , \12308 );
or \U$12073 ( \12326 , \12323 , \12324 , \12325 );
xor \U$12074 ( \12327 , \12322 , \12326 );
xor \U$12075 ( \12328 , \12313 , \12327 );
and \U$12076 ( \12329 , \12280 , \12296 );
and \U$12077 ( \12330 , \12296 , \12309 );
and \U$12078 ( \12331 , \12280 , \12309 );
or \U$12079 ( \12332 , \12329 , \12330 , \12331 );
and \U$12080 ( \12333 , \12252 , \12262 );
xor \U$12081 ( \12334 , \12332 , \12333 );
and \U$12082 ( \12335 , \6057 , \7099 );
and \U$12083 ( \12336 , \6029 , \7097 );
nor \U$12084 ( \12337 , \12335 , \12336 );
xnor \U$12085 ( \12338 , \12337 , \7105 );
and \U$12086 ( \12339 , \6065 , \7117 );
and \U$12087 ( \12340 , \6048 , \7115 );
nor \U$12088 ( \12341 , \12339 , \12340 );
xnor \U$12089 ( \12342 , \12341 , \7123 );
xor \U$12090 ( \12343 , \12338 , \12342 );
and \U$12091 ( \12344 , \5998 , \7043 );
and \U$12092 ( \12345 , \5967 , \7041 );
nor \U$12093 ( \12346 , \12344 , \12345 );
xnor \U$12094 ( \12347 , \12346 , \7049 );
and \U$12095 ( \12348 , \6018 , \7061 );
and \U$12096 ( \12349 , \5986 , \7059 );
nor \U$12097 ( \12350 , \12348 , \12349 );
xnor \U$12098 ( \12351 , \12350 , \7067 );
xor \U$12099 ( \12352 , \12347 , \12351 );
and \U$12100 ( \12353 , \6041 , \7082 );
and \U$12101 ( \12354 , \6006 , \7080 );
nor \U$12102 ( \12355 , \12353 , \12354 );
xnor \U$12103 ( \12356 , \12355 , \7088 );
xor \U$12104 ( \12357 , \12352 , \12356 );
xor \U$12105 ( \12358 , \12343 , \12357 );
and \U$12106 ( \12359 , \5937 , \6991 );
and \U$12107 ( \12360 , \5906 , \6988 );
nor \U$12108 ( \12361 , \12359 , \12360 );
xnor \U$12109 ( \12362 , \12361 , \6985 );
and \U$12110 ( \12363 , \5957 , \7006 );
and \U$12111 ( \12364 , \5925 , \7004 );
nor \U$12112 ( \12365 , \12363 , \12364 );
xnor \U$12113 ( \12366 , \12365 , \7012 );
xor \U$12114 ( \12367 , \12362 , \12366 );
and \U$12115 ( \12368 , \5979 , \7026 );
and \U$12116 ( \12369 , \5945 , \7024 );
nor \U$12117 ( \12370 , \12368 , \12369 );
xnor \U$12118 ( \12371 , \12370 , \7032 );
xor \U$12119 ( \12372 , \12367 , \12371 );
xor \U$12120 ( \12373 , \12358 , \12372 );
xor \U$12121 ( \12374 , \12334 , \12373 );
xor \U$12122 ( \12375 , \12328 , \12374 );
and \U$12123 ( \12376 , \5979 , \6991 );
and \U$12124 ( \12377 , \5945 , \6988 );
nor \U$12125 ( \12378 , \12376 , \12377 );
xnor \U$12126 ( \12379 , \12378 , \6985 );
and \U$12127 ( \12380 , \5998 , \7006 );
and \U$12128 ( \12381 , \5967 , \7004 );
nor \U$12129 ( \12382 , \12380 , \12381 );
xnor \U$12130 ( \12383 , \12382 , \7012 );
and \U$12131 ( \12384 , \12379 , \12383 );
and \U$12132 ( \12385 , \6018 , \7026 );
and \U$12133 ( \12386 , \5986 , \7024 );
nor \U$12134 ( \12387 , \12385 , \12386 );
xnor \U$12135 ( \12388 , \12387 , \7032 );
and \U$12136 ( \12389 , \12383 , \12388 );
and \U$12137 ( \12390 , \12379 , \12388 );
or \U$12138 ( \12391 , \12384 , \12389 , \12390 );
and \U$12139 ( \12392 , \6041 , \7043 );
and \U$12140 ( \12393 , \6006 , \7041 );
nor \U$12141 ( \12394 , \12392 , \12393 );
xnor \U$12142 ( \12395 , \12394 , \7049 );
and \U$12143 ( \12396 , \6057 , \7061 );
and \U$12144 ( \12397 , \6029 , \7059 );
nor \U$12145 ( \12398 , \12396 , \12397 );
xnor \U$12146 ( \12399 , \12398 , \7067 );
and \U$12147 ( \12400 , \12395 , \12399 );
and \U$12148 ( \12401 , \6065 , \7082 );
and \U$12149 ( \12402 , \6048 , \7080 );
nor \U$12150 ( \12403 , \12401 , \12402 );
xnor \U$12151 ( \12404 , \12403 , \7088 );
and \U$12152 ( \12405 , \12399 , \12404 );
and \U$12153 ( \12406 , \12395 , \12404 );
or \U$12154 ( \12407 , \12400 , \12405 , \12406 );
and \U$12155 ( \12408 , \12391 , \12407 );
and \U$12156 ( \12409 , \6048 , \7082 );
and \U$12157 ( \12410 , \6057 , \7080 );
nor \U$12158 ( \12411 , \12409 , \12410 );
xnor \U$12159 ( \12412 , \12411 , \7088 );
and \U$12160 ( \12413 , \12407 , \12412 );
and \U$12161 ( \12414 , \12391 , \12412 );
or \U$12162 ( \12415 , \12408 , \12413 , \12414 );
nand \U$12163 ( \12416 , \6065 , \7097 );
xnor \U$12164 ( \12417 , \12416 , \7105 );
xor \U$12165 ( \12418 , \12218 , \12222 );
xor \U$12166 ( \12419 , \12418 , \12227 );
and \U$12167 ( \12420 , \12417 , \12419 );
xor \U$12168 ( \12421 , \7105 , \12206 );
xor \U$12169 ( \12422 , \12421 , \12211 );
and \U$12170 ( \12423 , \12419 , \12422 );
and \U$12171 ( \12424 , \12417 , \12422 );
or \U$12172 ( \12425 , \12420 , \12423 , \12424 );
and \U$12173 ( \12426 , \12415 , \12425 );
xor \U$12174 ( \12427 , \12284 , \12288 );
xor \U$12175 ( \12428 , \12427 , \12293 );
and \U$12176 ( \12429 , \12425 , \12428 );
and \U$12177 ( \12430 , \12415 , \12428 );
or \U$12178 ( \12431 , \12426 , \12429 , \12430 );
xor \U$12179 ( \12432 , \12268 , \12272 );
xor \U$12180 ( \12433 , \12432 , \12277 );
xor \U$12181 ( \12434 , \12214 , \12230 );
xor \U$12182 ( \12435 , \12434 , \12235 );
and \U$12183 ( \12436 , \12433 , \12435 );
and \U$12184 ( \12437 , \12431 , \12436 );
xor \U$12185 ( \12438 , \12238 , \12263 );
xor \U$12186 ( \12439 , \12438 , \12310 );
and \U$12187 ( \12440 , \12436 , \12439 );
and \U$12188 ( \12441 , \12431 , \12439 );
or \U$12189 ( \12442 , \12437 , \12440 , \12441 );
nor \U$12190 ( \12443 , \12375 , \12442 );
and \U$12191 ( \12444 , \12332 , \12333 );
and \U$12192 ( \12445 , \12333 , \12373 );
and \U$12193 ( \12446 , \12332 , \12373 );
or \U$12194 ( \12447 , \12444 , \12445 , \12446 );
nand \U$12195 ( \12448 , \6065 , \7138 );
xnor \U$12196 ( \12449 , \12448 , \7146 );
and \U$12197 ( \12450 , \6006 , \7082 );
and \U$12198 ( \12451 , \6018 , \7080 );
nor \U$12199 ( \12452 , \12450 , \12451 );
xnor \U$12200 ( \12453 , \12452 , \7088 );
and \U$12201 ( \12454 , \6029 , \7099 );
and \U$12202 ( \12455 , \6041 , \7097 );
nor \U$12203 ( \12456 , \12454 , \12455 );
xnor \U$12204 ( \12457 , \12456 , \7105 );
xor \U$12205 ( \12458 , \12453 , \12457 );
and \U$12206 ( \12459 , \6048 , \7117 );
and \U$12207 ( \12460 , \6057 , \7115 );
nor \U$12208 ( \12461 , \12459 , \12460 );
xnor \U$12209 ( \12462 , \12461 , \7123 );
xor \U$12210 ( \12463 , \12458 , \12462 );
xor \U$12211 ( \12464 , \12449 , \12463 );
and \U$12212 ( \12465 , \5945 , \7026 );
and \U$12213 ( \12466 , \5957 , \7024 );
nor \U$12214 ( \12467 , \12465 , \12466 );
xnor \U$12215 ( \12468 , \12467 , \7032 );
and \U$12216 ( \12469 , \5967 , \7043 );
and \U$12217 ( \12470 , \5979 , \7041 );
nor \U$12218 ( \12471 , \12469 , \12470 );
xnor \U$12219 ( \12472 , \12471 , \7049 );
xor \U$12220 ( \12473 , \12468 , \12472 );
and \U$12221 ( \12474 , \5986 , \7061 );
and \U$12222 ( \12475 , \5998 , \7059 );
nor \U$12223 ( \12476 , \12474 , \12475 );
xnor \U$12224 ( \12477 , \12476 , \7067 );
xor \U$12225 ( \12478 , \12473 , \12477 );
xor \U$12226 ( \12479 , \12464 , \12478 );
and \U$12227 ( \12480 , \12362 , \12366 );
and \U$12228 ( \12481 , \12366 , \12371 );
and \U$12229 ( \12482 , \12362 , \12371 );
or \U$12230 ( \12483 , \12480 , \12481 , \12482 );
and \U$12231 ( \12484 , \12347 , \12351 );
and \U$12232 ( \12485 , \12351 , \12356 );
and \U$12233 ( \12486 , \12347 , \12356 );
or \U$12234 ( \12487 , \12484 , \12485 , \12486 );
xor \U$12235 ( \12488 , \12483 , \12487 );
and \U$12236 ( \12489 , \12338 , \12342 );
xor \U$12237 ( \12490 , \12488 , \12489 );
xor \U$12238 ( \12491 , \12479 , \12490 );
xor \U$12239 ( \12492 , \12447 , \12491 );
and \U$12240 ( \12493 , \12317 , \12321 );
and \U$12241 ( \12494 , \12321 , \12326 );
and \U$12242 ( \12495 , \12317 , \12326 );
or \U$12243 ( \12496 , \12493 , \12494 , \12495 );
and \U$12244 ( \12497 , \12343 , \12357 );
and \U$12245 ( \12498 , \12357 , \12372 );
and \U$12246 ( \12499 , \12343 , \12372 );
or \U$12247 ( \12500 , \12497 , \12498 , \12499 );
xor \U$12248 ( \12501 , \12496 , \12500 );
and \U$12249 ( \12502 , \5906 , \6991 );
and \U$12250 ( \12503 , \5918 , \6988 );
nor \U$12251 ( \12504 , \12502 , \12503 );
xnor \U$12252 ( \12505 , \12504 , \6985 );
xor \U$12253 ( \12506 , \7146 , \12505 );
and \U$12254 ( \12507 , \5925 , \7006 );
and \U$12255 ( \12508 , \5937 , \7004 );
nor \U$12256 ( \12509 , \12507 , \12508 );
xnor \U$12257 ( \12510 , \12509 , \7012 );
xor \U$12258 ( \12511 , \12506 , \12510 );
xor \U$12259 ( \12512 , \12501 , \12511 );
xor \U$12260 ( \12513 , \12492 , \12512 );
and \U$12261 ( \12514 , \12313 , \12327 );
and \U$12262 ( \12515 , \12327 , \12374 );
and \U$12263 ( \12516 , \12313 , \12374 );
or \U$12264 ( \12517 , \12514 , \12515 , \12516 );
nor \U$12265 ( \12518 , \12513 , \12517 );
nor \U$12266 ( \12519 , \12443 , \12518 );
and \U$12267 ( \12520 , \12483 , \12487 );
and \U$12268 ( \12521 , \12487 , \12489 );
and \U$12269 ( \12522 , \12483 , \12489 );
or \U$12270 ( \12523 , \12520 , \12521 , \12522 );
and \U$12271 ( \12524 , \12449 , \12463 );
and \U$12272 ( \12525 , \12463 , \12478 );
and \U$12273 ( \12526 , \12449 , \12478 );
or \U$12274 ( \12527 , \12524 , \12525 , \12526 );
xor \U$12275 ( \12528 , \12523 , \12527 );
and \U$12276 ( \12529 , \6041 , \7099 );
and \U$12277 ( \12530 , \6006 , \7097 );
nor \U$12278 ( \12531 , \12529 , \12530 );
xnor \U$12279 ( \12532 , \12531 , \7105 );
and \U$12280 ( \12533 , \6057 , \7117 );
and \U$12281 ( \12534 , \6029 , \7115 );
nor \U$12282 ( \12535 , \12533 , \12534 );
xnor \U$12283 ( \12536 , \12535 , \7123 );
xor \U$12284 ( \12537 , \12532 , \12536 );
and \U$12285 ( \12538 , \6065 , \7140 );
and \U$12286 ( \12539 , \6048 , \7138 );
nor \U$12287 ( \12540 , \12538 , \12539 );
xnor \U$12288 ( \12541 , \12540 , \7146 );
xor \U$12289 ( \12542 , \12537 , \12541 );
and \U$12290 ( \12543 , \5979 , \7043 );
and \U$12291 ( \12544 , \5945 , \7041 );
nor \U$12292 ( \12545 , \12543 , \12544 );
xnor \U$12293 ( \12546 , \12545 , \7049 );
and \U$12294 ( \12547 , \5998 , \7061 );
and \U$12295 ( \12548 , \5967 , \7059 );
nor \U$12296 ( \12549 , \12547 , \12548 );
xnor \U$12297 ( \12550 , \12549 , \7067 );
xor \U$12298 ( \12551 , \12546 , \12550 );
and \U$12299 ( \12552 , \6018 , \7082 );
and \U$12300 ( \12553 , \5986 , \7080 );
nor \U$12301 ( \12554 , \12552 , \12553 );
xnor \U$12302 ( \12555 , \12554 , \7088 );
xor \U$12303 ( \12556 , \12551 , \12555 );
xor \U$12304 ( \12557 , \12542 , \12556 );
and \U$12305 ( \12558 , \5918 , \6991 );
and \U$12306 ( \12559 , \5881 , \6988 );
nor \U$12307 ( \12560 , \12558 , \12559 );
xnor \U$12308 ( \12561 , \12560 , \6985 );
and \U$12309 ( \12562 , \5937 , \7006 );
and \U$12310 ( \12563 , \5906 , \7004 );
nor \U$12311 ( \12564 , \12562 , \12563 );
xnor \U$12312 ( \12565 , \12564 , \7012 );
xor \U$12313 ( \12566 , \12561 , \12565 );
and \U$12314 ( \12567 , \5957 , \7026 );
and \U$12315 ( \12568 , \5925 , \7024 );
nor \U$12316 ( \12569 , \12567 , \12568 );
xnor \U$12317 ( \12570 , \12569 , \7032 );
xor \U$12318 ( \12571 , \12566 , \12570 );
xor \U$12319 ( \12572 , \12557 , \12571 );
xor \U$12320 ( \12573 , \12528 , \12572 );
and \U$12321 ( \12574 , \12496 , \12500 );
and \U$12322 ( \12575 , \12500 , \12511 );
and \U$12323 ( \12576 , \12496 , \12511 );
or \U$12324 ( \12577 , \12574 , \12575 , \12576 );
and \U$12325 ( \12578 , \12479 , \12490 );
xor \U$12326 ( \12579 , \12577 , \12578 );
and \U$12327 ( \12580 , \7146 , \12505 );
and \U$12328 ( \12581 , \12505 , \12510 );
and \U$12329 ( \12582 , \7146 , \12510 );
or \U$12330 ( \12583 , \12580 , \12581 , \12582 );
and \U$12331 ( \12584 , \12468 , \12472 );
and \U$12332 ( \12585 , \12472 , \12477 );
and \U$12333 ( \12586 , \12468 , \12477 );
or \U$12334 ( \12587 , \12584 , \12585 , \12586 );
xor \U$12335 ( \12588 , \12583 , \12587 );
and \U$12336 ( \12589 , \12453 , \12457 );
and \U$12337 ( \12590 , \12457 , \12462 );
and \U$12338 ( \12591 , \12453 , \12462 );
or \U$12339 ( \12592 , \12589 , \12590 , \12591 );
xor \U$12340 ( \12593 , \12588 , \12592 );
xor \U$12341 ( \12594 , \12579 , \12593 );
xor \U$12342 ( \12595 , \12573 , \12594 );
and \U$12343 ( \12596 , \12447 , \12491 );
and \U$12344 ( \12597 , \12491 , \12512 );
and \U$12345 ( \12598 , \12447 , \12512 );
or \U$12346 ( \12599 , \12596 , \12597 , \12598 );
nor \U$12347 ( \12600 , \12595 , \12599 );
and \U$12348 ( \12601 , \12577 , \12578 );
and \U$12349 ( \12602 , \12578 , \12593 );
and \U$12350 ( \12603 , \12577 , \12593 );
or \U$12351 ( \12604 , \12601 , \12602 , \12603 );
and \U$12352 ( \12605 , \12523 , \12527 );
and \U$12353 ( \12606 , \12527 , \12572 );
and \U$12354 ( \12607 , \12523 , \12572 );
or \U$12355 ( \12608 , \12605 , \12606 , \12607 );
and \U$12356 ( \12609 , \5881 , \6991 );
and \U$12357 ( \12610 , \5893 , \6988 );
nor \U$12358 ( \12611 , \12609 , \12610 );
xnor \U$12359 ( \12612 , \12611 , \6985 );
xor \U$12360 ( \12613 , \7163 , \12612 );
and \U$12361 ( \12614 , \5906 , \7006 );
and \U$12362 ( \12615 , \5918 , \7004 );
nor \U$12363 ( \12616 , \12614 , \12615 );
xnor \U$12364 ( \12617 , \12616 , \7012 );
xor \U$12365 ( \12618 , \12613 , \12617 );
and \U$12366 ( \12619 , \6048 , \7140 );
and \U$12367 ( \12620 , \6057 , \7138 );
nor \U$12368 ( \12621 , \12619 , \12620 );
xnor \U$12369 ( \12622 , \12621 , \7146 );
nand \U$12370 ( \12623 , \6065 , \7155 );
xnor \U$12371 ( \12624 , \12623 , \7163 );
xor \U$12372 ( \12625 , \12622 , \12624 );
and \U$12373 ( \12626 , \5986 , \7082 );
and \U$12374 ( \12627 , \5998 , \7080 );
nor \U$12375 ( \12628 , \12626 , \12627 );
xnor \U$12376 ( \12629 , \12628 , \7088 );
and \U$12377 ( \12630 , \6006 , \7099 );
and \U$12378 ( \12631 , \6018 , \7097 );
nor \U$12379 ( \12632 , \12630 , \12631 );
xnor \U$12380 ( \12633 , \12632 , \7105 );
xor \U$12381 ( \12634 , \12629 , \12633 );
and \U$12382 ( \12635 , \6029 , \7117 );
and \U$12383 ( \12636 , \6041 , \7115 );
nor \U$12384 ( \12637 , \12635 , \12636 );
xnor \U$12385 ( \12638 , \12637 , \7123 );
xor \U$12386 ( \12639 , \12634 , \12638 );
xor \U$12387 ( \12640 , \12625 , \12639 );
xor \U$12388 ( \12641 , \12618 , \12640 );
and \U$12389 ( \12642 , \12561 , \12565 );
and \U$12390 ( \12643 , \12565 , \12570 );
and \U$12391 ( \12644 , \12561 , \12570 );
or \U$12392 ( \12645 , \12642 , \12643 , \12644 );
and \U$12393 ( \12646 , \12546 , \12550 );
and \U$12394 ( \12647 , \12550 , \12555 );
and \U$12395 ( \12648 , \12546 , \12555 );
or \U$12396 ( \12649 , \12646 , \12647 , \12648 );
xor \U$12397 ( \12650 , \12645 , \12649 );
and \U$12398 ( \12651 , \12532 , \12536 );
and \U$12399 ( \12652 , \12536 , \12541 );
and \U$12400 ( \12653 , \12532 , \12541 );
or \U$12401 ( \12654 , \12651 , \12652 , \12653 );
xor \U$12402 ( \12655 , \12650 , \12654 );
xor \U$12403 ( \12656 , \12641 , \12655 );
xor \U$12404 ( \12657 , \12608 , \12656 );
and \U$12405 ( \12658 , \12583 , \12587 );
and \U$12406 ( \12659 , \12587 , \12592 );
and \U$12407 ( \12660 , \12583 , \12592 );
or \U$12408 ( \12661 , \12658 , \12659 , \12660 );
and \U$12409 ( \12662 , \12542 , \12556 );
and \U$12410 ( \12663 , \12556 , \12571 );
and \U$12411 ( \12664 , \12542 , \12571 );
or \U$12412 ( \12665 , \12662 , \12663 , \12664 );
xor \U$12413 ( \12666 , \12661 , \12665 );
and \U$12414 ( \12667 , \5925 , \7026 );
and \U$12415 ( \12668 , \5937 , \7024 );
nor \U$12416 ( \12669 , \12667 , \12668 );
xnor \U$12417 ( \12670 , \12669 , \7032 );
and \U$12418 ( \12671 , \5945 , \7043 );
and \U$12419 ( \12672 , \5957 , \7041 );
nor \U$12420 ( \12673 , \12671 , \12672 );
xnor \U$12421 ( \12674 , \12673 , \7049 );
xor \U$12422 ( \12675 , \12670 , \12674 );
and \U$12423 ( \12676 , \5967 , \7061 );
and \U$12424 ( \12677 , \5979 , \7059 );
nor \U$12425 ( \12678 , \12676 , \12677 );
xnor \U$12426 ( \12679 , \12678 , \7067 );
xor \U$12427 ( \12680 , \12675 , \12679 );
xor \U$12428 ( \12681 , \12666 , \12680 );
xor \U$12429 ( \12682 , \12657 , \12681 );
xor \U$12430 ( \12683 , \12604 , \12682 );
and \U$12431 ( \12684 , \12573 , \12594 );
nor \U$12432 ( \12685 , \12683 , \12684 );
nor \U$12433 ( \12686 , \12600 , \12685 );
nand \U$12434 ( \12687 , \12519 , \12686 );
and \U$12435 ( \12688 , \12608 , \12656 );
and \U$12436 ( \12689 , \12656 , \12681 );
and \U$12437 ( \12690 , \12608 , \12681 );
or \U$12438 ( \12691 , \12688 , \12689 , \12690 );
and \U$12439 ( \12692 , \7163 , \12612 );
and \U$12440 ( \12693 , \12612 , \12617 );
and \U$12441 ( \12694 , \7163 , \12617 );
or \U$12442 ( \12695 , \12692 , \12693 , \12694 );
and \U$12443 ( \12696 , \12670 , \12674 );
and \U$12444 ( \12697 , \12674 , \12679 );
and \U$12445 ( \12698 , \12670 , \12679 );
or \U$12446 ( \12699 , \12696 , \12697 , \12698 );
xor \U$12447 ( \12700 , \12695 , \12699 );
and \U$12448 ( \12701 , \12629 , \12633 );
and \U$12449 ( \12702 , \12633 , \12638 );
and \U$12450 ( \12703 , \12629 , \12638 );
or \U$12451 ( \12704 , \12701 , \12702 , \12703 );
xor \U$12452 ( \12705 , \12700 , \12704 );
and \U$12453 ( \12706 , \12645 , \12649 );
and \U$12454 ( \12707 , \12649 , \12654 );
and \U$12455 ( \12708 , \12645 , \12654 );
or \U$12456 ( \12709 , \12706 , \12707 , \12708 );
and \U$12457 ( \12710 , \12622 , \12624 );
and \U$12458 ( \12711 , \12624 , \12639 );
and \U$12459 ( \12712 , \12622 , \12639 );
or \U$12460 ( \12713 , \12710 , \12711 , \12712 );
xor \U$12461 ( \12714 , \12709 , \12713 );
and \U$12462 ( \12715 , \5893 , \6991 );
and \U$12463 ( \12716 , \5861 , \6988 );
nor \U$12464 ( \12717 , \12715 , \12716 );
xnor \U$12465 ( \12718 , \12717 , \6985 );
and \U$12466 ( \12719 , \5918 , \7006 );
and \U$12467 ( \12720 , \5881 , \7004 );
nor \U$12468 ( \12721 , \12719 , \12720 );
xnor \U$12469 ( \12722 , \12721 , \7012 );
xor \U$12470 ( \12723 , \12718 , \12722 );
and \U$12471 ( \12724 , \5937 , \7026 );
and \U$12472 ( \12725 , \5906 , \7024 );
nor \U$12473 ( \12726 , \12724 , \12725 );
xnor \U$12474 ( \12727 , \12726 , \7032 );
xor \U$12475 ( \12728 , \12723 , \12727 );
xor \U$12476 ( \12729 , \12714 , \12728 );
xor \U$12477 ( \12730 , \12705 , \12729 );
xor \U$12478 ( \12731 , \12691 , \12730 );
and \U$12479 ( \12732 , \12661 , \12665 );
and \U$12480 ( \12733 , \12665 , \12680 );
and \U$12481 ( \12734 , \12661 , \12680 );
or \U$12482 ( \12735 , \12732 , \12733 , \12734 );
and \U$12483 ( \12736 , \12618 , \12640 );
and \U$12484 ( \12737 , \12640 , \12655 );
and \U$12485 ( \12738 , \12618 , \12655 );
or \U$12486 ( \12739 , \12736 , \12737 , \12738 );
xor \U$12487 ( \12740 , \12735 , \12739 );
and \U$12488 ( \12741 , \6065 , \7157 );
and \U$12489 ( \12742 , \6048 , \7155 );
nor \U$12490 ( \12743 , \12741 , \12742 );
xnor \U$12491 ( \12744 , \12743 , \7163 );
and \U$12492 ( \12745 , \6018 , \7099 );
and \U$12493 ( \12746 , \5986 , \7097 );
nor \U$12494 ( \12747 , \12745 , \12746 );
xnor \U$12495 ( \12748 , \12747 , \7105 );
and \U$12496 ( \12749 , \6041 , \7117 );
and \U$12497 ( \12750 , \6006 , \7115 );
nor \U$12498 ( \12751 , \12749 , \12750 );
xnor \U$12499 ( \12752 , \12751 , \7123 );
xor \U$12500 ( \12753 , \12748 , \12752 );
and \U$12501 ( \12754 , \6057 , \7140 );
and \U$12502 ( \12755 , \6029 , \7138 );
nor \U$12503 ( \12756 , \12754 , \12755 );
xnor \U$12504 ( \12757 , \12756 , \7146 );
xor \U$12505 ( \12758 , \12753 , \12757 );
xor \U$12506 ( \12759 , \12744 , \12758 );
and \U$12507 ( \12760 , \5957 , \7043 );
and \U$12508 ( \12761 , \5925 , \7041 );
nor \U$12509 ( \12762 , \12760 , \12761 );
xnor \U$12510 ( \12763 , \12762 , \7049 );
and \U$12511 ( \12764 , \5979 , \7061 );
and \U$12512 ( \12765 , \5945 , \7059 );
nor \U$12513 ( \12766 , \12764 , \12765 );
xnor \U$12514 ( \12767 , \12766 , \7067 );
xor \U$12515 ( \12768 , \12763 , \12767 );
and \U$12516 ( \12769 , \5998 , \7082 );
and \U$12517 ( \12770 , \5967 , \7080 );
nor \U$12518 ( \12771 , \12769 , \12770 );
xnor \U$12519 ( \12772 , \12771 , \7088 );
xor \U$12520 ( \12773 , \12768 , \12772 );
xor \U$12521 ( \12774 , \12759 , \12773 );
xor \U$12522 ( \12775 , \12740 , \12774 );
xor \U$12523 ( \12776 , \12731 , \12775 );
and \U$12524 ( \12777 , \12604 , \12682 );
nor \U$12525 ( \12778 , \12776 , \12777 );
and \U$12526 ( \12779 , \12735 , \12739 );
and \U$12527 ( \12780 , \12739 , \12774 );
and \U$12528 ( \12781 , \12735 , \12774 );
or \U$12529 ( \12782 , \12779 , \12780 , \12781 );
and \U$12530 ( \12783 , \12705 , \12729 );
xor \U$12531 ( \12784 , \12782 , \12783 );
and \U$12532 ( \12785 , \12709 , \12713 );
and \U$12533 ( \12786 , \12713 , \12728 );
and \U$12534 ( \12787 , \12709 , \12728 );
or \U$12535 ( \12788 , \12785 , \12786 , \12787 );
and \U$12536 ( \12789 , \6029 , \7140 );
and \U$12537 ( \12790 , \6041 , \7138 );
nor \U$12538 ( \12791 , \12789 , \12790 );
xnor \U$12539 ( \12792 , \12791 , \7146 );
and \U$12540 ( \12793 , \6048 , \7157 );
and \U$12541 ( \12794 , \6057 , \7155 );
nor \U$12542 ( \12795 , \12793 , \12794 );
xnor \U$12543 ( \12796 , \12795 , \7163 );
xor \U$12544 ( \12797 , \12792 , \12796 );
nand \U$12545 ( \12798 , \6065 , \7173 );
xnor \U$12546 ( \12799 , \12798 , \7181 );
xor \U$12547 ( \12800 , \12797 , \12799 );
and \U$12548 ( \12801 , \5967 , \7082 );
and \U$12549 ( \12802 , \5979 , \7080 );
nor \U$12550 ( \12803 , \12801 , \12802 );
xnor \U$12551 ( \12804 , \12803 , \7088 );
and \U$12552 ( \12805 , \5986 , \7099 );
and \U$12553 ( \12806 , \5998 , \7097 );
nor \U$12554 ( \12807 , \12805 , \12806 );
xnor \U$12555 ( \12808 , \12807 , \7105 );
xor \U$12556 ( \12809 , \12804 , \12808 );
and \U$12557 ( \12810 , \6006 , \7117 );
and \U$12558 ( \12811 , \6018 , \7115 );
nor \U$12559 ( \12812 , \12810 , \12811 );
xnor \U$12560 ( \12813 , \12812 , \7123 );
xor \U$12561 ( \12814 , \12809 , \12813 );
xor \U$12562 ( \12815 , \12800 , \12814 );
and \U$12563 ( \12816 , \5906 , \7026 );
and \U$12564 ( \12817 , \5918 , \7024 );
nor \U$12565 ( \12818 , \12816 , \12817 );
xnor \U$12566 ( \12819 , \12818 , \7032 );
and \U$12567 ( \12820 , \5925 , \7043 );
and \U$12568 ( \12821 , \5937 , \7041 );
nor \U$12569 ( \12822 , \12820 , \12821 );
xnor \U$12570 ( \12823 , \12822 , \7049 );
xor \U$12571 ( \12824 , \12819 , \12823 );
and \U$12572 ( \12825 , \5945 , \7061 );
and \U$12573 ( \12826 , \5957 , \7059 );
nor \U$12574 ( \12827 , \12825 , \12826 );
xnor \U$12575 ( \12828 , \12827 , \7067 );
xor \U$12576 ( \12829 , \12824 , \12828 );
xor \U$12577 ( \12830 , \12815 , \12829 );
and \U$12578 ( \12831 , \12718 , \12722 );
and \U$12579 ( \12832 , \12722 , \12727 );
and \U$12580 ( \12833 , \12718 , \12727 );
or \U$12581 ( \12834 , \12831 , \12832 , \12833 );
and \U$12582 ( \12835 , \12763 , \12767 );
and \U$12583 ( \12836 , \12767 , \12772 );
and \U$12584 ( \12837 , \12763 , \12772 );
or \U$12585 ( \12838 , \12835 , \12836 , \12837 );
xor \U$12586 ( \12839 , \12834 , \12838 );
and \U$12587 ( \12840 , \12748 , \12752 );
and \U$12588 ( \12841 , \12752 , \12757 );
and \U$12589 ( \12842 , \12748 , \12757 );
or \U$12590 ( \12843 , \12840 , \12841 , \12842 );
xor \U$12591 ( \12844 , \12839 , \12843 );
xor \U$12592 ( \12845 , \12830 , \12844 );
xor \U$12593 ( \12846 , \12788 , \12845 );
and \U$12594 ( \12847 , \12695 , \12699 );
and \U$12595 ( \12848 , \12699 , \12704 );
and \U$12596 ( \12849 , \12695 , \12704 );
or \U$12597 ( \12850 , \12847 , \12848 , \12849 );
and \U$12598 ( \12851 , \12744 , \12758 );
and \U$12599 ( \12852 , \12758 , \12773 );
and \U$12600 ( \12853 , \12744 , \12773 );
or \U$12601 ( \12854 , \12851 , \12852 , \12853 );
xor \U$12602 ( \12855 , \12850 , \12854 );
and \U$12603 ( \12856 , \5861 , \6991 );
and \U$12604 ( \12857 , \5873 , \6988 );
nor \U$12605 ( \12858 , \12856 , \12857 );
xnor \U$12606 ( \12859 , \12858 , \6985 );
xor \U$12607 ( \12860 , \7181 , \12859 );
and \U$12608 ( \12861 , \5881 , \7006 );
and \U$12609 ( \12862 , \5893 , \7004 );
nor \U$12610 ( \12863 , \12861 , \12862 );
xnor \U$12611 ( \12864 , \12863 , \7012 );
xor \U$12612 ( \12865 , \12860 , \12864 );
xor \U$12613 ( \12866 , \12855 , \12865 );
xor \U$12614 ( \12867 , \12846 , \12866 );
xor \U$12615 ( \12868 , \12784 , \12867 );
and \U$12616 ( \12869 , \12691 , \12730 );
and \U$12617 ( \12870 , \12730 , \12775 );
and \U$12618 ( \12871 , \12691 , \12775 );
or \U$12619 ( \12872 , \12869 , \12870 , \12871 );
nor \U$12620 ( \12873 , \12868 , \12872 );
nor \U$12621 ( \12874 , \12778 , \12873 );
and \U$12622 ( \12875 , \12788 , \12845 );
and \U$12623 ( \12876 , \12845 , \12866 );
and \U$12624 ( \12877 , \12788 , \12866 );
or \U$12625 ( \12878 , \12875 , \12876 , \12877 );
and \U$12626 ( \12879 , \7181 , \12859 );
and \U$12627 ( \12880 , \12859 , \12864 );
and \U$12628 ( \12881 , \7181 , \12864 );
or \U$12629 ( \12882 , \12879 , \12880 , \12881 );
and \U$12630 ( \12883 , \12819 , \12823 );
and \U$12631 ( \12884 , \12823 , \12828 );
and \U$12632 ( \12885 , \12819 , \12828 );
or \U$12633 ( \12886 , \12883 , \12884 , \12885 );
xor \U$12634 ( \12887 , \12882 , \12886 );
and \U$12635 ( \12888 , \12804 , \12808 );
and \U$12636 ( \12889 , \12808 , \12813 );
and \U$12637 ( \12890 , \12804 , \12813 );
or \U$12638 ( \12891 , \12888 , \12889 , \12890 );
xor \U$12639 ( \12892 , \12887 , \12891 );
and \U$12640 ( \12893 , \12834 , \12838 );
and \U$12641 ( \12894 , \12838 , \12843 );
and \U$12642 ( \12895 , \12834 , \12843 );
or \U$12643 ( \12896 , \12893 , \12894 , \12895 );
and \U$12644 ( \12897 , \12800 , \12814 );
and \U$12645 ( \12898 , \12814 , \12829 );
and \U$12646 ( \12899 , \12800 , \12829 );
or \U$12647 ( \12900 , \12897 , \12898 , \12899 );
xor \U$12648 ( \12901 , \12896 , \12900 );
and \U$12649 ( \12902 , \5998 , \7099 );
and \U$12650 ( \12903 , \5967 , \7097 );
nor \U$12651 ( \12904 , \12902 , \12903 );
xnor \U$12652 ( \12905 , \12904 , \7105 );
and \U$12653 ( \12906 , \6018 , \7117 );
and \U$12654 ( \12907 , \5986 , \7115 );
nor \U$12655 ( \12908 , \12906 , \12907 );
xnor \U$12656 ( \12909 , \12908 , \7123 );
xor \U$12657 ( \12910 , \12905 , \12909 );
and \U$12658 ( \12911 , \6041 , \7140 );
and \U$12659 ( \12912 , \6006 , \7138 );
nor \U$12660 ( \12913 , \12911 , \12912 );
xnor \U$12661 ( \12914 , \12913 , \7146 );
xor \U$12662 ( \12915 , \12910 , \12914 );
and \U$12663 ( \12916 , \5937 , \7043 );
and \U$12664 ( \12917 , \5906 , \7041 );
nor \U$12665 ( \12918 , \12916 , \12917 );
xnor \U$12666 ( \12919 , \12918 , \7049 );
and \U$12667 ( \12920 , \5957 , \7061 );
and \U$12668 ( \12921 , \5925 , \7059 );
nor \U$12669 ( \12922 , \12920 , \12921 );
xnor \U$12670 ( \12923 , \12922 , \7067 );
xor \U$12671 ( \12924 , \12919 , \12923 );
and \U$12672 ( \12925 , \5979 , \7082 );
and \U$12673 ( \12926 , \5945 , \7080 );
nor \U$12674 ( \12927 , \12925 , \12926 );
xnor \U$12675 ( \12928 , \12927 , \7088 );
xor \U$12676 ( \12929 , \12924 , \12928 );
xor \U$12677 ( \12930 , \12915 , \12929 );
and \U$12678 ( \12931 , \5873 , \6991 );
and \U$12679 ( \12932 , \5842 , \6988 );
nor \U$12680 ( \12933 , \12931 , \12932 );
xnor \U$12681 ( \12934 , \12933 , \6985 );
and \U$12682 ( \12935 , \5893 , \7006 );
and \U$12683 ( \12936 , \5861 , \7004 );
nor \U$12684 ( \12937 , \12935 , \12936 );
xnor \U$12685 ( \12938 , \12937 , \7012 );
xor \U$12686 ( \12939 , \12934 , \12938 );
and \U$12687 ( \12940 , \5918 , \7026 );
and \U$12688 ( \12941 , \5881 , \7024 );
nor \U$12689 ( \12942 , \12940 , \12941 );
xnor \U$12690 ( \12943 , \12942 , \7032 );
xor \U$12691 ( \12944 , \12939 , \12943 );
xor \U$12692 ( \12945 , \12930 , \12944 );
xor \U$12693 ( \12946 , \12901 , \12945 );
xor \U$12694 ( \12947 , \12892 , \12946 );
xor \U$12695 ( \12948 , \12878 , \12947 );
and \U$12696 ( \12949 , \12850 , \12854 );
and \U$12697 ( \12950 , \12854 , \12865 );
and \U$12698 ( \12951 , \12850 , \12865 );
or \U$12699 ( \12952 , \12949 , \12950 , \12951 );
and \U$12700 ( \12953 , \12830 , \12844 );
xor \U$12701 ( \12954 , \12952 , \12953 );
and \U$12702 ( \12955 , \12792 , \12796 );
and \U$12703 ( \12956 , \12796 , \12799 );
and \U$12704 ( \12957 , \12792 , \12799 );
or \U$12705 ( \12958 , \12955 , \12956 , \12957 );
and \U$12706 ( \12959 , \6057 , \7157 );
and \U$12707 ( \12960 , \6029 , \7155 );
nor \U$12708 ( \12961 , \12959 , \12960 );
xnor \U$12709 ( \12962 , \12961 , \7163 );
xor \U$12710 ( \12963 , \12958 , \12962 );
and \U$12711 ( \12964 , \6065 , \7175 );
and \U$12712 ( \12965 , \6048 , \7173 );
nor \U$12713 ( \12966 , \12964 , \12965 );
xnor \U$12714 ( \12967 , \12966 , \7181 );
xor \U$12715 ( \12968 , \12963 , \12967 );
xor \U$12716 ( \12969 , \12954 , \12968 );
xor \U$12717 ( \12970 , \12948 , \12969 );
and \U$12718 ( \12971 , \12782 , \12783 );
and \U$12719 ( \12972 , \12783 , \12867 );
and \U$12720 ( \12973 , \12782 , \12867 );
or \U$12721 ( \12974 , \12971 , \12972 , \12973 );
nor \U$12722 ( \12975 , \12970 , \12974 );
and \U$12723 ( \12976 , \12952 , \12953 );
and \U$12724 ( \12977 , \12953 , \12968 );
and \U$12725 ( \12978 , \12952 , \12968 );
or \U$12726 ( \12979 , \12976 , \12977 , \12978 );
and \U$12727 ( \12980 , \12892 , \12946 );
xor \U$12728 ( \12981 , \12979 , \12980 );
and \U$12729 ( \12982 , \12896 , \12900 );
and \U$12730 ( \12983 , \12900 , \12945 );
and \U$12731 ( \12984 , \12896 , \12945 );
or \U$12732 ( \12985 , \12982 , \12983 , \12984 );
and \U$12733 ( \12986 , \5881 , \7026 );
and \U$12734 ( \12987 , \5893 , \7024 );
nor \U$12735 ( \12988 , \12986 , \12987 );
xnor \U$12736 ( \12989 , \12988 , \7032 );
and \U$12737 ( \12990 , \5906 , \7043 );
and \U$12738 ( \12991 , \5918 , \7041 );
nor \U$12739 ( \12992 , \12990 , \12991 );
xnor \U$12740 ( \12993 , \12992 , \7049 );
xor \U$12741 ( \12994 , \12989 , \12993 );
and \U$12742 ( \12995 , \5925 , \7061 );
and \U$12743 ( \12996 , \5937 , \7059 );
nor \U$12744 ( \12997 , \12995 , \12996 );
xnor \U$12745 ( \12998 , \12997 , \7067 );
xor \U$12746 ( \12999 , \12994 , \12998 );
and \U$12747 ( \13000 , \5842 , \6991 );
and \U$12748 ( \13001 , \5854 , \6988 );
nor \U$12749 ( \13002 , \13000 , \13001 );
xnor \U$12750 ( \13003 , \13002 , \6985 );
xor \U$12751 ( \13004 , \7198 , \13003 );
and \U$12752 ( \13005 , \5861 , \7006 );
and \U$12753 ( \13006 , \5873 , \7004 );
nor \U$12754 ( \13007 , \13005 , \13006 );
xnor \U$12755 ( \13008 , \13007 , \7012 );
xor \U$12756 ( \13009 , \13004 , \13008 );
xor \U$12757 ( \13010 , \12999 , \13009 );
nand \U$12758 ( \13011 , \6065 , \7190 );
xnor \U$12759 ( \13012 , \13011 , \7198 );
and \U$12760 ( \13013 , \6006 , \7140 );
and \U$12761 ( \13014 , \6018 , \7138 );
nor \U$12762 ( \13015 , \13013 , \13014 );
xnor \U$12763 ( \13016 , \13015 , \7146 );
and \U$12764 ( \13017 , \6029 , \7157 );
and \U$12765 ( \13018 , \6041 , \7155 );
nor \U$12766 ( \13019 , \13017 , \13018 );
xnor \U$12767 ( \13020 , \13019 , \7163 );
xor \U$12768 ( \13021 , \13016 , \13020 );
and \U$12769 ( \13022 , \6048 , \7175 );
and \U$12770 ( \13023 , \6057 , \7173 );
nor \U$12771 ( \13024 , \13022 , \13023 );
xnor \U$12772 ( \13025 , \13024 , \7181 );
xor \U$12773 ( \13026 , \13021 , \13025 );
xor \U$12774 ( \13027 , \13012 , \13026 );
and \U$12775 ( \13028 , \5945 , \7082 );
and \U$12776 ( \13029 , \5957 , \7080 );
nor \U$12777 ( \13030 , \13028 , \13029 );
xnor \U$12778 ( \13031 , \13030 , \7088 );
and \U$12779 ( \13032 , \5967 , \7099 );
and \U$12780 ( \13033 , \5979 , \7097 );
nor \U$12781 ( \13034 , \13032 , \13033 );
xnor \U$12782 ( \13035 , \13034 , \7105 );
xor \U$12783 ( \13036 , \13031 , \13035 );
and \U$12784 ( \13037 , \5986 , \7117 );
and \U$12785 ( \13038 , \5998 , \7115 );
nor \U$12786 ( \13039 , \13037 , \13038 );
xnor \U$12787 ( \13040 , \13039 , \7123 );
xor \U$12788 ( \13041 , \13036 , \13040 );
xor \U$12789 ( \13042 , \13027 , \13041 );
xor \U$12790 ( \13043 , \13010 , \13042 );
and \U$12791 ( \13044 , \12934 , \12938 );
and \U$12792 ( \13045 , \12938 , \12943 );
and \U$12793 ( \13046 , \12934 , \12943 );
or \U$12794 ( \13047 , \13044 , \13045 , \13046 );
and \U$12795 ( \13048 , \12919 , \12923 );
and \U$12796 ( \13049 , \12923 , \12928 );
and \U$12797 ( \13050 , \12919 , \12928 );
or \U$12798 ( \13051 , \13048 , \13049 , \13050 );
xor \U$12799 ( \13052 , \13047 , \13051 );
and \U$12800 ( \13053 , \12905 , \12909 );
and \U$12801 ( \13054 , \12909 , \12914 );
and \U$12802 ( \13055 , \12905 , \12914 );
or \U$12803 ( \13056 , \13053 , \13054 , \13055 );
xor \U$12804 ( \13057 , \13052 , \13056 );
xor \U$12805 ( \13058 , \13043 , \13057 );
xor \U$12806 ( \13059 , \12985 , \13058 );
and \U$12807 ( \13060 , \12882 , \12886 );
and \U$12808 ( \13061 , \12886 , \12891 );
and \U$12809 ( \13062 , \12882 , \12891 );
or \U$12810 ( \13063 , \13060 , \13061 , \13062 );
and \U$12811 ( \13064 , \12958 , \12962 );
and \U$12812 ( \13065 , \12962 , \12967 );
and \U$12813 ( \13066 , \12958 , \12967 );
or \U$12814 ( \13067 , \13064 , \13065 , \13066 );
xor \U$12815 ( \13068 , \13063 , \13067 );
and \U$12816 ( \13069 , \12915 , \12929 );
and \U$12817 ( \13070 , \12929 , \12944 );
and \U$12818 ( \13071 , \12915 , \12944 );
or \U$12819 ( \13072 , \13069 , \13070 , \13071 );
xor \U$12820 ( \13073 , \13068 , \13072 );
xor \U$12821 ( \13074 , \13059 , \13073 );
xor \U$12822 ( \13075 , \12981 , \13074 );
and \U$12823 ( \13076 , \12878 , \12947 );
and \U$12824 ( \13077 , \12947 , \12969 );
and \U$12825 ( \13078 , \12878 , \12969 );
or \U$12826 ( \13079 , \13076 , \13077 , \13078 );
nor \U$12827 ( \13080 , \13075 , \13079 );
nor \U$12828 ( \13081 , \12975 , \13080 );
nand \U$12829 ( \13082 , \12874 , \13081 );
nor \U$12830 ( \13083 , \12687 , \13082 );
and \U$12831 ( \13084 , \12985 , \13058 );
and \U$12832 ( \13085 , \13058 , \13073 );
and \U$12833 ( \13086 , \12985 , \13073 );
or \U$12834 ( \13087 , \13084 , \13085 , \13086 );
and \U$12835 ( \13088 , \13047 , \13051 );
and \U$12836 ( \13089 , \13051 , \13056 );
and \U$12837 ( \13090 , \13047 , \13056 );
or \U$12838 ( \13091 , \13088 , \13089 , \13090 );
and \U$12839 ( \13092 , \13012 , \13026 );
and \U$12840 ( \13093 , \13026 , \13041 );
and \U$12841 ( \13094 , \13012 , \13041 );
or \U$12842 ( \13095 , \13092 , \13093 , \13094 );
xor \U$12843 ( \13096 , \13091 , \13095 );
and \U$12844 ( \13097 , \12999 , \13009 );
xor \U$12845 ( \13098 , \13096 , \13097 );
xor \U$12846 ( \13099 , \13087 , \13098 );
and \U$12847 ( \13100 , \13063 , \13067 );
and \U$12848 ( \13101 , \13067 , \13072 );
and \U$12849 ( \13102 , \13063 , \13072 );
or \U$12850 ( \13103 , \13100 , \13101 , \13102 );
and \U$12851 ( \13104 , \13010 , \13042 );
and \U$12852 ( \13105 , \13042 , \13057 );
and \U$12853 ( \13106 , \13010 , \13057 );
or \U$12854 ( \13107 , \13104 , \13105 , \13106 );
xor \U$12855 ( \13108 , \13103 , \13107 );
and \U$12856 ( \13109 , \5918 , \7043 );
and \U$12857 ( \13110 , \5881 , \7041 );
nor \U$12858 ( \13111 , \13109 , \13110 );
xnor \U$12859 ( \13112 , \13111 , \7049 );
and \U$12860 ( \13113 , \5937 , \7061 );
and \U$12861 ( \13114 , \5906 , \7059 );
nor \U$12862 ( \13115 , \13113 , \13114 );
xnor \U$12863 ( \13116 , \13115 , \7067 );
xor \U$12864 ( \13117 , \13112 , \13116 );
and \U$12865 ( \13118 , \5957 , \7082 );
and \U$12866 ( \13119 , \5925 , \7080 );
nor \U$12867 ( \13120 , \13118 , \13119 );
xnor \U$12868 ( \13121 , \13120 , \7088 );
xor \U$12869 ( \13122 , \13117 , \13121 );
and \U$12870 ( \13123 , \5854 , \6991 );
and \U$12871 ( \13124 , \5819 , \6988 );
nor \U$12872 ( \13125 , \13123 , \13124 );
xnor \U$12873 ( \13126 , \13125 , \6985 );
and \U$12874 ( \13127 , \5873 , \7006 );
and \U$12875 ( \13128 , \5842 , \7004 );
nor \U$12876 ( \13129 , \13127 , \13128 );
xnor \U$12877 ( \13130 , \13129 , \7012 );
xor \U$12878 ( \13131 , \13126 , \13130 );
and \U$12879 ( \13132 , \5893 , \7026 );
and \U$12880 ( \13133 , \5861 , \7024 );
nor \U$12881 ( \13134 , \13132 , \13133 );
xnor \U$12882 ( \13135 , \13134 , \7032 );
xor \U$12883 ( \13136 , \13131 , \13135 );
xor \U$12884 ( \13137 , \13122 , \13136 );
and \U$12885 ( \13138 , \13016 , \13020 );
and \U$12886 ( \13139 , \13020 , \13025 );
and \U$12887 ( \13140 , \13016 , \13025 );
or \U$12888 ( \13141 , \13138 , \13139 , \13140 );
and \U$12889 ( \13142 , \6041 , \7157 );
and \U$12890 ( \13143 , \6006 , \7155 );
nor \U$12891 ( \13144 , \13142 , \13143 );
xnor \U$12892 ( \13145 , \13144 , \7163 );
and \U$12893 ( \13146 , \6057 , \7175 );
and \U$12894 ( \13147 , \6029 , \7173 );
nor \U$12895 ( \13148 , \13146 , \13147 );
xnor \U$12896 ( \13149 , \13148 , \7181 );
xor \U$12897 ( \13150 , \13145 , \13149 );
and \U$12898 ( \13151 , \6065 , \7192 );
and \U$12899 ( \13152 , \6048 , \7190 );
nor \U$12900 ( \13153 , \13151 , \13152 );
xnor \U$12901 ( \13154 , \13153 , \7198 );
xor \U$12902 ( \13155 , \13150 , \13154 );
xor \U$12903 ( \13156 , \13141 , \13155 );
and \U$12904 ( \13157 , \5979 , \7099 );
and \U$12905 ( \13158 , \5945 , \7097 );
nor \U$12906 ( \13159 , \13157 , \13158 );
xnor \U$12907 ( \13160 , \13159 , \7105 );
and \U$12908 ( \13161 , \5998 , \7117 );
and \U$12909 ( \13162 , \5967 , \7115 );
nor \U$12910 ( \13163 , \13161 , \13162 );
xnor \U$12911 ( \13164 , \13163 , \7123 );
xor \U$12912 ( \13165 , \13160 , \13164 );
and \U$12913 ( \13166 , \6018 , \7140 );
and \U$12914 ( \13167 , \5986 , \7138 );
nor \U$12915 ( \13168 , \13166 , \13167 );
xnor \U$12916 ( \13169 , \13168 , \7146 );
xor \U$12917 ( \13170 , \13165 , \13169 );
xor \U$12918 ( \13171 , \13156 , \13170 );
xor \U$12919 ( \13172 , \13137 , \13171 );
and \U$12920 ( \13173 , \7198 , \13003 );
and \U$12921 ( \13174 , \13003 , \13008 );
and \U$12922 ( \13175 , \7198 , \13008 );
or \U$12923 ( \13176 , \13173 , \13174 , \13175 );
and \U$12924 ( \13177 , \12989 , \12993 );
and \U$12925 ( \13178 , \12993 , \12998 );
and \U$12926 ( \13179 , \12989 , \12998 );
or \U$12927 ( \13180 , \13177 , \13178 , \13179 );
xor \U$12928 ( \13181 , \13176 , \13180 );
and \U$12929 ( \13182 , \13031 , \13035 );
and \U$12930 ( \13183 , \13035 , \13040 );
and \U$12931 ( \13184 , \13031 , \13040 );
or \U$12932 ( \13185 , \13182 , \13183 , \13184 );
xor \U$12933 ( \13186 , \13181 , \13185 );
xor \U$12934 ( \13187 , \13172 , \13186 );
xor \U$12935 ( \13188 , \13108 , \13187 );
xor \U$12936 ( \13189 , \13099 , \13188 );
and \U$12937 ( \13190 , \12979 , \12980 );
and \U$12938 ( \13191 , \12980 , \13074 );
and \U$12939 ( \13192 , \12979 , \13074 );
or \U$12940 ( \13193 , \13190 , \13191 , \13192 );
nor \U$12941 ( \13194 , \13189 , \13193 );
and \U$12942 ( \13195 , \13103 , \13107 );
and \U$12943 ( \13196 , \13107 , \13187 );
and \U$12944 ( \13197 , \13103 , \13187 );
or \U$12945 ( \13198 , \13195 , \13196 , \13197 );
and \U$12946 ( \13199 , \13176 , \13180 );
and \U$12947 ( \13200 , \13180 , \13185 );
and \U$12948 ( \13201 , \13176 , \13185 );
or \U$12949 ( \13202 , \13199 , \13200 , \13201 );
and \U$12950 ( \13203 , \13141 , \13155 );
and \U$12951 ( \13204 , \13155 , \13170 );
and \U$12952 ( \13205 , \13141 , \13170 );
or \U$12953 ( \13206 , \13203 , \13204 , \13205 );
xor \U$12954 ( \13207 , \13202 , \13206 );
and \U$12955 ( \13208 , \13122 , \13136 );
xor \U$12956 ( \13209 , \13207 , \13208 );
xor \U$12957 ( \13210 , \13198 , \13209 );
and \U$12958 ( \13211 , \13091 , \13095 );
and \U$12959 ( \13212 , \13095 , \13097 );
and \U$12960 ( \13213 , \13091 , \13097 );
or \U$12961 ( \13214 , \13211 , \13212 , \13213 );
and \U$12962 ( \13215 , \13137 , \13171 );
and \U$12963 ( \13216 , \13171 , \13186 );
and \U$12964 ( \13217 , \13137 , \13186 );
or \U$12965 ( \13218 , \13215 , \13216 , \13217 );
xor \U$12966 ( \13219 , \13214 , \13218 );
and \U$12967 ( \13220 , \5925 , \7082 );
and \U$12968 ( \13221 , \5937 , \7080 );
nor \U$12969 ( \13222 , \13220 , \13221 );
xnor \U$12970 ( \13223 , \13222 , \7088 );
and \U$12971 ( \13224 , \5945 , \7099 );
and \U$12972 ( \13225 , \5957 , \7097 );
nor \U$12973 ( \13226 , \13224 , \13225 );
xnor \U$12974 ( \13227 , \13226 , \7105 );
xor \U$12975 ( \13228 , \13223 , \13227 );
and \U$12976 ( \13229 , \5967 , \7117 );
and \U$12977 ( \13230 , \5979 , \7115 );
nor \U$12978 ( \13231 , \13229 , \13230 );
xnor \U$12979 ( \13232 , \13231 , \7123 );
xor \U$12980 ( \13233 , \13228 , \13232 );
and \U$12981 ( \13234 , \5861 , \7026 );
and \U$12982 ( \13235 , \5873 , \7024 );
nor \U$12983 ( \13236 , \13234 , \13235 );
xnor \U$12984 ( \13237 , \13236 , \7032 );
and \U$12985 ( \13238 , \5881 , \7043 );
and \U$12986 ( \13239 , \5893 , \7041 );
nor \U$12987 ( \13240 , \13238 , \13239 );
xnor \U$12988 ( \13241 , \13240 , \7049 );
xor \U$12989 ( \13242 , \13237 , \13241 );
and \U$12990 ( \13243 , \5906 , \7061 );
and \U$12991 ( \13244 , \5918 , \7059 );
nor \U$12992 ( \13245 , \13243 , \13244 );
xnor \U$12993 ( \13246 , \13245 , \7067 );
xor \U$12994 ( \13247 , \13242 , \13246 );
xor \U$12995 ( \13248 , \13233 , \13247 );
and \U$12996 ( \13249 , \5819 , \6991 );
and \U$12997 ( \13250 , \5831 , \6988 );
nor \U$12998 ( \13251 , \13249 , \13250 );
xnor \U$12999 ( \13252 , \13251 , \6985 );
xor \U$13000 ( \13253 , \6824 , \13252 );
and \U$13001 ( \13254 , \5842 , \7006 );
and \U$13002 ( \13255 , \5854 , \7004 );
nor \U$13003 ( \13256 , \13254 , \13255 );
xnor \U$13004 ( \13257 , \13256 , \7012 );
xor \U$13005 ( \13258 , \13253 , \13257 );
xor \U$13006 ( \13259 , \13248 , \13258 );
and \U$13007 ( \13260 , \13145 , \13149 );
and \U$13008 ( \13261 , \13149 , \13154 );
and \U$13009 ( \13262 , \13145 , \13154 );
or \U$13010 ( \13263 , \13260 , \13261 , \13262 );
and \U$13011 ( \13264 , \6048 , \7192 );
and \U$13012 ( \13265 , \6057 , \7190 );
nor \U$13013 ( \13266 , \13264 , \13265 );
xnor \U$13014 ( \13267 , \13266 , \7198 );
nand \U$13015 ( \13268 , \6065 , \7201 );
xnor \U$13016 ( \13269 , \13268 , \6824 );
xor \U$13017 ( \13270 , \13267 , \13269 );
xor \U$13018 ( \13271 , \13263 , \13270 );
and \U$13019 ( \13272 , \5986 , \7140 );
and \U$13020 ( \13273 , \5998 , \7138 );
nor \U$13021 ( \13274 , \13272 , \13273 );
xnor \U$13022 ( \13275 , \13274 , \7146 );
and \U$13023 ( \13276 , \6006 , \7157 );
and \U$13024 ( \13277 , \6018 , \7155 );
nor \U$13025 ( \13278 , \13276 , \13277 );
xnor \U$13026 ( \13279 , \13278 , \7163 );
xor \U$13027 ( \13280 , \13275 , \13279 );
and \U$13028 ( \13281 , \6029 , \7175 );
and \U$13029 ( \13282 , \6041 , \7173 );
nor \U$13030 ( \13283 , \13281 , \13282 );
xnor \U$13031 ( \13284 , \13283 , \7181 );
xor \U$13032 ( \13285 , \13280 , \13284 );
xor \U$13033 ( \13286 , \13271 , \13285 );
xor \U$13034 ( \13287 , \13259 , \13286 );
and \U$13035 ( \13288 , \13126 , \13130 );
and \U$13036 ( \13289 , \13130 , \13135 );
and \U$13037 ( \13290 , \13126 , \13135 );
or \U$13038 ( \13291 , \13288 , \13289 , \13290 );
and \U$13039 ( \13292 , \13112 , \13116 );
and \U$13040 ( \13293 , \13116 , \13121 );
and \U$13041 ( \13294 , \13112 , \13121 );
or \U$13042 ( \13295 , \13292 , \13293 , \13294 );
xor \U$13043 ( \13296 , \13291 , \13295 );
and \U$13044 ( \13297 , \13160 , \13164 );
and \U$13045 ( \13298 , \13164 , \13169 );
and \U$13046 ( \13299 , \13160 , \13169 );
or \U$13047 ( \13300 , \13297 , \13298 , \13299 );
xor \U$13048 ( \13301 , \13296 , \13300 );
xor \U$13049 ( \13302 , \13287 , \13301 );
xor \U$13050 ( \13303 , \13219 , \13302 );
xor \U$13051 ( \13304 , \13210 , \13303 );
and \U$13052 ( \13305 , \13087 , \13098 );
and \U$13053 ( \13306 , \13098 , \13188 );
and \U$13054 ( \13307 , \13087 , \13188 );
or \U$13055 ( \13308 , \13305 , \13306 , \13307 );
nor \U$13056 ( \13309 , \13304 , \13308 );
nor \U$13057 ( \13310 , \13194 , \13309 );
and \U$13058 ( \13311 , \13214 , \13218 );
and \U$13059 ( \13312 , \13218 , \13302 );
and \U$13060 ( \13313 , \13214 , \13302 );
or \U$13061 ( \13314 , \13311 , \13312 , \13313 );
xor \U$13062 ( \13315 , \7770 , \7774 );
xor \U$13063 ( \13316 , \13315 , \7779 );
xor \U$13064 ( \13317 , \7822 , \7826 );
xor \U$13065 ( \13318 , \13317 , \7831 );
xor \U$13066 ( \13319 , \7803 , \7807 );
xor \U$13067 ( \13320 , \13319 , \7812 );
xor \U$13068 ( \13321 , \13318 , \13320 );
xor \U$13069 ( \13322 , \7786 , \7790 );
xor \U$13070 ( \13323 , \13322 , \7795 );
xor \U$13071 ( \13324 , \13321 , \13323 );
xor \U$13072 ( \13325 , \13316 , \13324 );
and \U$13073 ( \13326 , \13275 , \13279 );
and \U$13074 ( \13327 , \13279 , \13284 );
and \U$13075 ( \13328 , \13275 , \13284 );
or \U$13076 ( \13329 , \13326 , \13327 , \13328 );
and \U$13077 ( \13330 , \13267 , \13269 );
xor \U$13078 ( \13331 , \13329 , \13330 );
and \U$13079 ( \13332 , \6065 , \7203 );
and \U$13080 ( \13333 , \6048 , \7201 );
nor \U$13081 ( \13334 , \13332 , \13333 );
xnor \U$13082 ( \13335 , \13334 , \6824 );
xor \U$13083 ( \13336 , \13331 , \13335 );
xor \U$13084 ( \13337 , \13325 , \13336 );
and \U$13085 ( \13338 , \13291 , \13295 );
and \U$13086 ( \13339 , \13295 , \13300 );
and \U$13087 ( \13340 , \13291 , \13300 );
or \U$13088 ( \13341 , \13338 , \13339 , \13340 );
and \U$13089 ( \13342 , \13263 , \13270 );
and \U$13090 ( \13343 , \13270 , \13285 );
and \U$13091 ( \13344 , \13263 , \13285 );
or \U$13092 ( \13345 , \13342 , \13343 , \13344 );
xor \U$13093 ( \13346 , \13341 , \13345 );
and \U$13094 ( \13347 , \13233 , \13247 );
and \U$13095 ( \13348 , \13247 , \13258 );
and \U$13096 ( \13349 , \13233 , \13258 );
or \U$13097 ( \13350 , \13347 , \13348 , \13349 );
xor \U$13098 ( \13351 , \13346 , \13350 );
xor \U$13099 ( \13352 , \13337 , \13351 );
xor \U$13100 ( \13353 , \13314 , \13352 );
and \U$13101 ( \13354 , \13202 , \13206 );
and \U$13102 ( \13355 , \13206 , \13208 );
and \U$13103 ( \13356 , \13202 , \13208 );
or \U$13104 ( \13357 , \13354 , \13355 , \13356 );
and \U$13105 ( \13358 , \13259 , \13286 );
and \U$13106 ( \13359 , \13286 , \13301 );
and \U$13107 ( \13360 , \13259 , \13301 );
or \U$13108 ( \13361 , \13358 , \13359 , \13360 );
xor \U$13109 ( \13362 , \13357 , \13361 );
and \U$13110 ( \13363 , \6824 , \13252 );
and \U$13111 ( \13364 , \13252 , \13257 );
and \U$13112 ( \13365 , \6824 , \13257 );
or \U$13113 ( \13366 , \13363 , \13364 , \13365 );
and \U$13114 ( \13367 , \13237 , \13241 );
and \U$13115 ( \13368 , \13241 , \13246 );
and \U$13116 ( \13369 , \13237 , \13246 );
or \U$13117 ( \13370 , \13367 , \13368 , \13369 );
xor \U$13118 ( \13371 , \13366 , \13370 );
and \U$13119 ( \13372 , \13223 , \13227 );
and \U$13120 ( \13373 , \13227 , \13232 );
and \U$13121 ( \13374 , \13223 , \13232 );
or \U$13122 ( \13375 , \13372 , \13373 , \13374 );
xor \U$13123 ( \13376 , \13371 , \13375 );
xor \U$13124 ( \13377 , \13362 , \13376 );
xor \U$13125 ( \13378 , \13353 , \13377 );
and \U$13126 ( \13379 , \13198 , \13209 );
and \U$13127 ( \13380 , \13209 , \13303 );
and \U$13128 ( \13381 , \13198 , \13303 );
or \U$13129 ( \13382 , \13379 , \13380 , \13381 );
nor \U$13130 ( \13383 , \13378 , \13382 );
and \U$13131 ( \13384 , \13341 , \13345 );
and \U$13132 ( \13385 , \13345 , \13350 );
and \U$13133 ( \13386 , \13341 , \13350 );
or \U$13134 ( \13387 , \13384 , \13385 , \13386 );
and \U$13135 ( \13388 , \13316 , \13324 );
and \U$13136 ( \13389 , \13324 , \13336 );
and \U$13137 ( \13390 , \13316 , \13336 );
or \U$13138 ( \13391 , \13388 , \13389 , \13390 );
xor \U$13139 ( \13392 , \13387 , \13391 );
xor \U$13140 ( \13393 , \7845 , \7847 );
xor \U$13141 ( \13394 , \13393 , \7850 );
xor \U$13142 ( \13395 , \7834 , \7836 );
xor \U$13143 ( \13396 , \13395 , \7839 );
xor \U$13144 ( \13397 , \13394 , \13396 );
xor \U$13145 ( \13398 , \7782 , \7798 );
xor \U$13146 ( \13399 , \13398 , \7815 );
xor \U$13147 ( \13400 , \13397 , \13399 );
xor \U$13148 ( \13401 , \13392 , \13400 );
and \U$13149 ( \13402 , \13357 , \13361 );
and \U$13150 ( \13403 , \13361 , \13376 );
and \U$13151 ( \13404 , \13357 , \13376 );
or \U$13152 ( \13405 , \13402 , \13403 , \13404 );
and \U$13153 ( \13406 , \13337 , \13351 );
xor \U$13154 ( \13407 , \13405 , \13406 );
and \U$13155 ( \13408 , \13366 , \13370 );
and \U$13156 ( \13409 , \13370 , \13375 );
and \U$13157 ( \13410 , \13366 , \13375 );
or \U$13158 ( \13411 , \13408 , \13409 , \13410 );
and \U$13159 ( \13412 , \13329 , \13330 );
and \U$13160 ( \13413 , \13330 , \13335 );
and \U$13161 ( \13414 , \13329 , \13335 );
or \U$13162 ( \13415 , \13412 , \13413 , \13414 );
xor \U$13163 ( \13416 , \13411 , \13415 );
and \U$13164 ( \13417 , \13318 , \13320 );
and \U$13165 ( \13418 , \13320 , \13323 );
and \U$13166 ( \13419 , \13318 , \13323 );
or \U$13167 ( \13420 , \13417 , \13418 , \13419 );
xor \U$13168 ( \13421 , \13416 , \13420 );
xor \U$13169 ( \13422 , \13407 , \13421 );
xor \U$13170 ( \13423 , \13401 , \13422 );
and \U$13171 ( \13424 , \13314 , \13352 );
and \U$13172 ( \13425 , \13352 , \13377 );
and \U$13173 ( \13426 , \13314 , \13377 );
or \U$13174 ( \13427 , \13424 , \13425 , \13426 );
nor \U$13175 ( \13428 , \13423 , \13427 );
nor \U$13176 ( \13429 , \13383 , \13428 );
nand \U$13177 ( \13430 , \13310 , \13429 );
and \U$13178 ( \13431 , \13405 , \13406 );
and \U$13179 ( \13432 , \13406 , \13421 );
and \U$13180 ( \13433 , \13405 , \13421 );
or \U$13181 ( \13434 , \13431 , \13432 , \13433 );
and \U$13182 ( \13435 , \13387 , \13391 );
and \U$13183 ( \13436 , \13391 , \13400 );
and \U$13184 ( \13437 , \13387 , \13400 );
or \U$13185 ( \13438 , \13435 , \13436 , \13437 );
xor \U$13186 ( \13439 , \7016 , \7071 );
xor \U$13187 ( \13440 , \13439 , \7127 );
xor \U$13188 ( \13441 , \7858 , \7860 );
xor \U$13189 ( \13442 , \13441 , \7863 );
xor \U$13190 ( \13443 , \13440 , \13442 );
xor \U$13191 ( \13444 , \7818 , \7842 );
xor \U$13192 ( \13445 , \13444 , \7853 );
xor \U$13193 ( \13446 , \13443 , \13445 );
xor \U$13194 ( \13447 , \13438 , \13446 );
and \U$13195 ( \13448 , \13411 , \13415 );
and \U$13196 ( \13449 , \13415 , \13420 );
and \U$13197 ( \13450 , \13411 , \13420 );
or \U$13198 ( \13451 , \13448 , \13449 , \13450 );
and \U$13199 ( \13452 , \13394 , \13396 );
and \U$13200 ( \13453 , \13396 , \13399 );
and \U$13201 ( \13454 , \13394 , \13399 );
or \U$13202 ( \13455 , \13452 , \13453 , \13454 );
xor \U$13203 ( \13456 , \13451 , \13455 );
xor \U$13204 ( \13457 , \7185 , \7213 );
xor \U$13205 ( \13458 , \13457 , \7218 );
xor \U$13206 ( \13459 , \13456 , \13458 );
xor \U$13207 ( \13460 , \13447 , \13459 );
xor \U$13208 ( \13461 , \13434 , \13460 );
and \U$13209 ( \13462 , \13401 , \13422 );
nor \U$13210 ( \13463 , \13461 , \13462 );
and \U$13211 ( \13464 , \13438 , \13446 );
and \U$13212 ( \13465 , \13446 , \13459 );
and \U$13213 ( \13466 , \13438 , \13459 );
or \U$13214 ( \13467 , \13464 , \13465 , \13466 );
xor \U$13215 ( \13468 , \7130 , \7221 );
xor \U$13216 ( \13469 , \13468 , \7258 );
xor \U$13217 ( \13470 , \7856 , \7866 );
xor \U$13218 ( \13471 , \13470 , \7869 );
xor \U$13219 ( \13472 , \13469 , \13471 );
xor \U$13220 ( \13473 , \13467 , \13472 );
and \U$13221 ( \13474 , \13451 , \13455 );
and \U$13222 ( \13475 , \13455 , \13458 );
and \U$13223 ( \13476 , \13451 , \13458 );
or \U$13224 ( \13477 , \13474 , \13475 , \13476 );
and \U$13225 ( \13478 , \13440 , \13442 );
and \U$13226 ( \13479 , \13442 , \13445 );
and \U$13227 ( \13480 , \13440 , \13445 );
or \U$13228 ( \13481 , \13478 , \13479 , \13480 );
xor \U$13229 ( \13482 , \13477 , \13481 );
xor \U$13230 ( \13483 , \7271 , \7315 );
xor \U$13231 ( \13484 , \13483 , \7338 );
xor \U$13232 ( \13485 , \13482 , \13484 );
xor \U$13233 ( \13486 , \13473 , \13485 );
and \U$13234 ( \13487 , \13434 , \13460 );
nor \U$13235 ( \13488 , \13486 , \13487 );
nor \U$13236 ( \13489 , \13463 , \13488 );
and \U$13237 ( \13490 , \13477 , \13481 );
and \U$13238 ( \13491 , \13481 , \13484 );
and \U$13239 ( \13492 , \13477 , \13484 );
or \U$13240 ( \13493 , \13490 , \13491 , \13492 );
and \U$13241 ( \13494 , \13469 , \13471 );
xor \U$13242 ( \13495 , \13493 , \13494 );
xor \U$13243 ( \13496 , \7872 , \7873 );
xor \U$13244 ( \13497 , \13496 , \7876 );
xor \U$13245 ( \13498 , \13495 , \13497 );
and \U$13246 ( \13499 , \13467 , \13472 );
and \U$13247 ( \13500 , \13472 , \13485 );
and \U$13248 ( \13501 , \13467 , \13485 );
or \U$13249 ( \13502 , \13499 , \13500 , \13501 );
nor \U$13250 ( \13503 , \13498 , \13502 );
xor \U$13251 ( \13504 , \7879 , \7880 );
xor \U$13252 ( \13505 , \13504 , \7883 );
and \U$13253 ( \13506 , \13493 , \13494 );
and \U$13254 ( \13507 , \13494 , \13497 );
and \U$13255 ( \13508 , \13493 , \13497 );
or \U$13256 ( \13509 , \13506 , \13507 , \13508 );
nor \U$13257 ( \13510 , \13505 , \13509 );
nor \U$13258 ( \13511 , \13503 , \13510 );
nand \U$13259 ( \13512 , \13489 , \13511 );
nor \U$13260 ( \13513 , \13430 , \13512 );
nand \U$13261 ( \13514 , \13083 , \13513 );
and \U$13262 ( \13515 , \6018 , \6991 );
and \U$13263 ( \13516 , \5986 , \6988 );
nor \U$13264 ( \13517 , \13515 , \13516 );
xnor \U$13265 ( \13518 , \13517 , \6985 );
and \U$13266 ( \13519 , \6041 , \7006 );
and \U$13267 ( \13520 , \6006 , \7004 );
nor \U$13268 ( \13521 , \13519 , \13520 );
xnor \U$13269 ( \13522 , \13521 , \7012 );
xor \U$13270 ( \13523 , \13518 , \13522 );
and \U$13271 ( \13524 , \6057 , \7026 );
and \U$13272 ( \13525 , \6029 , \7024 );
nor \U$13273 ( \13526 , \13524 , \13525 );
xnor \U$13274 ( \13527 , \13526 , \7032 );
xor \U$13275 ( \13528 , \13523 , \13527 );
and \U$13276 ( \13529 , \6006 , \6991 );
and \U$13277 ( \13530 , \6018 , \6988 );
nor \U$13278 ( \13531 , \13529 , \13530 );
xnor \U$13279 ( \13532 , \13531 , \6985 );
and \U$13280 ( \13533 , \7049 , \13532 );
and \U$13281 ( \13534 , \6029 , \7006 );
and \U$13282 ( \13535 , \6041 , \7004 );
nor \U$13283 ( \13536 , \13534 , \13535 );
xnor \U$13284 ( \13537 , \13536 , \7012 );
and \U$13285 ( \13538 , \13532 , \13537 );
and \U$13286 ( \13539 , \7049 , \13537 );
or \U$13287 ( \13540 , \13533 , \13538 , \13539 );
and \U$13288 ( \13541 , \6048 , \7026 );
and \U$13289 ( \13542 , \6057 , \7024 );
nor \U$13290 ( \13543 , \13541 , \13542 );
xnor \U$13291 ( \13544 , \13543 , \7032 );
nand \U$13292 ( \13545 , \6065 , \7041 );
xnor \U$13293 ( \13546 , \13545 , \7049 );
and \U$13294 ( \13547 , \13544 , \13546 );
xor \U$13295 ( \13548 , \13540 , \13547 );
and \U$13296 ( \13549 , \6065 , \7043 );
and \U$13297 ( \13550 , \6048 , \7041 );
nor \U$13298 ( \13551 , \13549 , \13550 );
xnor \U$13299 ( \13552 , \13551 , \7049 );
xor \U$13300 ( \13553 , \13548 , \13552 );
xor \U$13301 ( \13554 , \13528 , \13553 );
and \U$13302 ( \13555 , \6041 , \6991 );
and \U$13303 ( \13556 , \6006 , \6988 );
nor \U$13304 ( \13557 , \13555 , \13556 );
xnor \U$13305 ( \13558 , \13557 , \6985 );
and \U$13306 ( \13559 , \6057 , \7006 );
and \U$13307 ( \13560 , \6029 , \7004 );
nor \U$13308 ( \13561 , \13559 , \13560 );
xnor \U$13309 ( \13562 , \13561 , \7012 );
and \U$13310 ( \13563 , \13558 , \13562 );
and \U$13311 ( \13564 , \6065 , \7026 );
and \U$13312 ( \13565 , \6048 , \7024 );
nor \U$13313 ( \13566 , \13564 , \13565 );
xnor \U$13314 ( \13567 , \13566 , \7032 );
and \U$13315 ( \13568 , \13562 , \13567 );
and \U$13316 ( \13569 , \13558 , \13567 );
or \U$13317 ( \13570 , \13563 , \13568 , \13569 );
xor \U$13318 ( \13571 , \13544 , \13546 );
and \U$13319 ( \13572 , \13570 , \13571 );
xor \U$13320 ( \13573 , \7049 , \13532 );
xor \U$13321 ( \13574 , \13573 , \13537 );
and \U$13322 ( \13575 , \13571 , \13574 );
and \U$13323 ( \13576 , \13570 , \13574 );
or \U$13324 ( \13577 , \13572 , \13575 , \13576 );
nor \U$13325 ( \13578 , \13554 , \13577 );
and \U$13326 ( \13579 , \13540 , \13547 );
and \U$13327 ( \13580 , \13547 , \13552 );
and \U$13328 ( \13581 , \13540 , \13552 );
or \U$13329 ( \13582 , \13579 , \13580 , \13581 );
and \U$13330 ( \13583 , \13518 , \13522 );
and \U$13331 ( \13584 , \13522 , \13527 );
and \U$13332 ( \13585 , \13518 , \13527 );
or \U$13333 ( \13586 , \13583 , \13584 , \13585 );
and \U$13334 ( \13587 , \6029 , \7026 );
and \U$13335 ( \13588 , \6041 , \7024 );
nor \U$13336 ( \13589 , \13587 , \13588 );
xnor \U$13337 ( \13590 , \13589 , \7032 );
and \U$13338 ( \13591 , \6048 , \7043 );
and \U$13339 ( \13592 , \6057 , \7041 );
nor \U$13340 ( \13593 , \13591 , \13592 );
xnor \U$13341 ( \13594 , \13593 , \7049 );
xor \U$13342 ( \13595 , \13590 , \13594 );
nand \U$13343 ( \13596 , \6065 , \7059 );
xnor \U$13344 ( \13597 , \13596 , \7067 );
xor \U$13345 ( \13598 , \13595 , \13597 );
xor \U$13346 ( \13599 , \13586 , \13598 );
and \U$13347 ( \13600 , \5986 , \6991 );
and \U$13348 ( \13601 , \5998 , \6988 );
nor \U$13349 ( \13602 , \13600 , \13601 );
xnor \U$13350 ( \13603 , \13602 , \6985 );
xor \U$13351 ( \13604 , \7067 , \13603 );
and \U$13352 ( \13605 , \6006 , \7006 );
and \U$13353 ( \13606 , \6018 , \7004 );
nor \U$13354 ( \13607 , \13605 , \13606 );
xnor \U$13355 ( \13608 , \13607 , \7012 );
xor \U$13356 ( \13609 , \13604 , \13608 );
xor \U$13357 ( \13610 , \13599 , \13609 );
xor \U$13358 ( \13611 , \13582 , \13610 );
and \U$13359 ( \13612 , \13528 , \13553 );
nor \U$13360 ( \13613 , \13611 , \13612 );
nor \U$13361 ( \13614 , \13578 , \13613 );
and \U$13362 ( \13615 , \13586 , \13598 );
and \U$13363 ( \13616 , \13598 , \13609 );
and \U$13364 ( \13617 , \13586 , \13609 );
or \U$13365 ( \13618 , \13615 , \13616 , \13617 );
and \U$13366 ( \13619 , \6065 , \7061 );
and \U$13367 ( \13620 , \6048 , \7059 );
nor \U$13368 ( \13621 , \13619 , \13620 );
xnor \U$13369 ( \13622 , \13621 , \7067 );
and \U$13370 ( \13623 , \5998 , \6991 );
and \U$13371 ( \13624 , \5967 , \6988 );
nor \U$13372 ( \13625 , \13623 , \13624 );
xnor \U$13373 ( \13626 , \13625 , \6985 );
and \U$13374 ( \13627 , \6018 , \7006 );
and \U$13375 ( \13628 , \5986 , \7004 );
nor \U$13376 ( \13629 , \13627 , \13628 );
xnor \U$13377 ( \13630 , \13629 , \7012 );
xor \U$13378 ( \13631 , \13626 , \13630 );
and \U$13379 ( \13632 , \6041 , \7026 );
and \U$13380 ( \13633 , \6006 , \7024 );
nor \U$13381 ( \13634 , \13632 , \13633 );
xnor \U$13382 ( \13635 , \13634 , \7032 );
xor \U$13383 ( \13636 , \13631 , \13635 );
xor \U$13384 ( \13637 , \13622 , \13636 );
xor \U$13385 ( \13638 , \13618 , \13637 );
and \U$13386 ( \13639 , \7067 , \13603 );
and \U$13387 ( \13640 , \13603 , \13608 );
and \U$13388 ( \13641 , \7067 , \13608 );
or \U$13389 ( \13642 , \13639 , \13640 , \13641 );
and \U$13390 ( \13643 , \13590 , \13594 );
and \U$13391 ( \13644 , \13594 , \13597 );
and \U$13392 ( \13645 , \13590 , \13597 );
or \U$13393 ( \13646 , \13643 , \13644 , \13645 );
xor \U$13394 ( \13647 , \13642 , \13646 );
and \U$13395 ( \13648 , \6057 , \7043 );
and \U$13396 ( \13649 , \6029 , \7041 );
nor \U$13397 ( \13650 , \13648 , \13649 );
xnor \U$13398 ( \13651 , \13650 , \7049 );
xor \U$13399 ( \13652 , \13647 , \13651 );
xor \U$13400 ( \13653 , \13638 , \13652 );
and \U$13401 ( \13654 , \13582 , \13610 );
nor \U$13402 ( \13655 , \13653 , \13654 );
and \U$13403 ( \13656 , \13626 , \13630 );
and \U$13404 ( \13657 , \13630 , \13635 );
and \U$13405 ( \13658 , \13626 , \13635 );
or \U$13406 ( \13659 , \13656 , \13657 , \13658 );
nand \U$13407 ( \13660 , \6065 , \7080 );
xnor \U$13408 ( \13661 , \13660 , \7088 );
xor \U$13409 ( \13662 , \13659 , \13661 );
and \U$13410 ( \13663 , \6006 , \7026 );
and \U$13411 ( \13664 , \6018 , \7024 );
nor \U$13412 ( \13665 , \13663 , \13664 );
xnor \U$13413 ( \13666 , \13665 , \7032 );
and \U$13414 ( \13667 , \6029 , \7043 );
and \U$13415 ( \13668 , \6041 , \7041 );
nor \U$13416 ( \13669 , \13667 , \13668 );
xnor \U$13417 ( \13670 , \13669 , \7049 );
xor \U$13418 ( \13671 , \13666 , \13670 );
and \U$13419 ( \13672 , \6048 , \7061 );
and \U$13420 ( \13673 , \6057 , \7059 );
nor \U$13421 ( \13674 , \13672 , \13673 );
xnor \U$13422 ( \13675 , \13674 , \7067 );
xor \U$13423 ( \13676 , \13671 , \13675 );
xor \U$13424 ( \13677 , \13662 , \13676 );
and \U$13425 ( \13678 , \13642 , \13646 );
and \U$13426 ( \13679 , \13646 , \13651 );
and \U$13427 ( \13680 , \13642 , \13651 );
or \U$13428 ( \13681 , \13678 , \13679 , \13680 );
and \U$13429 ( \13682 , \13622 , \13636 );
xor \U$13430 ( \13683 , \13681 , \13682 );
and \U$13431 ( \13684 , \5967 , \6991 );
and \U$13432 ( \13685 , \5979 , \6988 );
nor \U$13433 ( \13686 , \13684 , \13685 );
xnor \U$13434 ( \13687 , \13686 , \6985 );
xor \U$13435 ( \13688 , \7088 , \13687 );
and \U$13436 ( \13689 , \5986 , \7006 );
and \U$13437 ( \13690 , \5998 , \7004 );
nor \U$13438 ( \13691 , \13689 , \13690 );
xnor \U$13439 ( \13692 , \13691 , \7012 );
xor \U$13440 ( \13693 , \13688 , \13692 );
xor \U$13441 ( \13694 , \13683 , \13693 );
xor \U$13442 ( \13695 , \13677 , \13694 );
and \U$13443 ( \13696 , \13618 , \13637 );
and \U$13444 ( \13697 , \13637 , \13652 );
and \U$13445 ( \13698 , \13618 , \13652 );
or \U$13446 ( \13699 , \13696 , \13697 , \13698 );
nor \U$13447 ( \13700 , \13695 , \13699 );
nor \U$13448 ( \13701 , \13655 , \13700 );
nand \U$13449 ( \13702 , \13614 , \13701 );
and \U$13450 ( \13703 , \13681 , \13682 );
and \U$13451 ( \13704 , \13682 , \13693 );
and \U$13452 ( \13705 , \13681 , \13693 );
or \U$13453 ( \13706 , \13703 , \13704 , \13705 );
and \U$13454 ( \13707 , \13659 , \13661 );
and \U$13455 ( \13708 , \13661 , \13676 );
and \U$13456 ( \13709 , \13659 , \13676 );
or \U$13457 ( \13710 , \13707 , \13708 , \13709 );
xor \U$13458 ( \13711 , \12379 , \12383 );
xor \U$13459 ( \13712 , \13711 , \12388 );
xor \U$13460 ( \13713 , \13710 , \13712 );
and \U$13461 ( \13714 , \7088 , \13687 );
and \U$13462 ( \13715 , \13687 , \13692 );
and \U$13463 ( \13716 , \7088 , \13692 );
or \U$13464 ( \13717 , \13714 , \13715 , \13716 );
and \U$13465 ( \13718 , \13666 , \13670 );
and \U$13466 ( \13719 , \13670 , \13675 );
and \U$13467 ( \13720 , \13666 , \13675 );
or \U$13468 ( \13721 , \13718 , \13719 , \13720 );
xor \U$13469 ( \13722 , \13717 , \13721 );
xor \U$13470 ( \13723 , \12395 , \12399 );
xor \U$13471 ( \13724 , \13723 , \12404 );
xor \U$13472 ( \13725 , \13722 , \13724 );
xor \U$13473 ( \13726 , \13713 , \13725 );
xor \U$13474 ( \13727 , \13706 , \13726 );
and \U$13475 ( \13728 , \13677 , \13694 );
nor \U$13476 ( \13729 , \13727 , \13728 );
and \U$13477 ( \13730 , \13710 , \13712 );
and \U$13478 ( \13731 , \13712 , \13725 );
and \U$13479 ( \13732 , \13710 , \13725 );
or \U$13480 ( \13733 , \13730 , \13731 , \13732 );
and \U$13481 ( \13734 , \13717 , \13721 );
and \U$13482 ( \13735 , \13721 , \13724 );
and \U$13483 ( \13736 , \13717 , \13724 );
or \U$13484 ( \13737 , \13734 , \13735 , \13736 );
xor \U$13485 ( \13738 , \12417 , \12419 );
xor \U$13486 ( \13739 , \13738 , \12422 );
xor \U$13487 ( \13740 , \13737 , \13739 );
xor \U$13488 ( \13741 , \12391 , \12407 );
xor \U$13489 ( \13742 , \13741 , \12412 );
xor \U$13490 ( \13743 , \13740 , \13742 );
xor \U$13491 ( \13744 , \13733 , \13743 );
and \U$13492 ( \13745 , \13706 , \13726 );
nor \U$13493 ( \13746 , \13744 , \13745 );
nor \U$13494 ( \13747 , \13729 , \13746 );
and \U$13495 ( \13748 , \13737 , \13739 );
and \U$13496 ( \13749 , \13739 , \13742 );
and \U$13497 ( \13750 , \13737 , \13742 );
or \U$13498 ( \13751 , \13748 , \13749 , \13750 );
xor \U$13499 ( \13752 , \12433 , \12435 );
xor \U$13500 ( \13753 , \13751 , \13752 );
xor \U$13501 ( \13754 , \12415 , \12425 );
xor \U$13502 ( \13755 , \13754 , \12428 );
xor \U$13503 ( \13756 , \13753 , \13755 );
and \U$13504 ( \13757 , \13733 , \13743 );
nor \U$13505 ( \13758 , \13756 , \13757 );
xor \U$13506 ( \13759 , \12431 , \12436 );
xor \U$13507 ( \13760 , \13759 , \12439 );
and \U$13508 ( \13761 , \13751 , \13752 );
and \U$13509 ( \13762 , \13752 , \13755 );
and \U$13510 ( \13763 , \13751 , \13755 );
or \U$13511 ( \13764 , \13761 , \13762 , \13763 );
nor \U$13512 ( \13765 , \13760 , \13764 );
nor \U$13513 ( \13766 , \13758 , \13765 );
nand \U$13514 ( \13767 , \13747 , \13766 );
nor \U$13515 ( \13768 , \13702 , \13767 );
and \U$13516 ( \13769 , \6057 , \6991 );
and \U$13517 ( \13770 , \6029 , \6988 );
nor \U$13518 ( \13771 , \13769 , \13770 );
xnor \U$13519 ( \13772 , \13771 , \6985 );
and \U$13520 ( \13773 , \6065 , \7006 );
and \U$13521 ( \13774 , \6048 , \7004 );
nor \U$13522 ( \13775 , \13773 , \13774 );
xnor \U$13523 ( \13776 , \13775 , \7012 );
xor \U$13524 ( \13777 , \13772 , \13776 );
and \U$13525 ( \13778 , \6048 , \6991 );
and \U$13526 ( \13779 , \6057 , \6988 );
nor \U$13527 ( \13780 , \13778 , \13779 );
xnor \U$13528 ( \13781 , \13780 , \6985 );
and \U$13529 ( \13782 , \13781 , \7012 );
nor \U$13530 ( \13783 , \13777 , \13782 );
nand \U$13531 ( \13784 , \6065 , \7024 );
xnor \U$13532 ( \13785 , \13784 , \7032 );
and \U$13533 ( \13786 , \6029 , \6991 );
and \U$13534 ( \13787 , \6041 , \6988 );
nor \U$13535 ( \13788 , \13786 , \13787 );
xnor \U$13536 ( \13789 , \13788 , \6985 );
xor \U$13537 ( \13790 , \7032 , \13789 );
and \U$13538 ( \13791 , \6048 , \7006 );
and \U$13539 ( \13792 , \6057 , \7004 );
nor \U$13540 ( \13793 , \13791 , \13792 );
xnor \U$13541 ( \13794 , \13793 , \7012 );
xor \U$13542 ( \13795 , \13790 , \13794 );
xor \U$13543 ( \13796 , \13785 , \13795 );
and \U$13544 ( \13797 , \13772 , \13776 );
nor \U$13545 ( \13798 , \13796 , \13797 );
nor \U$13546 ( \13799 , \13783 , \13798 );
and \U$13547 ( \13800 , \7032 , \13789 );
and \U$13548 ( \13801 , \13789 , \13794 );
and \U$13549 ( \13802 , \7032 , \13794 );
or \U$13550 ( \13803 , \13800 , \13801 , \13802 );
xor \U$13551 ( \13804 , \13558 , \13562 );
xor \U$13552 ( \13805 , \13804 , \13567 );
xor \U$13553 ( \13806 , \13803 , \13805 );
and \U$13554 ( \13807 , \13785 , \13795 );
nor \U$13555 ( \13808 , \13806 , \13807 );
xor \U$13556 ( \13809 , \13570 , \13571 );
xor \U$13557 ( \13810 , \13809 , \13574 );
and \U$13558 ( \13811 , \13803 , \13805 );
nor \U$13559 ( \13812 , \13810 , \13811 );
nor \U$13560 ( \13813 , \13808 , \13812 );
nand \U$13561 ( \13814 , \13799 , \13813 );
xor \U$13562 ( \13815 , \13781 , \7012 );
nand \U$13563 ( \13816 , \6065 , \7004 );
xnor \U$13564 ( \13817 , \13816 , \7012 );
nor \U$13565 ( \13818 , \13815 , \13817 );
and \U$13566 ( \13819 , \6065 , \6991 );
and \U$13567 ( \13820 , \6048 , \6988 );
nor \U$13568 ( \13821 , \13819 , \13820 );
xnor \U$13569 ( \13822 , \13821 , \6985 );
nand \U$13570 ( \13823 , \6065 , \6988 );
xnor \U$13571 ( \13824 , \13823 , \6985 );
and \U$13572 ( \13825 , \13824 , \6985 );
nand \U$13573 ( \13826 , \13822 , \13825 );
or \U$13574 ( \13827 , \13818 , \13826 );
nand \U$13575 ( \13828 , \13815 , \13817 );
nand \U$13576 ( \13829 , \13827 , \13828 );
not \U$13577 ( \13830 , \13829 );
or \U$13578 ( \13831 , \13814 , \13830 );
nand \U$13579 ( \13832 , \13777 , \13782 );
or \U$13580 ( \13833 , \13798 , \13832 );
nand \U$13581 ( \13834 , \13796 , \13797 );
nand \U$13582 ( \13835 , \13833 , \13834 );
and \U$13583 ( \13836 , \13813 , \13835 );
nand \U$13584 ( \13837 , \13806 , \13807 );
or \U$13585 ( \13838 , \13812 , \13837 );
nand \U$13586 ( \13839 , \13810 , \13811 );
nand \U$13587 ( \13840 , \13838 , \13839 );
nor \U$13588 ( \13841 , \13836 , \13840 );
nand \U$13589 ( \13842 , \13831 , \13841 );
and \U$13590 ( \13843 , \13768 , \13842 );
nand \U$13591 ( \13844 , \13554 , \13577 );
or \U$13592 ( \13845 , \13613 , \13844 );
nand \U$13593 ( \13846 , \13611 , \13612 );
nand \U$13594 ( \13847 , \13845 , \13846 );
and \U$13595 ( \13848 , \13701 , \13847 );
nand \U$13596 ( \13849 , \13653 , \13654 );
or \U$13597 ( \13850 , \13700 , \13849 );
nand \U$13598 ( \13851 , \13695 , \13699 );
nand \U$13599 ( \13852 , \13850 , \13851 );
nor \U$13600 ( \13853 , \13848 , \13852 );
or \U$13601 ( \13854 , \13767 , \13853 );
nand \U$13602 ( \13855 , \13727 , \13728 );
or \U$13603 ( \13856 , \13746 , \13855 );
nand \U$13604 ( \13857 , \13744 , \13745 );
nand \U$13605 ( \13858 , \13856 , \13857 );
and \U$13606 ( \13859 , \13766 , \13858 );
nand \U$13607 ( \13860 , \13756 , \13757 );
or \U$13608 ( \13861 , \13765 , \13860 );
nand \U$13609 ( \13862 , \13760 , \13764 );
nand \U$13610 ( \13863 , \13861 , \13862 );
nor \U$13611 ( \13864 , \13859 , \13863 );
nand \U$13612 ( \13865 , \13854 , \13864 );
nor \U$13613 ( \13866 , \13843 , \13865 );
or \U$13614 ( \13867 , \13514 , \13866 );
nand \U$13615 ( \13868 , \12375 , \12442 );
or \U$13616 ( \13869 , \12518 , \13868 );
nand \U$13617 ( \13870 , \12513 , \12517 );
nand \U$13618 ( \13871 , \13869 , \13870 );
and \U$13619 ( \13872 , \12686 , \13871 );
nand \U$13620 ( \13873 , \12595 , \12599 );
or \U$13621 ( \13874 , \12685 , \13873 );
nand \U$13622 ( \13875 , \12683 , \12684 );
nand \U$13623 ( \13876 , \13874 , \13875 );
nor \U$13624 ( \13877 , \13872 , \13876 );
or \U$13625 ( \13878 , \13082 , \13877 );
nand \U$13626 ( \13879 , \12776 , \12777 );
or \U$13627 ( \13880 , \12873 , \13879 );
nand \U$13628 ( \13881 , \12868 , \12872 );
nand \U$13629 ( \13882 , \13880 , \13881 );
and \U$13630 ( \13883 , \13081 , \13882 );
nand \U$13631 ( \13884 , \12970 , \12974 );
or \U$13632 ( \13885 , \13080 , \13884 );
nand \U$13633 ( \13886 , \13075 , \13079 );
nand \U$13634 ( \13887 , \13885 , \13886 );
nor \U$13635 ( \13888 , \13883 , \13887 );
nand \U$13636 ( \13889 , \13878 , \13888 );
and \U$13637 ( \13890 , \13513 , \13889 );
nand \U$13638 ( \13891 , \13189 , \13193 );
or \U$13639 ( \13892 , \13309 , \13891 );
nand \U$13640 ( \13893 , \13304 , \13308 );
nand \U$13641 ( \13894 , \13892 , \13893 );
and \U$13642 ( \13895 , \13429 , \13894 );
nand \U$13643 ( \13896 , \13378 , \13382 );
or \U$13644 ( \13897 , \13428 , \13896 );
nand \U$13645 ( \13898 , \13423 , \13427 );
nand \U$13646 ( \13899 , \13897 , \13898 );
nor \U$13647 ( \13900 , \13895 , \13899 );
or \U$13648 ( \13901 , \13512 , \13900 );
nand \U$13649 ( \13902 , \13461 , \13462 );
or \U$13650 ( \13903 , \13488 , \13902 );
nand \U$13651 ( \13904 , \13486 , \13487 );
nand \U$13652 ( \13905 , \13903 , \13904 );
and \U$13653 ( \13906 , \13511 , \13905 );
nand \U$13654 ( \13907 , \13498 , \13502 );
or \U$13655 ( \13908 , \13510 , \13907 );
nand \U$13656 ( \13909 , \13505 , \13509 );
nand \U$13657 ( \13910 , \13908 , \13909 );
nor \U$13658 ( \13911 , \13906 , \13910 );
nand \U$13659 ( \13912 , \13901 , \13911 );
nor \U$13660 ( \13913 , \13890 , \13912 );
nand \U$13661 ( \13914 , \13867 , \13913 );
and \U$13662 ( \13915 , \12202 , \13914 );
nand \U$13663 ( \13916 , \7766 , \7886 );
or \U$13664 ( \13917 , \8041 , \13916 );
nand \U$13665 ( \13918 , \8036 , \8040 );
nand \U$13666 ( \13919 , \13917 , \13918 );
and \U$13667 ( \13920 , \8360 , \13919 );
nand \U$13668 ( \13921 , \8195 , \8199 );
or \U$13669 ( \13922 , \8359 , \13921 );
nand \U$13670 ( \13923 , \8354 , \8358 );
nand \U$13671 ( \13924 , \13922 , \13923 );
nor \U$13672 ( \13925 , \13920 , \13924 );
or \U$13673 ( \13926 , \9009 , \13925 );
nand \U$13674 ( \13927 , \8516 , \8520 );
or \U$13675 ( \13928 , \8682 , \13927 );
nand \U$13676 ( \13929 , \8677 , \8681 );
nand \U$13677 ( \13930 , \13928 , \13929 );
and \U$13678 ( \13931 , \9008 , \13930 );
nand \U$13679 ( \13932 , \8841 , \8845 );
or \U$13680 ( \13933 , \9007 , \13932 );
nand \U$13681 ( \13934 , \9002 , \9006 );
nand \U$13682 ( \13935 , \13933 , \13934 );
nor \U$13683 ( \13936 , \13931 , \13935 );
nand \U$13684 ( \13937 , \13926 , \13936 );
and \U$13685 ( \13938 , \10313 , \13937 );
nand \U$13686 ( \13939 , \9168 , \9172 );
or \U$13687 ( \13940 , \9334 , \13939 );
nand \U$13688 ( \13941 , \9329 , \9333 );
nand \U$13689 ( \13942 , \13940 , \13941 );
and \U$13690 ( \13943 , \9660 , \13942 );
nand \U$13691 ( \13944 , \9493 , \9497 );
or \U$13692 ( \13945 , \9659 , \13944 );
nand \U$13693 ( \13946 , \9654 , \9658 );
nand \U$13694 ( \13947 , \13945 , \13946 );
nor \U$13695 ( \13948 , \13943 , \13947 );
or \U$13696 ( \13949 , \10312 , \13948 );
nand \U$13697 ( \13950 , \9819 , \9823 );
or \U$13698 ( \13951 , \9985 , \13950 );
nand \U$13699 ( \13952 , \9980 , \9984 );
nand \U$13700 ( \13953 , \13951 , \13952 );
and \U$13701 ( \13954 , \10311 , \13953 );
nand \U$13702 ( \13955 , \10144 , \10148 );
or \U$13703 ( \13956 , \10310 , \13955 );
nand \U$13704 ( \13957 , \10305 , \10309 );
nand \U$13705 ( \13958 , \13956 , \13957 );
nor \U$13706 ( \13959 , \13954 , \13958 );
nand \U$13707 ( \13960 , \13949 , \13959 );
nor \U$13708 ( \13961 , \13938 , \13960 );
or \U$13709 ( \13962 , \12201 , \13961 );
nand \U$13710 ( \13963 , \10472 , \10476 );
or \U$13711 ( \13964 , \10638 , \13963 );
nand \U$13712 ( \13965 , \10633 , \10637 );
nand \U$13713 ( \13966 , \13964 , \13965 );
and \U$13714 ( \13967 , \10964 , \13966 );
nand \U$13715 ( \13968 , \10797 , \10801 );
or \U$13716 ( \13969 , \10963 , \13968 );
nand \U$13717 ( \13970 , \10958 , \10962 );
nand \U$13718 ( \13971 , \13969 , \13970 );
nor \U$13719 ( \13972 , \13967 , \13971 );
or \U$13720 ( \13973 , \11616 , \13972 );
nand \U$13721 ( \13974 , \11123 , \11127 );
or \U$13722 ( \13975 , \11289 , \13974 );
nand \U$13723 ( \13976 , \11284 , \11288 );
nand \U$13724 ( \13977 , \13975 , \13976 );
and \U$13725 ( \13978 , \11615 , \13977 );
nand \U$13726 ( \13979 , \11448 , \11452 );
or \U$13727 ( \13980 , \11614 , \13979 );
nand \U$13728 ( \13981 , \11609 , \11613 );
nand \U$13729 ( \13982 , \13980 , \13981 );
nor \U$13730 ( \13983 , \13978 , \13982 );
nand \U$13731 ( \13984 , \13973 , \13983 );
and \U$13732 ( \13985 , \12200 , \13984 );
nand \U$13733 ( \13986 , \11775 , \11779 );
or \U$13734 ( \13987 , \11941 , \13986 );
nand \U$13735 ( \13988 , \11936 , \11940 );
nand \U$13736 ( \13989 , \13987 , \13988 );
and \U$13737 ( \13990 , \12106 , \13989 );
nand \U$13738 ( \13991 , \12035 , \12039 );
or \U$13739 ( \13992 , \12105 , \13991 );
nand \U$13740 ( \13993 , \12100 , \12104 );
nand \U$13741 ( \13994 , \13992 , \13993 );
nor \U$13742 ( \13995 , \13990 , \13994 );
or \U$13743 ( \13996 , \12199 , \13995 );
nand \U$13744 ( \13997 , \12144 , \12148 );
or \U$13745 ( \13998 , \12174 , \13997 );
nand \U$13746 ( \13999 , \12169 , \12173 );
nand \U$13747 ( \14000 , \13998 , \13999 );
and \U$13748 ( \14001 , \12198 , \14000 );
nand \U$13749 ( \14002 , \12185 , \12189 );
or \U$13750 ( \14003 , \12197 , \14002 );
nand \U$13751 ( \14004 , \12192 , \12196 );
nand \U$13752 ( \14005 , \14003 , \14004 );
nor \U$13753 ( \14006 , \14001 , \14005 );
nand \U$13754 ( \14007 , \13996 , \14006 );
nor \U$13755 ( \14008 , \13985 , \14007 );
nand \U$13756 ( \14009 , \13962 , \14008 );
nor \U$13757 ( \14010 , \13915 , \14009 );
not \U$13758 ( \14011 , \14010 );
xnor \U$13759 ( \14012 , \6982 , \14011 );
buf g36c1_GF_PartitionCandidate( \14013_nG36c1 , \14012 );
buf \U$13760 ( \14014 , \14013_nG36c1 );
not \U$13761 ( \14015 , \12197 );
nand \U$13762 ( \14016 , \14004 , \14015 );
nor \U$13763 ( \14017 , \13510 , \7887 );
nor \U$13764 ( \14018 , \8041 , \8200 );
nand \U$13765 ( \14019 , \14017 , \14018 );
nor \U$13766 ( \14020 , \8359 , \8521 );
nor \U$13767 ( \14021 , \8682 , \8846 );
nand \U$13768 ( \14022 , \14020 , \14021 );
nor \U$13769 ( \14023 , \14019 , \14022 );
nor \U$13770 ( \14024 , \9007 , \9173 );
nor \U$13771 ( \14025 , \9334 , \9498 );
nand \U$13772 ( \14026 , \14024 , \14025 );
nor \U$13773 ( \14027 , \9659 , \9824 );
nor \U$13774 ( \14028 , \9985 , \10149 );
nand \U$13775 ( \14029 , \14027 , \14028 );
nor \U$13776 ( \14030 , \14026 , \14029 );
nand \U$13777 ( \14031 , \14023 , \14030 );
nor \U$13778 ( \14032 , \10310 , \10477 );
nor \U$13779 ( \14033 , \10638 , \10802 );
nand \U$13780 ( \14034 , \14032 , \14033 );
nor \U$13781 ( \14035 , \10963 , \11128 );
nor \U$13782 ( \14036 , \11289 , \11453 );
nand \U$13783 ( \14037 , \14035 , \14036 );
nor \U$13784 ( \14038 , \14034 , \14037 );
nor \U$13785 ( \14039 , \11614 , \11780 );
nor \U$13786 ( \14040 , \11941 , \12040 );
nand \U$13787 ( \14041 , \14039 , \14040 );
nor \U$13788 ( \14042 , \12105 , \12149 );
nor \U$13789 ( \14043 , \12174 , \12190 );
nand \U$13790 ( \14044 , \14042 , \14043 );
nor \U$13791 ( \14045 , \14041 , \14044 );
nand \U$13792 ( \14046 , \14038 , \14045 );
nor \U$13793 ( \14047 , \14031 , \14046 );
nor \U$13794 ( \14048 , \13765 , \12443 );
nor \U$13795 ( \14049 , \12518 , \12600 );
nand \U$13796 ( \14050 , \14048 , \14049 );
nor \U$13797 ( \14051 , \12685 , \12778 );
nor \U$13798 ( \14052 , \12873 , \12975 );
nand \U$13799 ( \14053 , \14051 , \14052 );
nor \U$13800 ( \14054 , \14050 , \14053 );
nor \U$13801 ( \14055 , \13080 , \13194 );
nor \U$13802 ( \14056 , \13309 , \13383 );
nand \U$13803 ( \14057 , \14055 , \14056 );
nor \U$13804 ( \14058 , \13428 , \13463 );
nor \U$13805 ( \14059 , \13488 , \13503 );
nand \U$13806 ( \14060 , \14058 , \14059 );
nor \U$13807 ( \14061 , \14057 , \14060 );
nand \U$13808 ( \14062 , \14054 , \14061 );
nor \U$13809 ( \14063 , \13812 , \13578 );
nor \U$13810 ( \14064 , \13613 , \13655 );
nand \U$13811 ( \14065 , \14063 , \14064 );
nor \U$13812 ( \14066 , \13700 , \13729 );
nor \U$13813 ( \14067 , \13746 , \13758 );
nand \U$13814 ( \14068 , \14066 , \14067 );
nor \U$13815 ( \14069 , \14065 , \14068 );
nor \U$13816 ( \14070 , \13818 , \13783 );
nor \U$13817 ( \14071 , \13798 , \13808 );
nand \U$13818 ( \14072 , \14070 , \14071 );
or \U$13819 ( \14073 , \14072 , \13826 );
or \U$13820 ( \14074 , \13783 , \13828 );
nand \U$13821 ( \14075 , \14074 , \13832 );
and \U$13822 ( \14076 , \14071 , \14075 );
or \U$13823 ( \14077 , \13808 , \13834 );
nand \U$13824 ( \14078 , \14077 , \13837 );
nor \U$13825 ( \14079 , \14076 , \14078 );
nand \U$13826 ( \14080 , \14073 , \14079 );
and \U$13827 ( \14081 , \14069 , \14080 );
or \U$13828 ( \14082 , \13578 , \13839 );
nand \U$13829 ( \14083 , \14082 , \13844 );
and \U$13830 ( \14084 , \14064 , \14083 );
or \U$13831 ( \14085 , \13655 , \13846 );
nand \U$13832 ( \14086 , \14085 , \13849 );
nor \U$13833 ( \14087 , \14084 , \14086 );
or \U$13834 ( \14088 , \14068 , \14087 );
or \U$13835 ( \14089 , \13729 , \13851 );
nand \U$13836 ( \14090 , \14089 , \13855 );
and \U$13837 ( \14091 , \14067 , \14090 );
or \U$13838 ( \14092 , \13758 , \13857 );
nand \U$13839 ( \14093 , \14092 , \13860 );
nor \U$13840 ( \14094 , \14091 , \14093 );
nand \U$13841 ( \14095 , \14088 , \14094 );
nor \U$13842 ( \14096 , \14081 , \14095 );
or \U$13843 ( \14097 , \14062 , \14096 );
or \U$13844 ( \14098 , \12443 , \13862 );
nand \U$13845 ( \14099 , \14098 , \13868 );
and \U$13846 ( \14100 , \14049 , \14099 );
or \U$13847 ( \14101 , \12600 , \13870 );
nand \U$13848 ( \14102 , \14101 , \13873 );
nor \U$13849 ( \14103 , \14100 , \14102 );
or \U$13850 ( \14104 , \14053 , \14103 );
or \U$13851 ( \14105 , \12778 , \13875 );
nand \U$13852 ( \14106 , \14105 , \13879 );
and \U$13853 ( \14107 , \14052 , \14106 );
or \U$13854 ( \14108 , \12975 , \13881 );
nand \U$13855 ( \14109 , \14108 , \13884 );
nor \U$13856 ( \14110 , \14107 , \14109 );
nand \U$13857 ( \14111 , \14104 , \14110 );
and \U$13858 ( \14112 , \14061 , \14111 );
or \U$13859 ( \14113 , \13194 , \13886 );
nand \U$13860 ( \14114 , \14113 , \13891 );
and \U$13861 ( \14115 , \14056 , \14114 );
or \U$13862 ( \14116 , \13383 , \13893 );
nand \U$13863 ( \14117 , \14116 , \13896 );
nor \U$13864 ( \14118 , \14115 , \14117 );
or \U$13865 ( \14119 , \14060 , \14118 );
or \U$13866 ( \14120 , \13463 , \13898 );
nand \U$13867 ( \14121 , \14120 , \13902 );
and \U$13868 ( \14122 , \14059 , \14121 );
or \U$13869 ( \14123 , \13503 , \13904 );
nand \U$13870 ( \14124 , \14123 , \13907 );
nor \U$13871 ( \14125 , \14122 , \14124 );
nand \U$13872 ( \14126 , \14119 , \14125 );
nor \U$13873 ( \14127 , \14112 , \14126 );
nand \U$13874 ( \14128 , \14097 , \14127 );
and \U$13875 ( \14129 , \14047 , \14128 );
or \U$13876 ( \14130 , \7887 , \13909 );
nand \U$13877 ( \14131 , \14130 , \13916 );
and \U$13878 ( \14132 , \14018 , \14131 );
or \U$13879 ( \14133 , \8200 , \13918 );
nand \U$13880 ( \14134 , \14133 , \13921 );
nor \U$13881 ( \14135 , \14132 , \14134 );
or \U$13882 ( \14136 , \14022 , \14135 );
or \U$13883 ( \14137 , \8521 , \13923 );
nand \U$13884 ( \14138 , \14137 , \13927 );
and \U$13885 ( \14139 , \14021 , \14138 );
or \U$13886 ( \14140 , \8846 , \13929 );
nand \U$13887 ( \14141 , \14140 , \13932 );
nor \U$13888 ( \14142 , \14139 , \14141 );
nand \U$13889 ( \14143 , \14136 , \14142 );
and \U$13890 ( \14144 , \14030 , \14143 );
or \U$13891 ( \14145 , \9173 , \13934 );
nand \U$13892 ( \14146 , \14145 , \13939 );
and \U$13893 ( \14147 , \14025 , \14146 );
or \U$13894 ( \14148 , \9498 , \13941 );
nand \U$13895 ( \14149 , \14148 , \13944 );
nor \U$13896 ( \14150 , \14147 , \14149 );
or \U$13897 ( \14151 , \14029 , \14150 );
or \U$13898 ( \14152 , \9824 , \13946 );
nand \U$13899 ( \14153 , \14152 , \13950 );
and \U$13900 ( \14154 , \14028 , \14153 );
or \U$13901 ( \14155 , \10149 , \13952 );
nand \U$13902 ( \14156 , \14155 , \13955 );
nor \U$13903 ( \14157 , \14154 , \14156 );
nand \U$13904 ( \14158 , \14151 , \14157 );
nor \U$13905 ( \14159 , \14144 , \14158 );
or \U$13906 ( \14160 , \14046 , \14159 );
or \U$13907 ( \14161 , \10477 , \13957 );
nand \U$13908 ( \14162 , \14161 , \13963 );
and \U$13909 ( \14163 , \14033 , \14162 );
or \U$13910 ( \14164 , \10802 , \13965 );
nand \U$13911 ( \14165 , \14164 , \13968 );
nor \U$13912 ( \14166 , \14163 , \14165 );
or \U$13913 ( \14167 , \14037 , \14166 );
or \U$13914 ( \14168 , \11128 , \13970 );
nand \U$13915 ( \14169 , \14168 , \13974 );
and \U$13916 ( \14170 , \14036 , \14169 );
or \U$13917 ( \14171 , \11453 , \13976 );
nand \U$13918 ( \14172 , \14171 , \13979 );
nor \U$13919 ( \14173 , \14170 , \14172 );
nand \U$13920 ( \14174 , \14167 , \14173 );
and \U$13921 ( \14175 , \14045 , \14174 );
or \U$13922 ( \14176 , \11780 , \13981 );
nand \U$13923 ( \14177 , \14176 , \13986 );
and \U$13924 ( \14178 , \14040 , \14177 );
or \U$13925 ( \14179 , \12040 , \13988 );
nand \U$13926 ( \14180 , \14179 , \13991 );
nor \U$13927 ( \14181 , \14178 , \14180 );
or \U$13928 ( \14182 , \14044 , \14181 );
or \U$13929 ( \14183 , \12149 , \13993 );
nand \U$13930 ( \14184 , \14183 , \13997 );
and \U$13931 ( \14185 , \14043 , \14184 );
or \U$13932 ( \14186 , \12190 , \13999 );
nand \U$13933 ( \14187 , \14186 , \14002 );
nor \U$13934 ( \14188 , \14185 , \14187 );
nand \U$13935 ( \14189 , \14182 , \14188 );
nor \U$13936 ( \14190 , \14175 , \14189 );
nand \U$13937 ( \14191 , \14160 , \14190 );
nor \U$13938 ( \14192 , \14129 , \14191 );
not \U$13939 ( \14193 , \14192 );
xnor \U$13940 ( \14194 , \14016 , \14193 );
buf g3776_GF_PartitionCandidate( \14195_nG3776 , \14194 );
buf \U$13941 ( \14196 , \14195_nG3776 );
not \U$13942 ( \14197 , \12190 );
nand \U$13943 ( \14198 , \14002 , \14197 );
nand \U$13944 ( \14199 , \13511 , \8042 );
nand \U$13945 ( \14200 , \8360 , \8683 );
nor \U$13946 ( \14201 , \14199 , \14200 );
nand \U$13947 ( \14202 , \9008 , \9335 );
nand \U$13948 ( \14203 , \9660 , \9986 );
nor \U$13949 ( \14204 , \14202 , \14203 );
nand \U$13950 ( \14205 , \14201 , \14204 );
nand \U$13951 ( \14206 , \10311 , \10639 );
nand \U$13952 ( \14207 , \10964 , \11290 );
nor \U$13953 ( \14208 , \14206 , \14207 );
nand \U$13954 ( \14209 , \11615 , \11942 );
nand \U$13955 ( \14210 , \12106 , \12175 );
nor \U$13956 ( \14211 , \14209 , \14210 );
nand \U$13957 ( \14212 , \14208 , \14211 );
nor \U$13958 ( \14213 , \14205 , \14212 );
nand \U$13959 ( \14214 , \13766 , \12519 );
nand \U$13960 ( \14215 , \12686 , \12874 );
nor \U$13961 ( \14216 , \14214 , \14215 );
nand \U$13962 ( \14217 , \13081 , \13310 );
nand \U$13963 ( \14218 , \13429 , \13489 );
nor \U$13964 ( \14219 , \14217 , \14218 );
nand \U$13965 ( \14220 , \14216 , \14219 );
nand \U$13966 ( \14221 , \13813 , \13614 );
nand \U$13967 ( \14222 , \13701 , \13747 );
nor \U$13968 ( \14223 , \14221 , \14222 );
and \U$13969 ( \14224 , \13799 , \13829 );
nor \U$13970 ( \14225 , \14224 , \13835 );
not \U$13971 ( \14226 , \14225 );
and \U$13972 ( \14227 , \14223 , \14226 );
and \U$13973 ( \14228 , \13614 , \13840 );
nor \U$13974 ( \14229 , \14228 , \13847 );
or \U$13975 ( \14230 , \14222 , \14229 );
and \U$13976 ( \14231 , \13747 , \13852 );
nor \U$13977 ( \14232 , \14231 , \13858 );
nand \U$13978 ( \14233 , \14230 , \14232 );
nor \U$13979 ( \14234 , \14227 , \14233 );
or \U$13980 ( \14235 , \14220 , \14234 );
and \U$13981 ( \14236 , \12519 , \13863 );
nor \U$13982 ( \14237 , \14236 , \13871 );
or \U$13983 ( \14238 , \14215 , \14237 );
and \U$13984 ( \14239 , \12874 , \13876 );
nor \U$13985 ( \14240 , \14239 , \13882 );
nand \U$13986 ( \14241 , \14238 , \14240 );
and \U$13987 ( \14242 , \14219 , \14241 );
and \U$13988 ( \14243 , \13310 , \13887 );
nor \U$13989 ( \14244 , \14243 , \13894 );
or \U$13990 ( \14245 , \14218 , \14244 );
and \U$13991 ( \14246 , \13489 , \13899 );
nor \U$13992 ( \14247 , \14246 , \13905 );
nand \U$13993 ( \14248 , \14245 , \14247 );
nor \U$13994 ( \14249 , \14242 , \14248 );
nand \U$13995 ( \14250 , \14235 , \14249 );
and \U$13996 ( \14251 , \14213 , \14250 );
and \U$13997 ( \14252 , \8042 , \13910 );
nor \U$13998 ( \14253 , \14252 , \13919 );
or \U$13999 ( \14254 , \14200 , \14253 );
and \U$14000 ( \14255 , \8683 , \13924 );
nor \U$14001 ( \14256 , \14255 , \13930 );
nand \U$14002 ( \14257 , \14254 , \14256 );
and \U$14003 ( \14258 , \14204 , \14257 );
and \U$14004 ( \14259 , \9335 , \13935 );
nor \U$14005 ( \14260 , \14259 , \13942 );
or \U$14006 ( \14261 , \14203 , \14260 );
and \U$14007 ( \14262 , \9986 , \13947 );
nor \U$14008 ( \14263 , \14262 , \13953 );
nand \U$14009 ( \14264 , \14261 , \14263 );
nor \U$14010 ( \14265 , \14258 , \14264 );
or \U$14011 ( \14266 , \14212 , \14265 );
and \U$14012 ( \14267 , \10639 , \13958 );
nor \U$14013 ( \14268 , \14267 , \13966 );
or \U$14014 ( \14269 , \14207 , \14268 );
and \U$14015 ( \14270 , \11290 , \13971 );
nor \U$14016 ( \14271 , \14270 , \13977 );
nand \U$14017 ( \14272 , \14269 , \14271 );
and \U$14018 ( \14273 , \14211 , \14272 );
and \U$14019 ( \14274 , \11942 , \13982 );
nor \U$14020 ( \14275 , \14274 , \13989 );
or \U$14021 ( \14276 , \14210 , \14275 );
and \U$14022 ( \14277 , \12175 , \13994 );
nor \U$14023 ( \14278 , \14277 , \14000 );
nand \U$14024 ( \14279 , \14276 , \14278 );
nor \U$14025 ( \14280 , \14273 , \14279 );
nand \U$14026 ( \14281 , \14266 , \14280 );
nor \U$14027 ( \14282 , \14251 , \14281 );
not \U$14028 ( \14283 , \14282 );
xnor \U$14029 ( \14284 , \14198 , \14283 );
buf g37cf_GF_PartitionCandidate( \14285_nG37cf , \14284 );
buf \U$14030 ( \14286 , \14285_nG37cf );
not \U$14031 ( \14287 , \12174 );
nand \U$14032 ( \14288 , \13999 , \14287 );
nand \U$14033 ( \14289 , \14059 , \14017 );
nand \U$14034 ( \14290 , \14018 , \14020 );
nor \U$14035 ( \14291 , \14289 , \14290 );
nand \U$14036 ( \14292 , \14021 , \14024 );
nand \U$14037 ( \14293 , \14025 , \14027 );
nor \U$14038 ( \14294 , \14292 , \14293 );
nand \U$14039 ( \14295 , \14291 , \14294 );
nand \U$14040 ( \14296 , \14028 , \14032 );
nand \U$14041 ( \14297 , \14033 , \14035 );
nor \U$14042 ( \14298 , \14296 , \14297 );
nand \U$14043 ( \14299 , \14036 , \14039 );
nand \U$14044 ( \14300 , \14040 , \14042 );
nor \U$14045 ( \14301 , \14299 , \14300 );
nand \U$14046 ( \14302 , \14298 , \14301 );
nor \U$14047 ( \14303 , \14295 , \14302 );
nand \U$14048 ( \14304 , \14067 , \14048 );
nand \U$14049 ( \14305 , \14049 , \14051 );
nor \U$14050 ( \14306 , \14304 , \14305 );
nand \U$14051 ( \14307 , \14052 , \14055 );
nand \U$14052 ( \14308 , \14056 , \14058 );
nor \U$14053 ( \14309 , \14307 , \14308 );
nand \U$14054 ( \14310 , \14306 , \14309 );
nand \U$14055 ( \14311 , \14071 , \14063 );
nand \U$14056 ( \14312 , \14064 , \14066 );
nor \U$14057 ( \14313 , \14311 , \14312 );
not \U$14058 ( \14314 , \13826 );
and \U$14059 ( \14315 , \14070 , \14314 );
nor \U$14060 ( \14316 , \14315 , \14075 );
not \U$14061 ( \14317 , \14316 );
and \U$14062 ( \14318 , \14313 , \14317 );
and \U$14063 ( \14319 , \14063 , \14078 );
nor \U$14064 ( \14320 , \14319 , \14083 );
or \U$14065 ( \14321 , \14312 , \14320 );
and \U$14066 ( \14322 , \14066 , \14086 );
nor \U$14067 ( \14323 , \14322 , \14090 );
nand \U$14068 ( \14324 , \14321 , \14323 );
nor \U$14069 ( \14325 , \14318 , \14324 );
or \U$14070 ( \14326 , \14310 , \14325 );
and \U$14071 ( \14327 , \14048 , \14093 );
nor \U$14072 ( \14328 , \14327 , \14099 );
or \U$14073 ( \14329 , \14305 , \14328 );
and \U$14074 ( \14330 , \14051 , \14102 );
nor \U$14075 ( \14331 , \14330 , \14106 );
nand \U$14076 ( \14332 , \14329 , \14331 );
and \U$14077 ( \14333 , \14309 , \14332 );
and \U$14078 ( \14334 , \14055 , \14109 );
nor \U$14079 ( \14335 , \14334 , \14114 );
or \U$14080 ( \14336 , \14308 , \14335 );
and \U$14081 ( \14337 , \14058 , \14117 );
nor \U$14082 ( \14338 , \14337 , \14121 );
nand \U$14083 ( \14339 , \14336 , \14338 );
nor \U$14084 ( \14340 , \14333 , \14339 );
nand \U$14085 ( \14341 , \14326 , \14340 );
and \U$14086 ( \14342 , \14303 , \14341 );
and \U$14087 ( \14343 , \14017 , \14124 );
nor \U$14088 ( \14344 , \14343 , \14131 );
or \U$14089 ( \14345 , \14290 , \14344 );
and \U$14090 ( \14346 , \14020 , \14134 );
nor \U$14091 ( \14347 , \14346 , \14138 );
nand \U$14092 ( \14348 , \14345 , \14347 );
and \U$14093 ( \14349 , \14294 , \14348 );
and \U$14094 ( \14350 , \14024 , \14141 );
nor \U$14095 ( \14351 , \14350 , \14146 );
or \U$14096 ( \14352 , \14293 , \14351 );
and \U$14097 ( \14353 , \14027 , \14149 );
nor \U$14098 ( \14354 , \14353 , \14153 );
nand \U$14099 ( \14355 , \14352 , \14354 );
nor \U$14100 ( \14356 , \14349 , \14355 );
or \U$14101 ( \14357 , \14302 , \14356 );
and \U$14102 ( \14358 , \14032 , \14156 );
nor \U$14103 ( \14359 , \14358 , \14162 );
or \U$14104 ( \14360 , \14297 , \14359 );
and \U$14105 ( \14361 , \14035 , \14165 );
nor \U$14106 ( \14362 , \14361 , \14169 );
nand \U$14107 ( \14363 , \14360 , \14362 );
and \U$14108 ( \14364 , \14301 , \14363 );
and \U$14109 ( \14365 , \14039 , \14172 );
nor \U$14110 ( \14366 , \14365 , \14177 );
or \U$14111 ( \14367 , \14300 , \14366 );
and \U$14112 ( \14368 , \14042 , \14180 );
nor \U$14113 ( \14369 , \14368 , \14184 );
nand \U$14114 ( \14370 , \14367 , \14369 );
nor \U$14115 ( \14371 , \14364 , \14370 );
nand \U$14116 ( \14372 , \14357 , \14371 );
nor \U$14117 ( \14373 , \14342 , \14372 );
not \U$14118 ( \14374 , \14373 );
xnor \U$14119 ( \14375 , \14288 , \14374 );
buf g3829_GF_PartitionCandidate( \14376_nG3829 , \14375 );
buf \U$14120 ( \14377 , \14376_nG3829 );
not \U$14121 ( \14378 , \12149 );
nand \U$14122 ( \14379 , \13997 , \14378 );
nor \U$14123 ( \14380 , \13512 , \8361 );
nor \U$14124 ( \14381 , \9009 , \9661 );
nand \U$14125 ( \14382 , \14380 , \14381 );
nor \U$14126 ( \14383 , \10312 , \10965 );
nor \U$14127 ( \14384 , \11616 , \12107 );
nand \U$14128 ( \14385 , \14383 , \14384 );
nor \U$14129 ( \14386 , \14382 , \14385 );
nor \U$14130 ( \14387 , \13767 , \12687 );
nor \U$14131 ( \14388 , \13082 , \13430 );
nand \U$14132 ( \14389 , \14387 , \14388 );
nor \U$14133 ( \14390 , \13814 , \13702 );
and \U$14134 ( \14391 , \14390 , \13829 );
or \U$14135 ( \14392 , \13702 , \13841 );
nand \U$14136 ( \14393 , \14392 , \13853 );
nor \U$14137 ( \14394 , \14391 , \14393 );
or \U$14138 ( \14395 , \14389 , \14394 );
or \U$14139 ( \14396 , \12687 , \13864 );
nand \U$14140 ( \14397 , \14396 , \13877 );
and \U$14141 ( \14398 , \14388 , \14397 );
or \U$14142 ( \14399 , \13430 , \13888 );
nand \U$14143 ( \14400 , \14399 , \13900 );
nor \U$14144 ( \14401 , \14398 , \14400 );
nand \U$14145 ( \14402 , \14395 , \14401 );
and \U$14146 ( \14403 , \14386 , \14402 );
or \U$14147 ( \14404 , \8361 , \13911 );
nand \U$14148 ( \14405 , \14404 , \13925 );
and \U$14149 ( \14406 , \14381 , \14405 );
or \U$14150 ( \14407 , \9661 , \13936 );
nand \U$14151 ( \14408 , \14407 , \13948 );
nor \U$14152 ( \14409 , \14406 , \14408 );
or \U$14153 ( \14410 , \14385 , \14409 );
or \U$14154 ( \14411 , \10965 , \13959 );
nand \U$14155 ( \14412 , \14411 , \13972 );
and \U$14156 ( \14413 , \14384 , \14412 );
or \U$14157 ( \14414 , \12107 , \13983 );
nand \U$14158 ( \14415 , \14414 , \13995 );
nor \U$14159 ( \14416 , \14413 , \14415 );
nand \U$14160 ( \14417 , \14410 , \14416 );
nor \U$14161 ( \14418 , \14403 , \14417 );
not \U$14162 ( \14419 , \14418 );
xnor \U$14163 ( \14420 , \14379 , \14419 );
buf g3855_GF_PartitionCandidate( \14421_nG3855 , \14420 );
buf \U$14164 ( \14422 , \14421_nG3855 );
not \U$14165 ( \14423 , \12105 );
nand \U$14166 ( \14424 , \13993 , \14423 );
nor \U$14167 ( \14425 , \14060 , \14019 );
nor \U$14168 ( \14426 , \14022 , \14026 );
nand \U$14169 ( \14427 , \14425 , \14426 );
nor \U$14170 ( \14428 , \14029 , \14034 );
nor \U$14171 ( \14429 , \14037 , \14041 );
nand \U$14172 ( \14430 , \14428 , \14429 );
nor \U$14173 ( \14431 , \14427 , \14430 );
nor \U$14174 ( \14432 , \14068 , \14050 );
nor \U$14175 ( \14433 , \14053 , \14057 );
nand \U$14176 ( \14434 , \14432 , \14433 );
nor \U$14177 ( \14435 , \14072 , \14065 );
and \U$14178 ( \14436 , \14435 , \14314 );
or \U$14179 ( \14437 , \14065 , \14079 );
nand \U$14180 ( \14438 , \14437 , \14087 );
nor \U$14181 ( \14439 , \14436 , \14438 );
or \U$14182 ( \14440 , \14434 , \14439 );
or \U$14183 ( \14441 , \14050 , \14094 );
nand \U$14184 ( \14442 , \14441 , \14103 );
and \U$14185 ( \14443 , \14433 , \14442 );
or \U$14186 ( \14444 , \14057 , \14110 );
nand \U$14187 ( \14445 , \14444 , \14118 );
nor \U$14188 ( \14446 , \14443 , \14445 );
nand \U$14189 ( \14447 , \14440 , \14446 );
and \U$14190 ( \14448 , \14431 , \14447 );
or \U$14191 ( \14449 , \14019 , \14125 );
nand \U$14192 ( \14450 , \14449 , \14135 );
and \U$14193 ( \14451 , \14426 , \14450 );
or \U$14194 ( \14452 , \14026 , \14142 );
nand \U$14195 ( \14453 , \14452 , \14150 );
nor \U$14196 ( \14454 , \14451 , \14453 );
or \U$14197 ( \14455 , \14430 , \14454 );
or \U$14198 ( \14456 , \14034 , \14157 );
nand \U$14199 ( \14457 , \14456 , \14166 );
and \U$14200 ( \14458 , \14429 , \14457 );
or \U$14201 ( \14459 , \14041 , \14173 );
nand \U$14202 ( \14460 , \14459 , \14181 );
nor \U$14203 ( \14461 , \14458 , \14460 );
nand \U$14204 ( \14462 , \14455 , \14461 );
nor \U$14205 ( \14463 , \14448 , \14462 );
not \U$14206 ( \14464 , \14463 );
xnor \U$14207 ( \14465 , \14424 , \14464 );
buf g3881_GF_PartitionCandidate( \14466_nG3881 , \14465 );
buf \U$14208 ( \14467 , \14466_nG3881 );
not \U$14209 ( \14468 , \12040 );
nand \U$14210 ( \14469 , \13991 , \14468 );
nor \U$14211 ( \14470 , \14218 , \14199 );
nor \U$14212 ( \14471 , \14200 , \14202 );
nand \U$14213 ( \14472 , \14470 , \14471 );
nor \U$14214 ( \14473 , \14203 , \14206 );
nor \U$14215 ( \14474 , \14207 , \14209 );
nand \U$14216 ( \14475 , \14473 , \14474 );
nor \U$14217 ( \14476 , \14472 , \14475 );
nor \U$14218 ( \14477 , \14222 , \14214 );
nor \U$14219 ( \14478 , \14215 , \14217 );
nand \U$14220 ( \14479 , \14477 , \14478 );
or \U$14221 ( \14480 , \14221 , \14225 );
nand \U$14222 ( \14481 , \14480 , \14229 );
not \U$14223 ( \14482 , \14481 );
or \U$14224 ( \14483 , \14479 , \14482 );
or \U$14225 ( \14484 , \14214 , \14232 );
nand \U$14226 ( \14485 , \14484 , \14237 );
and \U$14227 ( \14486 , \14478 , \14485 );
or \U$14228 ( \14487 , \14217 , \14240 );
nand \U$14229 ( \14488 , \14487 , \14244 );
nor \U$14230 ( \14489 , \14486 , \14488 );
nand \U$14231 ( \14490 , \14483 , \14489 );
and \U$14232 ( \14491 , \14476 , \14490 );
or \U$14233 ( \14492 , \14199 , \14247 );
nand \U$14234 ( \14493 , \14492 , \14253 );
and \U$14235 ( \14494 , \14471 , \14493 );
or \U$14236 ( \14495 , \14202 , \14256 );
nand \U$14237 ( \14496 , \14495 , \14260 );
nor \U$14238 ( \14497 , \14494 , \14496 );
or \U$14239 ( \14498 , \14475 , \14497 );
or \U$14240 ( \14499 , \14206 , \14263 );
nand \U$14241 ( \14500 , \14499 , \14268 );
and \U$14242 ( \14501 , \14474 , \14500 );
or \U$14243 ( \14502 , \14209 , \14271 );
nand \U$14244 ( \14503 , \14502 , \14275 );
nor \U$14245 ( \14504 , \14501 , \14503 );
nand \U$14246 ( \14505 , \14498 , \14504 );
nor \U$14247 ( \14506 , \14491 , \14505 );
not \U$14248 ( \14507 , \14506 );
xnor \U$14249 ( \14508 , \14469 , \14507 );
buf g38ab_GF_PartitionCandidate( \14509_nG38ab , \14508 );
buf \U$14250 ( \14510 , \14509_nG38ab );
not \U$14251 ( \14511 , \11941 );
nand \U$14252 ( \14512 , \13988 , \14511 );
nor \U$14253 ( \14513 , \14308 , \14289 );
nor \U$14254 ( \14514 , \14290 , \14292 );
nand \U$14255 ( \14515 , \14513 , \14514 );
nor \U$14256 ( \14516 , \14293 , \14296 );
nor \U$14257 ( \14517 , \14297 , \14299 );
nand \U$14258 ( \14518 , \14516 , \14517 );
nor \U$14259 ( \14519 , \14515 , \14518 );
nor \U$14260 ( \14520 , \14312 , \14304 );
nor \U$14261 ( \14521 , \14305 , \14307 );
nand \U$14262 ( \14522 , \14520 , \14521 );
or \U$14263 ( \14523 , \14311 , \14316 );
nand \U$14264 ( \14524 , \14523 , \14320 );
not \U$14265 ( \14525 , \14524 );
or \U$14266 ( \14526 , \14522 , \14525 );
or \U$14267 ( \14527 , \14304 , \14323 );
nand \U$14268 ( \14528 , \14527 , \14328 );
and \U$14269 ( \14529 , \14521 , \14528 );
or \U$14270 ( \14530 , \14307 , \14331 );
nand \U$14271 ( \14531 , \14530 , \14335 );
nor \U$14272 ( \14532 , \14529 , \14531 );
nand \U$14273 ( \14533 , \14526 , \14532 );
and \U$14274 ( \14534 , \14519 , \14533 );
or \U$14275 ( \14535 , \14289 , \14338 );
nand \U$14276 ( \14536 , \14535 , \14344 );
and \U$14277 ( \14537 , \14514 , \14536 );
or \U$14278 ( \14538 , \14292 , \14347 );
nand \U$14279 ( \14539 , \14538 , \14351 );
nor \U$14280 ( \14540 , \14537 , \14539 );
or \U$14281 ( \14541 , \14518 , \14540 );
or \U$14282 ( \14542 , \14296 , \14354 );
nand \U$14283 ( \14543 , \14542 , \14359 );
and \U$14284 ( \14544 , \14517 , \14543 );
or \U$14285 ( \14545 , \14299 , \14362 );
nand \U$14286 ( \14546 , \14545 , \14366 );
nor \U$14287 ( \14547 , \14544 , \14546 );
nand \U$14288 ( \14548 , \14541 , \14547 );
nor \U$14289 ( \14549 , \14534 , \14548 );
not \U$14290 ( \14550 , \14549 );
xnor \U$14291 ( \14551 , \14512 , \14550 );
buf g38d5_GF_PartitionCandidate( \14552_nG38d5 , \14551 );
buf \U$14292 ( \14553 , \14552_nG38d5 );
not \U$14293 ( \14554 , \11780 );
nand \U$14294 ( \14555 , \13986 , \14554 );
nand \U$14295 ( \14556 , \13513 , \9010 );
nand \U$14296 ( \14557 , \10313 , \11617 );
nor \U$14297 ( \14558 , \14556 , \14557 );
nand \U$14298 ( \14559 , \13768 , \13083 );
not \U$14299 ( \14560 , \13842 );
or \U$14300 ( \14561 , \14559 , \14560 );
and \U$14301 ( \14562 , \13083 , \13865 );
nor \U$14302 ( \14563 , \14562 , \13889 );
nand \U$14303 ( \14564 , \14561 , \14563 );
and \U$14304 ( \14565 , \14558 , \14564 );
and \U$14305 ( \14566 , \9010 , \13912 );
nor \U$14306 ( \14567 , \14566 , \13937 );
or \U$14307 ( \14568 , \14557 , \14567 );
and \U$14308 ( \14569 , \11617 , \13960 );
nor \U$14309 ( \14570 , \14569 , \13984 );
nand \U$14310 ( \14571 , \14568 , \14570 );
nor \U$14311 ( \14572 , \14565 , \14571 );
not \U$14312 ( \14573 , \14572 );
xnor \U$14313 ( \14574 , \14555 , \14573 );
buf g38eb_GF_PartitionCandidate( \14575_nG38eb , \14574 );
buf \U$14314 ( \14576 , \14575_nG38eb );
not \U$14315 ( \14577 , \11614 );
nand \U$14316 ( \14578 , \13981 , \14577 );
nand \U$14317 ( \14579 , \14061 , \14023 );
nand \U$14318 ( \14580 , \14030 , \14038 );
nor \U$14319 ( \14581 , \14579 , \14580 );
nand \U$14320 ( \14582 , \14069 , \14054 );
not \U$14321 ( \14583 , \14080 );
or \U$14322 ( \14584 , \14582 , \14583 );
and \U$14323 ( \14585 , \14054 , \14095 );
nor \U$14324 ( \14586 , \14585 , \14111 );
nand \U$14325 ( \14587 , \14584 , \14586 );
and \U$14326 ( \14588 , \14581 , \14587 );
and \U$14327 ( \14589 , \14023 , \14126 );
nor \U$14328 ( \14590 , \14589 , \14143 );
or \U$14329 ( \14591 , \14580 , \14590 );
and \U$14330 ( \14592 , \14038 , \14158 );
nor \U$14331 ( \14593 , \14592 , \14174 );
nand \U$14332 ( \14594 , \14591 , \14593 );
nor \U$14333 ( \14595 , \14588 , \14594 );
not \U$14334 ( \14596 , \14595 );
xnor \U$14335 ( \14597 , \14578 , \14596 );
buf g3901_GF_PartitionCandidate( \14598_nG3901 , \14597 );
buf \U$14336 ( \14599 , \14598_nG3901 );
not \U$14337 ( \14600 , \11453 );
nand \U$14338 ( \14601 , \13979 , \14600 );
nand \U$14339 ( \14602 , \14219 , \14201 );
nand \U$14340 ( \14603 , \14204 , \14208 );
nor \U$14341 ( \14604 , \14602 , \14603 );
nand \U$14342 ( \14605 , \14223 , \14216 );
or \U$14343 ( \14606 , \14605 , \14225 );
and \U$14344 ( \14607 , \14216 , \14233 );
nor \U$14345 ( \14608 , \14607 , \14241 );
nand \U$14346 ( \14609 , \14606 , \14608 );
and \U$14347 ( \14610 , \14604 , \14609 );
and \U$14348 ( \14611 , \14201 , \14248 );
nor \U$14349 ( \14612 , \14611 , \14257 );
or \U$14350 ( \14613 , \14603 , \14612 );
and \U$14351 ( \14614 , \14208 , \14264 );
nor \U$14352 ( \14615 , \14614 , \14272 );
nand \U$14353 ( \14616 , \14613 , \14615 );
nor \U$14354 ( \14617 , \14610 , \14616 );
not \U$14355 ( \14618 , \14617 );
xnor \U$14356 ( \14619 , \14601 , \14618 );
buf g3916_GF_PartitionCandidate( \14620_nG3916 , \14619 );
buf \U$14357 ( \14621 , \14620_nG3916 );
not \U$14358 ( \14622 , \11289 );
nand \U$14359 ( \14623 , \13976 , \14622 );
nand \U$14360 ( \14624 , \14309 , \14291 );
nand \U$14361 ( \14625 , \14294 , \14298 );
nor \U$14362 ( \14626 , \14624 , \14625 );
nand \U$14363 ( \14627 , \14313 , \14306 );
or \U$14364 ( \14628 , \14627 , \14316 );
and \U$14365 ( \14629 , \14306 , \14324 );
nor \U$14366 ( \14630 , \14629 , \14332 );
nand \U$14367 ( \14631 , \14628 , \14630 );
and \U$14368 ( \14632 , \14626 , \14631 );
and \U$14369 ( \14633 , \14291 , \14339 );
nor \U$14370 ( \14634 , \14633 , \14348 );
or \U$14371 ( \14635 , \14625 , \14634 );
and \U$14372 ( \14636 , \14298 , \14355 );
nor \U$14373 ( \14637 , \14636 , \14363 );
nand \U$14374 ( \14638 , \14635 , \14637 );
nor \U$14375 ( \14639 , \14632 , \14638 );
not \U$14376 ( \14640 , \14639 );
xnor \U$14377 ( \14641 , \14623 , \14640 );
buf g392b_GF_PartitionCandidate( \14642_nG392b , \14641 );
buf \U$14378 ( \14643 , \14642_nG392b );
not \U$14379 ( \14644 , \11128 );
nand \U$14380 ( \14645 , \13974 , \14644 );
nand \U$14381 ( \14646 , \14388 , \14380 );
nand \U$14382 ( \14647 , \14381 , \14383 );
nor \U$14383 ( \14648 , \14646 , \14647 );
nand \U$14384 ( \14649 , \14390 , \14387 );
or \U$14385 ( \14650 , \14649 , \13830 );
and \U$14386 ( \14651 , \14387 , \14393 );
nor \U$14387 ( \14652 , \14651 , \14397 );
nand \U$14388 ( \14653 , \14650 , \14652 );
and \U$14389 ( \14654 , \14648 , \14653 );
and \U$14390 ( \14655 , \14380 , \14400 );
nor \U$14391 ( \14656 , \14655 , \14405 );
or \U$14392 ( \14657 , \14647 , \14656 );
and \U$14393 ( \14658 , \14383 , \14408 );
nor \U$14394 ( \14659 , \14658 , \14412 );
nand \U$14395 ( \14660 , \14657 , \14659 );
nor \U$14396 ( \14661 , \14654 , \14660 );
not \U$14397 ( \14662 , \14661 );
xnor \U$14398 ( \14663 , \14645 , \14662 );
buf g3940_GF_PartitionCandidate( \14664_nG3940 , \14663 );
buf \U$14399 ( \14665 , \14664_nG3940 );
not \U$14400 ( \14666 , \10963 );
nand \U$14401 ( \14667 , \13970 , \14666 );
nand \U$14402 ( \14668 , \14433 , \14425 );
nand \U$14403 ( \14669 , \14426 , \14428 );
nor \U$14404 ( \14670 , \14668 , \14669 );
nand \U$14405 ( \14671 , \14435 , \14432 );
or \U$14406 ( \14672 , \14671 , \13826 );
and \U$14407 ( \14673 , \14432 , \14438 );
nor \U$14408 ( \14674 , \14673 , \14442 );
nand \U$14409 ( \14675 , \14672 , \14674 );
and \U$14410 ( \14676 , \14670 , \14675 );
and \U$14411 ( \14677 , \14425 , \14445 );
nor \U$14412 ( \14678 , \14677 , \14450 );
or \U$14413 ( \14679 , \14669 , \14678 );
and \U$14414 ( \14680 , \14428 , \14453 );
nor \U$14415 ( \14681 , \14680 , \14457 );
nand \U$14416 ( \14682 , \14679 , \14681 );
nor \U$14417 ( \14683 , \14676 , \14682 );
not \U$14418 ( \14684 , \14683 );
xnor \U$14419 ( \14685 , \14667 , \14684 );
buf g3955_GF_PartitionCandidate( \14686_nG3955 , \14685 );
buf \U$14420 ( \14687 , \14686_nG3955 );
not \U$14421 ( \14688 , \10802 );
nand \U$14422 ( \14689 , \13968 , \14688 );
nand \U$14423 ( \14690 , \14478 , \14470 );
nand \U$14424 ( \14691 , \14471 , \14473 );
nor \U$14425 ( \14692 , \14690 , \14691 );
and \U$14426 ( \14693 , \14477 , \14481 );
nor \U$14427 ( \14694 , \14693 , \14485 );
not \U$14428 ( \14695 , \14694 );
and \U$14429 ( \14696 , \14692 , \14695 );
and \U$14430 ( \14697 , \14470 , \14488 );
nor \U$14431 ( \14698 , \14697 , \14493 );
or \U$14432 ( \14699 , \14691 , \14698 );
and \U$14433 ( \14700 , \14473 , \14496 );
nor \U$14434 ( \14701 , \14700 , \14500 );
nand \U$14435 ( \14702 , \14699 , \14701 );
nor \U$14436 ( \14703 , \14696 , \14702 );
not \U$14437 ( \14704 , \14703 );
xnor \U$14438 ( \14705 , \14689 , \14704 );
buf g3968_GF_PartitionCandidate( \14706_nG3968 , \14705 );
buf \U$14439 ( \14707 , \14706_nG3968 );
not \U$14440 ( \14708 , \10638 );
nand \U$14441 ( \14709 , \13965 , \14708 );
nand \U$14442 ( \14710 , \14521 , \14513 );
nand \U$14443 ( \14711 , \14514 , \14516 );
nor \U$14444 ( \14712 , \14710 , \14711 );
and \U$14445 ( \14713 , \14520 , \14524 );
nor \U$14446 ( \14714 , \14713 , \14528 );
not \U$14447 ( \14715 , \14714 );
and \U$14448 ( \14716 , \14712 , \14715 );
and \U$14449 ( \14717 , \14513 , \14531 );
nor \U$14450 ( \14718 , \14717 , \14536 );
or \U$14451 ( \14719 , \14711 , \14718 );
and \U$14452 ( \14720 , \14516 , \14539 );
nor \U$14453 ( \14721 , \14720 , \14543 );
nand \U$14454 ( \14722 , \14719 , \14721 );
nor \U$14455 ( \14723 , \14716 , \14722 );
not \U$14456 ( \14724 , \14723 );
xnor \U$14457 ( \14725 , \14709 , \14724 );
buf g397b_GF_PartitionCandidate( \14726_nG397b , \14725 );
buf \U$14458 ( \14727 , \14726_nG397b );
not \U$14459 ( \14728 , \10477 );
nand \U$14460 ( \14729 , \13963 , \14728 );
nor \U$14461 ( \14730 , \13514 , \10314 );
not \U$14462 ( \14731 , \13866 );
and \U$14463 ( \14732 , \14730 , \14731 );
or \U$14464 ( \14733 , \10314 , \13913 );
nand \U$14465 ( \14734 , \14733 , \13961 );
nor \U$14466 ( \14735 , \14732 , \14734 );
not \U$14467 ( \14736 , \14735 );
xnor \U$14468 ( \14737 , \14729 , \14736 );
buf g3986_GF_PartitionCandidate( \14738_nG3986 , \14737 );
buf \U$14469 ( \14739 , \14738_nG3986 );
not \U$14470 ( \14740 , \10310 );
nand \U$14471 ( \14741 , \13957 , \14740 );
nor \U$14472 ( \14742 , \14062 , \14031 );
not \U$14473 ( \14743 , \14096 );
and \U$14474 ( \14744 , \14742 , \14743 );
or \U$14475 ( \14745 , \14031 , \14127 );
nand \U$14476 ( \14746 , \14745 , \14159 );
nor \U$14477 ( \14747 , \14744 , \14746 );
not \U$14478 ( \14748 , \14747 );
xnor \U$14479 ( \14749 , \14741 , \14748 );
buf g3991_GF_PartitionCandidate( \14750_nG3991 , \14749 );
buf \U$14480 ( \14751 , \14750_nG3991 );
not \U$14481 ( \14752 , \10149 );
nand \U$14482 ( \14753 , \13955 , \14752 );
nor \U$14483 ( \14754 , \14220 , \14205 );
not \U$14484 ( \14755 , \14234 );
and \U$14485 ( \14756 , \14754 , \14755 );
or \U$14486 ( \14757 , \14205 , \14249 );
nand \U$14487 ( \14758 , \14757 , \14265 );
nor \U$14488 ( \14759 , \14756 , \14758 );
not \U$14489 ( \14760 , \14759 );
xnor \U$14490 ( \14761 , \14753 , \14760 );
buf g399c_GF_PartitionCandidate( \14762_nG399c , \14761 );
buf \U$14491 ( \14763 , \14762_nG399c );
not \U$14492 ( \14764 , \9985 );
nand \U$14493 ( \14765 , \13952 , \14764 );
nor \U$14494 ( \14766 , \14310 , \14295 );
not \U$14495 ( \14767 , \14325 );
and \U$14496 ( \14768 , \14766 , \14767 );
or \U$14497 ( \14769 , \14295 , \14340 );
nand \U$14498 ( \14770 , \14769 , \14356 );
nor \U$14499 ( \14771 , \14768 , \14770 );
not \U$14500 ( \14772 , \14771 );
xnor \U$14501 ( \14773 , \14765 , \14772 );
buf g39a7_GF_PartitionCandidate( \14774_nG39a7 , \14773 );
buf \U$14502 ( \14775 , \14774_nG39a7 );
not \U$14503 ( \14776 , \9824 );
nand \U$14504 ( \14777 , \13950 , \14776 );
nor \U$14505 ( \14778 , \14389 , \14382 );
not \U$14506 ( \14779 , \14394 );
and \U$14507 ( \14780 , \14778 , \14779 );
or \U$14508 ( \14781 , \14382 , \14401 );
nand \U$14509 ( \14782 , \14781 , \14409 );
nor \U$14510 ( \14783 , \14780 , \14782 );
not \U$14511 ( \14784 , \14783 );
xnor \U$14512 ( \14785 , \14777 , \14784 );
buf g39b2_GF_PartitionCandidate( \14786_nG39b2 , \14785 );
buf \U$14513 ( \14787 , \14786_nG39b2 );
not \U$14514 ( \14788 , \9659 );
nand \U$14515 ( \14789 , \13946 , \14788 );
nor \U$14516 ( \14790 , \14434 , \14427 );
not \U$14517 ( \14791 , \14439 );
and \U$14518 ( \14792 , \14790 , \14791 );
or \U$14519 ( \14793 , \14427 , \14446 );
nand \U$14520 ( \14794 , \14793 , \14454 );
nor \U$14521 ( \14795 , \14792 , \14794 );
not \U$14522 ( \14796 , \14795 );
xnor \U$14523 ( \14797 , \14789 , \14796 );
buf g39bd_GF_PartitionCandidate( \14798_nG39bd , \14797 );
buf \U$14524 ( \14799 , \14798_nG39bd );
not \U$14525 ( \14800 , \9498 );
nand \U$14526 ( \14801 , \13944 , \14800 );
nor \U$14527 ( \14802 , \14479 , \14472 );
and \U$14528 ( \14803 , \14802 , \14481 );
or \U$14529 ( \14804 , \14472 , \14489 );
nand \U$14530 ( \14805 , \14804 , \14497 );
nor \U$14531 ( \14806 , \14803 , \14805 );
not \U$14532 ( \14807 , \14806 );
xnor \U$14533 ( \14808 , \14801 , \14807 );
buf g39c7_GF_PartitionCandidate( \14809_nG39c7 , \14808 );
buf \U$14534 ( \14810 , \14809_nG39c7 );
not \U$14535 ( \14811 , \9334 );
nand \U$14536 ( \14812 , \13941 , \14811 );
nor \U$14537 ( \14813 , \14522 , \14515 );
and \U$14538 ( \14814 , \14813 , \14524 );
or \U$14539 ( \14815 , \14515 , \14532 );
nand \U$14540 ( \14816 , \14815 , \14540 );
nor \U$14541 ( \14817 , \14814 , \14816 );
not \U$14542 ( \14818 , \14817 );
xnor \U$14543 ( \14819 , \14812 , \14818 );
buf g39d1_GF_PartitionCandidate( \14820_nG39d1 , \14819 );
buf \U$14544 ( \14821 , \14820_nG39d1 );
not \U$14545 ( \14822 , \9173 );
nand \U$14546 ( \14823 , \13939 , \14822 );
nor \U$14547 ( \14824 , \14559 , \14556 );
and \U$14548 ( \14825 , \14824 , \13842 );
or \U$14549 ( \14826 , \14556 , \14563 );
nand \U$14550 ( \14827 , \14826 , \14567 );
nor \U$14551 ( \14828 , \14825 , \14827 );
not \U$14552 ( \14829 , \14828 );
xnor \U$14553 ( \14830 , \14823 , \14829 );
buf g39db_GF_PartitionCandidate( \14831_nG39db , \14830 );
buf \U$14554 ( \14832 , \14831_nG39db );
not \U$14555 ( \14833 , \9007 );
nand \U$14556 ( \14834 , \13934 , \14833 );
nor \U$14557 ( \14835 , \14582 , \14579 );
and \U$14558 ( \14836 , \14835 , \14080 );
or \U$14559 ( \14837 , \14579 , \14586 );
nand \U$14560 ( \14838 , \14837 , \14590 );
nor \U$14561 ( \14839 , \14836 , \14838 );
not \U$14562 ( \14840 , \14839 );
xnor \U$14563 ( \14841 , \14834 , \14840 );
buf g39e5_GF_PartitionCandidate( \14842_nG39e5 , \14841 );
buf \U$14564 ( \14843 , \14842_nG39e5 );
not \U$14565 ( \14844 , \8846 );
nand \U$14566 ( \14845 , \13932 , \14844 );
nor \U$14567 ( \14846 , \14605 , \14602 );
and \U$14568 ( \14847 , \14846 , \14226 );
or \U$14569 ( \14848 , \14602 , \14608 );
nand \U$14570 ( \14849 , \14848 , \14612 );
nor \U$14571 ( \14850 , \14847 , \14849 );
not \U$14572 ( \14851 , \14850 );
xnor \U$14573 ( \14852 , \14845 , \14851 );
buf g39ef_GF_PartitionCandidate( \14853_nG39ef , \14852 );
buf \U$14574 ( \14854 , \14853_nG39ef );
not \U$14575 ( \14855 , \8682 );
nand \U$14576 ( \14856 , \13929 , \14855 );
nor \U$14577 ( \14857 , \14627 , \14624 );
and \U$14578 ( \14858 , \14857 , \14317 );
or \U$14579 ( \14859 , \14624 , \14630 );
nand \U$14580 ( \14860 , \14859 , \14634 );
nor \U$14581 ( \14861 , \14858 , \14860 );
not \U$14582 ( \14862 , \14861 );
xnor \U$14583 ( \14863 , \14856 , \14862 );
buf g39f9_GF_PartitionCandidate( \14864_nG39f9 , \14863 );
buf \U$14584 ( \14865 , \14864_nG39f9 );
not \U$14585 ( \14866 , \8521 );
nand \U$14586 ( \14867 , \13927 , \14866 );
nor \U$14587 ( \14868 , \14649 , \14646 );
and \U$14588 ( \14869 , \14868 , \13829 );
or \U$14589 ( \14870 , \14646 , \14652 );
nand \U$14590 ( \14871 , \14870 , \14656 );
nor \U$14591 ( \14872 , \14869 , \14871 );
not \U$14592 ( \14873 , \14872 );
xnor \U$14593 ( \14874 , \14867 , \14873 );
buf g3a03_GF_PartitionCandidate( \14875_nG3a03 , \14874 );
buf \U$14594 ( \14876 , \14875_nG3a03 );
not \U$14595 ( \14877 , \8359 );
nand \U$14596 ( \14878 , \13923 , \14877 );
nor \U$14597 ( \14879 , \14671 , \14668 );
and \U$14598 ( \14880 , \14879 , \14314 );
or \U$14599 ( \14881 , \14668 , \14674 );
nand \U$14600 ( \14882 , \14881 , \14678 );
nor \U$14601 ( \14883 , \14880 , \14882 );
not \U$14602 ( \14884 , \14883 );
xnor \U$14603 ( \14885 , \14878 , \14884 );
buf g3a0d_GF_PartitionCandidate( \14886_nG3a0d , \14885 );
buf \U$14604 ( \14887 , \14886_nG3a0d );
not \U$14605 ( \14888 , \8200 );
nand \U$14606 ( \14889 , \13921 , \14888 );
or \U$14607 ( \14890 , \14690 , \14694 );
nand \U$14608 ( \14891 , \14890 , \14698 );
xnor \U$14609 ( \14892 , \14889 , \14891 );
buf g3a13_GF_PartitionCandidate( \14893_nG3a13 , \14892 );
buf \U$14610 ( \14894 , \14893_nG3a13 );
not \U$14611 ( \14895 , \8041 );
nand \U$14612 ( \14896 , \13918 , \14895 );
or \U$14613 ( \14897 , \14710 , \14714 );
nand \U$14614 ( \14898 , \14897 , \14718 );
xnor \U$14615 ( \14899 , \14896 , \14898 );
buf g3a19_GF_PartitionCandidate( \14900_nG3a19 , \14899 );
buf \U$14616 ( \14901 , \14900_nG3a19 );
not \U$14617 ( \14902 , \7887 );
nand \U$14618 ( \14903 , \13916 , \14902 );
xnor \U$14619 ( \14904 , \14903 , \13914 );
buf g3a1d_GF_PartitionCandidate( \14905_nG3a1d , \14904 );
buf \U$14620 ( \14906 , \14905_nG3a1d );
not \U$14621 ( \14907 , \13510 );
nand \U$14622 ( \14908 , \13909 , \14907 );
xnor \U$14623 ( \14909 , \14908 , \14128 );
buf g3a21_GF_PartitionCandidate( \14910_nG3a21 , \14909 );
buf \U$14624 ( \14911 , \14910_nG3a21 );
not \U$14625 ( \14912 , \13503 );
nand \U$14626 ( \14913 , \13907 , \14912 );
xnor \U$14627 ( \14914 , \14913 , \14250 );
buf g3a25_GF_PartitionCandidate( \14915_nG3a25 , \14914 );
buf \U$14628 ( \14916 , \14915_nG3a25 );
not \U$14629 ( \14917 , \13488 );
nand \U$14630 ( \14918 , \13904 , \14917 );
xnor \U$14631 ( \14919 , \14918 , \14341 );
buf g3a29_GF_PartitionCandidate( \14920_nG3a29 , \14919 );
buf \U$14632 ( \14921 , \14920_nG3a29 );
not \U$14633 ( \14922 , \13463 );
nand \U$14634 ( \14923 , \13902 , \14922 );
xnor \U$14635 ( \14924 , \14923 , \14402 );
buf g3a2d_GF_PartitionCandidate( \14925_nG3a2d , \14924 );
buf \U$14636 ( \14926 , \14925_nG3a2d );
not \U$14637 ( \14927 , \13428 );
nand \U$14638 ( \14928 , \13898 , \14927 );
xnor \U$14639 ( \14929 , \14928 , \14447 );
buf g3a31_GF_PartitionCandidate( \14930_nG3a31 , \14929 );
buf \U$14640 ( \14931 , \14930_nG3a31 );
not \U$14641 ( \14932 , \13383 );
nand \U$14642 ( \14933 , \13896 , \14932 );
xnor \U$14643 ( \14934 , \14933 , \14490 );
buf g3a35_GF_PartitionCandidate( \14935_nG3a35 , \14934 );
buf \U$14644 ( \14936 , \14935_nG3a35 );
not \U$14645 ( \14937 , \13309 );
nand \U$14646 ( \14938 , \13893 , \14937 );
xnor \U$14647 ( \14939 , \14938 , \14533 );
buf g3a39_GF_PartitionCandidate( \14940_nG3a39 , \14939 );
buf \U$14648 ( \14941 , \14940_nG3a39 );
not \U$14649 ( \14942 , \13194 );
nand \U$14650 ( \14943 , \13891 , \14942 );
xnor \U$14651 ( \14944 , \14943 , \14564 );
buf g3a3d_GF_PartitionCandidate( \14945_nG3a3d , \14944 );
buf \U$14652 ( \14946 , \14945_nG3a3d );
not \U$14653 ( \14947 , \13080 );
nand \U$14654 ( \14948 , \13886 , \14947 );
xnor \U$14655 ( \14949 , \14948 , \14587 );
buf g3a41_GF_PartitionCandidate( \14950_nG3a41 , \14949 );
buf \U$14656 ( \14951 , \14950_nG3a41 );
not \U$14657 ( \14952 , \12975 );
nand \U$14658 ( \14953 , \13884 , \14952 );
xnor \U$14659 ( \14954 , \14953 , \14609 );
buf g3a45_GF_PartitionCandidate( \14955_nG3a45 , \14954 );
buf \U$14660 ( \14956 , \14955_nG3a45 );
not \U$14661 ( \14957 , \12873 );
nand \U$14662 ( \14958 , \13881 , \14957 );
xnor \U$14663 ( \14959 , \14958 , \14631 );
buf g3a49_GF_PartitionCandidate( \14960_nG3a49 , \14959 );
buf \U$14664 ( \14961 , \14960_nG3a49 );
not \U$14665 ( \14962 , \12778 );
nand \U$14666 ( \14963 , \13879 , \14962 );
xnor \U$14667 ( \14964 , \14963 , \14653 );
buf g3a4d_GF_PartitionCandidate( \14965_nG3a4d , \14964 );
buf \U$14668 ( \14966 , \14965_nG3a4d );
not \U$14669 ( \14967 , \12685 );
nand \U$14670 ( \14968 , \13875 , \14967 );
xnor \U$14671 ( \14969 , \14968 , \14675 );
buf g3a51_GF_PartitionCandidate( \14970_nG3a51 , \14969 );
buf \U$14672 ( \14971 , \14970_nG3a51 );
not \U$14673 ( \14972 , \12600 );
nand \U$14674 ( \14973 , \13873 , \14972 );
xnor \U$14675 ( \14974 , \14973 , \14695 );
buf g3a55_GF_PartitionCandidate( \14975_nG3a55 , \14974 );
buf \U$14676 ( \14976 , \14975_nG3a55 );
not \U$14677 ( \14977 , \12518 );
nand \U$14678 ( \14978 , \13870 , \14977 );
xnor \U$14679 ( \14979 , \14978 , \14715 );
buf g3a59_GF_PartitionCandidate( \14980_nG3a59 , \14979 );
buf \U$14680 ( \14981 , \14980_nG3a59 );
not \U$14681 ( \14982 , \12443 );
nand \U$14682 ( \14983 , \13868 , \14982 );
xnor \U$14683 ( \14984 , \14983 , \14731 );
buf g3a5d_GF_PartitionCandidate( \14985_nG3a5d , \14984 );
buf \U$14684 ( \14986 , \14985_nG3a5d );
not \U$14685 ( \14987 , \13765 );
nand \U$14686 ( \14988 , \13862 , \14987 );
xnor \U$14687 ( \14989 , \14988 , \14743 );
buf g3a61_GF_PartitionCandidate( \14990_nG3a61 , \14989 );
buf \U$14688 ( \14991 , \14990_nG3a61 );
not \U$14689 ( \14992 , \13758 );
nand \U$14690 ( \14993 , \13860 , \14992 );
xnor \U$14691 ( \14994 , \14993 , \14755 );
buf g3a65_GF_PartitionCandidate( \14995_nG3a65 , \14994 );
buf \U$14692 ( \14996 , \14995_nG3a65 );
not \U$14693 ( \14997 , \13746 );
nand \U$14694 ( \14998 , \13857 , \14997 );
xnor \U$14695 ( \14999 , \14998 , \14767 );
buf g3a69_GF_PartitionCandidate( \15000_nG3a69 , \14999 );
buf \U$14696 ( \15001 , \15000_nG3a69 );
not \U$14697 ( \15002 , \13729 );
nand \U$14698 ( \15003 , \13855 , \15002 );
xnor \U$14699 ( \15004 , \15003 , \14779 );
buf g3a6d_GF_PartitionCandidate( \15005_nG3a6d , \15004 );
buf \U$14700 ( \15006 , \15005_nG3a6d );
not \U$14701 ( \15007 , \13700 );
nand \U$14702 ( \15008 , \13851 , \15007 );
xnor \U$14703 ( \15009 , \15008 , \14791 );
buf g3a71_GF_PartitionCandidate( \15010_nG3a71 , \15009 );
buf \U$14704 ( \15011 , \15010_nG3a71 );
not \U$14705 ( \15012 , \13655 );
nand \U$14706 ( \15013 , \13849 , \15012 );
xnor \U$14707 ( \15014 , \15013 , \14481 );
buf g3a75_GF_PartitionCandidate( \15015_nG3a75 , \15014 );
buf \U$14708 ( \15016 , \15015_nG3a75 );
not \U$14709 ( \15017 , \13613 );
nand \U$14710 ( \15018 , \13846 , \15017 );
xnor \U$14711 ( \15019 , \15018 , \14524 );
buf g3a79_GF_PartitionCandidate( \15020_nG3a79 , \15019 );
buf \U$14712 ( \15021 , \15020_nG3a79 );
not \U$14713 ( \15022 , \13578 );
nand \U$14714 ( \15023 , \13844 , \15022 );
xnor \U$14715 ( \15024 , \15023 , \13842 );
buf g3a7d_GF_PartitionCandidate( \15025_nG3a7d , \15024 );
buf \U$14716 ( \15026 , \15025_nG3a7d );
not \U$14717 ( \15027 , \13812 );
nand \U$14718 ( \15028 , \13839 , \15027 );
xnor \U$14719 ( \15029 , \15028 , \14080 );
buf g3a81_GF_PartitionCandidate( \15030_nG3a81 , \15029 );
buf \U$14720 ( \15031 , \15030_nG3a81 );
endmodule

